VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_devinatkin_dual_oscillator
  CLASS BLOCK ;
  FOREIGN tt_um_devinatkin_dual_oscillator ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 93.243820 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 19.610 12.575 23.390 143.370 ;
      LAYER nwell ;
        RECT 23.390 53.000 32.290 143.370 ;
      LAYER pwell ;
        RECT 32.290 53.000 36.070 143.370 ;
      LAYER nwell ;
        RECT 23.390 12.575 27.840 53.000 ;
      LAYER li1 ;
        RECT 23.680 143.190 24.480 143.200 ;
        RECT 31.200 143.190 32.000 143.200 ;
        RECT 19.720 143.020 23.220 143.190 ;
        RECT 19.710 143.010 23.220 143.020 ;
        RECT 19.710 141.910 19.890 143.010 ;
        RECT 19.720 139.190 19.890 141.910 ;
        RECT 20.290 141.720 21.290 141.890 ;
        RECT 21.580 141.720 22.580 141.890 ;
        RECT 20.060 140.510 20.230 141.550 ;
        RECT 21.350 140.510 21.520 141.550 ;
        RECT 22.640 140.510 22.810 141.550 ;
        RECT 20.290 140.170 21.290 140.340 ;
        RECT 21.580 140.170 22.580 140.340 ;
        RECT 23.050 139.190 23.220 143.010 ;
        RECT 19.720 139.020 23.220 139.190 ;
        RECT 19.710 138.920 23.220 139.020 ;
        RECT 19.710 137.910 19.890 138.920 ;
        RECT 19.720 135.130 19.890 137.910 ;
        RECT 20.290 137.720 21.290 137.890 ;
        RECT 21.580 137.720 22.580 137.890 ;
        RECT 20.060 136.510 20.230 137.550 ;
        RECT 21.350 136.510 21.520 137.550 ;
        RECT 22.640 136.510 22.810 137.550 ;
        RECT 20.290 136.170 21.290 136.340 ;
        RECT 21.580 136.170 22.580 136.340 ;
        RECT 23.050 135.130 23.220 138.920 ;
        RECT 19.720 134.920 23.220 135.130 ;
        RECT 19.710 134.910 23.220 134.920 ;
        RECT 19.710 133.810 19.890 134.910 ;
        RECT 19.720 131.040 19.890 133.810 ;
        RECT 20.290 133.620 21.290 133.790 ;
        RECT 21.580 133.620 22.580 133.790 ;
        RECT 20.060 132.410 20.230 133.450 ;
        RECT 21.350 132.410 21.520 133.450 ;
        RECT 22.640 132.410 22.810 133.450 ;
        RECT 20.290 132.070 21.290 132.240 ;
        RECT 21.580 132.070 22.580 132.240 ;
        RECT 23.050 131.040 23.220 134.910 ;
        RECT 19.720 130.870 23.220 131.040 ;
        RECT 19.710 130.820 23.220 130.870 ;
        RECT 19.710 129.760 19.890 130.820 ;
        RECT 19.720 126.990 19.890 129.760 ;
        RECT 20.290 129.570 21.290 129.740 ;
        RECT 21.580 129.570 22.580 129.740 ;
        RECT 20.060 128.360 20.230 129.400 ;
        RECT 21.350 128.360 21.520 129.400 ;
        RECT 22.640 128.360 22.810 129.400 ;
        RECT 20.290 128.020 21.290 128.190 ;
        RECT 21.580 128.020 22.580 128.190 ;
        RECT 23.050 126.990 23.220 130.820 ;
        RECT 19.720 126.820 23.220 126.990 ;
        RECT 19.710 126.770 23.220 126.820 ;
        RECT 19.710 125.710 19.890 126.770 ;
        RECT 19.720 122.940 19.890 125.710 ;
        RECT 20.290 125.520 21.290 125.690 ;
        RECT 21.580 125.520 22.580 125.690 ;
        RECT 20.060 124.310 20.230 125.350 ;
        RECT 21.350 124.310 21.520 125.350 ;
        RECT 22.640 124.310 22.810 125.350 ;
        RECT 20.290 123.970 21.290 124.140 ;
        RECT 21.580 123.970 22.580 124.140 ;
        RECT 23.050 122.940 23.220 126.770 ;
        RECT 19.720 122.770 23.220 122.940 ;
        RECT 19.710 122.720 23.220 122.770 ;
        RECT 19.710 121.660 19.890 122.720 ;
        RECT 19.720 118.890 19.890 121.660 ;
        RECT 20.290 121.470 21.290 121.640 ;
        RECT 21.580 121.470 22.580 121.640 ;
        RECT 20.060 120.260 20.230 121.300 ;
        RECT 21.350 120.260 21.520 121.300 ;
        RECT 22.640 120.260 22.810 121.300 ;
        RECT 20.290 119.920 21.290 120.090 ;
        RECT 21.580 119.920 22.580 120.090 ;
        RECT 23.050 118.890 23.220 122.720 ;
        RECT 19.720 118.720 23.220 118.890 ;
        RECT 19.710 118.670 23.220 118.720 ;
        RECT 19.710 117.610 19.890 118.670 ;
        RECT 19.720 114.840 19.890 117.610 ;
        RECT 20.290 117.420 21.290 117.590 ;
        RECT 21.580 117.420 22.580 117.590 ;
        RECT 20.060 116.210 20.230 117.250 ;
        RECT 21.350 116.210 21.520 117.250 ;
        RECT 22.640 116.210 22.810 117.250 ;
        RECT 20.290 115.870 21.290 116.040 ;
        RECT 21.580 115.870 22.580 116.040 ;
        RECT 23.050 114.840 23.220 118.670 ;
        RECT 19.720 114.670 23.220 114.840 ;
        RECT 19.710 114.620 23.220 114.670 ;
        RECT 19.710 113.560 19.890 114.620 ;
        RECT 19.720 110.790 19.890 113.560 ;
        RECT 20.290 113.370 21.290 113.540 ;
        RECT 21.580 113.370 22.580 113.540 ;
        RECT 20.060 112.160 20.230 113.200 ;
        RECT 21.350 112.160 21.520 113.200 ;
        RECT 22.640 112.160 22.810 113.200 ;
        RECT 20.290 111.820 21.290 111.990 ;
        RECT 21.580 111.820 22.580 111.990 ;
        RECT 23.050 110.790 23.220 114.620 ;
        RECT 19.720 110.620 23.220 110.790 ;
        RECT 19.710 110.570 23.220 110.620 ;
        RECT 19.710 109.510 19.890 110.570 ;
        RECT 19.720 106.740 19.890 109.510 ;
        RECT 20.290 109.320 21.290 109.490 ;
        RECT 21.580 109.320 22.580 109.490 ;
        RECT 20.060 108.110 20.230 109.150 ;
        RECT 21.350 108.110 21.520 109.150 ;
        RECT 22.640 108.110 22.810 109.150 ;
        RECT 20.290 107.770 21.290 107.940 ;
        RECT 21.580 107.770 22.580 107.940 ;
        RECT 23.050 106.740 23.220 110.570 ;
        RECT 19.720 106.570 23.220 106.740 ;
        RECT 19.710 106.520 23.220 106.570 ;
        RECT 19.710 105.460 19.890 106.520 ;
        RECT 19.720 102.690 19.890 105.460 ;
        RECT 20.290 105.270 21.290 105.440 ;
        RECT 21.580 105.270 22.580 105.440 ;
        RECT 20.060 104.060 20.230 105.100 ;
        RECT 21.350 104.060 21.520 105.100 ;
        RECT 22.640 104.060 22.810 105.100 ;
        RECT 20.290 103.720 21.290 103.890 ;
        RECT 21.580 103.720 22.580 103.890 ;
        RECT 23.050 102.690 23.220 106.520 ;
        RECT 19.720 102.520 23.220 102.690 ;
        RECT 19.710 102.470 23.220 102.520 ;
        RECT 19.710 101.410 19.890 102.470 ;
        RECT 19.720 98.640 19.890 101.410 ;
        RECT 20.290 101.220 21.290 101.390 ;
        RECT 21.580 101.220 22.580 101.390 ;
        RECT 20.060 100.010 20.230 101.050 ;
        RECT 21.350 100.010 21.520 101.050 ;
        RECT 22.640 100.010 22.810 101.050 ;
        RECT 20.290 99.670 21.290 99.840 ;
        RECT 21.580 99.670 22.580 99.840 ;
        RECT 23.050 98.640 23.220 102.470 ;
        RECT 19.720 98.470 23.220 98.640 ;
        RECT 19.710 98.420 23.220 98.470 ;
        RECT 19.710 97.360 19.890 98.420 ;
        RECT 19.720 94.590 19.890 97.360 ;
        RECT 20.290 97.170 21.290 97.340 ;
        RECT 21.580 97.170 22.580 97.340 ;
        RECT 20.060 95.960 20.230 97.000 ;
        RECT 21.350 95.960 21.520 97.000 ;
        RECT 22.640 95.960 22.810 97.000 ;
        RECT 20.290 95.620 21.290 95.790 ;
        RECT 21.580 95.620 22.580 95.790 ;
        RECT 23.050 94.590 23.220 98.420 ;
        RECT 19.720 94.420 23.220 94.590 ;
        RECT 19.710 94.370 23.220 94.420 ;
        RECT 19.710 93.310 19.890 94.370 ;
        RECT 19.720 90.540 19.890 93.310 ;
        RECT 20.290 93.120 21.290 93.290 ;
        RECT 21.580 93.120 22.580 93.290 ;
        RECT 20.060 91.910 20.230 92.950 ;
        RECT 21.350 91.910 21.520 92.950 ;
        RECT 22.640 91.910 22.810 92.950 ;
        RECT 20.290 91.570 21.290 91.740 ;
        RECT 21.580 91.570 22.580 91.740 ;
        RECT 23.050 90.540 23.220 94.370 ;
        RECT 19.720 90.370 23.220 90.540 ;
        RECT 19.710 90.320 23.220 90.370 ;
        RECT 19.710 89.260 19.890 90.320 ;
        RECT 19.720 86.490 19.890 89.260 ;
        RECT 20.290 89.070 21.290 89.240 ;
        RECT 21.580 89.070 22.580 89.240 ;
        RECT 20.060 87.860 20.230 88.900 ;
        RECT 21.350 87.860 21.520 88.900 ;
        RECT 22.640 87.860 22.810 88.900 ;
        RECT 20.290 87.520 21.290 87.690 ;
        RECT 21.580 87.520 22.580 87.690 ;
        RECT 23.050 86.490 23.220 90.320 ;
        RECT 19.720 86.320 23.220 86.490 ;
        RECT 19.710 86.270 23.220 86.320 ;
        RECT 19.710 85.210 19.890 86.270 ;
        RECT 19.720 82.440 19.890 85.210 ;
        RECT 20.290 85.020 21.290 85.190 ;
        RECT 21.580 85.020 22.580 85.190 ;
        RECT 20.060 83.810 20.230 84.850 ;
        RECT 21.350 83.810 21.520 84.850 ;
        RECT 22.640 83.810 22.810 84.850 ;
        RECT 20.290 83.470 21.290 83.640 ;
        RECT 21.580 83.470 22.580 83.640 ;
        RECT 23.050 82.440 23.220 86.270 ;
        RECT 19.720 82.270 23.220 82.440 ;
        RECT 19.710 82.220 23.220 82.270 ;
        RECT 19.710 81.160 19.890 82.220 ;
        RECT 19.720 78.390 19.890 81.160 ;
        RECT 20.290 80.970 21.290 81.140 ;
        RECT 21.580 80.970 22.580 81.140 ;
        RECT 20.060 79.760 20.230 80.800 ;
        RECT 21.350 79.760 21.520 80.800 ;
        RECT 22.640 79.760 22.810 80.800 ;
        RECT 20.290 79.420 21.290 79.590 ;
        RECT 21.580 79.420 22.580 79.590 ;
        RECT 23.050 78.390 23.220 82.220 ;
        RECT 19.720 78.220 23.220 78.390 ;
        RECT 19.710 78.170 23.220 78.220 ;
        RECT 19.710 77.110 19.890 78.170 ;
        RECT 19.720 74.340 19.890 77.110 ;
        RECT 20.290 76.920 21.290 77.090 ;
        RECT 21.580 76.920 22.580 77.090 ;
        RECT 20.060 75.710 20.230 76.750 ;
        RECT 21.350 75.710 21.520 76.750 ;
        RECT 22.640 75.710 22.810 76.750 ;
        RECT 20.290 75.370 21.290 75.540 ;
        RECT 21.580 75.370 22.580 75.540 ;
        RECT 23.050 74.340 23.220 78.170 ;
        RECT 19.720 74.170 23.220 74.340 ;
        RECT 19.710 74.120 23.220 74.170 ;
        RECT 19.710 73.060 19.890 74.120 ;
        RECT 19.720 70.290 19.890 73.060 ;
        RECT 20.290 72.870 21.290 73.040 ;
        RECT 21.580 72.870 22.580 73.040 ;
        RECT 20.060 71.660 20.230 72.700 ;
        RECT 21.350 71.660 21.520 72.700 ;
        RECT 22.640 71.660 22.810 72.700 ;
        RECT 20.290 71.320 21.290 71.490 ;
        RECT 21.580 71.320 22.580 71.490 ;
        RECT 23.050 70.290 23.220 74.120 ;
        RECT 19.720 70.120 23.220 70.290 ;
        RECT 19.710 70.070 23.220 70.120 ;
        RECT 19.710 69.010 19.890 70.070 ;
        RECT 19.720 66.240 19.890 69.010 ;
        RECT 20.290 68.820 21.290 68.990 ;
        RECT 21.580 68.820 22.580 68.990 ;
        RECT 20.060 67.610 20.230 68.650 ;
        RECT 21.350 67.610 21.520 68.650 ;
        RECT 22.640 67.610 22.810 68.650 ;
        RECT 20.290 67.270 21.290 67.440 ;
        RECT 21.580 67.270 22.580 67.440 ;
        RECT 23.050 66.240 23.220 70.070 ;
        RECT 19.720 66.070 23.220 66.240 ;
        RECT 19.710 66.020 23.220 66.070 ;
        RECT 19.710 64.960 19.890 66.020 ;
        RECT 19.720 62.190 19.890 64.960 ;
        RECT 20.290 64.770 21.290 64.940 ;
        RECT 21.580 64.770 22.580 64.940 ;
        RECT 20.060 63.560 20.230 64.600 ;
        RECT 21.350 63.560 21.520 64.600 ;
        RECT 22.640 63.560 22.810 64.600 ;
        RECT 20.290 63.220 21.290 63.390 ;
        RECT 21.580 63.220 22.580 63.390 ;
        RECT 23.050 62.190 23.220 66.020 ;
        RECT 19.720 62.020 23.220 62.190 ;
        RECT 19.710 61.970 23.220 62.020 ;
        RECT 19.710 60.910 19.890 61.970 ;
        RECT 19.720 58.140 19.890 60.910 ;
        RECT 20.290 60.720 21.290 60.890 ;
        RECT 21.580 60.720 22.580 60.890 ;
        RECT 20.060 59.510 20.230 60.550 ;
        RECT 21.350 59.510 21.520 60.550 ;
        RECT 22.640 59.510 22.810 60.550 ;
        RECT 20.290 59.170 21.290 59.340 ;
        RECT 21.580 59.170 22.580 59.340 ;
        RECT 23.050 58.140 23.220 61.970 ;
        RECT 19.720 57.970 23.220 58.140 ;
        RECT 19.710 57.920 23.220 57.970 ;
        RECT 19.710 56.860 19.890 57.920 ;
        RECT 19.720 54.090 19.890 56.860 ;
        RECT 20.290 56.670 21.290 56.840 ;
        RECT 21.580 56.670 22.580 56.840 ;
        RECT 20.060 55.460 20.230 56.500 ;
        RECT 21.350 55.460 21.520 56.500 ;
        RECT 22.640 55.460 22.810 56.500 ;
        RECT 20.290 55.120 21.290 55.290 ;
        RECT 21.580 55.120 22.580 55.290 ;
        RECT 23.050 54.090 23.220 57.920 ;
        RECT 19.720 53.920 23.220 54.090 ;
        RECT 19.710 53.870 23.220 53.920 ;
        RECT 19.710 52.810 19.890 53.870 ;
        RECT 19.720 50.040 19.890 52.810 ;
        RECT 20.290 52.620 21.290 52.790 ;
        RECT 21.580 52.620 22.580 52.790 ;
        RECT 20.060 51.410 20.230 52.450 ;
        RECT 21.350 51.410 21.520 52.450 ;
        RECT 22.640 51.410 22.810 52.450 ;
        RECT 20.290 51.070 21.290 51.240 ;
        RECT 21.580 51.070 22.580 51.240 ;
        RECT 23.050 50.040 23.220 53.870 ;
        RECT 19.720 49.870 23.220 50.040 ;
        RECT 19.710 49.820 23.220 49.870 ;
        RECT 19.710 48.760 19.890 49.820 ;
        RECT 19.720 45.990 19.890 48.760 ;
        RECT 20.290 48.570 21.290 48.740 ;
        RECT 21.580 48.570 22.580 48.740 ;
        RECT 20.060 47.360 20.230 48.400 ;
        RECT 21.350 47.360 21.520 48.400 ;
        RECT 22.640 47.360 22.810 48.400 ;
        RECT 20.290 47.020 21.290 47.190 ;
        RECT 21.580 47.020 22.580 47.190 ;
        RECT 23.050 45.990 23.220 49.820 ;
        RECT 19.720 45.820 23.220 45.990 ;
        RECT 19.710 45.770 23.220 45.820 ;
        RECT 19.710 44.710 19.890 45.770 ;
        RECT 19.720 41.940 19.890 44.710 ;
        RECT 20.290 44.520 21.290 44.690 ;
        RECT 21.580 44.520 22.580 44.690 ;
        RECT 20.060 43.310 20.230 44.350 ;
        RECT 21.350 43.310 21.520 44.350 ;
        RECT 22.640 43.310 22.810 44.350 ;
        RECT 20.290 42.970 21.290 43.140 ;
        RECT 21.580 42.970 22.580 43.140 ;
        RECT 23.050 41.940 23.220 45.770 ;
        RECT 19.720 41.770 23.220 41.940 ;
        RECT 19.710 41.720 23.220 41.770 ;
        RECT 19.710 40.660 19.890 41.720 ;
        RECT 19.720 37.890 19.890 40.660 ;
        RECT 20.290 40.470 21.290 40.640 ;
        RECT 21.580 40.470 22.580 40.640 ;
        RECT 20.060 39.260 20.230 40.300 ;
        RECT 21.350 39.260 21.520 40.300 ;
        RECT 22.640 39.260 22.810 40.300 ;
        RECT 20.290 38.920 21.290 39.090 ;
        RECT 21.580 38.920 22.580 39.090 ;
        RECT 23.050 37.890 23.220 41.720 ;
        RECT 19.720 37.720 23.220 37.890 ;
        RECT 19.710 37.670 23.220 37.720 ;
        RECT 19.710 36.610 19.890 37.670 ;
        RECT 19.720 33.840 19.890 36.610 ;
        RECT 20.290 36.420 21.290 36.590 ;
        RECT 21.580 36.420 22.580 36.590 ;
        RECT 20.060 35.210 20.230 36.250 ;
        RECT 21.350 35.210 21.520 36.250 ;
        RECT 22.640 35.210 22.810 36.250 ;
        RECT 20.290 34.870 21.290 35.040 ;
        RECT 21.580 34.870 22.580 35.040 ;
        RECT 23.050 33.840 23.220 37.670 ;
        RECT 19.720 33.670 23.220 33.840 ;
        RECT 19.710 33.620 23.220 33.670 ;
        RECT 19.710 32.560 19.890 33.620 ;
        RECT 19.720 29.790 19.890 32.560 ;
        RECT 20.290 32.370 21.290 32.540 ;
        RECT 21.580 32.370 22.580 32.540 ;
        RECT 20.060 31.160 20.230 32.200 ;
        RECT 21.350 31.160 21.520 32.200 ;
        RECT 22.640 31.160 22.810 32.200 ;
        RECT 20.290 30.820 21.290 30.990 ;
        RECT 21.580 30.820 22.580 30.990 ;
        RECT 23.050 29.790 23.220 33.620 ;
        RECT 19.720 29.620 23.220 29.790 ;
        RECT 19.710 29.570 23.220 29.620 ;
        RECT 19.710 28.510 19.890 29.570 ;
        RECT 19.720 25.730 19.890 28.510 ;
        RECT 20.290 28.320 21.290 28.490 ;
        RECT 21.580 28.320 22.580 28.490 ;
        RECT 20.060 27.110 20.230 28.150 ;
        RECT 21.350 27.110 21.520 28.150 ;
        RECT 22.640 27.110 22.810 28.150 ;
        RECT 20.290 26.770 21.290 26.940 ;
        RECT 21.580 26.770 22.580 26.940 ;
        RECT 23.050 25.730 23.220 29.570 ;
        RECT 19.720 25.535 23.220 25.730 ;
        RECT 19.710 25.520 23.220 25.535 ;
        RECT 19.710 24.425 19.890 25.520 ;
        RECT 19.720 21.645 19.890 24.425 ;
        RECT 20.290 24.235 21.290 24.405 ;
        RECT 21.580 24.235 22.580 24.405 ;
        RECT 20.060 23.025 20.230 24.065 ;
        RECT 21.350 23.025 21.520 24.065 ;
        RECT 22.640 23.025 22.810 24.065 ;
        RECT 20.290 22.685 21.290 22.855 ;
        RECT 21.580 22.685 22.580 22.855 ;
        RECT 23.050 21.645 23.220 25.520 ;
        RECT 19.720 21.410 23.220 21.645 ;
        RECT 19.710 21.400 23.220 21.410 ;
        RECT 19.710 20.300 19.890 21.400 ;
        RECT 19.720 17.520 19.890 20.300 ;
        RECT 20.290 20.110 21.290 20.280 ;
        RECT 21.580 20.110 22.580 20.280 ;
        RECT 20.060 18.900 20.230 19.940 ;
        RECT 21.350 18.900 21.520 19.940 ;
        RECT 22.640 18.900 22.810 19.940 ;
        RECT 20.290 18.560 21.290 18.730 ;
        RECT 21.580 18.560 22.580 18.730 ;
        RECT 23.050 17.520 23.220 21.400 ;
        RECT 19.720 17.310 23.220 17.520 ;
        RECT 23.570 143.020 27.670 143.190 ;
        RECT 23.570 139.200 23.740 143.020 ;
        RECT 24.480 142.195 25.480 142.365 ;
        RECT 25.770 142.195 26.770 142.365 ;
        RECT 24.250 139.940 24.420 141.980 ;
        RECT 25.540 139.940 25.710 141.980 ;
        RECT 26.830 139.940 27.000 141.980 ;
        RECT 24.480 139.555 25.480 139.725 ;
        RECT 25.770 139.555 26.770 139.725 ;
        RECT 23.570 139.190 24.480 139.200 ;
        RECT 27.490 139.190 27.670 143.020 ;
        RECT 23.570 138.920 27.670 139.190 ;
        RECT 23.570 135.130 23.740 138.920 ;
        RECT 24.480 138.195 25.480 138.365 ;
        RECT 25.770 138.195 26.770 138.365 ;
        RECT 24.250 135.940 24.420 137.980 ;
        RECT 25.540 135.940 25.710 137.980 ;
        RECT 26.830 135.940 27.000 137.980 ;
        RECT 24.480 135.555 25.480 135.725 ;
        RECT 25.770 135.555 26.770 135.725 ;
        RECT 27.490 135.130 27.670 138.920 ;
        RECT 23.570 134.920 27.670 135.130 ;
        RECT 23.570 131.050 23.740 134.920 ;
        RECT 24.480 134.095 25.480 134.265 ;
        RECT 25.770 134.095 26.770 134.265 ;
        RECT 24.250 131.840 24.420 133.880 ;
        RECT 25.540 131.840 25.710 133.880 ;
        RECT 26.830 131.840 27.000 133.880 ;
        RECT 24.480 131.455 25.480 131.625 ;
        RECT 25.770 131.455 26.770 131.625 ;
        RECT 23.570 131.040 24.480 131.050 ;
        RECT 27.490 131.040 27.670 134.920 ;
        RECT 23.570 130.820 27.670 131.040 ;
        RECT 23.570 127.000 23.740 130.820 ;
        RECT 24.480 130.045 25.480 130.215 ;
        RECT 25.770 130.045 26.770 130.215 ;
        RECT 24.250 127.790 24.420 129.830 ;
        RECT 25.540 127.790 25.710 129.830 ;
        RECT 26.830 127.790 27.000 129.830 ;
        RECT 24.480 127.405 25.480 127.575 ;
        RECT 25.770 127.405 26.770 127.575 ;
        RECT 23.570 126.990 24.480 127.000 ;
        RECT 27.490 126.990 27.670 130.820 ;
        RECT 23.570 126.770 27.670 126.990 ;
        RECT 23.570 122.950 23.740 126.770 ;
        RECT 24.480 125.995 25.480 126.165 ;
        RECT 25.770 125.995 26.770 126.165 ;
        RECT 24.250 123.740 24.420 125.780 ;
        RECT 25.540 123.740 25.710 125.780 ;
        RECT 26.830 123.740 27.000 125.780 ;
        RECT 24.480 123.355 25.480 123.525 ;
        RECT 25.770 123.355 26.770 123.525 ;
        RECT 23.570 122.940 24.480 122.950 ;
        RECT 27.490 122.940 27.670 126.770 ;
        RECT 23.570 122.720 27.670 122.940 ;
        RECT 23.570 118.900 23.740 122.720 ;
        RECT 24.480 121.945 25.480 122.115 ;
        RECT 25.770 121.945 26.770 122.115 ;
        RECT 24.250 119.690 24.420 121.730 ;
        RECT 25.540 119.690 25.710 121.730 ;
        RECT 26.830 119.690 27.000 121.730 ;
        RECT 24.480 119.305 25.480 119.475 ;
        RECT 25.770 119.305 26.770 119.475 ;
        RECT 23.570 118.890 24.480 118.900 ;
        RECT 27.490 118.890 27.670 122.720 ;
        RECT 23.570 118.670 27.670 118.890 ;
        RECT 23.570 114.850 23.740 118.670 ;
        RECT 24.480 117.895 25.480 118.065 ;
        RECT 25.770 117.895 26.770 118.065 ;
        RECT 24.250 115.640 24.420 117.680 ;
        RECT 25.540 115.640 25.710 117.680 ;
        RECT 26.830 115.640 27.000 117.680 ;
        RECT 24.480 115.255 25.480 115.425 ;
        RECT 25.770 115.255 26.770 115.425 ;
        RECT 23.570 114.840 24.480 114.850 ;
        RECT 27.490 114.840 27.670 118.670 ;
        RECT 23.570 114.620 27.670 114.840 ;
        RECT 23.570 110.800 23.740 114.620 ;
        RECT 24.480 113.845 25.480 114.015 ;
        RECT 25.770 113.845 26.770 114.015 ;
        RECT 24.250 111.590 24.420 113.630 ;
        RECT 25.540 111.590 25.710 113.630 ;
        RECT 26.830 111.590 27.000 113.630 ;
        RECT 24.480 111.205 25.480 111.375 ;
        RECT 25.770 111.205 26.770 111.375 ;
        RECT 23.570 110.790 24.480 110.800 ;
        RECT 27.490 110.790 27.670 114.620 ;
        RECT 23.570 110.570 27.670 110.790 ;
        RECT 23.570 106.750 23.740 110.570 ;
        RECT 24.480 109.795 25.480 109.965 ;
        RECT 25.770 109.795 26.770 109.965 ;
        RECT 24.250 107.540 24.420 109.580 ;
        RECT 25.540 107.540 25.710 109.580 ;
        RECT 26.830 107.540 27.000 109.580 ;
        RECT 24.480 107.155 25.480 107.325 ;
        RECT 25.770 107.155 26.770 107.325 ;
        RECT 23.570 106.740 24.480 106.750 ;
        RECT 27.490 106.740 27.670 110.570 ;
        RECT 23.570 106.520 27.670 106.740 ;
        RECT 23.570 102.700 23.740 106.520 ;
        RECT 24.480 105.745 25.480 105.915 ;
        RECT 25.770 105.745 26.770 105.915 ;
        RECT 24.250 103.490 24.420 105.530 ;
        RECT 25.540 103.490 25.710 105.530 ;
        RECT 26.830 103.490 27.000 105.530 ;
        RECT 24.480 103.105 25.480 103.275 ;
        RECT 25.770 103.105 26.770 103.275 ;
        RECT 23.570 102.690 24.480 102.700 ;
        RECT 27.490 102.690 27.670 106.520 ;
        RECT 23.570 102.470 27.670 102.690 ;
        RECT 23.570 98.650 23.740 102.470 ;
        RECT 24.480 101.695 25.480 101.865 ;
        RECT 25.770 101.695 26.770 101.865 ;
        RECT 24.250 99.440 24.420 101.480 ;
        RECT 25.540 99.440 25.710 101.480 ;
        RECT 26.830 99.440 27.000 101.480 ;
        RECT 24.480 99.055 25.480 99.225 ;
        RECT 25.770 99.055 26.770 99.225 ;
        RECT 23.570 98.640 24.480 98.650 ;
        RECT 27.490 98.640 27.670 102.470 ;
        RECT 23.570 98.420 27.670 98.640 ;
        RECT 23.570 94.600 23.740 98.420 ;
        RECT 24.480 97.645 25.480 97.815 ;
        RECT 25.770 97.645 26.770 97.815 ;
        RECT 24.250 95.390 24.420 97.430 ;
        RECT 25.540 95.390 25.710 97.430 ;
        RECT 26.830 95.390 27.000 97.430 ;
        RECT 24.480 95.005 25.480 95.175 ;
        RECT 25.770 95.005 26.770 95.175 ;
        RECT 23.570 94.590 24.480 94.600 ;
        RECT 27.490 94.590 27.670 98.420 ;
        RECT 23.570 94.370 27.670 94.590 ;
        RECT 23.570 90.550 23.740 94.370 ;
        RECT 24.480 93.595 25.480 93.765 ;
        RECT 25.770 93.595 26.770 93.765 ;
        RECT 24.250 91.340 24.420 93.380 ;
        RECT 25.540 91.340 25.710 93.380 ;
        RECT 26.830 91.340 27.000 93.380 ;
        RECT 24.480 90.955 25.480 91.125 ;
        RECT 25.770 90.955 26.770 91.125 ;
        RECT 23.570 90.540 24.480 90.550 ;
        RECT 27.490 90.540 27.670 94.370 ;
        RECT 23.570 90.320 27.670 90.540 ;
        RECT 23.570 86.500 23.740 90.320 ;
        RECT 24.480 89.545 25.480 89.715 ;
        RECT 25.770 89.545 26.770 89.715 ;
        RECT 24.250 87.290 24.420 89.330 ;
        RECT 25.540 87.290 25.710 89.330 ;
        RECT 26.830 87.290 27.000 89.330 ;
        RECT 24.480 86.905 25.480 87.075 ;
        RECT 25.770 86.905 26.770 87.075 ;
        RECT 23.570 86.490 24.480 86.500 ;
        RECT 27.490 86.490 27.670 90.320 ;
        RECT 23.570 86.270 27.670 86.490 ;
        RECT 23.570 82.450 23.740 86.270 ;
        RECT 24.480 85.495 25.480 85.665 ;
        RECT 25.770 85.495 26.770 85.665 ;
        RECT 24.250 83.240 24.420 85.280 ;
        RECT 25.540 83.240 25.710 85.280 ;
        RECT 26.830 83.240 27.000 85.280 ;
        RECT 24.480 82.855 25.480 83.025 ;
        RECT 25.770 82.855 26.770 83.025 ;
        RECT 23.570 82.440 24.480 82.450 ;
        RECT 27.490 82.440 27.670 86.270 ;
        RECT 23.570 82.220 27.670 82.440 ;
        RECT 23.570 78.400 23.740 82.220 ;
        RECT 24.480 81.445 25.480 81.615 ;
        RECT 25.770 81.445 26.770 81.615 ;
        RECT 24.250 79.190 24.420 81.230 ;
        RECT 25.540 79.190 25.710 81.230 ;
        RECT 26.830 79.190 27.000 81.230 ;
        RECT 24.480 78.805 25.480 78.975 ;
        RECT 25.770 78.805 26.770 78.975 ;
        RECT 23.570 78.390 24.480 78.400 ;
        RECT 27.490 78.390 27.670 82.220 ;
        RECT 23.570 78.170 27.670 78.390 ;
        RECT 23.570 74.350 23.740 78.170 ;
        RECT 24.480 77.395 25.480 77.565 ;
        RECT 25.770 77.395 26.770 77.565 ;
        RECT 24.250 75.140 24.420 77.180 ;
        RECT 25.540 75.140 25.710 77.180 ;
        RECT 26.830 75.140 27.000 77.180 ;
        RECT 24.480 74.755 25.480 74.925 ;
        RECT 25.770 74.755 26.770 74.925 ;
        RECT 23.570 74.340 24.480 74.350 ;
        RECT 27.490 74.340 27.670 78.170 ;
        RECT 23.570 74.120 27.670 74.340 ;
        RECT 23.570 70.300 23.740 74.120 ;
        RECT 24.480 73.345 25.480 73.515 ;
        RECT 25.770 73.345 26.770 73.515 ;
        RECT 24.250 71.090 24.420 73.130 ;
        RECT 25.540 71.090 25.710 73.130 ;
        RECT 26.830 71.090 27.000 73.130 ;
        RECT 24.480 70.705 25.480 70.875 ;
        RECT 25.770 70.705 26.770 70.875 ;
        RECT 23.570 70.290 24.480 70.300 ;
        RECT 27.490 70.290 27.670 74.120 ;
        RECT 23.570 70.070 27.670 70.290 ;
        RECT 23.570 66.250 23.740 70.070 ;
        RECT 24.480 69.295 25.480 69.465 ;
        RECT 25.770 69.295 26.770 69.465 ;
        RECT 24.250 67.040 24.420 69.080 ;
        RECT 25.540 67.040 25.710 69.080 ;
        RECT 26.830 67.040 27.000 69.080 ;
        RECT 24.480 66.655 25.480 66.825 ;
        RECT 25.770 66.655 26.770 66.825 ;
        RECT 23.570 66.240 24.480 66.250 ;
        RECT 27.490 66.240 27.670 70.070 ;
        RECT 23.570 66.020 27.670 66.240 ;
        RECT 23.570 62.200 23.740 66.020 ;
        RECT 24.480 65.245 25.480 65.415 ;
        RECT 25.770 65.245 26.770 65.415 ;
        RECT 24.250 62.990 24.420 65.030 ;
        RECT 25.540 62.990 25.710 65.030 ;
        RECT 26.830 62.990 27.000 65.030 ;
        RECT 24.480 62.605 25.480 62.775 ;
        RECT 25.770 62.605 26.770 62.775 ;
        RECT 23.570 62.190 24.480 62.200 ;
        RECT 27.490 62.190 27.670 66.020 ;
        RECT 23.570 61.970 27.670 62.190 ;
        RECT 23.570 58.150 23.740 61.970 ;
        RECT 24.480 61.195 25.480 61.365 ;
        RECT 25.770 61.195 26.770 61.365 ;
        RECT 24.250 58.940 24.420 60.980 ;
        RECT 25.540 58.940 25.710 60.980 ;
        RECT 26.830 58.940 27.000 60.980 ;
        RECT 24.480 58.555 25.480 58.725 ;
        RECT 25.770 58.555 26.770 58.725 ;
        RECT 23.570 58.140 24.480 58.150 ;
        RECT 27.490 58.140 27.670 61.970 ;
        RECT 23.570 57.920 27.670 58.140 ;
        RECT 23.570 54.100 23.740 57.920 ;
        RECT 24.480 57.145 25.480 57.315 ;
        RECT 25.770 57.145 26.770 57.315 ;
        RECT 24.250 54.890 24.420 56.930 ;
        RECT 25.540 54.890 25.710 56.930 ;
        RECT 26.830 54.890 27.000 56.930 ;
        RECT 24.480 54.505 25.480 54.675 ;
        RECT 25.770 54.505 26.770 54.675 ;
        RECT 23.570 54.090 24.480 54.100 ;
        RECT 27.490 54.090 27.670 57.920 ;
        RECT 28.010 143.020 32.110 143.190 ;
        RECT 28.010 139.130 28.190 143.020 ;
        RECT 28.910 142.195 29.910 142.365 ;
        RECT 30.200 142.195 31.200 142.365 ;
        RECT 28.680 139.940 28.850 141.980 ;
        RECT 29.970 139.940 30.140 141.980 ;
        RECT 31.260 139.940 31.430 141.980 ;
        RECT 28.910 139.555 29.910 139.725 ;
        RECT 30.200 139.555 31.200 139.725 ;
        RECT 31.940 139.140 32.110 143.020 ;
        RECT 31.200 139.130 32.110 139.140 ;
        RECT 28.010 138.920 32.110 139.130 ;
        RECT 28.010 135.070 28.190 138.920 ;
        RECT 28.910 138.135 29.910 138.305 ;
        RECT 30.200 138.135 31.200 138.305 ;
        RECT 28.680 135.880 28.850 137.920 ;
        RECT 29.970 135.880 30.140 137.920 ;
        RECT 31.260 135.880 31.430 137.920 ;
        RECT 28.910 135.495 29.910 135.665 ;
        RECT 30.200 135.495 31.200 135.665 ;
        RECT 31.940 135.080 32.110 138.920 ;
        RECT 31.200 135.070 32.110 135.080 ;
        RECT 28.010 134.860 32.110 135.070 ;
        RECT 28.010 131.010 28.190 134.860 ;
        RECT 28.910 134.075 29.910 134.245 ;
        RECT 30.200 134.075 31.200 134.245 ;
        RECT 28.680 131.820 28.850 133.860 ;
        RECT 29.970 131.820 30.140 133.860 ;
        RECT 31.260 131.820 31.430 133.860 ;
        RECT 28.910 131.435 29.910 131.605 ;
        RECT 30.200 131.435 31.200 131.605 ;
        RECT 31.940 131.020 32.110 134.860 ;
        RECT 31.200 131.010 32.110 131.020 ;
        RECT 28.010 130.800 32.110 131.010 ;
        RECT 28.010 126.950 28.190 130.800 ;
        RECT 28.910 130.015 29.910 130.185 ;
        RECT 30.200 130.015 31.200 130.185 ;
        RECT 28.680 127.760 28.850 129.800 ;
        RECT 29.970 127.760 30.140 129.800 ;
        RECT 31.260 127.760 31.430 129.800 ;
        RECT 28.910 127.375 29.910 127.545 ;
        RECT 30.200 127.375 31.200 127.545 ;
        RECT 31.940 126.960 32.110 130.800 ;
        RECT 31.200 126.950 32.110 126.960 ;
        RECT 28.010 126.740 32.110 126.950 ;
        RECT 28.010 122.890 28.190 126.740 ;
        RECT 28.910 125.955 29.910 126.125 ;
        RECT 30.200 125.955 31.200 126.125 ;
        RECT 28.680 123.700 28.850 125.740 ;
        RECT 29.970 123.700 30.140 125.740 ;
        RECT 31.260 123.700 31.430 125.740 ;
        RECT 28.910 123.315 29.910 123.485 ;
        RECT 30.200 123.315 31.200 123.485 ;
        RECT 31.940 122.900 32.110 126.740 ;
        RECT 31.200 122.890 32.110 122.900 ;
        RECT 28.010 122.680 32.110 122.890 ;
        RECT 28.010 118.830 28.190 122.680 ;
        RECT 28.910 121.895 29.910 122.065 ;
        RECT 30.200 121.895 31.200 122.065 ;
        RECT 28.680 119.640 28.850 121.680 ;
        RECT 29.970 119.640 30.140 121.680 ;
        RECT 31.260 119.640 31.430 121.680 ;
        RECT 28.910 119.255 29.910 119.425 ;
        RECT 30.200 119.255 31.200 119.425 ;
        RECT 31.940 118.840 32.110 122.680 ;
        RECT 31.200 118.830 32.110 118.840 ;
        RECT 28.010 118.620 32.110 118.830 ;
        RECT 28.010 114.770 28.190 118.620 ;
        RECT 28.910 117.835 29.910 118.005 ;
        RECT 30.200 117.835 31.200 118.005 ;
        RECT 28.680 115.580 28.850 117.620 ;
        RECT 29.970 115.580 30.140 117.620 ;
        RECT 31.260 115.580 31.430 117.620 ;
        RECT 28.910 115.195 29.910 115.365 ;
        RECT 30.200 115.195 31.200 115.365 ;
        RECT 31.940 114.780 32.110 118.620 ;
        RECT 31.200 114.770 32.110 114.780 ;
        RECT 28.010 114.560 32.110 114.770 ;
        RECT 28.010 110.710 28.190 114.560 ;
        RECT 28.910 113.775 29.910 113.945 ;
        RECT 30.200 113.775 31.200 113.945 ;
        RECT 28.680 111.520 28.850 113.560 ;
        RECT 29.970 111.520 30.140 113.560 ;
        RECT 31.260 111.520 31.430 113.560 ;
        RECT 28.910 111.135 29.910 111.305 ;
        RECT 30.200 111.135 31.200 111.305 ;
        RECT 31.940 110.720 32.110 114.560 ;
        RECT 31.200 110.710 32.110 110.720 ;
        RECT 28.010 110.500 32.110 110.710 ;
        RECT 28.010 106.650 28.190 110.500 ;
        RECT 28.910 109.715 29.910 109.885 ;
        RECT 30.200 109.715 31.200 109.885 ;
        RECT 28.680 107.460 28.850 109.500 ;
        RECT 29.970 107.460 30.140 109.500 ;
        RECT 31.260 107.460 31.430 109.500 ;
        RECT 28.910 107.075 29.910 107.245 ;
        RECT 30.200 107.075 31.200 107.245 ;
        RECT 31.940 106.660 32.110 110.500 ;
        RECT 31.200 106.650 32.110 106.660 ;
        RECT 28.010 106.440 32.110 106.650 ;
        RECT 28.010 102.590 28.190 106.440 ;
        RECT 28.910 105.655 29.910 105.825 ;
        RECT 30.200 105.655 31.200 105.825 ;
        RECT 28.680 103.400 28.850 105.440 ;
        RECT 29.970 103.400 30.140 105.440 ;
        RECT 31.260 103.400 31.430 105.440 ;
        RECT 28.910 103.015 29.910 103.185 ;
        RECT 30.200 103.015 31.200 103.185 ;
        RECT 31.940 102.600 32.110 106.440 ;
        RECT 31.200 102.590 32.110 102.600 ;
        RECT 28.010 102.380 32.110 102.590 ;
        RECT 28.010 98.530 28.190 102.380 ;
        RECT 28.910 101.595 29.910 101.765 ;
        RECT 30.200 101.595 31.200 101.765 ;
        RECT 28.680 99.340 28.850 101.380 ;
        RECT 29.970 99.340 30.140 101.380 ;
        RECT 31.260 99.340 31.430 101.380 ;
        RECT 28.910 98.955 29.910 99.125 ;
        RECT 30.200 98.955 31.200 99.125 ;
        RECT 31.940 98.540 32.110 102.380 ;
        RECT 31.200 98.530 32.110 98.540 ;
        RECT 28.010 98.320 32.110 98.530 ;
        RECT 28.010 94.470 28.190 98.320 ;
        RECT 28.910 97.535 29.910 97.705 ;
        RECT 30.200 97.535 31.200 97.705 ;
        RECT 28.680 95.280 28.850 97.320 ;
        RECT 29.970 95.280 30.140 97.320 ;
        RECT 31.260 95.280 31.430 97.320 ;
        RECT 28.910 94.895 29.910 95.065 ;
        RECT 30.200 94.895 31.200 95.065 ;
        RECT 31.940 94.480 32.110 98.320 ;
        RECT 31.200 94.470 32.110 94.480 ;
        RECT 28.010 94.260 32.110 94.470 ;
        RECT 28.010 90.410 28.190 94.260 ;
        RECT 28.910 93.475 29.910 93.645 ;
        RECT 30.200 93.475 31.200 93.645 ;
        RECT 28.680 91.220 28.850 93.260 ;
        RECT 29.970 91.220 30.140 93.260 ;
        RECT 31.260 91.220 31.430 93.260 ;
        RECT 28.910 90.835 29.910 91.005 ;
        RECT 30.200 90.835 31.200 91.005 ;
        RECT 31.940 90.420 32.110 94.260 ;
        RECT 31.200 90.410 32.110 90.420 ;
        RECT 28.010 90.200 32.110 90.410 ;
        RECT 28.010 86.350 28.190 90.200 ;
        RECT 28.910 89.415 29.910 89.585 ;
        RECT 30.200 89.415 31.200 89.585 ;
        RECT 28.680 87.160 28.850 89.200 ;
        RECT 29.970 87.160 30.140 89.200 ;
        RECT 31.260 87.160 31.430 89.200 ;
        RECT 28.910 86.775 29.910 86.945 ;
        RECT 30.200 86.775 31.200 86.945 ;
        RECT 31.940 86.360 32.110 90.200 ;
        RECT 31.200 86.350 32.110 86.360 ;
        RECT 28.010 86.140 32.110 86.350 ;
        RECT 28.010 82.290 28.190 86.140 ;
        RECT 28.910 85.355 29.910 85.525 ;
        RECT 30.200 85.355 31.200 85.525 ;
        RECT 28.680 83.100 28.850 85.140 ;
        RECT 29.970 83.100 30.140 85.140 ;
        RECT 31.260 83.100 31.430 85.140 ;
        RECT 28.910 82.715 29.910 82.885 ;
        RECT 30.200 82.715 31.200 82.885 ;
        RECT 31.940 82.300 32.110 86.140 ;
        RECT 31.200 82.290 32.110 82.300 ;
        RECT 28.010 82.080 32.110 82.290 ;
        RECT 28.010 78.230 28.190 82.080 ;
        RECT 28.910 81.295 29.910 81.465 ;
        RECT 30.200 81.295 31.200 81.465 ;
        RECT 28.680 79.040 28.850 81.080 ;
        RECT 29.970 79.040 30.140 81.080 ;
        RECT 31.260 79.040 31.430 81.080 ;
        RECT 28.910 78.655 29.910 78.825 ;
        RECT 30.200 78.655 31.200 78.825 ;
        RECT 31.940 78.240 32.110 82.080 ;
        RECT 31.200 78.230 32.110 78.240 ;
        RECT 28.010 78.020 32.110 78.230 ;
        RECT 28.010 74.170 28.190 78.020 ;
        RECT 28.910 77.235 29.910 77.405 ;
        RECT 30.200 77.235 31.200 77.405 ;
        RECT 28.680 74.980 28.850 77.020 ;
        RECT 29.970 74.980 30.140 77.020 ;
        RECT 31.260 74.980 31.430 77.020 ;
        RECT 28.910 74.595 29.910 74.765 ;
        RECT 30.200 74.595 31.200 74.765 ;
        RECT 31.940 74.180 32.110 78.020 ;
        RECT 31.200 74.170 32.110 74.180 ;
        RECT 28.010 73.960 32.110 74.170 ;
        RECT 28.010 70.110 28.190 73.960 ;
        RECT 28.910 73.175 29.910 73.345 ;
        RECT 30.200 73.175 31.200 73.345 ;
        RECT 28.680 70.920 28.850 72.960 ;
        RECT 29.970 70.920 30.140 72.960 ;
        RECT 31.260 70.920 31.430 72.960 ;
        RECT 28.910 70.535 29.910 70.705 ;
        RECT 30.200 70.535 31.200 70.705 ;
        RECT 31.940 70.120 32.110 73.960 ;
        RECT 31.200 70.110 32.110 70.120 ;
        RECT 28.010 69.900 32.110 70.110 ;
        RECT 28.010 66.050 28.190 69.900 ;
        RECT 28.910 69.115 29.910 69.285 ;
        RECT 30.200 69.115 31.200 69.285 ;
        RECT 28.680 66.860 28.850 68.900 ;
        RECT 29.970 66.860 30.140 68.900 ;
        RECT 31.260 66.860 31.430 68.900 ;
        RECT 28.910 66.475 29.910 66.645 ;
        RECT 30.200 66.475 31.200 66.645 ;
        RECT 31.940 66.060 32.110 69.900 ;
        RECT 31.200 66.050 32.110 66.060 ;
        RECT 28.010 65.840 32.110 66.050 ;
        RECT 28.010 61.990 28.190 65.840 ;
        RECT 28.910 65.055 29.910 65.225 ;
        RECT 30.200 65.055 31.200 65.225 ;
        RECT 28.680 62.800 28.850 64.840 ;
        RECT 29.970 62.800 30.140 64.840 ;
        RECT 31.260 62.800 31.430 64.840 ;
        RECT 28.910 62.415 29.910 62.585 ;
        RECT 30.200 62.415 31.200 62.585 ;
        RECT 31.940 62.000 32.110 65.840 ;
        RECT 31.200 61.990 32.110 62.000 ;
        RECT 28.010 61.780 32.110 61.990 ;
        RECT 28.010 57.930 28.190 61.780 ;
        RECT 28.910 60.995 29.910 61.165 ;
        RECT 30.200 60.995 31.200 61.165 ;
        RECT 28.680 58.740 28.850 60.780 ;
        RECT 29.970 58.740 30.140 60.780 ;
        RECT 31.260 58.740 31.430 60.780 ;
        RECT 28.910 58.355 29.910 58.525 ;
        RECT 30.200 58.355 31.200 58.525 ;
        RECT 31.940 57.930 32.110 61.780 ;
        RECT 28.010 57.720 32.110 57.930 ;
        RECT 32.460 143.020 35.960 143.190 ;
        RECT 32.460 143.010 35.970 143.020 ;
        RECT 32.460 139.130 32.630 143.010 ;
        RECT 35.790 141.910 35.970 143.010 ;
        RECT 33.100 141.720 34.100 141.890 ;
        RECT 34.390 141.720 35.390 141.890 ;
        RECT 32.870 140.510 33.040 141.550 ;
        RECT 34.160 140.510 34.330 141.550 ;
        RECT 35.450 140.510 35.620 141.550 ;
        RECT 33.100 140.170 34.100 140.340 ;
        RECT 34.390 140.170 35.390 140.340 ;
        RECT 35.790 139.130 35.960 141.910 ;
        RECT 32.460 138.960 35.960 139.130 ;
        RECT 32.460 138.920 35.970 138.960 ;
        RECT 32.460 135.070 32.630 138.920 ;
        RECT 35.790 137.850 35.970 138.920 ;
        RECT 33.100 137.660 34.100 137.830 ;
        RECT 34.390 137.660 35.390 137.830 ;
        RECT 32.870 136.450 33.040 137.490 ;
        RECT 34.160 136.450 34.330 137.490 ;
        RECT 35.450 136.450 35.620 137.490 ;
        RECT 33.100 136.110 34.100 136.280 ;
        RECT 34.390 136.110 35.390 136.280 ;
        RECT 35.790 135.070 35.960 137.850 ;
        RECT 32.460 134.900 35.960 135.070 ;
        RECT 32.460 134.860 35.970 134.900 ;
        RECT 32.460 131.010 32.630 134.860 ;
        RECT 35.790 133.790 35.970 134.860 ;
        RECT 33.100 133.600 34.100 133.770 ;
        RECT 34.390 133.600 35.390 133.770 ;
        RECT 32.870 132.390 33.040 133.430 ;
        RECT 34.160 132.390 34.330 133.430 ;
        RECT 35.450 132.390 35.620 133.430 ;
        RECT 33.100 132.050 34.100 132.220 ;
        RECT 34.390 132.050 35.390 132.220 ;
        RECT 35.790 131.010 35.960 133.790 ;
        RECT 32.460 130.840 35.960 131.010 ;
        RECT 32.460 130.800 35.970 130.840 ;
        RECT 32.460 126.950 32.630 130.800 ;
        RECT 35.790 129.730 35.970 130.800 ;
        RECT 33.100 129.540 34.100 129.710 ;
        RECT 34.390 129.540 35.390 129.710 ;
        RECT 32.870 128.330 33.040 129.370 ;
        RECT 34.160 128.330 34.330 129.370 ;
        RECT 35.450 128.330 35.620 129.370 ;
        RECT 33.100 127.990 34.100 128.160 ;
        RECT 34.390 127.990 35.390 128.160 ;
        RECT 35.790 126.950 35.960 129.730 ;
        RECT 32.460 126.780 35.960 126.950 ;
        RECT 32.460 126.740 35.970 126.780 ;
        RECT 32.460 122.890 32.630 126.740 ;
        RECT 35.790 125.670 35.970 126.740 ;
        RECT 33.100 125.480 34.100 125.650 ;
        RECT 34.390 125.480 35.390 125.650 ;
        RECT 32.870 124.270 33.040 125.310 ;
        RECT 34.160 124.270 34.330 125.310 ;
        RECT 35.450 124.270 35.620 125.310 ;
        RECT 33.100 123.930 34.100 124.100 ;
        RECT 34.390 123.930 35.390 124.100 ;
        RECT 35.790 122.890 35.960 125.670 ;
        RECT 32.460 122.720 35.960 122.890 ;
        RECT 32.460 122.680 35.970 122.720 ;
        RECT 32.460 118.830 32.630 122.680 ;
        RECT 35.790 121.610 35.970 122.680 ;
        RECT 33.100 121.420 34.100 121.590 ;
        RECT 34.390 121.420 35.390 121.590 ;
        RECT 32.870 120.210 33.040 121.250 ;
        RECT 34.160 120.210 34.330 121.250 ;
        RECT 35.450 120.210 35.620 121.250 ;
        RECT 33.100 119.870 34.100 120.040 ;
        RECT 34.390 119.870 35.390 120.040 ;
        RECT 35.790 118.830 35.960 121.610 ;
        RECT 32.460 118.660 35.960 118.830 ;
        RECT 32.460 118.620 35.970 118.660 ;
        RECT 32.460 114.770 32.630 118.620 ;
        RECT 35.790 117.550 35.970 118.620 ;
        RECT 33.100 117.360 34.100 117.530 ;
        RECT 34.390 117.360 35.390 117.530 ;
        RECT 32.870 116.150 33.040 117.190 ;
        RECT 34.160 116.150 34.330 117.190 ;
        RECT 35.450 116.150 35.620 117.190 ;
        RECT 33.100 115.810 34.100 115.980 ;
        RECT 34.390 115.810 35.390 115.980 ;
        RECT 35.790 114.770 35.960 117.550 ;
        RECT 32.460 114.600 35.960 114.770 ;
        RECT 32.460 114.560 35.970 114.600 ;
        RECT 32.460 110.710 32.630 114.560 ;
        RECT 35.790 113.490 35.970 114.560 ;
        RECT 33.100 113.300 34.100 113.470 ;
        RECT 34.390 113.300 35.390 113.470 ;
        RECT 32.870 112.090 33.040 113.130 ;
        RECT 34.160 112.090 34.330 113.130 ;
        RECT 35.450 112.090 35.620 113.130 ;
        RECT 33.100 111.750 34.100 111.920 ;
        RECT 34.390 111.750 35.390 111.920 ;
        RECT 35.790 110.710 35.960 113.490 ;
        RECT 32.460 110.540 35.960 110.710 ;
        RECT 32.460 110.500 35.970 110.540 ;
        RECT 32.460 106.650 32.630 110.500 ;
        RECT 35.790 109.430 35.970 110.500 ;
        RECT 33.100 109.240 34.100 109.410 ;
        RECT 34.390 109.240 35.390 109.410 ;
        RECT 32.870 108.030 33.040 109.070 ;
        RECT 34.160 108.030 34.330 109.070 ;
        RECT 35.450 108.030 35.620 109.070 ;
        RECT 33.100 107.690 34.100 107.860 ;
        RECT 34.390 107.690 35.390 107.860 ;
        RECT 35.790 106.650 35.960 109.430 ;
        RECT 32.460 106.480 35.960 106.650 ;
        RECT 32.460 106.440 35.970 106.480 ;
        RECT 32.460 102.590 32.630 106.440 ;
        RECT 35.790 105.370 35.970 106.440 ;
        RECT 33.100 105.180 34.100 105.350 ;
        RECT 34.390 105.180 35.390 105.350 ;
        RECT 32.870 103.970 33.040 105.010 ;
        RECT 34.160 103.970 34.330 105.010 ;
        RECT 35.450 103.970 35.620 105.010 ;
        RECT 33.100 103.630 34.100 103.800 ;
        RECT 34.390 103.630 35.390 103.800 ;
        RECT 35.790 102.590 35.960 105.370 ;
        RECT 32.460 102.420 35.960 102.590 ;
        RECT 32.460 102.380 35.970 102.420 ;
        RECT 32.460 98.530 32.630 102.380 ;
        RECT 35.790 101.310 35.970 102.380 ;
        RECT 33.100 101.120 34.100 101.290 ;
        RECT 34.390 101.120 35.390 101.290 ;
        RECT 32.870 99.910 33.040 100.950 ;
        RECT 34.160 99.910 34.330 100.950 ;
        RECT 35.450 99.910 35.620 100.950 ;
        RECT 33.100 99.570 34.100 99.740 ;
        RECT 34.390 99.570 35.390 99.740 ;
        RECT 35.790 98.530 35.960 101.310 ;
        RECT 32.460 98.360 35.960 98.530 ;
        RECT 32.460 98.320 35.970 98.360 ;
        RECT 32.460 94.470 32.630 98.320 ;
        RECT 35.790 97.250 35.970 98.320 ;
        RECT 33.100 97.060 34.100 97.230 ;
        RECT 34.390 97.060 35.390 97.230 ;
        RECT 32.870 95.850 33.040 96.890 ;
        RECT 34.160 95.850 34.330 96.890 ;
        RECT 35.450 95.850 35.620 96.890 ;
        RECT 33.100 95.510 34.100 95.680 ;
        RECT 34.390 95.510 35.390 95.680 ;
        RECT 35.790 94.470 35.960 97.250 ;
        RECT 32.460 94.300 35.960 94.470 ;
        RECT 32.460 94.260 35.970 94.300 ;
        RECT 32.460 90.410 32.630 94.260 ;
        RECT 35.790 93.190 35.970 94.260 ;
        RECT 33.100 93.000 34.100 93.170 ;
        RECT 34.390 93.000 35.390 93.170 ;
        RECT 32.870 91.790 33.040 92.830 ;
        RECT 34.160 91.790 34.330 92.830 ;
        RECT 35.450 91.790 35.620 92.830 ;
        RECT 33.100 91.450 34.100 91.620 ;
        RECT 34.390 91.450 35.390 91.620 ;
        RECT 35.790 90.410 35.960 93.190 ;
        RECT 32.460 90.240 35.960 90.410 ;
        RECT 32.460 90.200 35.970 90.240 ;
        RECT 32.460 86.350 32.630 90.200 ;
        RECT 35.790 89.130 35.970 90.200 ;
        RECT 33.100 88.940 34.100 89.110 ;
        RECT 34.390 88.940 35.390 89.110 ;
        RECT 32.870 87.730 33.040 88.770 ;
        RECT 34.160 87.730 34.330 88.770 ;
        RECT 35.450 87.730 35.620 88.770 ;
        RECT 33.100 87.390 34.100 87.560 ;
        RECT 34.390 87.390 35.390 87.560 ;
        RECT 35.790 86.350 35.960 89.130 ;
        RECT 32.460 86.180 35.960 86.350 ;
        RECT 32.460 86.140 35.970 86.180 ;
        RECT 32.460 82.290 32.630 86.140 ;
        RECT 35.790 85.070 35.970 86.140 ;
        RECT 33.100 84.880 34.100 85.050 ;
        RECT 34.390 84.880 35.390 85.050 ;
        RECT 32.870 83.670 33.040 84.710 ;
        RECT 34.160 83.670 34.330 84.710 ;
        RECT 35.450 83.670 35.620 84.710 ;
        RECT 33.100 83.330 34.100 83.500 ;
        RECT 34.390 83.330 35.390 83.500 ;
        RECT 35.790 82.290 35.960 85.070 ;
        RECT 32.460 82.120 35.960 82.290 ;
        RECT 32.460 82.080 35.970 82.120 ;
        RECT 32.460 78.230 32.630 82.080 ;
        RECT 35.790 81.010 35.970 82.080 ;
        RECT 33.100 80.820 34.100 80.990 ;
        RECT 34.390 80.820 35.390 80.990 ;
        RECT 32.870 79.610 33.040 80.650 ;
        RECT 34.160 79.610 34.330 80.650 ;
        RECT 35.450 79.610 35.620 80.650 ;
        RECT 33.100 79.270 34.100 79.440 ;
        RECT 34.390 79.270 35.390 79.440 ;
        RECT 35.790 78.230 35.960 81.010 ;
        RECT 32.460 78.060 35.960 78.230 ;
        RECT 32.460 78.020 35.970 78.060 ;
        RECT 32.460 74.170 32.630 78.020 ;
        RECT 35.790 76.950 35.970 78.020 ;
        RECT 33.100 76.760 34.100 76.930 ;
        RECT 34.390 76.760 35.390 76.930 ;
        RECT 32.870 75.550 33.040 76.590 ;
        RECT 34.160 75.550 34.330 76.590 ;
        RECT 35.450 75.550 35.620 76.590 ;
        RECT 33.100 75.210 34.100 75.380 ;
        RECT 34.390 75.210 35.390 75.380 ;
        RECT 35.790 74.170 35.960 76.950 ;
        RECT 32.460 74.000 35.960 74.170 ;
        RECT 32.460 73.960 35.970 74.000 ;
        RECT 32.460 70.110 32.630 73.960 ;
        RECT 35.790 72.890 35.970 73.960 ;
        RECT 33.100 72.700 34.100 72.870 ;
        RECT 34.390 72.700 35.390 72.870 ;
        RECT 32.870 71.490 33.040 72.530 ;
        RECT 34.160 71.490 34.330 72.530 ;
        RECT 35.450 71.490 35.620 72.530 ;
        RECT 33.100 71.150 34.100 71.320 ;
        RECT 34.390 71.150 35.390 71.320 ;
        RECT 35.790 70.110 35.960 72.890 ;
        RECT 32.460 69.940 35.960 70.110 ;
        RECT 32.460 69.900 35.970 69.940 ;
        RECT 32.460 66.050 32.630 69.900 ;
        RECT 35.790 68.830 35.970 69.900 ;
        RECT 33.100 68.640 34.100 68.810 ;
        RECT 34.390 68.640 35.390 68.810 ;
        RECT 32.870 67.430 33.040 68.470 ;
        RECT 34.160 67.430 34.330 68.470 ;
        RECT 35.450 67.430 35.620 68.470 ;
        RECT 33.100 67.090 34.100 67.260 ;
        RECT 34.390 67.090 35.390 67.260 ;
        RECT 35.790 66.050 35.960 68.830 ;
        RECT 32.460 65.880 35.960 66.050 ;
        RECT 32.460 65.840 35.970 65.880 ;
        RECT 32.460 61.990 32.630 65.840 ;
        RECT 35.790 64.770 35.970 65.840 ;
        RECT 33.100 64.580 34.100 64.750 ;
        RECT 34.390 64.580 35.390 64.750 ;
        RECT 32.870 63.370 33.040 64.410 ;
        RECT 34.160 63.370 34.330 64.410 ;
        RECT 35.450 63.370 35.620 64.410 ;
        RECT 33.100 63.030 34.100 63.200 ;
        RECT 34.390 63.030 35.390 63.200 ;
        RECT 35.790 61.990 35.960 64.770 ;
        RECT 32.460 61.820 35.960 61.990 ;
        RECT 32.460 61.780 35.970 61.820 ;
        RECT 32.460 57.930 32.630 61.780 ;
        RECT 35.790 60.710 35.970 61.780 ;
        RECT 33.100 60.520 34.100 60.690 ;
        RECT 34.390 60.520 35.390 60.690 ;
        RECT 32.870 59.310 33.040 60.350 ;
        RECT 34.160 59.310 34.330 60.350 ;
        RECT 35.450 59.310 35.620 60.350 ;
        RECT 33.100 58.970 34.100 59.140 ;
        RECT 34.390 58.970 35.390 59.140 ;
        RECT 35.790 57.930 35.960 60.710 ;
        RECT 32.460 57.720 35.960 57.930 ;
        RECT 31.200 57.450 32.000 57.460 ;
        RECT 23.570 53.870 27.670 54.090 ;
        RECT 23.570 50.050 23.740 53.870 ;
        RECT 24.480 53.095 25.480 53.265 ;
        RECT 25.770 53.095 26.770 53.265 ;
        RECT 24.250 50.840 24.420 52.880 ;
        RECT 25.540 50.840 25.710 52.880 ;
        RECT 26.830 50.840 27.000 52.880 ;
        RECT 24.480 50.455 25.480 50.625 ;
        RECT 25.770 50.455 26.770 50.625 ;
        RECT 23.570 50.040 24.480 50.050 ;
        RECT 27.490 50.040 27.670 53.870 ;
        RECT 28.010 57.280 32.110 57.450 ;
        RECT 28.010 53.390 28.190 57.280 ;
        RECT 28.910 56.455 29.910 56.625 ;
        RECT 30.200 56.455 31.200 56.625 ;
        RECT 28.680 54.200 28.850 56.240 ;
        RECT 29.970 54.200 30.140 56.240 ;
        RECT 31.260 54.200 31.430 56.240 ;
        RECT 28.910 53.815 29.910 53.985 ;
        RECT 30.200 53.815 31.200 53.985 ;
        RECT 31.940 53.390 32.110 57.280 ;
        RECT 28.010 53.180 32.110 53.390 ;
        RECT 32.460 57.280 35.960 57.450 ;
        RECT 32.460 57.270 35.970 57.280 ;
        RECT 32.460 53.390 32.630 57.270 ;
        RECT 35.790 56.170 35.970 57.270 ;
        RECT 33.100 55.980 34.100 56.150 ;
        RECT 34.390 55.980 35.390 56.150 ;
        RECT 32.870 54.770 33.040 55.810 ;
        RECT 34.160 54.770 34.330 55.810 ;
        RECT 35.450 54.770 35.620 55.810 ;
        RECT 33.100 54.430 34.100 54.600 ;
        RECT 34.390 54.430 35.390 54.600 ;
        RECT 35.790 53.390 35.960 56.170 ;
        RECT 32.460 53.180 35.960 53.390 ;
        RECT 23.570 49.820 27.670 50.040 ;
        RECT 23.570 46.000 23.740 49.820 ;
        RECT 24.480 49.045 25.480 49.215 ;
        RECT 25.770 49.045 26.770 49.215 ;
        RECT 24.250 46.790 24.420 48.830 ;
        RECT 25.540 46.790 25.710 48.830 ;
        RECT 26.830 46.790 27.000 48.830 ;
        RECT 24.480 46.405 25.480 46.575 ;
        RECT 25.770 46.405 26.770 46.575 ;
        RECT 23.570 45.990 24.480 46.000 ;
        RECT 27.490 45.990 27.670 49.820 ;
        RECT 23.570 45.770 27.670 45.990 ;
        RECT 23.570 41.950 23.740 45.770 ;
        RECT 24.480 44.995 25.480 45.165 ;
        RECT 25.770 44.995 26.770 45.165 ;
        RECT 24.250 42.740 24.420 44.780 ;
        RECT 25.540 42.740 25.710 44.780 ;
        RECT 26.830 42.740 27.000 44.780 ;
        RECT 24.480 42.355 25.480 42.525 ;
        RECT 25.770 42.355 26.770 42.525 ;
        RECT 23.570 41.940 24.480 41.950 ;
        RECT 27.490 41.940 27.670 45.770 ;
        RECT 23.570 41.720 27.670 41.940 ;
        RECT 23.570 37.900 23.740 41.720 ;
        RECT 24.480 40.945 25.480 41.115 ;
        RECT 25.770 40.945 26.770 41.115 ;
        RECT 24.250 38.690 24.420 40.730 ;
        RECT 25.540 38.690 25.710 40.730 ;
        RECT 26.830 38.690 27.000 40.730 ;
        RECT 24.480 38.305 25.480 38.475 ;
        RECT 25.770 38.305 26.770 38.475 ;
        RECT 23.570 37.890 24.480 37.900 ;
        RECT 27.490 37.890 27.670 41.720 ;
        RECT 23.570 37.670 27.670 37.890 ;
        RECT 23.570 33.850 23.740 37.670 ;
        RECT 24.480 36.895 25.480 37.065 ;
        RECT 25.770 36.895 26.770 37.065 ;
        RECT 24.250 34.640 24.420 36.680 ;
        RECT 25.540 34.640 25.710 36.680 ;
        RECT 26.830 34.640 27.000 36.680 ;
        RECT 24.480 34.255 25.480 34.425 ;
        RECT 25.770 34.255 26.770 34.425 ;
        RECT 23.570 33.840 24.480 33.850 ;
        RECT 27.490 33.840 27.670 37.670 ;
        RECT 23.570 33.620 27.670 33.840 ;
        RECT 23.570 29.800 23.740 33.620 ;
        RECT 24.480 32.845 25.480 33.015 ;
        RECT 25.770 32.845 26.770 33.015 ;
        RECT 24.250 30.590 24.420 32.630 ;
        RECT 25.540 30.590 25.710 32.630 ;
        RECT 26.830 30.590 27.000 32.630 ;
        RECT 24.480 30.205 25.480 30.375 ;
        RECT 25.770 30.205 26.770 30.375 ;
        RECT 23.570 29.790 24.480 29.800 ;
        RECT 27.490 29.790 27.670 33.620 ;
        RECT 23.570 29.570 27.670 29.790 ;
        RECT 23.570 25.730 23.740 29.570 ;
        RECT 24.480 28.795 25.480 28.965 ;
        RECT 25.770 28.795 26.770 28.965 ;
        RECT 24.250 26.540 24.420 28.580 ;
        RECT 25.540 26.540 25.710 28.580 ;
        RECT 26.830 26.540 27.000 28.580 ;
        RECT 24.480 26.155 25.480 26.325 ;
        RECT 25.770 26.155 26.770 26.325 ;
        RECT 27.490 25.730 27.670 29.570 ;
        RECT 23.570 25.520 27.670 25.730 ;
        RECT 23.570 21.645 23.740 25.520 ;
        RECT 24.480 24.710 25.480 24.880 ;
        RECT 25.770 24.710 26.770 24.880 ;
        RECT 24.250 22.455 24.420 24.495 ;
        RECT 25.540 22.455 25.710 24.495 ;
        RECT 26.830 22.455 27.000 24.495 ;
        RECT 24.480 22.070 25.480 22.240 ;
        RECT 25.770 22.070 26.770 22.240 ;
        RECT 27.490 21.645 27.670 25.520 ;
        RECT 23.570 21.410 27.670 21.645 ;
        RECT 23.570 17.520 23.740 21.410 ;
        RECT 24.480 20.585 25.480 20.755 ;
        RECT 25.770 20.585 26.770 20.755 ;
        RECT 24.250 18.330 24.420 20.370 ;
        RECT 25.540 18.330 25.710 20.370 ;
        RECT 26.830 18.330 27.000 20.370 ;
        RECT 24.480 17.945 25.480 18.115 ;
        RECT 25.770 17.945 26.770 18.115 ;
        RECT 27.490 17.520 27.670 21.410 ;
        RECT 23.570 17.310 27.670 17.520 ;
        RECT 23.680 17.025 24.480 17.035 ;
        RECT 19.720 16.855 23.220 17.025 ;
        RECT 19.710 16.845 23.220 16.855 ;
        RECT 19.710 15.745 19.890 16.845 ;
        RECT 19.720 12.965 19.890 15.745 ;
        RECT 20.290 15.555 21.290 15.725 ;
        RECT 21.580 15.555 22.580 15.725 ;
        RECT 20.060 14.345 20.230 15.385 ;
        RECT 21.350 14.345 21.520 15.385 ;
        RECT 22.640 14.345 22.810 15.385 ;
        RECT 20.290 14.005 21.290 14.175 ;
        RECT 21.580 14.005 22.580 14.175 ;
        RECT 23.050 12.965 23.220 16.845 ;
        RECT 19.720 12.755 23.220 12.965 ;
        RECT 23.570 16.855 27.670 17.025 ;
        RECT 23.570 12.965 23.740 16.855 ;
        RECT 24.480 16.030 25.480 16.200 ;
        RECT 25.770 16.030 26.770 16.200 ;
        RECT 24.250 13.775 24.420 15.815 ;
        RECT 25.540 13.775 25.710 15.815 ;
        RECT 26.830 13.775 27.000 15.815 ;
        RECT 24.480 13.390 25.480 13.560 ;
        RECT 25.770 13.390 26.770 13.560 ;
        RECT 27.490 12.965 27.670 16.855 ;
        RECT 23.570 12.755 27.670 12.965 ;
      LAYER mcon ;
        RECT 20.370 141.720 21.210 141.890 ;
        RECT 21.660 141.720 22.500 141.890 ;
        RECT 20.060 140.590 20.230 141.470 ;
        RECT 21.350 140.590 21.520 141.470 ;
        RECT 22.640 140.590 22.810 141.470 ;
        RECT 20.370 140.170 21.210 140.340 ;
        RECT 21.660 140.170 22.500 140.340 ;
        RECT 19.720 139.260 19.890 139.700 ;
        RECT 20.370 137.720 21.210 137.890 ;
        RECT 21.660 137.720 22.500 137.890 ;
        RECT 20.060 136.590 20.230 137.470 ;
        RECT 21.350 136.590 21.520 137.470 ;
        RECT 22.640 136.590 22.810 137.470 ;
        RECT 20.370 136.170 21.210 136.340 ;
        RECT 21.660 136.170 22.500 136.340 ;
        RECT 19.720 135.260 19.890 135.700 ;
        RECT 20.370 133.620 21.210 133.790 ;
        RECT 21.660 133.620 22.500 133.790 ;
        RECT 20.060 132.490 20.230 133.370 ;
        RECT 21.350 132.490 21.520 133.370 ;
        RECT 22.640 132.490 22.810 133.370 ;
        RECT 20.370 132.070 21.210 132.240 ;
        RECT 21.660 132.070 22.500 132.240 ;
        RECT 19.720 131.160 19.890 131.600 ;
        RECT 20.370 129.570 21.210 129.740 ;
        RECT 21.660 129.570 22.500 129.740 ;
        RECT 20.060 128.440 20.230 129.320 ;
        RECT 21.350 128.440 21.520 129.320 ;
        RECT 22.640 128.440 22.810 129.320 ;
        RECT 20.370 128.020 21.210 128.190 ;
        RECT 21.660 128.020 22.500 128.190 ;
        RECT 19.720 127.110 19.890 127.550 ;
        RECT 20.370 125.520 21.210 125.690 ;
        RECT 21.660 125.520 22.500 125.690 ;
        RECT 20.060 124.390 20.230 125.270 ;
        RECT 21.350 124.390 21.520 125.270 ;
        RECT 22.640 124.390 22.810 125.270 ;
        RECT 20.370 123.970 21.210 124.140 ;
        RECT 21.660 123.970 22.500 124.140 ;
        RECT 19.720 123.060 19.890 123.500 ;
        RECT 20.370 121.470 21.210 121.640 ;
        RECT 21.660 121.470 22.500 121.640 ;
        RECT 20.060 120.340 20.230 121.220 ;
        RECT 21.350 120.340 21.520 121.220 ;
        RECT 22.640 120.340 22.810 121.220 ;
        RECT 20.370 119.920 21.210 120.090 ;
        RECT 21.660 119.920 22.500 120.090 ;
        RECT 19.720 119.010 19.890 119.450 ;
        RECT 20.370 117.420 21.210 117.590 ;
        RECT 21.660 117.420 22.500 117.590 ;
        RECT 20.060 116.290 20.230 117.170 ;
        RECT 21.350 116.290 21.520 117.170 ;
        RECT 22.640 116.290 22.810 117.170 ;
        RECT 20.370 115.870 21.210 116.040 ;
        RECT 21.660 115.870 22.500 116.040 ;
        RECT 19.720 114.960 19.890 115.400 ;
        RECT 20.370 113.370 21.210 113.540 ;
        RECT 21.660 113.370 22.500 113.540 ;
        RECT 20.060 112.240 20.230 113.120 ;
        RECT 21.350 112.240 21.520 113.120 ;
        RECT 22.640 112.240 22.810 113.120 ;
        RECT 20.370 111.820 21.210 111.990 ;
        RECT 21.660 111.820 22.500 111.990 ;
        RECT 19.720 110.910 19.890 111.350 ;
        RECT 20.370 109.320 21.210 109.490 ;
        RECT 21.660 109.320 22.500 109.490 ;
        RECT 20.060 108.190 20.230 109.070 ;
        RECT 21.350 108.190 21.520 109.070 ;
        RECT 22.640 108.190 22.810 109.070 ;
        RECT 20.370 107.770 21.210 107.940 ;
        RECT 21.660 107.770 22.500 107.940 ;
        RECT 19.720 106.860 19.890 107.300 ;
        RECT 20.370 105.270 21.210 105.440 ;
        RECT 21.660 105.270 22.500 105.440 ;
        RECT 20.060 104.140 20.230 105.020 ;
        RECT 21.350 104.140 21.520 105.020 ;
        RECT 22.640 104.140 22.810 105.020 ;
        RECT 20.370 103.720 21.210 103.890 ;
        RECT 21.660 103.720 22.500 103.890 ;
        RECT 19.720 102.810 19.890 103.250 ;
        RECT 20.370 101.220 21.210 101.390 ;
        RECT 21.660 101.220 22.500 101.390 ;
        RECT 20.060 100.090 20.230 100.970 ;
        RECT 21.350 100.090 21.520 100.970 ;
        RECT 22.640 100.090 22.810 100.970 ;
        RECT 20.370 99.670 21.210 99.840 ;
        RECT 21.660 99.670 22.500 99.840 ;
        RECT 19.720 98.760 19.890 99.200 ;
        RECT 20.370 97.170 21.210 97.340 ;
        RECT 21.660 97.170 22.500 97.340 ;
        RECT 20.060 96.040 20.230 96.920 ;
        RECT 21.350 96.040 21.520 96.920 ;
        RECT 22.640 96.040 22.810 96.920 ;
        RECT 20.370 95.620 21.210 95.790 ;
        RECT 21.660 95.620 22.500 95.790 ;
        RECT 19.720 94.710 19.890 95.150 ;
        RECT 20.370 93.120 21.210 93.290 ;
        RECT 21.660 93.120 22.500 93.290 ;
        RECT 20.060 91.990 20.230 92.870 ;
        RECT 21.350 91.990 21.520 92.870 ;
        RECT 22.640 91.990 22.810 92.870 ;
        RECT 20.370 91.570 21.210 91.740 ;
        RECT 21.660 91.570 22.500 91.740 ;
        RECT 19.720 90.660 19.890 91.100 ;
        RECT 20.370 89.070 21.210 89.240 ;
        RECT 21.660 89.070 22.500 89.240 ;
        RECT 20.060 87.940 20.230 88.820 ;
        RECT 21.350 87.940 21.520 88.820 ;
        RECT 22.640 87.940 22.810 88.820 ;
        RECT 20.370 87.520 21.210 87.690 ;
        RECT 21.660 87.520 22.500 87.690 ;
        RECT 19.720 86.610 19.890 87.050 ;
        RECT 20.370 85.020 21.210 85.190 ;
        RECT 21.660 85.020 22.500 85.190 ;
        RECT 20.060 83.890 20.230 84.770 ;
        RECT 21.350 83.890 21.520 84.770 ;
        RECT 22.640 83.890 22.810 84.770 ;
        RECT 20.370 83.470 21.210 83.640 ;
        RECT 21.660 83.470 22.500 83.640 ;
        RECT 19.720 82.560 19.890 83.000 ;
        RECT 20.370 80.970 21.210 81.140 ;
        RECT 21.660 80.970 22.500 81.140 ;
        RECT 20.060 79.840 20.230 80.720 ;
        RECT 21.350 79.840 21.520 80.720 ;
        RECT 22.640 79.840 22.810 80.720 ;
        RECT 20.370 79.420 21.210 79.590 ;
        RECT 21.660 79.420 22.500 79.590 ;
        RECT 19.720 78.510 19.890 78.950 ;
        RECT 20.370 76.920 21.210 77.090 ;
        RECT 21.660 76.920 22.500 77.090 ;
        RECT 20.060 75.790 20.230 76.670 ;
        RECT 21.350 75.790 21.520 76.670 ;
        RECT 22.640 75.790 22.810 76.670 ;
        RECT 20.370 75.370 21.210 75.540 ;
        RECT 21.660 75.370 22.500 75.540 ;
        RECT 19.720 74.460 19.890 74.900 ;
        RECT 20.370 72.870 21.210 73.040 ;
        RECT 21.660 72.870 22.500 73.040 ;
        RECT 20.060 71.740 20.230 72.620 ;
        RECT 21.350 71.740 21.520 72.620 ;
        RECT 22.640 71.740 22.810 72.620 ;
        RECT 20.370 71.320 21.210 71.490 ;
        RECT 21.660 71.320 22.500 71.490 ;
        RECT 19.720 70.410 19.890 70.850 ;
        RECT 20.370 68.820 21.210 68.990 ;
        RECT 21.660 68.820 22.500 68.990 ;
        RECT 20.060 67.690 20.230 68.570 ;
        RECT 21.350 67.690 21.520 68.570 ;
        RECT 22.640 67.690 22.810 68.570 ;
        RECT 20.370 67.270 21.210 67.440 ;
        RECT 21.660 67.270 22.500 67.440 ;
        RECT 19.720 66.360 19.890 66.800 ;
        RECT 20.370 64.770 21.210 64.940 ;
        RECT 21.660 64.770 22.500 64.940 ;
        RECT 20.060 63.640 20.230 64.520 ;
        RECT 21.350 63.640 21.520 64.520 ;
        RECT 22.640 63.640 22.810 64.520 ;
        RECT 20.370 63.220 21.210 63.390 ;
        RECT 21.660 63.220 22.500 63.390 ;
        RECT 19.720 62.310 19.890 62.750 ;
        RECT 20.370 60.720 21.210 60.890 ;
        RECT 21.660 60.720 22.500 60.890 ;
        RECT 20.060 59.590 20.230 60.470 ;
        RECT 21.350 59.590 21.520 60.470 ;
        RECT 22.640 59.590 22.810 60.470 ;
        RECT 20.370 59.170 21.210 59.340 ;
        RECT 21.660 59.170 22.500 59.340 ;
        RECT 19.720 58.260 19.890 58.700 ;
        RECT 20.370 56.670 21.210 56.840 ;
        RECT 21.660 56.670 22.500 56.840 ;
        RECT 20.060 55.540 20.230 56.420 ;
        RECT 21.350 55.540 21.520 56.420 ;
        RECT 22.640 55.540 22.810 56.420 ;
        RECT 20.370 55.120 21.210 55.290 ;
        RECT 21.660 55.120 22.500 55.290 ;
        RECT 19.720 54.210 19.890 54.650 ;
        RECT 20.370 52.620 21.210 52.790 ;
        RECT 21.660 52.620 22.500 52.790 ;
        RECT 20.060 51.490 20.230 52.370 ;
        RECT 21.350 51.490 21.520 52.370 ;
        RECT 22.640 51.490 22.810 52.370 ;
        RECT 20.370 51.070 21.210 51.240 ;
        RECT 21.660 51.070 22.500 51.240 ;
        RECT 19.720 50.160 19.890 50.600 ;
        RECT 20.370 48.570 21.210 48.740 ;
        RECT 21.660 48.570 22.500 48.740 ;
        RECT 20.060 47.440 20.230 48.320 ;
        RECT 21.350 47.440 21.520 48.320 ;
        RECT 22.640 47.440 22.810 48.320 ;
        RECT 20.370 47.020 21.210 47.190 ;
        RECT 21.660 47.020 22.500 47.190 ;
        RECT 19.720 46.110 19.890 46.550 ;
        RECT 20.370 44.520 21.210 44.690 ;
        RECT 21.660 44.520 22.500 44.690 ;
        RECT 20.060 43.390 20.230 44.270 ;
        RECT 21.350 43.390 21.520 44.270 ;
        RECT 22.640 43.390 22.810 44.270 ;
        RECT 20.370 42.970 21.210 43.140 ;
        RECT 21.660 42.970 22.500 43.140 ;
        RECT 19.720 42.060 19.890 42.500 ;
        RECT 20.370 40.470 21.210 40.640 ;
        RECT 21.660 40.470 22.500 40.640 ;
        RECT 20.060 39.340 20.230 40.220 ;
        RECT 21.350 39.340 21.520 40.220 ;
        RECT 22.640 39.340 22.810 40.220 ;
        RECT 20.370 38.920 21.210 39.090 ;
        RECT 21.660 38.920 22.500 39.090 ;
        RECT 19.720 38.010 19.890 38.450 ;
        RECT 20.370 36.420 21.210 36.590 ;
        RECT 21.660 36.420 22.500 36.590 ;
        RECT 20.060 35.290 20.230 36.170 ;
        RECT 21.350 35.290 21.520 36.170 ;
        RECT 22.640 35.290 22.810 36.170 ;
        RECT 20.370 34.870 21.210 35.040 ;
        RECT 21.660 34.870 22.500 35.040 ;
        RECT 19.720 33.960 19.890 34.400 ;
        RECT 20.370 32.370 21.210 32.540 ;
        RECT 21.660 32.370 22.500 32.540 ;
        RECT 20.060 31.240 20.230 32.120 ;
        RECT 21.350 31.240 21.520 32.120 ;
        RECT 22.640 31.240 22.810 32.120 ;
        RECT 20.370 30.820 21.210 30.990 ;
        RECT 21.660 30.820 22.500 30.990 ;
        RECT 19.720 29.910 19.890 30.350 ;
        RECT 20.370 28.320 21.210 28.490 ;
        RECT 21.660 28.320 22.500 28.490 ;
        RECT 20.060 27.190 20.230 28.070 ;
        RECT 21.350 27.190 21.520 28.070 ;
        RECT 22.640 27.190 22.810 28.070 ;
        RECT 20.370 26.770 21.210 26.940 ;
        RECT 21.660 26.770 22.500 26.940 ;
        RECT 19.720 25.860 19.890 26.300 ;
        RECT 20.370 24.235 21.210 24.405 ;
        RECT 21.660 24.235 22.500 24.405 ;
        RECT 20.060 23.105 20.230 23.985 ;
        RECT 21.350 23.105 21.520 23.985 ;
        RECT 22.640 23.105 22.810 23.985 ;
        RECT 20.370 22.685 21.210 22.855 ;
        RECT 21.660 22.685 22.500 22.855 ;
        RECT 19.720 21.775 19.890 22.215 ;
        RECT 20.370 20.110 21.210 20.280 ;
        RECT 21.660 20.110 22.500 20.280 ;
        RECT 20.060 18.980 20.230 19.860 ;
        RECT 21.350 18.980 21.520 19.860 ;
        RECT 22.640 18.980 22.810 19.860 ;
        RECT 20.370 18.560 21.210 18.730 ;
        RECT 21.660 18.560 22.500 18.730 ;
        RECT 19.720 17.650 19.890 18.090 ;
        RECT 24.560 142.195 25.400 142.365 ;
        RECT 25.850 142.195 26.690 142.365 ;
        RECT 24.250 140.020 24.420 141.900 ;
        RECT 25.540 140.020 25.710 141.900 ;
        RECT 26.830 140.020 27.000 141.900 ;
        RECT 24.560 139.555 25.400 139.725 ;
        RECT 25.850 139.555 26.690 139.725 ;
        RECT 27.490 139.220 27.670 142.890 ;
        RECT 24.560 138.195 25.400 138.365 ;
        RECT 25.850 138.195 26.690 138.365 ;
        RECT 24.250 136.020 24.420 137.900 ;
        RECT 25.540 136.020 25.710 137.900 ;
        RECT 26.830 136.020 27.000 137.900 ;
        RECT 24.560 135.555 25.400 135.725 ;
        RECT 25.850 135.555 26.690 135.725 ;
        RECT 27.490 135.220 27.670 138.890 ;
        RECT 24.560 134.095 25.400 134.265 ;
        RECT 25.850 134.095 26.690 134.265 ;
        RECT 24.250 131.920 24.420 133.800 ;
        RECT 25.540 131.920 25.710 133.800 ;
        RECT 26.830 131.920 27.000 133.800 ;
        RECT 24.560 131.455 25.400 131.625 ;
        RECT 25.850 131.455 26.690 131.625 ;
        RECT 27.490 131.120 27.670 134.790 ;
        RECT 24.560 130.045 25.400 130.215 ;
        RECT 25.850 130.045 26.690 130.215 ;
        RECT 24.250 127.870 24.420 129.750 ;
        RECT 25.540 127.870 25.710 129.750 ;
        RECT 26.830 127.870 27.000 129.750 ;
        RECT 24.560 127.405 25.400 127.575 ;
        RECT 25.850 127.405 26.690 127.575 ;
        RECT 27.490 127.070 27.670 130.740 ;
        RECT 24.560 125.995 25.400 126.165 ;
        RECT 25.850 125.995 26.690 126.165 ;
        RECT 24.250 123.820 24.420 125.700 ;
        RECT 25.540 123.820 25.710 125.700 ;
        RECT 26.830 123.820 27.000 125.700 ;
        RECT 24.560 123.355 25.400 123.525 ;
        RECT 25.850 123.355 26.690 123.525 ;
        RECT 27.490 123.020 27.670 126.690 ;
        RECT 24.560 121.945 25.400 122.115 ;
        RECT 25.850 121.945 26.690 122.115 ;
        RECT 24.250 119.770 24.420 121.650 ;
        RECT 25.540 119.770 25.710 121.650 ;
        RECT 26.830 119.770 27.000 121.650 ;
        RECT 24.560 119.305 25.400 119.475 ;
        RECT 25.850 119.305 26.690 119.475 ;
        RECT 27.490 118.970 27.670 122.640 ;
        RECT 24.560 117.895 25.400 118.065 ;
        RECT 25.850 117.895 26.690 118.065 ;
        RECT 24.250 115.720 24.420 117.600 ;
        RECT 25.540 115.720 25.710 117.600 ;
        RECT 26.830 115.720 27.000 117.600 ;
        RECT 24.560 115.255 25.400 115.425 ;
        RECT 25.850 115.255 26.690 115.425 ;
        RECT 27.490 114.920 27.670 118.590 ;
        RECT 24.560 113.845 25.400 114.015 ;
        RECT 25.850 113.845 26.690 114.015 ;
        RECT 24.250 111.670 24.420 113.550 ;
        RECT 25.540 111.670 25.710 113.550 ;
        RECT 26.830 111.670 27.000 113.550 ;
        RECT 24.560 111.205 25.400 111.375 ;
        RECT 25.850 111.205 26.690 111.375 ;
        RECT 27.490 110.870 27.670 114.540 ;
        RECT 24.560 109.795 25.400 109.965 ;
        RECT 25.850 109.795 26.690 109.965 ;
        RECT 24.250 107.620 24.420 109.500 ;
        RECT 25.540 107.620 25.710 109.500 ;
        RECT 26.830 107.620 27.000 109.500 ;
        RECT 24.560 107.155 25.400 107.325 ;
        RECT 25.850 107.155 26.690 107.325 ;
        RECT 27.490 106.820 27.670 110.490 ;
        RECT 24.560 105.745 25.400 105.915 ;
        RECT 25.850 105.745 26.690 105.915 ;
        RECT 24.250 103.570 24.420 105.450 ;
        RECT 25.540 103.570 25.710 105.450 ;
        RECT 26.830 103.570 27.000 105.450 ;
        RECT 24.560 103.105 25.400 103.275 ;
        RECT 25.850 103.105 26.690 103.275 ;
        RECT 27.490 102.770 27.670 106.440 ;
        RECT 24.560 101.695 25.400 101.865 ;
        RECT 25.850 101.695 26.690 101.865 ;
        RECT 24.250 99.520 24.420 101.400 ;
        RECT 25.540 99.520 25.710 101.400 ;
        RECT 26.830 99.520 27.000 101.400 ;
        RECT 24.560 99.055 25.400 99.225 ;
        RECT 25.850 99.055 26.690 99.225 ;
        RECT 27.490 98.720 27.670 102.390 ;
        RECT 24.560 97.645 25.400 97.815 ;
        RECT 25.850 97.645 26.690 97.815 ;
        RECT 24.250 95.470 24.420 97.350 ;
        RECT 25.540 95.470 25.710 97.350 ;
        RECT 26.830 95.470 27.000 97.350 ;
        RECT 24.560 95.005 25.400 95.175 ;
        RECT 25.850 95.005 26.690 95.175 ;
        RECT 27.490 94.670 27.670 98.340 ;
        RECT 24.560 93.595 25.400 93.765 ;
        RECT 25.850 93.595 26.690 93.765 ;
        RECT 24.250 91.420 24.420 93.300 ;
        RECT 25.540 91.420 25.710 93.300 ;
        RECT 26.830 91.420 27.000 93.300 ;
        RECT 24.560 90.955 25.400 91.125 ;
        RECT 25.850 90.955 26.690 91.125 ;
        RECT 27.490 90.620 27.670 94.290 ;
        RECT 24.560 89.545 25.400 89.715 ;
        RECT 25.850 89.545 26.690 89.715 ;
        RECT 24.250 87.370 24.420 89.250 ;
        RECT 25.540 87.370 25.710 89.250 ;
        RECT 26.830 87.370 27.000 89.250 ;
        RECT 24.560 86.905 25.400 87.075 ;
        RECT 25.850 86.905 26.690 87.075 ;
        RECT 27.490 86.570 27.670 90.240 ;
        RECT 24.560 85.495 25.400 85.665 ;
        RECT 25.850 85.495 26.690 85.665 ;
        RECT 24.250 83.320 24.420 85.200 ;
        RECT 25.540 83.320 25.710 85.200 ;
        RECT 26.830 83.320 27.000 85.200 ;
        RECT 24.560 82.855 25.400 83.025 ;
        RECT 25.850 82.855 26.690 83.025 ;
        RECT 27.490 82.520 27.670 86.190 ;
        RECT 24.560 81.445 25.400 81.615 ;
        RECT 25.850 81.445 26.690 81.615 ;
        RECT 24.250 79.270 24.420 81.150 ;
        RECT 25.540 79.270 25.710 81.150 ;
        RECT 26.830 79.270 27.000 81.150 ;
        RECT 24.560 78.805 25.400 78.975 ;
        RECT 25.850 78.805 26.690 78.975 ;
        RECT 27.490 78.470 27.670 82.140 ;
        RECT 24.560 77.395 25.400 77.565 ;
        RECT 25.850 77.395 26.690 77.565 ;
        RECT 24.250 75.220 24.420 77.100 ;
        RECT 25.540 75.220 25.710 77.100 ;
        RECT 26.830 75.220 27.000 77.100 ;
        RECT 24.560 74.755 25.400 74.925 ;
        RECT 25.850 74.755 26.690 74.925 ;
        RECT 27.490 74.420 27.670 78.090 ;
        RECT 24.560 73.345 25.400 73.515 ;
        RECT 25.850 73.345 26.690 73.515 ;
        RECT 24.250 71.170 24.420 73.050 ;
        RECT 25.540 71.170 25.710 73.050 ;
        RECT 26.830 71.170 27.000 73.050 ;
        RECT 24.560 70.705 25.400 70.875 ;
        RECT 25.850 70.705 26.690 70.875 ;
        RECT 27.490 70.370 27.670 74.040 ;
        RECT 24.560 69.295 25.400 69.465 ;
        RECT 25.850 69.295 26.690 69.465 ;
        RECT 24.250 67.120 24.420 69.000 ;
        RECT 25.540 67.120 25.710 69.000 ;
        RECT 26.830 67.120 27.000 69.000 ;
        RECT 24.560 66.655 25.400 66.825 ;
        RECT 25.850 66.655 26.690 66.825 ;
        RECT 27.490 66.320 27.670 69.990 ;
        RECT 24.560 65.245 25.400 65.415 ;
        RECT 25.850 65.245 26.690 65.415 ;
        RECT 24.250 63.070 24.420 64.950 ;
        RECT 25.540 63.070 25.710 64.950 ;
        RECT 26.830 63.070 27.000 64.950 ;
        RECT 24.560 62.605 25.400 62.775 ;
        RECT 25.850 62.605 26.690 62.775 ;
        RECT 27.490 62.270 27.670 65.940 ;
        RECT 24.560 61.195 25.400 61.365 ;
        RECT 25.850 61.195 26.690 61.365 ;
        RECT 24.250 59.020 24.420 60.900 ;
        RECT 25.540 59.020 25.710 60.900 ;
        RECT 26.830 59.020 27.000 60.900 ;
        RECT 24.560 58.555 25.400 58.725 ;
        RECT 25.850 58.555 26.690 58.725 ;
        RECT 27.490 58.220 27.670 61.890 ;
        RECT 24.560 57.145 25.400 57.315 ;
        RECT 25.850 57.145 26.690 57.315 ;
        RECT 24.250 54.970 24.420 56.850 ;
        RECT 25.540 54.970 25.710 56.850 ;
        RECT 26.830 54.970 27.000 56.850 ;
        RECT 24.560 54.505 25.400 54.675 ;
        RECT 25.850 54.505 26.690 54.675 ;
        RECT 27.490 54.170 27.670 57.840 ;
        RECT 28.010 139.220 28.190 142.890 ;
        RECT 28.990 142.195 29.830 142.365 ;
        RECT 30.280 142.195 31.120 142.365 ;
        RECT 28.680 140.020 28.850 141.900 ;
        RECT 29.970 140.020 30.140 141.900 ;
        RECT 31.260 140.020 31.430 141.900 ;
        RECT 28.990 139.555 29.830 139.725 ;
        RECT 30.280 139.555 31.120 139.725 ;
        RECT 28.010 135.160 28.190 138.830 ;
        RECT 28.990 138.135 29.830 138.305 ;
        RECT 30.280 138.135 31.120 138.305 ;
        RECT 28.680 135.960 28.850 137.840 ;
        RECT 29.970 135.960 30.140 137.840 ;
        RECT 31.260 135.960 31.430 137.840 ;
        RECT 28.990 135.495 29.830 135.665 ;
        RECT 30.280 135.495 31.120 135.665 ;
        RECT 28.010 131.100 28.190 134.770 ;
        RECT 28.990 134.075 29.830 134.245 ;
        RECT 30.280 134.075 31.120 134.245 ;
        RECT 28.680 131.900 28.850 133.780 ;
        RECT 29.970 131.900 30.140 133.780 ;
        RECT 31.260 131.900 31.430 133.780 ;
        RECT 28.990 131.435 29.830 131.605 ;
        RECT 30.280 131.435 31.120 131.605 ;
        RECT 28.010 127.040 28.190 130.710 ;
        RECT 28.990 130.015 29.830 130.185 ;
        RECT 30.280 130.015 31.120 130.185 ;
        RECT 28.680 127.840 28.850 129.720 ;
        RECT 29.970 127.840 30.140 129.720 ;
        RECT 31.260 127.840 31.430 129.720 ;
        RECT 28.990 127.375 29.830 127.545 ;
        RECT 30.280 127.375 31.120 127.545 ;
        RECT 28.010 122.980 28.190 126.650 ;
        RECT 28.990 125.955 29.830 126.125 ;
        RECT 30.280 125.955 31.120 126.125 ;
        RECT 28.680 123.780 28.850 125.660 ;
        RECT 29.970 123.780 30.140 125.660 ;
        RECT 31.260 123.780 31.430 125.660 ;
        RECT 28.990 123.315 29.830 123.485 ;
        RECT 30.280 123.315 31.120 123.485 ;
        RECT 28.010 118.920 28.190 122.590 ;
        RECT 28.990 121.895 29.830 122.065 ;
        RECT 30.280 121.895 31.120 122.065 ;
        RECT 28.680 119.720 28.850 121.600 ;
        RECT 29.970 119.720 30.140 121.600 ;
        RECT 31.260 119.720 31.430 121.600 ;
        RECT 28.990 119.255 29.830 119.425 ;
        RECT 30.280 119.255 31.120 119.425 ;
        RECT 28.010 114.860 28.190 118.530 ;
        RECT 28.990 117.835 29.830 118.005 ;
        RECT 30.280 117.835 31.120 118.005 ;
        RECT 28.680 115.660 28.850 117.540 ;
        RECT 29.970 115.660 30.140 117.540 ;
        RECT 31.260 115.660 31.430 117.540 ;
        RECT 28.990 115.195 29.830 115.365 ;
        RECT 30.280 115.195 31.120 115.365 ;
        RECT 28.010 110.800 28.190 114.470 ;
        RECT 28.990 113.775 29.830 113.945 ;
        RECT 30.280 113.775 31.120 113.945 ;
        RECT 28.680 111.600 28.850 113.480 ;
        RECT 29.970 111.600 30.140 113.480 ;
        RECT 31.260 111.600 31.430 113.480 ;
        RECT 28.990 111.135 29.830 111.305 ;
        RECT 30.280 111.135 31.120 111.305 ;
        RECT 28.010 106.740 28.190 110.410 ;
        RECT 28.990 109.715 29.830 109.885 ;
        RECT 30.280 109.715 31.120 109.885 ;
        RECT 28.680 107.540 28.850 109.420 ;
        RECT 29.970 107.540 30.140 109.420 ;
        RECT 31.260 107.540 31.430 109.420 ;
        RECT 28.990 107.075 29.830 107.245 ;
        RECT 30.280 107.075 31.120 107.245 ;
        RECT 28.010 102.680 28.190 106.350 ;
        RECT 28.990 105.655 29.830 105.825 ;
        RECT 30.280 105.655 31.120 105.825 ;
        RECT 28.680 103.480 28.850 105.360 ;
        RECT 29.970 103.480 30.140 105.360 ;
        RECT 31.260 103.480 31.430 105.360 ;
        RECT 28.990 103.015 29.830 103.185 ;
        RECT 30.280 103.015 31.120 103.185 ;
        RECT 28.010 98.620 28.190 102.290 ;
        RECT 28.990 101.595 29.830 101.765 ;
        RECT 30.280 101.595 31.120 101.765 ;
        RECT 28.680 99.420 28.850 101.300 ;
        RECT 29.970 99.420 30.140 101.300 ;
        RECT 31.260 99.420 31.430 101.300 ;
        RECT 28.990 98.955 29.830 99.125 ;
        RECT 30.280 98.955 31.120 99.125 ;
        RECT 28.010 94.560 28.190 98.230 ;
        RECT 28.990 97.535 29.830 97.705 ;
        RECT 30.280 97.535 31.120 97.705 ;
        RECT 28.680 95.360 28.850 97.240 ;
        RECT 29.970 95.360 30.140 97.240 ;
        RECT 31.260 95.360 31.430 97.240 ;
        RECT 28.990 94.895 29.830 95.065 ;
        RECT 30.280 94.895 31.120 95.065 ;
        RECT 28.010 90.500 28.190 94.170 ;
        RECT 28.990 93.475 29.830 93.645 ;
        RECT 30.280 93.475 31.120 93.645 ;
        RECT 28.680 91.300 28.850 93.180 ;
        RECT 29.970 91.300 30.140 93.180 ;
        RECT 31.260 91.300 31.430 93.180 ;
        RECT 28.990 90.835 29.830 91.005 ;
        RECT 30.280 90.835 31.120 91.005 ;
        RECT 28.010 86.440 28.190 90.110 ;
        RECT 28.990 89.415 29.830 89.585 ;
        RECT 30.280 89.415 31.120 89.585 ;
        RECT 28.680 87.240 28.850 89.120 ;
        RECT 29.970 87.240 30.140 89.120 ;
        RECT 31.260 87.240 31.430 89.120 ;
        RECT 28.990 86.775 29.830 86.945 ;
        RECT 30.280 86.775 31.120 86.945 ;
        RECT 28.010 82.380 28.190 86.050 ;
        RECT 28.990 85.355 29.830 85.525 ;
        RECT 30.280 85.355 31.120 85.525 ;
        RECT 28.680 83.180 28.850 85.060 ;
        RECT 29.970 83.180 30.140 85.060 ;
        RECT 31.260 83.180 31.430 85.060 ;
        RECT 28.990 82.715 29.830 82.885 ;
        RECT 30.280 82.715 31.120 82.885 ;
        RECT 28.010 78.320 28.190 81.990 ;
        RECT 28.990 81.295 29.830 81.465 ;
        RECT 30.280 81.295 31.120 81.465 ;
        RECT 28.680 79.120 28.850 81.000 ;
        RECT 29.970 79.120 30.140 81.000 ;
        RECT 31.260 79.120 31.430 81.000 ;
        RECT 28.990 78.655 29.830 78.825 ;
        RECT 30.280 78.655 31.120 78.825 ;
        RECT 28.010 74.260 28.190 77.930 ;
        RECT 28.990 77.235 29.830 77.405 ;
        RECT 30.280 77.235 31.120 77.405 ;
        RECT 28.680 75.060 28.850 76.940 ;
        RECT 29.970 75.060 30.140 76.940 ;
        RECT 31.260 75.060 31.430 76.940 ;
        RECT 28.990 74.595 29.830 74.765 ;
        RECT 30.280 74.595 31.120 74.765 ;
        RECT 28.010 70.200 28.190 73.870 ;
        RECT 28.990 73.175 29.830 73.345 ;
        RECT 30.280 73.175 31.120 73.345 ;
        RECT 28.680 71.000 28.850 72.880 ;
        RECT 29.970 71.000 30.140 72.880 ;
        RECT 31.260 71.000 31.430 72.880 ;
        RECT 28.990 70.535 29.830 70.705 ;
        RECT 30.280 70.535 31.120 70.705 ;
        RECT 28.010 66.140 28.190 69.810 ;
        RECT 28.990 69.115 29.830 69.285 ;
        RECT 30.280 69.115 31.120 69.285 ;
        RECT 28.680 66.940 28.850 68.820 ;
        RECT 29.970 66.940 30.140 68.820 ;
        RECT 31.260 66.940 31.430 68.820 ;
        RECT 28.990 66.475 29.830 66.645 ;
        RECT 30.280 66.475 31.120 66.645 ;
        RECT 28.010 62.080 28.190 65.750 ;
        RECT 28.990 65.055 29.830 65.225 ;
        RECT 30.280 65.055 31.120 65.225 ;
        RECT 28.680 62.880 28.850 64.760 ;
        RECT 29.970 62.880 30.140 64.760 ;
        RECT 31.260 62.880 31.430 64.760 ;
        RECT 28.990 62.415 29.830 62.585 ;
        RECT 30.280 62.415 31.120 62.585 ;
        RECT 28.010 58.020 28.190 61.690 ;
        RECT 28.990 60.995 29.830 61.165 ;
        RECT 30.280 60.995 31.120 61.165 ;
        RECT 28.680 58.820 28.850 60.700 ;
        RECT 29.970 58.820 30.140 60.700 ;
        RECT 31.260 58.820 31.430 60.700 ;
        RECT 28.990 58.355 29.830 58.525 ;
        RECT 30.280 58.355 31.120 58.525 ;
        RECT 33.180 141.720 34.020 141.890 ;
        RECT 34.470 141.720 35.310 141.890 ;
        RECT 32.870 140.590 33.040 141.470 ;
        RECT 34.160 140.590 34.330 141.470 ;
        RECT 35.450 140.590 35.620 141.470 ;
        RECT 33.180 140.170 34.020 140.340 ;
        RECT 34.470 140.170 35.310 140.340 ;
        RECT 35.790 139.260 35.960 139.700 ;
        RECT 33.180 137.660 34.020 137.830 ;
        RECT 34.470 137.660 35.310 137.830 ;
        RECT 32.870 136.530 33.040 137.410 ;
        RECT 34.160 136.530 34.330 137.410 ;
        RECT 35.450 136.530 35.620 137.410 ;
        RECT 33.180 136.110 34.020 136.280 ;
        RECT 34.470 136.110 35.310 136.280 ;
        RECT 35.790 135.200 35.960 135.640 ;
        RECT 33.180 133.600 34.020 133.770 ;
        RECT 34.470 133.600 35.310 133.770 ;
        RECT 32.870 132.470 33.040 133.350 ;
        RECT 34.160 132.470 34.330 133.350 ;
        RECT 35.450 132.470 35.620 133.350 ;
        RECT 33.180 132.050 34.020 132.220 ;
        RECT 34.470 132.050 35.310 132.220 ;
        RECT 35.790 131.140 35.960 131.580 ;
        RECT 33.180 129.540 34.020 129.710 ;
        RECT 34.470 129.540 35.310 129.710 ;
        RECT 32.870 128.410 33.040 129.290 ;
        RECT 34.160 128.410 34.330 129.290 ;
        RECT 35.450 128.410 35.620 129.290 ;
        RECT 33.180 127.990 34.020 128.160 ;
        RECT 34.470 127.990 35.310 128.160 ;
        RECT 35.790 127.080 35.960 127.520 ;
        RECT 33.180 125.480 34.020 125.650 ;
        RECT 34.470 125.480 35.310 125.650 ;
        RECT 32.870 124.350 33.040 125.230 ;
        RECT 34.160 124.350 34.330 125.230 ;
        RECT 35.450 124.350 35.620 125.230 ;
        RECT 33.180 123.930 34.020 124.100 ;
        RECT 34.470 123.930 35.310 124.100 ;
        RECT 35.790 123.020 35.960 123.460 ;
        RECT 33.180 121.420 34.020 121.590 ;
        RECT 34.470 121.420 35.310 121.590 ;
        RECT 32.870 120.290 33.040 121.170 ;
        RECT 34.160 120.290 34.330 121.170 ;
        RECT 35.450 120.290 35.620 121.170 ;
        RECT 33.180 119.870 34.020 120.040 ;
        RECT 34.470 119.870 35.310 120.040 ;
        RECT 35.790 118.960 35.960 119.400 ;
        RECT 33.180 117.360 34.020 117.530 ;
        RECT 34.470 117.360 35.310 117.530 ;
        RECT 32.870 116.230 33.040 117.110 ;
        RECT 34.160 116.230 34.330 117.110 ;
        RECT 35.450 116.230 35.620 117.110 ;
        RECT 33.180 115.810 34.020 115.980 ;
        RECT 34.470 115.810 35.310 115.980 ;
        RECT 35.790 114.900 35.960 115.340 ;
        RECT 33.180 113.300 34.020 113.470 ;
        RECT 34.470 113.300 35.310 113.470 ;
        RECT 32.870 112.170 33.040 113.050 ;
        RECT 34.160 112.170 34.330 113.050 ;
        RECT 35.450 112.170 35.620 113.050 ;
        RECT 33.180 111.750 34.020 111.920 ;
        RECT 34.470 111.750 35.310 111.920 ;
        RECT 35.790 110.840 35.960 111.280 ;
        RECT 33.180 109.240 34.020 109.410 ;
        RECT 34.470 109.240 35.310 109.410 ;
        RECT 32.870 108.110 33.040 108.990 ;
        RECT 34.160 108.110 34.330 108.990 ;
        RECT 35.450 108.110 35.620 108.990 ;
        RECT 33.180 107.690 34.020 107.860 ;
        RECT 34.470 107.690 35.310 107.860 ;
        RECT 35.790 106.780 35.960 107.220 ;
        RECT 33.180 105.180 34.020 105.350 ;
        RECT 34.470 105.180 35.310 105.350 ;
        RECT 32.870 104.050 33.040 104.930 ;
        RECT 34.160 104.050 34.330 104.930 ;
        RECT 35.450 104.050 35.620 104.930 ;
        RECT 33.180 103.630 34.020 103.800 ;
        RECT 34.470 103.630 35.310 103.800 ;
        RECT 35.790 102.720 35.960 103.160 ;
        RECT 33.180 101.120 34.020 101.290 ;
        RECT 34.470 101.120 35.310 101.290 ;
        RECT 32.870 99.990 33.040 100.870 ;
        RECT 34.160 99.990 34.330 100.870 ;
        RECT 35.450 99.990 35.620 100.870 ;
        RECT 33.180 99.570 34.020 99.740 ;
        RECT 34.470 99.570 35.310 99.740 ;
        RECT 35.790 98.660 35.960 99.100 ;
        RECT 33.180 97.060 34.020 97.230 ;
        RECT 34.470 97.060 35.310 97.230 ;
        RECT 32.870 95.930 33.040 96.810 ;
        RECT 34.160 95.930 34.330 96.810 ;
        RECT 35.450 95.930 35.620 96.810 ;
        RECT 33.180 95.510 34.020 95.680 ;
        RECT 34.470 95.510 35.310 95.680 ;
        RECT 35.790 94.600 35.960 95.040 ;
        RECT 33.180 93.000 34.020 93.170 ;
        RECT 34.470 93.000 35.310 93.170 ;
        RECT 32.870 91.870 33.040 92.750 ;
        RECT 34.160 91.870 34.330 92.750 ;
        RECT 35.450 91.870 35.620 92.750 ;
        RECT 33.180 91.450 34.020 91.620 ;
        RECT 34.470 91.450 35.310 91.620 ;
        RECT 35.790 90.540 35.960 90.980 ;
        RECT 33.180 88.940 34.020 89.110 ;
        RECT 34.470 88.940 35.310 89.110 ;
        RECT 32.870 87.810 33.040 88.690 ;
        RECT 34.160 87.810 34.330 88.690 ;
        RECT 35.450 87.810 35.620 88.690 ;
        RECT 33.180 87.390 34.020 87.560 ;
        RECT 34.470 87.390 35.310 87.560 ;
        RECT 35.790 86.480 35.960 86.920 ;
        RECT 33.180 84.880 34.020 85.050 ;
        RECT 34.470 84.880 35.310 85.050 ;
        RECT 32.870 83.750 33.040 84.630 ;
        RECT 34.160 83.750 34.330 84.630 ;
        RECT 35.450 83.750 35.620 84.630 ;
        RECT 33.180 83.330 34.020 83.500 ;
        RECT 34.470 83.330 35.310 83.500 ;
        RECT 35.790 82.420 35.960 82.860 ;
        RECT 33.180 80.820 34.020 80.990 ;
        RECT 34.470 80.820 35.310 80.990 ;
        RECT 32.870 79.690 33.040 80.570 ;
        RECT 34.160 79.690 34.330 80.570 ;
        RECT 35.450 79.690 35.620 80.570 ;
        RECT 33.180 79.270 34.020 79.440 ;
        RECT 34.470 79.270 35.310 79.440 ;
        RECT 35.790 78.360 35.960 78.800 ;
        RECT 33.180 76.760 34.020 76.930 ;
        RECT 34.470 76.760 35.310 76.930 ;
        RECT 32.870 75.630 33.040 76.510 ;
        RECT 34.160 75.630 34.330 76.510 ;
        RECT 35.450 75.630 35.620 76.510 ;
        RECT 33.180 75.210 34.020 75.380 ;
        RECT 34.470 75.210 35.310 75.380 ;
        RECT 35.790 74.300 35.960 74.740 ;
        RECT 33.180 72.700 34.020 72.870 ;
        RECT 34.470 72.700 35.310 72.870 ;
        RECT 32.870 71.570 33.040 72.450 ;
        RECT 34.160 71.570 34.330 72.450 ;
        RECT 35.450 71.570 35.620 72.450 ;
        RECT 33.180 71.150 34.020 71.320 ;
        RECT 34.470 71.150 35.310 71.320 ;
        RECT 35.790 70.240 35.960 70.680 ;
        RECT 33.180 68.640 34.020 68.810 ;
        RECT 34.470 68.640 35.310 68.810 ;
        RECT 32.870 67.510 33.040 68.390 ;
        RECT 34.160 67.510 34.330 68.390 ;
        RECT 35.450 67.510 35.620 68.390 ;
        RECT 33.180 67.090 34.020 67.260 ;
        RECT 34.470 67.090 35.310 67.260 ;
        RECT 35.790 66.180 35.960 66.620 ;
        RECT 33.180 64.580 34.020 64.750 ;
        RECT 34.470 64.580 35.310 64.750 ;
        RECT 32.870 63.450 33.040 64.330 ;
        RECT 34.160 63.450 34.330 64.330 ;
        RECT 35.450 63.450 35.620 64.330 ;
        RECT 33.180 63.030 34.020 63.200 ;
        RECT 34.470 63.030 35.310 63.200 ;
        RECT 35.790 62.120 35.960 62.560 ;
        RECT 33.180 60.520 34.020 60.690 ;
        RECT 34.470 60.520 35.310 60.690 ;
        RECT 32.870 59.390 33.040 60.270 ;
        RECT 34.160 59.390 34.330 60.270 ;
        RECT 35.450 59.390 35.620 60.270 ;
        RECT 33.180 58.970 34.020 59.140 ;
        RECT 34.470 58.970 35.310 59.140 ;
        RECT 35.790 58.060 35.960 58.500 ;
        RECT 24.560 53.095 25.400 53.265 ;
        RECT 25.850 53.095 26.690 53.265 ;
        RECT 24.250 50.920 24.420 52.800 ;
        RECT 25.540 50.920 25.710 52.800 ;
        RECT 26.830 50.920 27.000 52.800 ;
        RECT 24.560 50.455 25.400 50.625 ;
        RECT 25.850 50.455 26.690 50.625 ;
        RECT 27.490 50.120 27.670 53.790 ;
        RECT 28.010 53.480 28.190 57.150 ;
        RECT 28.990 56.455 29.830 56.625 ;
        RECT 30.280 56.455 31.120 56.625 ;
        RECT 28.680 54.280 28.850 56.160 ;
        RECT 29.970 54.280 30.140 56.160 ;
        RECT 31.260 54.280 31.430 56.160 ;
        RECT 28.990 53.815 29.830 53.985 ;
        RECT 30.280 53.815 31.120 53.985 ;
        RECT 33.180 55.980 34.020 56.150 ;
        RECT 34.470 55.980 35.310 56.150 ;
        RECT 32.870 54.850 33.040 55.730 ;
        RECT 34.160 54.850 34.330 55.730 ;
        RECT 35.450 54.850 35.620 55.730 ;
        RECT 33.180 54.430 34.020 54.600 ;
        RECT 34.470 54.430 35.310 54.600 ;
        RECT 35.790 53.520 35.960 53.960 ;
        RECT 24.560 49.045 25.400 49.215 ;
        RECT 25.850 49.045 26.690 49.215 ;
        RECT 24.250 46.870 24.420 48.750 ;
        RECT 25.540 46.870 25.710 48.750 ;
        RECT 26.830 46.870 27.000 48.750 ;
        RECT 24.560 46.405 25.400 46.575 ;
        RECT 25.850 46.405 26.690 46.575 ;
        RECT 27.490 46.070 27.670 49.740 ;
        RECT 24.560 44.995 25.400 45.165 ;
        RECT 25.850 44.995 26.690 45.165 ;
        RECT 24.250 42.820 24.420 44.700 ;
        RECT 25.540 42.820 25.710 44.700 ;
        RECT 26.830 42.820 27.000 44.700 ;
        RECT 24.560 42.355 25.400 42.525 ;
        RECT 25.850 42.355 26.690 42.525 ;
        RECT 27.490 42.020 27.670 45.690 ;
        RECT 24.560 40.945 25.400 41.115 ;
        RECT 25.850 40.945 26.690 41.115 ;
        RECT 24.250 38.770 24.420 40.650 ;
        RECT 25.540 38.770 25.710 40.650 ;
        RECT 26.830 38.770 27.000 40.650 ;
        RECT 24.560 38.305 25.400 38.475 ;
        RECT 25.850 38.305 26.690 38.475 ;
        RECT 27.490 37.970 27.670 41.640 ;
        RECT 24.560 36.895 25.400 37.065 ;
        RECT 25.850 36.895 26.690 37.065 ;
        RECT 24.250 34.720 24.420 36.600 ;
        RECT 25.540 34.720 25.710 36.600 ;
        RECT 26.830 34.720 27.000 36.600 ;
        RECT 24.560 34.255 25.400 34.425 ;
        RECT 25.850 34.255 26.690 34.425 ;
        RECT 27.490 33.920 27.670 37.590 ;
        RECT 24.560 32.845 25.400 33.015 ;
        RECT 25.850 32.845 26.690 33.015 ;
        RECT 24.250 30.670 24.420 32.550 ;
        RECT 25.540 30.670 25.710 32.550 ;
        RECT 26.830 30.670 27.000 32.550 ;
        RECT 24.560 30.205 25.400 30.375 ;
        RECT 25.850 30.205 26.690 30.375 ;
        RECT 27.490 29.870 27.670 33.540 ;
        RECT 24.560 28.795 25.400 28.965 ;
        RECT 25.850 28.795 26.690 28.965 ;
        RECT 24.250 26.620 24.420 28.500 ;
        RECT 25.540 26.620 25.710 28.500 ;
        RECT 26.830 26.620 27.000 28.500 ;
        RECT 24.560 26.155 25.400 26.325 ;
        RECT 25.850 26.155 26.690 26.325 ;
        RECT 27.490 25.820 27.670 29.490 ;
        RECT 24.560 24.710 25.400 24.880 ;
        RECT 25.850 24.710 26.690 24.880 ;
        RECT 24.250 22.535 24.420 24.415 ;
        RECT 25.540 22.535 25.710 24.415 ;
        RECT 26.830 22.535 27.000 24.415 ;
        RECT 24.560 22.070 25.400 22.240 ;
        RECT 25.850 22.070 26.690 22.240 ;
        RECT 27.490 21.735 27.670 25.405 ;
        RECT 24.560 20.585 25.400 20.755 ;
        RECT 25.850 20.585 26.690 20.755 ;
        RECT 24.250 18.410 24.420 20.290 ;
        RECT 25.540 18.410 25.710 20.290 ;
        RECT 26.830 18.410 27.000 20.290 ;
        RECT 24.560 17.945 25.400 18.115 ;
        RECT 25.850 17.945 26.690 18.115 ;
        RECT 27.490 17.610 27.670 21.280 ;
        RECT 20.370 15.555 21.210 15.725 ;
        RECT 21.660 15.555 22.500 15.725 ;
        RECT 20.060 14.425 20.230 15.305 ;
        RECT 21.350 14.425 21.520 15.305 ;
        RECT 22.640 14.425 22.810 15.305 ;
        RECT 20.370 14.005 21.210 14.175 ;
        RECT 21.660 14.005 22.500 14.175 ;
        RECT 19.720 13.095 19.890 13.535 ;
        RECT 24.560 16.030 25.400 16.200 ;
        RECT 25.850 16.030 26.690 16.200 ;
        RECT 24.250 13.855 24.420 15.735 ;
        RECT 25.540 13.855 25.710 15.735 ;
        RECT 26.830 13.855 27.000 15.735 ;
        RECT 24.560 13.390 25.400 13.560 ;
        RECT 25.850 13.390 26.690 13.560 ;
        RECT 27.490 13.055 27.670 16.725 ;
      LAYER met1 ;
        RECT 19.610 141.530 20.150 143.370 ;
        RECT 23.050 142.370 23.740 143.150 ;
        RECT 24.500 142.370 25.460 142.395 ;
        RECT 21.660 142.200 25.460 142.370 ;
        RECT 21.660 141.920 22.500 142.200 ;
        RECT 24.500 142.165 25.460 142.200 ;
        RECT 25.790 142.165 26.750 142.395 ;
        RECT 22.710 141.960 24.430 141.980 ;
        RECT 20.310 141.690 21.270 141.920 ;
        RECT 21.600 141.690 22.560 141.920 ;
        RECT 19.610 140.530 20.260 141.530 ;
        RECT 19.610 140.000 20.150 140.530 ;
        RECT 20.530 140.370 21.050 141.690 ;
        RECT 21.320 140.530 21.550 141.530 ;
        RECT 21.800 140.370 22.320 141.690 ;
        RECT 22.710 141.530 24.450 141.960 ;
        RECT 22.610 140.530 24.450 141.530 ;
        RECT 20.310 140.140 21.270 140.370 ;
        RECT 21.600 140.140 22.560 140.370 ;
        RECT 19.610 139.880 20.160 140.000 ;
        RECT 22.710 139.960 24.450 140.530 ;
        RECT 22.710 139.940 24.430 139.960 ;
        RECT 19.610 138.740 20.170 139.880 ;
        RECT 23.050 139.530 23.740 139.940 ;
        RECT 24.730 139.755 25.250 142.165 ;
        RECT 25.510 139.960 25.740 141.960 ;
        RECT 26.060 139.755 26.580 142.165 ;
        RECT 26.940 141.960 28.740 143.370 ;
        RECT 35.530 143.365 36.070 143.370 ;
        RECT 28.930 142.165 29.890 142.395 ;
        RECT 30.220 142.370 31.180 142.395 ;
        RECT 31.940 142.370 32.630 143.150 ;
        RECT 30.220 142.200 34.020 142.370 ;
        RECT 30.220 142.165 31.180 142.200 ;
        RECT 26.800 139.960 28.880 141.960 ;
        RECT 23.050 138.910 23.750 139.530 ;
        RECT 24.500 139.525 25.460 139.755 ;
        RECT 25.790 139.525 26.750 139.755 ;
        RECT 19.610 137.530 20.150 138.740 ;
        RECT 23.050 138.370 23.740 138.910 ;
        RECT 24.500 138.370 25.460 138.395 ;
        RECT 21.660 138.200 25.460 138.370 ;
        RECT 21.660 137.920 22.500 138.200 ;
        RECT 24.500 138.165 25.460 138.200 ;
        RECT 25.790 138.165 26.750 138.395 ;
        RECT 22.710 137.960 24.430 137.980 ;
        RECT 20.310 137.690 21.270 137.920 ;
        RECT 21.600 137.690 22.560 137.920 ;
        RECT 19.610 136.530 20.260 137.530 ;
        RECT 19.610 136.000 20.150 136.530 ;
        RECT 20.530 136.370 21.050 137.690 ;
        RECT 21.320 136.530 21.550 137.530 ;
        RECT 21.800 136.370 22.320 137.690 ;
        RECT 22.710 137.530 24.450 137.960 ;
        RECT 22.610 136.530 24.450 137.530 ;
        RECT 20.310 136.140 21.270 136.370 ;
        RECT 21.600 136.140 22.560 136.370 ;
        RECT 19.610 135.880 20.160 136.000 ;
        RECT 22.710 135.960 24.450 136.530 ;
        RECT 22.710 135.940 24.430 135.960 ;
        RECT 19.610 134.740 20.170 135.880 ;
        RECT 23.050 135.530 23.740 135.940 ;
        RECT 24.730 135.755 25.250 138.165 ;
        RECT 25.510 135.960 25.740 137.960 ;
        RECT 26.060 135.755 26.580 138.165 ;
        RECT 26.940 137.960 28.740 139.960 ;
        RECT 29.100 139.755 29.620 142.165 ;
        RECT 29.940 139.960 30.170 141.960 ;
        RECT 30.430 139.755 30.950 142.165 ;
        RECT 31.250 141.960 32.970 141.980 ;
        RECT 31.230 141.530 32.970 141.960 ;
        RECT 33.180 141.920 34.020 142.200 ;
        RECT 33.120 141.690 34.080 141.920 ;
        RECT 34.410 141.690 35.370 141.920 ;
        RECT 35.530 141.695 38.100 143.365 ;
        RECT 31.230 140.530 33.070 141.530 ;
        RECT 31.230 139.960 32.970 140.530 ;
        RECT 33.360 140.370 33.880 141.690 ;
        RECT 34.130 140.530 34.360 141.530 ;
        RECT 34.630 140.370 35.150 141.690 ;
        RECT 35.530 141.530 36.070 141.695 ;
        RECT 35.420 140.530 36.070 141.530 ;
        RECT 33.120 140.140 34.080 140.370 ;
        RECT 34.410 140.140 35.370 140.370 ;
        RECT 35.530 140.000 36.070 140.530 ;
        RECT 31.250 139.940 32.970 139.960 ;
        RECT 28.930 139.525 29.890 139.755 ;
        RECT 30.220 139.525 31.180 139.755 ;
        RECT 31.940 139.530 32.630 139.940 ;
        RECT 35.520 139.880 36.070 140.000 ;
        RECT 31.930 138.910 32.630 139.530 ;
        RECT 28.930 138.105 29.890 138.335 ;
        RECT 30.220 138.310 31.180 138.335 ;
        RECT 31.940 138.310 32.630 138.910 ;
        RECT 35.510 138.740 36.070 139.880 ;
        RECT 35.520 138.310 36.070 138.740 ;
        RECT 30.220 138.140 34.020 138.310 ;
        RECT 30.220 138.105 31.180 138.140 ;
        RECT 26.800 137.900 28.740 137.960 ;
        RECT 26.800 135.960 28.880 137.900 ;
        RECT 26.940 135.900 28.880 135.960 ;
        RECT 23.050 134.910 23.750 135.530 ;
        RECT 24.500 135.525 25.460 135.755 ;
        RECT 25.790 135.525 26.750 135.755 ;
        RECT 19.610 133.430 20.150 134.740 ;
        RECT 23.050 134.270 23.740 134.910 ;
        RECT 24.500 134.270 25.460 134.295 ;
        RECT 21.660 134.100 25.460 134.270 ;
        RECT 21.660 133.820 22.500 134.100 ;
        RECT 24.500 134.065 25.460 134.100 ;
        RECT 25.790 134.065 26.750 134.295 ;
        RECT 22.710 133.860 24.430 133.880 ;
        RECT 20.310 133.590 21.270 133.820 ;
        RECT 21.600 133.590 22.560 133.820 ;
        RECT 19.610 132.430 20.260 133.430 ;
        RECT 19.610 131.900 20.150 132.430 ;
        RECT 20.530 132.270 21.050 133.590 ;
        RECT 21.320 132.430 21.550 133.430 ;
        RECT 21.800 132.270 22.320 133.590 ;
        RECT 22.710 133.430 24.450 133.860 ;
        RECT 22.610 132.430 24.450 133.430 ;
        RECT 20.310 132.040 21.270 132.270 ;
        RECT 21.600 132.040 22.560 132.270 ;
        RECT 19.610 131.780 20.160 131.900 ;
        RECT 22.710 131.860 24.450 132.430 ;
        RECT 22.710 131.840 24.430 131.860 ;
        RECT 19.610 130.640 20.170 131.780 ;
        RECT 23.050 131.430 23.740 131.840 ;
        RECT 24.730 131.655 25.250 134.065 ;
        RECT 25.510 131.860 25.740 133.860 ;
        RECT 26.060 131.655 26.580 134.065 ;
        RECT 26.940 133.860 28.740 135.900 ;
        RECT 29.100 135.695 29.620 138.105 ;
        RECT 29.940 135.900 30.170 137.900 ;
        RECT 30.430 135.695 30.950 138.105 ;
        RECT 31.250 137.900 32.970 137.920 ;
        RECT 31.230 137.470 32.970 137.900 ;
        RECT 33.180 137.860 34.020 138.140 ;
        RECT 33.120 137.630 34.080 137.860 ;
        RECT 34.410 137.630 35.370 137.860 ;
        RECT 31.230 136.470 33.070 137.470 ;
        RECT 31.230 135.900 32.970 136.470 ;
        RECT 33.360 136.310 33.880 137.630 ;
        RECT 34.130 136.470 34.360 137.470 ;
        RECT 34.630 136.310 35.150 137.630 ;
        RECT 35.530 137.470 36.070 138.310 ;
        RECT 35.420 136.470 36.070 137.470 ;
        RECT 33.120 136.080 34.080 136.310 ;
        RECT 34.410 136.080 35.370 136.310 ;
        RECT 35.530 135.940 36.070 136.470 ;
        RECT 31.250 135.880 32.970 135.900 ;
        RECT 28.930 135.465 29.890 135.695 ;
        RECT 30.220 135.465 31.180 135.695 ;
        RECT 31.940 135.470 32.630 135.880 ;
        RECT 35.520 135.820 36.070 135.940 ;
        RECT 31.930 134.850 32.630 135.470 ;
        RECT 28.930 134.045 29.890 134.275 ;
        RECT 30.220 134.250 31.180 134.275 ;
        RECT 31.940 134.250 32.630 134.850 ;
        RECT 35.510 134.680 36.070 135.820 ;
        RECT 30.220 134.080 34.020 134.250 ;
        RECT 30.220 134.045 31.180 134.080 ;
        RECT 26.800 133.840 28.740 133.860 ;
        RECT 26.800 131.860 28.880 133.840 ;
        RECT 26.940 131.840 28.880 131.860 ;
        RECT 23.050 130.810 23.750 131.430 ;
        RECT 24.500 131.425 25.460 131.655 ;
        RECT 25.790 131.425 26.750 131.655 ;
        RECT 19.610 129.380 20.150 130.640 ;
        RECT 23.050 130.220 23.740 130.810 ;
        RECT 24.500 130.220 25.460 130.245 ;
        RECT 21.660 130.050 25.460 130.220 ;
        RECT 21.660 129.770 22.500 130.050 ;
        RECT 24.500 130.015 25.460 130.050 ;
        RECT 25.790 130.015 26.750 130.245 ;
        RECT 22.710 129.810 24.430 129.830 ;
        RECT 20.310 129.540 21.270 129.770 ;
        RECT 21.600 129.540 22.560 129.770 ;
        RECT 19.610 128.380 20.260 129.380 ;
        RECT 19.610 127.850 20.150 128.380 ;
        RECT 20.530 128.220 21.050 129.540 ;
        RECT 21.320 128.380 21.550 129.380 ;
        RECT 21.800 128.220 22.320 129.540 ;
        RECT 22.710 129.380 24.450 129.810 ;
        RECT 22.610 128.380 24.450 129.380 ;
        RECT 20.310 127.990 21.270 128.220 ;
        RECT 21.600 127.990 22.560 128.220 ;
        RECT 19.610 127.730 20.160 127.850 ;
        RECT 22.710 127.810 24.450 128.380 ;
        RECT 22.710 127.790 24.430 127.810 ;
        RECT 19.610 126.590 20.170 127.730 ;
        RECT 23.050 127.380 23.740 127.790 ;
        RECT 24.730 127.605 25.250 130.015 ;
        RECT 25.510 127.810 25.740 129.810 ;
        RECT 26.060 127.605 26.580 130.015 ;
        RECT 26.940 129.810 28.740 131.840 ;
        RECT 29.100 131.635 29.620 134.045 ;
        RECT 29.940 131.840 30.170 133.840 ;
        RECT 30.430 131.635 30.950 134.045 ;
        RECT 31.250 133.840 32.970 133.860 ;
        RECT 31.230 133.410 32.970 133.840 ;
        RECT 33.180 133.800 34.020 134.080 ;
        RECT 33.120 133.570 34.080 133.800 ;
        RECT 34.410 133.570 35.370 133.800 ;
        RECT 31.230 132.410 33.070 133.410 ;
        RECT 31.230 131.840 32.970 132.410 ;
        RECT 33.360 132.250 33.880 133.570 ;
        RECT 34.130 132.410 34.360 133.410 ;
        RECT 34.630 132.250 35.150 133.570 ;
        RECT 35.530 133.410 36.070 134.680 ;
        RECT 35.420 132.410 36.070 133.410 ;
        RECT 33.120 132.020 34.080 132.250 ;
        RECT 34.410 132.020 35.370 132.250 ;
        RECT 35.530 131.880 36.070 132.410 ;
        RECT 31.250 131.820 32.970 131.840 ;
        RECT 28.930 131.405 29.890 131.635 ;
        RECT 30.220 131.405 31.180 131.635 ;
        RECT 31.940 131.410 32.630 131.820 ;
        RECT 35.520 131.760 36.070 131.880 ;
        RECT 31.930 130.790 32.630 131.410 ;
        RECT 28.930 129.985 29.890 130.215 ;
        RECT 30.220 130.190 31.180 130.215 ;
        RECT 31.940 130.190 32.630 130.790 ;
        RECT 35.510 130.620 36.070 131.760 ;
        RECT 30.220 130.020 34.020 130.190 ;
        RECT 30.220 129.985 31.180 130.020 ;
        RECT 26.800 129.780 28.740 129.810 ;
        RECT 26.800 127.810 28.880 129.780 ;
        RECT 26.940 127.780 28.880 127.810 ;
        RECT 23.050 126.760 23.750 127.380 ;
        RECT 24.500 127.375 25.460 127.605 ;
        RECT 25.790 127.375 26.750 127.605 ;
        RECT 19.610 125.330 20.150 126.590 ;
        RECT 23.050 126.170 23.740 126.760 ;
        RECT 24.500 126.170 25.460 126.195 ;
        RECT 21.660 126.000 25.460 126.170 ;
        RECT 21.660 125.720 22.500 126.000 ;
        RECT 24.500 125.965 25.460 126.000 ;
        RECT 25.790 125.965 26.750 126.195 ;
        RECT 22.710 125.760 24.430 125.780 ;
        RECT 20.310 125.490 21.270 125.720 ;
        RECT 21.600 125.490 22.560 125.720 ;
        RECT 19.610 124.330 20.260 125.330 ;
        RECT 19.610 123.800 20.150 124.330 ;
        RECT 20.530 124.170 21.050 125.490 ;
        RECT 21.320 124.330 21.550 125.330 ;
        RECT 21.800 124.170 22.320 125.490 ;
        RECT 22.710 125.330 24.450 125.760 ;
        RECT 22.610 124.330 24.450 125.330 ;
        RECT 20.310 123.940 21.270 124.170 ;
        RECT 21.600 123.940 22.560 124.170 ;
        RECT 19.610 123.680 20.160 123.800 ;
        RECT 22.710 123.760 24.450 124.330 ;
        RECT 22.710 123.740 24.430 123.760 ;
        RECT 19.610 122.540 20.170 123.680 ;
        RECT 23.050 123.330 23.740 123.740 ;
        RECT 24.730 123.555 25.250 125.965 ;
        RECT 25.510 123.760 25.740 125.760 ;
        RECT 26.060 123.555 26.580 125.965 ;
        RECT 26.940 125.760 28.740 127.780 ;
        RECT 29.100 127.575 29.620 129.985 ;
        RECT 29.940 127.780 30.170 129.780 ;
        RECT 30.430 127.575 30.950 129.985 ;
        RECT 31.250 129.780 32.970 129.800 ;
        RECT 31.230 129.350 32.970 129.780 ;
        RECT 33.180 129.740 34.020 130.020 ;
        RECT 33.120 129.510 34.080 129.740 ;
        RECT 34.410 129.510 35.370 129.740 ;
        RECT 31.230 128.350 33.070 129.350 ;
        RECT 31.230 127.780 32.970 128.350 ;
        RECT 33.360 128.190 33.880 129.510 ;
        RECT 34.130 128.350 34.360 129.350 ;
        RECT 34.630 128.190 35.150 129.510 ;
        RECT 35.530 129.350 36.070 130.620 ;
        RECT 35.420 128.350 36.070 129.350 ;
        RECT 33.120 127.960 34.080 128.190 ;
        RECT 34.410 127.960 35.370 128.190 ;
        RECT 35.530 127.820 36.070 128.350 ;
        RECT 31.250 127.760 32.970 127.780 ;
        RECT 28.930 127.345 29.890 127.575 ;
        RECT 30.220 127.345 31.180 127.575 ;
        RECT 31.940 127.350 32.630 127.760 ;
        RECT 35.520 127.700 36.070 127.820 ;
        RECT 31.930 126.730 32.630 127.350 ;
        RECT 28.930 125.925 29.890 126.155 ;
        RECT 30.220 126.130 31.180 126.155 ;
        RECT 31.940 126.130 32.630 126.730 ;
        RECT 35.510 126.560 36.070 127.700 ;
        RECT 30.220 125.960 34.020 126.130 ;
        RECT 30.220 125.925 31.180 125.960 ;
        RECT 26.800 125.720 28.740 125.760 ;
        RECT 26.800 123.760 28.880 125.720 ;
        RECT 26.940 123.720 28.880 123.760 ;
        RECT 23.050 122.710 23.750 123.330 ;
        RECT 24.500 123.325 25.460 123.555 ;
        RECT 25.790 123.325 26.750 123.555 ;
        RECT 19.610 121.280 20.150 122.540 ;
        RECT 23.050 122.120 23.740 122.710 ;
        RECT 24.500 122.120 25.460 122.145 ;
        RECT 21.660 121.950 25.460 122.120 ;
        RECT 21.660 121.670 22.500 121.950 ;
        RECT 24.500 121.915 25.460 121.950 ;
        RECT 25.790 121.915 26.750 122.145 ;
        RECT 22.710 121.710 24.430 121.730 ;
        RECT 20.310 121.440 21.270 121.670 ;
        RECT 21.600 121.440 22.560 121.670 ;
        RECT 19.610 120.280 20.260 121.280 ;
        RECT 19.610 119.750 20.150 120.280 ;
        RECT 20.530 120.120 21.050 121.440 ;
        RECT 21.320 120.280 21.550 121.280 ;
        RECT 21.800 120.120 22.320 121.440 ;
        RECT 22.710 121.280 24.450 121.710 ;
        RECT 22.610 120.280 24.450 121.280 ;
        RECT 20.310 119.890 21.270 120.120 ;
        RECT 21.600 119.890 22.560 120.120 ;
        RECT 19.610 119.630 20.160 119.750 ;
        RECT 22.710 119.710 24.450 120.280 ;
        RECT 22.710 119.690 24.430 119.710 ;
        RECT 19.610 118.490 20.170 119.630 ;
        RECT 23.050 119.280 23.740 119.690 ;
        RECT 24.730 119.505 25.250 121.915 ;
        RECT 25.510 119.710 25.740 121.710 ;
        RECT 26.060 119.505 26.580 121.915 ;
        RECT 26.940 121.710 28.740 123.720 ;
        RECT 29.100 123.515 29.620 125.925 ;
        RECT 29.940 123.720 30.170 125.720 ;
        RECT 30.430 123.515 30.950 125.925 ;
        RECT 31.250 125.720 32.970 125.740 ;
        RECT 31.230 125.290 32.970 125.720 ;
        RECT 33.180 125.680 34.020 125.960 ;
        RECT 33.120 125.450 34.080 125.680 ;
        RECT 34.410 125.450 35.370 125.680 ;
        RECT 31.230 124.290 33.070 125.290 ;
        RECT 31.230 123.720 32.970 124.290 ;
        RECT 33.360 124.130 33.880 125.450 ;
        RECT 34.130 124.290 34.360 125.290 ;
        RECT 34.630 124.130 35.150 125.450 ;
        RECT 35.530 125.290 36.070 126.560 ;
        RECT 35.420 124.290 36.070 125.290 ;
        RECT 33.120 123.900 34.080 124.130 ;
        RECT 34.410 123.900 35.370 124.130 ;
        RECT 35.530 123.760 36.070 124.290 ;
        RECT 31.250 123.700 32.970 123.720 ;
        RECT 28.930 123.285 29.890 123.515 ;
        RECT 30.220 123.285 31.180 123.515 ;
        RECT 31.940 123.290 32.630 123.700 ;
        RECT 35.520 123.640 36.070 123.760 ;
        RECT 31.930 122.670 32.630 123.290 ;
        RECT 28.930 121.865 29.890 122.095 ;
        RECT 30.220 122.070 31.180 122.095 ;
        RECT 31.940 122.070 32.630 122.670 ;
        RECT 35.510 122.500 36.070 123.640 ;
        RECT 30.220 121.900 34.020 122.070 ;
        RECT 30.220 121.865 31.180 121.900 ;
        RECT 26.800 121.660 28.740 121.710 ;
        RECT 26.800 119.710 28.880 121.660 ;
        RECT 26.940 119.660 28.880 119.710 ;
        RECT 23.050 118.660 23.750 119.280 ;
        RECT 24.500 119.275 25.460 119.505 ;
        RECT 25.790 119.275 26.750 119.505 ;
        RECT 19.610 117.230 20.150 118.490 ;
        RECT 23.050 118.070 23.740 118.660 ;
        RECT 24.500 118.070 25.460 118.095 ;
        RECT 21.660 117.900 25.460 118.070 ;
        RECT 21.660 117.620 22.500 117.900 ;
        RECT 24.500 117.865 25.460 117.900 ;
        RECT 25.790 117.865 26.750 118.095 ;
        RECT 22.710 117.660 24.430 117.680 ;
        RECT 20.310 117.390 21.270 117.620 ;
        RECT 21.600 117.390 22.560 117.620 ;
        RECT 19.610 116.230 20.260 117.230 ;
        RECT 19.610 115.700 20.150 116.230 ;
        RECT 20.530 116.070 21.050 117.390 ;
        RECT 21.320 116.230 21.550 117.230 ;
        RECT 21.800 116.070 22.320 117.390 ;
        RECT 22.710 117.230 24.450 117.660 ;
        RECT 22.610 116.230 24.450 117.230 ;
        RECT 20.310 115.840 21.270 116.070 ;
        RECT 21.600 115.840 22.560 116.070 ;
        RECT 19.610 115.580 20.160 115.700 ;
        RECT 22.710 115.660 24.450 116.230 ;
        RECT 22.710 115.640 24.430 115.660 ;
        RECT 19.610 114.440 20.170 115.580 ;
        RECT 23.050 115.230 23.740 115.640 ;
        RECT 24.730 115.455 25.250 117.865 ;
        RECT 25.510 115.660 25.740 117.660 ;
        RECT 26.060 115.455 26.580 117.865 ;
        RECT 26.940 117.660 28.740 119.660 ;
        RECT 29.100 119.455 29.620 121.865 ;
        RECT 29.940 119.660 30.170 121.660 ;
        RECT 30.430 119.455 30.950 121.865 ;
        RECT 31.250 121.660 32.970 121.680 ;
        RECT 31.230 121.230 32.970 121.660 ;
        RECT 33.180 121.620 34.020 121.900 ;
        RECT 33.120 121.390 34.080 121.620 ;
        RECT 34.410 121.390 35.370 121.620 ;
        RECT 31.230 120.230 33.070 121.230 ;
        RECT 31.230 119.660 32.970 120.230 ;
        RECT 33.360 120.070 33.880 121.390 ;
        RECT 34.130 120.230 34.360 121.230 ;
        RECT 34.630 120.070 35.150 121.390 ;
        RECT 35.530 121.230 36.070 122.500 ;
        RECT 35.420 120.230 36.070 121.230 ;
        RECT 33.120 119.840 34.080 120.070 ;
        RECT 34.410 119.840 35.370 120.070 ;
        RECT 35.530 119.700 36.070 120.230 ;
        RECT 31.250 119.640 32.970 119.660 ;
        RECT 28.930 119.225 29.890 119.455 ;
        RECT 30.220 119.225 31.180 119.455 ;
        RECT 31.940 119.230 32.630 119.640 ;
        RECT 35.520 119.580 36.070 119.700 ;
        RECT 31.930 118.610 32.630 119.230 ;
        RECT 28.930 117.805 29.890 118.035 ;
        RECT 30.220 118.010 31.180 118.035 ;
        RECT 31.940 118.010 32.630 118.610 ;
        RECT 35.510 118.440 36.070 119.580 ;
        RECT 30.220 117.840 34.020 118.010 ;
        RECT 30.220 117.805 31.180 117.840 ;
        RECT 26.800 117.600 28.740 117.660 ;
        RECT 26.800 115.660 28.880 117.600 ;
        RECT 26.940 115.600 28.880 115.660 ;
        RECT 23.050 114.610 23.750 115.230 ;
        RECT 24.500 115.225 25.460 115.455 ;
        RECT 25.790 115.225 26.750 115.455 ;
        RECT 19.610 113.180 20.150 114.440 ;
        RECT 23.050 114.020 23.740 114.610 ;
        RECT 24.500 114.020 25.460 114.045 ;
        RECT 21.660 113.850 25.460 114.020 ;
        RECT 21.660 113.570 22.500 113.850 ;
        RECT 24.500 113.815 25.460 113.850 ;
        RECT 25.790 113.815 26.750 114.045 ;
        RECT 22.710 113.610 24.430 113.630 ;
        RECT 20.310 113.340 21.270 113.570 ;
        RECT 21.600 113.340 22.560 113.570 ;
        RECT 19.610 112.180 20.260 113.180 ;
        RECT 19.610 111.650 20.150 112.180 ;
        RECT 20.530 112.020 21.050 113.340 ;
        RECT 21.320 112.180 21.550 113.180 ;
        RECT 21.800 112.020 22.320 113.340 ;
        RECT 22.710 113.180 24.450 113.610 ;
        RECT 22.610 112.180 24.450 113.180 ;
        RECT 20.310 111.790 21.270 112.020 ;
        RECT 21.600 111.790 22.560 112.020 ;
        RECT 19.610 111.530 20.160 111.650 ;
        RECT 22.710 111.610 24.450 112.180 ;
        RECT 22.710 111.590 24.430 111.610 ;
        RECT 19.610 110.390 20.170 111.530 ;
        RECT 23.050 111.180 23.740 111.590 ;
        RECT 24.730 111.405 25.250 113.815 ;
        RECT 25.510 111.610 25.740 113.610 ;
        RECT 26.060 111.405 26.580 113.815 ;
        RECT 26.940 113.610 28.740 115.600 ;
        RECT 29.100 115.395 29.620 117.805 ;
        RECT 29.940 115.600 30.170 117.600 ;
        RECT 30.430 115.395 30.950 117.805 ;
        RECT 31.250 117.600 32.970 117.620 ;
        RECT 31.230 117.170 32.970 117.600 ;
        RECT 33.180 117.560 34.020 117.840 ;
        RECT 33.120 117.330 34.080 117.560 ;
        RECT 34.410 117.330 35.370 117.560 ;
        RECT 31.230 116.170 33.070 117.170 ;
        RECT 31.230 115.600 32.970 116.170 ;
        RECT 33.360 116.010 33.880 117.330 ;
        RECT 34.130 116.170 34.360 117.170 ;
        RECT 34.630 116.010 35.150 117.330 ;
        RECT 35.530 117.170 36.070 118.440 ;
        RECT 35.420 116.170 36.070 117.170 ;
        RECT 33.120 115.780 34.080 116.010 ;
        RECT 34.410 115.780 35.370 116.010 ;
        RECT 35.530 115.640 36.070 116.170 ;
        RECT 31.250 115.580 32.970 115.600 ;
        RECT 28.930 115.165 29.890 115.395 ;
        RECT 30.220 115.165 31.180 115.395 ;
        RECT 31.940 115.170 32.630 115.580 ;
        RECT 35.520 115.520 36.070 115.640 ;
        RECT 31.930 114.550 32.630 115.170 ;
        RECT 28.930 113.745 29.890 113.975 ;
        RECT 30.220 113.950 31.180 113.975 ;
        RECT 31.940 113.950 32.630 114.550 ;
        RECT 35.510 114.380 36.070 115.520 ;
        RECT 30.220 113.780 34.020 113.950 ;
        RECT 30.220 113.745 31.180 113.780 ;
        RECT 26.800 113.540 28.740 113.610 ;
        RECT 26.800 111.610 28.880 113.540 ;
        RECT 26.940 111.540 28.880 111.610 ;
        RECT 23.050 110.560 23.750 111.180 ;
        RECT 24.500 111.175 25.460 111.405 ;
        RECT 25.790 111.175 26.750 111.405 ;
        RECT 19.610 109.130 20.150 110.390 ;
        RECT 23.050 109.970 23.740 110.560 ;
        RECT 24.500 109.970 25.460 109.995 ;
        RECT 21.660 109.800 25.460 109.970 ;
        RECT 21.660 109.520 22.500 109.800 ;
        RECT 24.500 109.765 25.460 109.800 ;
        RECT 25.790 109.765 26.750 109.995 ;
        RECT 22.710 109.560 24.430 109.580 ;
        RECT 20.310 109.290 21.270 109.520 ;
        RECT 21.600 109.290 22.560 109.520 ;
        RECT 19.610 108.130 20.260 109.130 ;
        RECT 19.610 107.600 20.150 108.130 ;
        RECT 20.530 107.970 21.050 109.290 ;
        RECT 21.320 108.130 21.550 109.130 ;
        RECT 21.800 107.970 22.320 109.290 ;
        RECT 22.710 109.130 24.450 109.560 ;
        RECT 22.610 108.130 24.450 109.130 ;
        RECT 20.310 107.740 21.270 107.970 ;
        RECT 21.600 107.740 22.560 107.970 ;
        RECT 19.610 107.480 20.160 107.600 ;
        RECT 22.710 107.560 24.450 108.130 ;
        RECT 22.710 107.540 24.430 107.560 ;
        RECT 19.610 106.340 20.170 107.480 ;
        RECT 23.050 107.130 23.740 107.540 ;
        RECT 24.730 107.355 25.250 109.765 ;
        RECT 25.510 107.560 25.740 109.560 ;
        RECT 26.060 107.355 26.580 109.765 ;
        RECT 26.940 109.560 28.740 111.540 ;
        RECT 29.100 111.335 29.620 113.745 ;
        RECT 29.940 111.540 30.170 113.540 ;
        RECT 30.430 111.335 30.950 113.745 ;
        RECT 31.250 113.540 32.970 113.560 ;
        RECT 31.230 113.110 32.970 113.540 ;
        RECT 33.180 113.500 34.020 113.780 ;
        RECT 33.120 113.270 34.080 113.500 ;
        RECT 34.410 113.270 35.370 113.500 ;
        RECT 31.230 112.110 33.070 113.110 ;
        RECT 31.230 111.540 32.970 112.110 ;
        RECT 33.360 111.950 33.880 113.270 ;
        RECT 34.130 112.110 34.360 113.110 ;
        RECT 34.630 111.950 35.150 113.270 ;
        RECT 35.530 113.110 36.070 114.380 ;
        RECT 35.420 112.110 36.070 113.110 ;
        RECT 33.120 111.720 34.080 111.950 ;
        RECT 34.410 111.720 35.370 111.950 ;
        RECT 35.530 111.580 36.070 112.110 ;
        RECT 31.250 111.520 32.970 111.540 ;
        RECT 28.930 111.105 29.890 111.335 ;
        RECT 30.220 111.105 31.180 111.335 ;
        RECT 31.940 111.110 32.630 111.520 ;
        RECT 35.520 111.460 36.070 111.580 ;
        RECT 31.930 110.490 32.630 111.110 ;
        RECT 28.930 109.685 29.890 109.915 ;
        RECT 30.220 109.890 31.180 109.915 ;
        RECT 31.940 109.890 32.630 110.490 ;
        RECT 35.510 110.320 36.070 111.460 ;
        RECT 30.220 109.720 34.020 109.890 ;
        RECT 30.220 109.685 31.180 109.720 ;
        RECT 26.800 109.480 28.740 109.560 ;
        RECT 26.800 107.560 28.880 109.480 ;
        RECT 26.940 107.480 28.880 107.560 ;
        RECT 23.050 106.510 23.750 107.130 ;
        RECT 24.500 107.125 25.460 107.355 ;
        RECT 25.790 107.125 26.750 107.355 ;
        RECT 19.610 105.080 20.150 106.340 ;
        RECT 23.050 105.920 23.740 106.510 ;
        RECT 24.500 105.920 25.460 105.945 ;
        RECT 21.660 105.750 25.460 105.920 ;
        RECT 21.660 105.470 22.500 105.750 ;
        RECT 24.500 105.715 25.460 105.750 ;
        RECT 25.790 105.715 26.750 105.945 ;
        RECT 22.710 105.510 24.430 105.530 ;
        RECT 20.310 105.240 21.270 105.470 ;
        RECT 21.600 105.240 22.560 105.470 ;
        RECT 19.610 104.080 20.260 105.080 ;
        RECT 19.610 103.550 20.150 104.080 ;
        RECT 20.530 103.920 21.050 105.240 ;
        RECT 21.320 104.080 21.550 105.080 ;
        RECT 21.800 103.920 22.320 105.240 ;
        RECT 22.710 105.080 24.450 105.510 ;
        RECT 22.610 104.080 24.450 105.080 ;
        RECT 20.310 103.690 21.270 103.920 ;
        RECT 21.600 103.690 22.560 103.920 ;
        RECT 19.610 103.430 20.160 103.550 ;
        RECT 22.710 103.510 24.450 104.080 ;
        RECT 22.710 103.490 24.430 103.510 ;
        RECT 19.610 102.290 20.170 103.430 ;
        RECT 23.050 103.080 23.740 103.490 ;
        RECT 24.730 103.305 25.250 105.715 ;
        RECT 25.510 103.510 25.740 105.510 ;
        RECT 26.060 103.305 26.580 105.715 ;
        RECT 26.940 105.510 28.740 107.480 ;
        RECT 29.100 107.275 29.620 109.685 ;
        RECT 29.940 107.480 30.170 109.480 ;
        RECT 30.430 107.275 30.950 109.685 ;
        RECT 31.250 109.480 32.970 109.500 ;
        RECT 31.230 109.050 32.970 109.480 ;
        RECT 33.180 109.440 34.020 109.720 ;
        RECT 33.120 109.210 34.080 109.440 ;
        RECT 34.410 109.210 35.370 109.440 ;
        RECT 31.230 108.050 33.070 109.050 ;
        RECT 31.230 107.480 32.970 108.050 ;
        RECT 33.360 107.890 33.880 109.210 ;
        RECT 34.130 108.050 34.360 109.050 ;
        RECT 34.630 107.890 35.150 109.210 ;
        RECT 35.530 109.050 36.070 110.320 ;
        RECT 35.420 108.050 36.070 109.050 ;
        RECT 33.120 107.660 34.080 107.890 ;
        RECT 34.410 107.660 35.370 107.890 ;
        RECT 35.530 107.520 36.070 108.050 ;
        RECT 31.250 107.460 32.970 107.480 ;
        RECT 28.930 107.045 29.890 107.275 ;
        RECT 30.220 107.045 31.180 107.275 ;
        RECT 31.940 107.050 32.630 107.460 ;
        RECT 35.520 107.400 36.070 107.520 ;
        RECT 31.930 106.430 32.630 107.050 ;
        RECT 28.930 105.625 29.890 105.855 ;
        RECT 30.220 105.830 31.180 105.855 ;
        RECT 31.940 105.830 32.630 106.430 ;
        RECT 35.510 106.260 36.070 107.400 ;
        RECT 30.220 105.660 34.020 105.830 ;
        RECT 30.220 105.625 31.180 105.660 ;
        RECT 26.800 105.420 28.740 105.510 ;
        RECT 26.800 103.510 28.880 105.420 ;
        RECT 26.940 103.420 28.880 103.510 ;
        RECT 23.050 102.460 23.750 103.080 ;
        RECT 24.500 103.075 25.460 103.305 ;
        RECT 25.790 103.075 26.750 103.305 ;
        RECT 19.610 101.030 20.150 102.290 ;
        RECT 23.050 101.870 23.740 102.460 ;
        RECT 24.500 101.870 25.460 101.895 ;
        RECT 21.660 101.700 25.460 101.870 ;
        RECT 21.660 101.420 22.500 101.700 ;
        RECT 24.500 101.665 25.460 101.700 ;
        RECT 25.790 101.665 26.750 101.895 ;
        RECT 22.710 101.460 24.430 101.480 ;
        RECT 20.310 101.190 21.270 101.420 ;
        RECT 21.600 101.190 22.560 101.420 ;
        RECT 19.610 100.030 20.260 101.030 ;
        RECT 19.610 99.500 20.150 100.030 ;
        RECT 20.530 99.870 21.050 101.190 ;
        RECT 21.320 100.030 21.550 101.030 ;
        RECT 21.800 99.870 22.320 101.190 ;
        RECT 22.710 101.030 24.450 101.460 ;
        RECT 22.610 100.030 24.450 101.030 ;
        RECT 20.310 99.640 21.270 99.870 ;
        RECT 21.600 99.640 22.560 99.870 ;
        RECT 19.610 99.380 20.160 99.500 ;
        RECT 22.710 99.460 24.450 100.030 ;
        RECT 22.710 99.440 24.430 99.460 ;
        RECT 19.610 98.240 20.170 99.380 ;
        RECT 23.050 99.030 23.740 99.440 ;
        RECT 24.730 99.255 25.250 101.665 ;
        RECT 25.510 99.460 25.740 101.460 ;
        RECT 26.060 99.255 26.580 101.665 ;
        RECT 26.940 101.460 28.740 103.420 ;
        RECT 29.100 103.215 29.620 105.625 ;
        RECT 29.940 103.420 30.170 105.420 ;
        RECT 30.430 103.215 30.950 105.625 ;
        RECT 31.250 105.420 32.970 105.440 ;
        RECT 31.230 104.990 32.970 105.420 ;
        RECT 33.180 105.380 34.020 105.660 ;
        RECT 33.120 105.150 34.080 105.380 ;
        RECT 34.410 105.150 35.370 105.380 ;
        RECT 31.230 103.990 33.070 104.990 ;
        RECT 31.230 103.420 32.970 103.990 ;
        RECT 33.360 103.830 33.880 105.150 ;
        RECT 34.130 103.990 34.360 104.990 ;
        RECT 34.630 103.830 35.150 105.150 ;
        RECT 35.530 104.990 36.070 106.260 ;
        RECT 35.420 103.990 36.070 104.990 ;
        RECT 33.120 103.600 34.080 103.830 ;
        RECT 34.410 103.600 35.370 103.830 ;
        RECT 35.530 103.460 36.070 103.990 ;
        RECT 31.250 103.400 32.970 103.420 ;
        RECT 28.930 102.985 29.890 103.215 ;
        RECT 30.220 102.985 31.180 103.215 ;
        RECT 31.940 102.990 32.630 103.400 ;
        RECT 35.520 103.340 36.070 103.460 ;
        RECT 31.930 102.370 32.630 102.990 ;
        RECT 28.930 101.565 29.890 101.795 ;
        RECT 30.220 101.770 31.180 101.795 ;
        RECT 31.940 101.770 32.630 102.370 ;
        RECT 35.510 102.200 36.070 103.340 ;
        RECT 30.220 101.600 34.020 101.770 ;
        RECT 30.220 101.565 31.180 101.600 ;
        RECT 26.800 101.360 28.740 101.460 ;
        RECT 26.800 99.460 28.880 101.360 ;
        RECT 26.940 99.360 28.880 99.460 ;
        RECT 23.050 98.410 23.750 99.030 ;
        RECT 24.500 99.025 25.460 99.255 ;
        RECT 25.790 99.025 26.750 99.255 ;
        RECT 19.610 96.980 20.150 98.240 ;
        RECT 23.050 97.820 23.740 98.410 ;
        RECT 24.500 97.820 25.460 97.845 ;
        RECT 21.660 97.650 25.460 97.820 ;
        RECT 21.660 97.370 22.500 97.650 ;
        RECT 24.500 97.615 25.460 97.650 ;
        RECT 25.790 97.615 26.750 97.845 ;
        RECT 22.710 97.410 24.430 97.430 ;
        RECT 20.310 97.140 21.270 97.370 ;
        RECT 21.600 97.140 22.560 97.370 ;
        RECT 19.610 95.980 20.260 96.980 ;
        RECT 19.610 95.450 20.150 95.980 ;
        RECT 20.530 95.820 21.050 97.140 ;
        RECT 21.320 95.980 21.550 96.980 ;
        RECT 21.800 95.820 22.320 97.140 ;
        RECT 22.710 96.980 24.450 97.410 ;
        RECT 22.610 95.980 24.450 96.980 ;
        RECT 20.310 95.590 21.270 95.820 ;
        RECT 21.600 95.590 22.560 95.820 ;
        RECT 19.610 95.330 20.160 95.450 ;
        RECT 22.710 95.410 24.450 95.980 ;
        RECT 22.710 95.390 24.430 95.410 ;
        RECT 19.610 94.190 20.170 95.330 ;
        RECT 23.050 94.980 23.740 95.390 ;
        RECT 24.730 95.205 25.250 97.615 ;
        RECT 25.510 95.410 25.740 97.410 ;
        RECT 26.060 95.205 26.580 97.615 ;
        RECT 26.940 97.410 28.740 99.360 ;
        RECT 29.100 99.155 29.620 101.565 ;
        RECT 29.940 99.360 30.170 101.360 ;
        RECT 30.430 99.155 30.950 101.565 ;
        RECT 31.250 101.360 32.970 101.380 ;
        RECT 31.230 100.930 32.970 101.360 ;
        RECT 33.180 101.320 34.020 101.600 ;
        RECT 33.120 101.090 34.080 101.320 ;
        RECT 34.410 101.090 35.370 101.320 ;
        RECT 31.230 99.930 33.070 100.930 ;
        RECT 31.230 99.360 32.970 99.930 ;
        RECT 33.360 99.770 33.880 101.090 ;
        RECT 34.130 99.930 34.360 100.930 ;
        RECT 34.630 99.770 35.150 101.090 ;
        RECT 35.530 100.930 36.070 102.200 ;
        RECT 35.420 99.930 36.070 100.930 ;
        RECT 33.120 99.540 34.080 99.770 ;
        RECT 34.410 99.540 35.370 99.770 ;
        RECT 35.530 99.400 36.070 99.930 ;
        RECT 31.250 99.340 32.970 99.360 ;
        RECT 28.930 98.925 29.890 99.155 ;
        RECT 30.220 98.925 31.180 99.155 ;
        RECT 31.940 98.930 32.630 99.340 ;
        RECT 35.520 99.280 36.070 99.400 ;
        RECT 31.930 98.310 32.630 98.930 ;
        RECT 28.930 97.505 29.890 97.735 ;
        RECT 30.220 97.710 31.180 97.735 ;
        RECT 31.940 97.710 32.630 98.310 ;
        RECT 35.510 98.140 36.070 99.280 ;
        RECT 30.220 97.540 34.020 97.710 ;
        RECT 30.220 97.505 31.180 97.540 ;
        RECT 26.800 97.300 28.740 97.410 ;
        RECT 26.800 95.410 28.880 97.300 ;
        RECT 26.940 95.300 28.880 95.410 ;
        RECT 23.050 94.360 23.750 94.980 ;
        RECT 24.500 94.975 25.460 95.205 ;
        RECT 25.790 94.975 26.750 95.205 ;
        RECT 19.610 92.930 20.150 94.190 ;
        RECT 23.050 93.770 23.740 94.360 ;
        RECT 24.500 93.770 25.460 93.795 ;
        RECT 21.660 93.600 25.460 93.770 ;
        RECT 21.660 93.320 22.500 93.600 ;
        RECT 24.500 93.565 25.460 93.600 ;
        RECT 25.790 93.565 26.750 93.795 ;
        RECT 22.710 93.360 24.430 93.380 ;
        RECT 20.310 93.090 21.270 93.320 ;
        RECT 21.600 93.090 22.560 93.320 ;
        RECT 19.610 91.930 20.260 92.930 ;
        RECT 19.610 91.400 20.150 91.930 ;
        RECT 20.530 91.770 21.050 93.090 ;
        RECT 21.320 91.930 21.550 92.930 ;
        RECT 21.800 91.770 22.320 93.090 ;
        RECT 22.710 92.930 24.450 93.360 ;
        RECT 22.610 91.930 24.450 92.930 ;
        RECT 20.310 91.540 21.270 91.770 ;
        RECT 21.600 91.540 22.560 91.770 ;
        RECT 19.610 91.280 20.160 91.400 ;
        RECT 22.710 91.360 24.450 91.930 ;
        RECT 22.710 91.340 24.430 91.360 ;
        RECT 19.610 90.140 20.170 91.280 ;
        RECT 23.050 90.930 23.740 91.340 ;
        RECT 24.730 91.155 25.250 93.565 ;
        RECT 25.510 91.360 25.740 93.360 ;
        RECT 26.060 91.155 26.580 93.565 ;
        RECT 26.940 93.360 28.740 95.300 ;
        RECT 29.100 95.095 29.620 97.505 ;
        RECT 29.940 95.300 30.170 97.300 ;
        RECT 30.430 95.095 30.950 97.505 ;
        RECT 31.250 97.300 32.970 97.320 ;
        RECT 31.230 96.870 32.970 97.300 ;
        RECT 33.180 97.260 34.020 97.540 ;
        RECT 33.120 97.030 34.080 97.260 ;
        RECT 34.410 97.030 35.370 97.260 ;
        RECT 31.230 95.870 33.070 96.870 ;
        RECT 31.230 95.300 32.970 95.870 ;
        RECT 33.360 95.710 33.880 97.030 ;
        RECT 34.130 95.870 34.360 96.870 ;
        RECT 34.630 95.710 35.150 97.030 ;
        RECT 35.530 96.870 36.070 98.140 ;
        RECT 35.420 95.870 36.070 96.870 ;
        RECT 33.120 95.480 34.080 95.710 ;
        RECT 34.410 95.480 35.370 95.710 ;
        RECT 35.530 95.340 36.070 95.870 ;
        RECT 31.250 95.280 32.970 95.300 ;
        RECT 28.930 94.865 29.890 95.095 ;
        RECT 30.220 94.865 31.180 95.095 ;
        RECT 31.940 94.870 32.630 95.280 ;
        RECT 35.520 95.220 36.070 95.340 ;
        RECT 31.930 94.250 32.630 94.870 ;
        RECT 28.930 93.445 29.890 93.675 ;
        RECT 30.220 93.650 31.180 93.675 ;
        RECT 31.940 93.650 32.630 94.250 ;
        RECT 35.510 94.080 36.070 95.220 ;
        RECT 30.220 93.480 34.020 93.650 ;
        RECT 30.220 93.445 31.180 93.480 ;
        RECT 26.800 93.240 28.740 93.360 ;
        RECT 26.800 91.360 28.880 93.240 ;
        RECT 26.940 91.240 28.880 91.360 ;
        RECT 23.050 90.310 23.750 90.930 ;
        RECT 24.500 90.925 25.460 91.155 ;
        RECT 25.790 90.925 26.750 91.155 ;
        RECT 19.610 88.880 20.150 90.140 ;
        RECT 23.050 89.720 23.740 90.310 ;
        RECT 24.500 89.720 25.460 89.745 ;
        RECT 21.660 89.550 25.460 89.720 ;
        RECT 21.660 89.270 22.500 89.550 ;
        RECT 24.500 89.515 25.460 89.550 ;
        RECT 25.790 89.515 26.750 89.745 ;
        RECT 22.710 89.310 24.430 89.330 ;
        RECT 20.310 89.040 21.270 89.270 ;
        RECT 21.600 89.040 22.560 89.270 ;
        RECT 19.610 87.880 20.260 88.880 ;
        RECT 19.610 87.350 20.150 87.880 ;
        RECT 20.530 87.720 21.050 89.040 ;
        RECT 21.320 87.880 21.550 88.880 ;
        RECT 21.800 87.720 22.320 89.040 ;
        RECT 22.710 88.880 24.450 89.310 ;
        RECT 22.610 87.880 24.450 88.880 ;
        RECT 20.310 87.490 21.270 87.720 ;
        RECT 21.600 87.490 22.560 87.720 ;
        RECT 19.610 87.230 20.160 87.350 ;
        RECT 22.710 87.310 24.450 87.880 ;
        RECT 22.710 87.290 24.430 87.310 ;
        RECT 19.610 86.090 20.170 87.230 ;
        RECT 23.050 86.880 23.740 87.290 ;
        RECT 24.730 87.105 25.250 89.515 ;
        RECT 25.510 87.310 25.740 89.310 ;
        RECT 26.060 87.105 26.580 89.515 ;
        RECT 26.940 89.310 28.740 91.240 ;
        RECT 29.100 91.035 29.620 93.445 ;
        RECT 29.940 91.240 30.170 93.240 ;
        RECT 30.430 91.035 30.950 93.445 ;
        RECT 31.250 93.240 32.970 93.260 ;
        RECT 31.230 92.810 32.970 93.240 ;
        RECT 33.180 93.200 34.020 93.480 ;
        RECT 33.120 92.970 34.080 93.200 ;
        RECT 34.410 92.970 35.370 93.200 ;
        RECT 31.230 91.810 33.070 92.810 ;
        RECT 31.230 91.240 32.970 91.810 ;
        RECT 33.360 91.650 33.880 92.970 ;
        RECT 34.130 91.810 34.360 92.810 ;
        RECT 34.630 91.650 35.150 92.970 ;
        RECT 35.530 92.810 36.070 94.080 ;
        RECT 35.420 91.810 36.070 92.810 ;
        RECT 33.120 91.420 34.080 91.650 ;
        RECT 34.410 91.420 35.370 91.650 ;
        RECT 35.530 91.280 36.070 91.810 ;
        RECT 31.250 91.220 32.970 91.240 ;
        RECT 28.930 90.805 29.890 91.035 ;
        RECT 30.220 90.805 31.180 91.035 ;
        RECT 31.940 90.810 32.630 91.220 ;
        RECT 35.520 91.160 36.070 91.280 ;
        RECT 31.930 90.190 32.630 90.810 ;
        RECT 28.930 89.385 29.890 89.615 ;
        RECT 30.220 89.590 31.180 89.615 ;
        RECT 31.940 89.590 32.630 90.190 ;
        RECT 35.510 90.020 36.070 91.160 ;
        RECT 30.220 89.420 34.020 89.590 ;
        RECT 30.220 89.385 31.180 89.420 ;
        RECT 26.800 89.180 28.740 89.310 ;
        RECT 26.800 87.310 28.880 89.180 ;
        RECT 26.940 87.180 28.880 87.310 ;
        RECT 23.050 86.260 23.750 86.880 ;
        RECT 24.500 86.875 25.460 87.105 ;
        RECT 25.790 86.875 26.750 87.105 ;
        RECT 19.610 84.830 20.150 86.090 ;
        RECT 23.050 85.670 23.740 86.260 ;
        RECT 24.500 85.670 25.460 85.695 ;
        RECT 21.660 85.500 25.460 85.670 ;
        RECT 21.660 85.220 22.500 85.500 ;
        RECT 24.500 85.465 25.460 85.500 ;
        RECT 25.790 85.465 26.750 85.695 ;
        RECT 22.710 85.260 24.430 85.280 ;
        RECT 20.310 84.990 21.270 85.220 ;
        RECT 21.600 84.990 22.560 85.220 ;
        RECT 19.610 83.830 20.260 84.830 ;
        RECT 19.610 83.300 20.150 83.830 ;
        RECT 20.530 83.670 21.050 84.990 ;
        RECT 21.320 83.830 21.550 84.830 ;
        RECT 21.800 83.670 22.320 84.990 ;
        RECT 22.710 84.830 24.450 85.260 ;
        RECT 22.610 83.830 24.450 84.830 ;
        RECT 20.310 83.440 21.270 83.670 ;
        RECT 21.600 83.440 22.560 83.670 ;
        RECT 19.610 83.180 20.160 83.300 ;
        RECT 22.710 83.260 24.450 83.830 ;
        RECT 22.710 83.240 24.430 83.260 ;
        RECT 19.610 82.040 20.170 83.180 ;
        RECT 23.050 82.830 23.740 83.240 ;
        RECT 24.730 83.055 25.250 85.465 ;
        RECT 25.510 83.260 25.740 85.260 ;
        RECT 26.060 83.055 26.580 85.465 ;
        RECT 26.940 85.260 28.740 87.180 ;
        RECT 29.100 86.975 29.620 89.385 ;
        RECT 29.940 87.180 30.170 89.180 ;
        RECT 30.430 86.975 30.950 89.385 ;
        RECT 31.250 89.180 32.970 89.200 ;
        RECT 31.230 88.750 32.970 89.180 ;
        RECT 33.180 89.140 34.020 89.420 ;
        RECT 33.120 88.910 34.080 89.140 ;
        RECT 34.410 88.910 35.370 89.140 ;
        RECT 31.230 87.750 33.070 88.750 ;
        RECT 31.230 87.180 32.970 87.750 ;
        RECT 33.360 87.590 33.880 88.910 ;
        RECT 34.130 87.750 34.360 88.750 ;
        RECT 34.630 87.590 35.150 88.910 ;
        RECT 35.530 88.750 36.070 90.020 ;
        RECT 35.420 87.750 36.070 88.750 ;
        RECT 33.120 87.360 34.080 87.590 ;
        RECT 34.410 87.360 35.370 87.590 ;
        RECT 35.530 87.220 36.070 87.750 ;
        RECT 31.250 87.160 32.970 87.180 ;
        RECT 28.930 86.745 29.890 86.975 ;
        RECT 30.220 86.745 31.180 86.975 ;
        RECT 31.940 86.750 32.630 87.160 ;
        RECT 35.520 87.100 36.070 87.220 ;
        RECT 31.930 86.130 32.630 86.750 ;
        RECT 28.930 85.325 29.890 85.555 ;
        RECT 30.220 85.530 31.180 85.555 ;
        RECT 31.940 85.530 32.630 86.130 ;
        RECT 35.510 85.960 36.070 87.100 ;
        RECT 30.220 85.360 34.020 85.530 ;
        RECT 30.220 85.325 31.180 85.360 ;
        RECT 26.800 85.120 28.740 85.260 ;
        RECT 26.800 83.260 28.880 85.120 ;
        RECT 26.940 83.120 28.880 83.260 ;
        RECT 23.050 82.210 23.750 82.830 ;
        RECT 24.500 82.825 25.460 83.055 ;
        RECT 25.790 82.825 26.750 83.055 ;
        RECT 19.610 80.780 20.150 82.040 ;
        RECT 23.050 81.620 23.740 82.210 ;
        RECT 24.500 81.620 25.460 81.645 ;
        RECT 21.660 81.450 25.460 81.620 ;
        RECT 21.660 81.170 22.500 81.450 ;
        RECT 24.500 81.415 25.460 81.450 ;
        RECT 25.790 81.415 26.750 81.645 ;
        RECT 22.710 81.210 24.430 81.230 ;
        RECT 20.310 80.940 21.270 81.170 ;
        RECT 21.600 80.940 22.560 81.170 ;
        RECT 19.610 79.780 20.260 80.780 ;
        RECT 19.610 79.250 20.150 79.780 ;
        RECT 20.530 79.620 21.050 80.940 ;
        RECT 21.320 79.780 21.550 80.780 ;
        RECT 21.800 79.620 22.320 80.940 ;
        RECT 22.710 80.780 24.450 81.210 ;
        RECT 22.610 79.780 24.450 80.780 ;
        RECT 20.310 79.390 21.270 79.620 ;
        RECT 21.600 79.390 22.560 79.620 ;
        RECT 19.610 79.130 20.160 79.250 ;
        RECT 22.710 79.210 24.450 79.780 ;
        RECT 22.710 79.190 24.430 79.210 ;
        RECT 19.610 77.990 20.170 79.130 ;
        RECT 23.050 78.780 23.740 79.190 ;
        RECT 24.730 79.005 25.250 81.415 ;
        RECT 25.510 79.210 25.740 81.210 ;
        RECT 26.060 79.005 26.580 81.415 ;
        RECT 26.940 81.210 28.740 83.120 ;
        RECT 29.100 82.915 29.620 85.325 ;
        RECT 29.940 83.120 30.170 85.120 ;
        RECT 30.430 82.915 30.950 85.325 ;
        RECT 31.250 85.120 32.970 85.140 ;
        RECT 31.230 84.690 32.970 85.120 ;
        RECT 33.180 85.080 34.020 85.360 ;
        RECT 33.120 84.850 34.080 85.080 ;
        RECT 34.410 84.850 35.370 85.080 ;
        RECT 31.230 83.690 33.070 84.690 ;
        RECT 31.230 83.120 32.970 83.690 ;
        RECT 33.360 83.530 33.880 84.850 ;
        RECT 34.130 83.690 34.360 84.690 ;
        RECT 34.630 83.530 35.150 84.850 ;
        RECT 35.530 84.690 36.070 85.960 ;
        RECT 35.420 83.690 36.070 84.690 ;
        RECT 33.120 83.300 34.080 83.530 ;
        RECT 34.410 83.300 35.370 83.530 ;
        RECT 35.530 83.160 36.070 83.690 ;
        RECT 31.250 83.100 32.970 83.120 ;
        RECT 28.930 82.685 29.890 82.915 ;
        RECT 30.220 82.685 31.180 82.915 ;
        RECT 31.940 82.690 32.630 83.100 ;
        RECT 35.520 83.040 36.070 83.160 ;
        RECT 31.930 82.070 32.630 82.690 ;
        RECT 28.930 81.265 29.890 81.495 ;
        RECT 30.220 81.470 31.180 81.495 ;
        RECT 31.940 81.470 32.630 82.070 ;
        RECT 35.510 81.900 36.070 83.040 ;
        RECT 30.220 81.300 34.020 81.470 ;
        RECT 30.220 81.265 31.180 81.300 ;
        RECT 26.800 81.060 28.740 81.210 ;
        RECT 26.800 79.210 28.880 81.060 ;
        RECT 26.940 79.060 28.880 79.210 ;
        RECT 23.050 78.160 23.750 78.780 ;
        RECT 24.500 78.775 25.460 79.005 ;
        RECT 25.790 78.775 26.750 79.005 ;
        RECT 19.610 76.730 20.150 77.990 ;
        RECT 23.050 77.570 23.740 78.160 ;
        RECT 24.500 77.570 25.460 77.595 ;
        RECT 21.660 77.400 25.460 77.570 ;
        RECT 21.660 77.120 22.500 77.400 ;
        RECT 24.500 77.365 25.460 77.400 ;
        RECT 25.790 77.365 26.750 77.595 ;
        RECT 22.710 77.160 24.430 77.180 ;
        RECT 20.310 76.890 21.270 77.120 ;
        RECT 21.600 76.890 22.560 77.120 ;
        RECT 19.610 75.730 20.260 76.730 ;
        RECT 19.610 75.200 20.150 75.730 ;
        RECT 20.530 75.570 21.050 76.890 ;
        RECT 21.320 75.730 21.550 76.730 ;
        RECT 21.800 75.570 22.320 76.890 ;
        RECT 22.710 76.730 24.450 77.160 ;
        RECT 22.610 75.730 24.450 76.730 ;
        RECT 20.310 75.340 21.270 75.570 ;
        RECT 21.600 75.340 22.560 75.570 ;
        RECT 19.610 75.080 20.160 75.200 ;
        RECT 22.710 75.160 24.450 75.730 ;
        RECT 22.710 75.140 24.430 75.160 ;
        RECT 19.610 73.940 20.170 75.080 ;
        RECT 23.050 74.730 23.740 75.140 ;
        RECT 24.730 74.955 25.250 77.365 ;
        RECT 25.510 75.160 25.740 77.160 ;
        RECT 26.060 74.955 26.580 77.365 ;
        RECT 26.940 77.160 28.740 79.060 ;
        RECT 29.100 78.855 29.620 81.265 ;
        RECT 29.940 79.060 30.170 81.060 ;
        RECT 30.430 78.855 30.950 81.265 ;
        RECT 31.250 81.060 32.970 81.080 ;
        RECT 31.230 80.630 32.970 81.060 ;
        RECT 33.180 81.020 34.020 81.300 ;
        RECT 33.120 80.790 34.080 81.020 ;
        RECT 34.410 80.790 35.370 81.020 ;
        RECT 31.230 79.630 33.070 80.630 ;
        RECT 31.230 79.060 32.970 79.630 ;
        RECT 33.360 79.470 33.880 80.790 ;
        RECT 34.130 79.630 34.360 80.630 ;
        RECT 34.630 79.470 35.150 80.790 ;
        RECT 35.530 80.630 36.070 81.900 ;
        RECT 35.420 79.630 36.070 80.630 ;
        RECT 33.120 79.240 34.080 79.470 ;
        RECT 34.410 79.240 35.370 79.470 ;
        RECT 35.530 79.100 36.070 79.630 ;
        RECT 31.250 79.040 32.970 79.060 ;
        RECT 28.930 78.625 29.890 78.855 ;
        RECT 30.220 78.625 31.180 78.855 ;
        RECT 31.940 78.630 32.630 79.040 ;
        RECT 35.520 78.980 36.070 79.100 ;
        RECT 31.930 78.010 32.630 78.630 ;
        RECT 28.930 77.205 29.890 77.435 ;
        RECT 30.220 77.410 31.180 77.435 ;
        RECT 31.940 77.410 32.630 78.010 ;
        RECT 35.510 77.840 36.070 78.980 ;
        RECT 30.220 77.240 34.020 77.410 ;
        RECT 30.220 77.205 31.180 77.240 ;
        RECT 26.800 77.000 28.740 77.160 ;
        RECT 26.800 75.160 28.880 77.000 ;
        RECT 26.940 75.000 28.880 75.160 ;
        RECT 23.050 74.110 23.750 74.730 ;
        RECT 24.500 74.725 25.460 74.955 ;
        RECT 25.790 74.725 26.750 74.955 ;
        RECT 19.610 72.680 20.150 73.940 ;
        RECT 23.050 73.520 23.740 74.110 ;
        RECT 24.500 73.520 25.460 73.545 ;
        RECT 21.660 73.350 25.460 73.520 ;
        RECT 21.660 73.070 22.500 73.350 ;
        RECT 24.500 73.315 25.460 73.350 ;
        RECT 25.790 73.315 26.750 73.545 ;
        RECT 22.710 73.110 24.430 73.130 ;
        RECT 20.310 72.840 21.270 73.070 ;
        RECT 21.600 72.840 22.560 73.070 ;
        RECT 19.610 71.680 20.260 72.680 ;
        RECT 19.610 71.150 20.150 71.680 ;
        RECT 20.530 71.520 21.050 72.840 ;
        RECT 21.320 71.680 21.550 72.680 ;
        RECT 21.800 71.520 22.320 72.840 ;
        RECT 22.710 72.680 24.450 73.110 ;
        RECT 22.610 71.680 24.450 72.680 ;
        RECT 20.310 71.290 21.270 71.520 ;
        RECT 21.600 71.290 22.560 71.520 ;
        RECT 19.610 71.030 20.160 71.150 ;
        RECT 22.710 71.110 24.450 71.680 ;
        RECT 22.710 71.090 24.430 71.110 ;
        RECT 19.610 69.890 20.170 71.030 ;
        RECT 23.050 70.680 23.740 71.090 ;
        RECT 24.730 70.905 25.250 73.315 ;
        RECT 25.510 71.110 25.740 73.110 ;
        RECT 26.060 70.905 26.580 73.315 ;
        RECT 26.940 73.110 28.740 75.000 ;
        RECT 29.100 74.795 29.620 77.205 ;
        RECT 29.940 75.000 30.170 77.000 ;
        RECT 30.430 74.795 30.950 77.205 ;
        RECT 31.250 77.000 32.970 77.020 ;
        RECT 31.230 76.570 32.970 77.000 ;
        RECT 33.180 76.960 34.020 77.240 ;
        RECT 33.120 76.730 34.080 76.960 ;
        RECT 34.410 76.730 35.370 76.960 ;
        RECT 31.230 75.570 33.070 76.570 ;
        RECT 31.230 75.000 32.970 75.570 ;
        RECT 33.360 75.410 33.880 76.730 ;
        RECT 34.130 75.570 34.360 76.570 ;
        RECT 34.630 75.410 35.150 76.730 ;
        RECT 35.530 76.570 36.070 77.840 ;
        RECT 35.420 75.570 36.070 76.570 ;
        RECT 33.120 75.180 34.080 75.410 ;
        RECT 34.410 75.180 35.370 75.410 ;
        RECT 35.530 75.040 36.070 75.570 ;
        RECT 31.250 74.980 32.970 75.000 ;
        RECT 28.930 74.565 29.890 74.795 ;
        RECT 30.220 74.565 31.180 74.795 ;
        RECT 31.940 74.570 32.630 74.980 ;
        RECT 35.520 74.920 36.070 75.040 ;
        RECT 31.930 73.950 32.630 74.570 ;
        RECT 28.930 73.145 29.890 73.375 ;
        RECT 30.220 73.350 31.180 73.375 ;
        RECT 31.940 73.350 32.630 73.950 ;
        RECT 35.510 73.780 36.070 74.920 ;
        RECT 30.220 73.180 34.020 73.350 ;
        RECT 30.220 73.145 31.180 73.180 ;
        RECT 26.800 72.940 28.740 73.110 ;
        RECT 26.800 71.110 28.880 72.940 ;
        RECT 26.940 70.940 28.880 71.110 ;
        RECT 23.050 70.060 23.750 70.680 ;
        RECT 24.500 70.675 25.460 70.905 ;
        RECT 25.790 70.675 26.750 70.905 ;
        RECT 19.610 68.630 20.150 69.890 ;
        RECT 23.050 69.470 23.740 70.060 ;
        RECT 24.500 69.470 25.460 69.495 ;
        RECT 21.660 69.300 25.460 69.470 ;
        RECT 21.660 69.020 22.500 69.300 ;
        RECT 24.500 69.265 25.460 69.300 ;
        RECT 25.790 69.265 26.750 69.495 ;
        RECT 22.710 69.060 24.430 69.080 ;
        RECT 20.310 68.790 21.270 69.020 ;
        RECT 21.600 68.790 22.560 69.020 ;
        RECT 19.610 67.630 20.260 68.630 ;
        RECT 19.610 67.100 20.150 67.630 ;
        RECT 20.530 67.470 21.050 68.790 ;
        RECT 21.320 67.630 21.550 68.630 ;
        RECT 21.800 67.470 22.320 68.790 ;
        RECT 22.710 68.630 24.450 69.060 ;
        RECT 22.610 67.630 24.450 68.630 ;
        RECT 20.310 67.240 21.270 67.470 ;
        RECT 21.600 67.240 22.560 67.470 ;
        RECT 19.610 66.980 20.160 67.100 ;
        RECT 22.710 67.060 24.450 67.630 ;
        RECT 22.710 67.040 24.430 67.060 ;
        RECT 19.610 65.840 20.170 66.980 ;
        RECT 23.050 66.630 23.740 67.040 ;
        RECT 24.730 66.855 25.250 69.265 ;
        RECT 25.510 67.060 25.740 69.060 ;
        RECT 26.060 66.855 26.580 69.265 ;
        RECT 26.940 69.060 28.740 70.940 ;
        RECT 29.100 70.735 29.620 73.145 ;
        RECT 29.940 70.940 30.170 72.940 ;
        RECT 30.430 70.735 30.950 73.145 ;
        RECT 31.250 72.940 32.970 72.960 ;
        RECT 31.230 72.510 32.970 72.940 ;
        RECT 33.180 72.900 34.020 73.180 ;
        RECT 33.120 72.670 34.080 72.900 ;
        RECT 34.410 72.670 35.370 72.900 ;
        RECT 31.230 71.510 33.070 72.510 ;
        RECT 31.230 70.940 32.970 71.510 ;
        RECT 33.360 71.350 33.880 72.670 ;
        RECT 34.130 71.510 34.360 72.510 ;
        RECT 34.630 71.350 35.150 72.670 ;
        RECT 35.530 72.510 36.070 73.780 ;
        RECT 35.420 71.510 36.070 72.510 ;
        RECT 33.120 71.120 34.080 71.350 ;
        RECT 34.410 71.120 35.370 71.350 ;
        RECT 35.530 70.980 36.070 71.510 ;
        RECT 31.250 70.920 32.970 70.940 ;
        RECT 28.930 70.505 29.890 70.735 ;
        RECT 30.220 70.505 31.180 70.735 ;
        RECT 31.940 70.510 32.630 70.920 ;
        RECT 35.520 70.860 36.070 70.980 ;
        RECT 31.930 69.890 32.630 70.510 ;
        RECT 28.930 69.085 29.890 69.315 ;
        RECT 30.220 69.290 31.180 69.315 ;
        RECT 31.940 69.290 32.630 69.890 ;
        RECT 35.510 69.720 36.070 70.860 ;
        RECT 30.220 69.120 34.020 69.290 ;
        RECT 30.220 69.085 31.180 69.120 ;
        RECT 26.800 68.880 28.740 69.060 ;
        RECT 26.800 67.060 28.880 68.880 ;
        RECT 26.940 66.880 28.880 67.060 ;
        RECT 23.050 66.010 23.750 66.630 ;
        RECT 24.500 66.625 25.460 66.855 ;
        RECT 25.790 66.625 26.750 66.855 ;
        RECT 19.610 64.580 20.150 65.840 ;
        RECT 23.050 65.420 23.740 66.010 ;
        RECT 24.500 65.420 25.460 65.445 ;
        RECT 21.660 65.250 25.460 65.420 ;
        RECT 21.660 64.970 22.500 65.250 ;
        RECT 24.500 65.215 25.460 65.250 ;
        RECT 25.790 65.215 26.750 65.445 ;
        RECT 22.710 65.010 24.430 65.030 ;
        RECT 20.310 64.740 21.270 64.970 ;
        RECT 21.600 64.740 22.560 64.970 ;
        RECT 19.610 63.580 20.260 64.580 ;
        RECT 19.610 63.050 20.150 63.580 ;
        RECT 20.530 63.420 21.050 64.740 ;
        RECT 21.320 63.580 21.550 64.580 ;
        RECT 21.800 63.420 22.320 64.740 ;
        RECT 22.710 64.580 24.450 65.010 ;
        RECT 22.610 63.580 24.450 64.580 ;
        RECT 20.310 63.190 21.270 63.420 ;
        RECT 21.600 63.190 22.560 63.420 ;
        RECT 19.610 62.930 20.160 63.050 ;
        RECT 22.710 63.010 24.450 63.580 ;
        RECT 22.710 62.990 24.430 63.010 ;
        RECT 19.610 61.790 20.170 62.930 ;
        RECT 23.050 62.580 23.740 62.990 ;
        RECT 24.730 62.805 25.250 65.215 ;
        RECT 25.510 63.010 25.740 65.010 ;
        RECT 26.060 62.805 26.580 65.215 ;
        RECT 26.940 65.010 28.740 66.880 ;
        RECT 29.100 66.675 29.620 69.085 ;
        RECT 29.940 66.880 30.170 68.880 ;
        RECT 30.430 66.675 30.950 69.085 ;
        RECT 31.250 68.880 32.970 68.900 ;
        RECT 31.230 68.450 32.970 68.880 ;
        RECT 33.180 68.840 34.020 69.120 ;
        RECT 33.120 68.610 34.080 68.840 ;
        RECT 34.410 68.610 35.370 68.840 ;
        RECT 31.230 67.450 33.070 68.450 ;
        RECT 31.230 66.880 32.970 67.450 ;
        RECT 33.360 67.290 33.880 68.610 ;
        RECT 34.130 67.450 34.360 68.450 ;
        RECT 34.630 67.290 35.150 68.610 ;
        RECT 35.530 68.450 36.070 69.720 ;
        RECT 35.420 67.450 36.070 68.450 ;
        RECT 33.120 67.060 34.080 67.290 ;
        RECT 34.410 67.060 35.370 67.290 ;
        RECT 35.530 66.920 36.070 67.450 ;
        RECT 31.250 66.860 32.970 66.880 ;
        RECT 28.930 66.445 29.890 66.675 ;
        RECT 30.220 66.445 31.180 66.675 ;
        RECT 31.940 66.450 32.630 66.860 ;
        RECT 35.520 66.800 36.070 66.920 ;
        RECT 31.930 65.830 32.630 66.450 ;
        RECT 28.930 65.025 29.890 65.255 ;
        RECT 30.220 65.230 31.180 65.255 ;
        RECT 31.940 65.230 32.630 65.830 ;
        RECT 35.510 65.660 36.070 66.800 ;
        RECT 30.220 65.060 34.020 65.230 ;
        RECT 30.220 65.025 31.180 65.060 ;
        RECT 26.800 64.820 28.740 65.010 ;
        RECT 26.800 63.010 28.880 64.820 ;
        RECT 26.940 62.820 28.880 63.010 ;
        RECT 23.050 61.960 23.750 62.580 ;
        RECT 24.500 62.575 25.460 62.805 ;
        RECT 25.790 62.575 26.750 62.805 ;
        RECT 19.610 60.530 20.150 61.790 ;
        RECT 23.050 61.370 23.740 61.960 ;
        RECT 24.500 61.370 25.460 61.395 ;
        RECT 21.660 61.200 25.460 61.370 ;
        RECT 21.660 60.920 22.500 61.200 ;
        RECT 24.500 61.165 25.460 61.200 ;
        RECT 25.790 61.165 26.750 61.395 ;
        RECT 22.710 60.960 24.430 60.980 ;
        RECT 20.310 60.690 21.270 60.920 ;
        RECT 21.600 60.690 22.560 60.920 ;
        RECT 19.610 59.530 20.260 60.530 ;
        RECT 19.610 59.000 20.150 59.530 ;
        RECT 20.530 59.370 21.050 60.690 ;
        RECT 21.320 59.530 21.550 60.530 ;
        RECT 21.800 59.370 22.320 60.690 ;
        RECT 22.710 60.530 24.450 60.960 ;
        RECT 22.610 59.530 24.450 60.530 ;
        RECT 20.310 59.140 21.270 59.370 ;
        RECT 21.600 59.140 22.560 59.370 ;
        RECT 19.610 58.880 20.160 59.000 ;
        RECT 22.710 58.960 24.450 59.530 ;
        RECT 22.710 58.940 24.430 58.960 ;
        RECT 19.610 57.740 20.170 58.880 ;
        RECT 23.050 58.530 23.740 58.940 ;
        RECT 24.730 58.755 25.250 61.165 ;
        RECT 25.510 58.960 25.740 60.960 ;
        RECT 26.060 58.755 26.580 61.165 ;
        RECT 26.940 60.960 28.740 62.820 ;
        RECT 29.100 62.615 29.620 65.025 ;
        RECT 29.940 62.820 30.170 64.820 ;
        RECT 30.430 62.615 30.950 65.025 ;
        RECT 31.250 64.820 32.970 64.840 ;
        RECT 31.230 64.390 32.970 64.820 ;
        RECT 33.180 64.780 34.020 65.060 ;
        RECT 33.120 64.550 34.080 64.780 ;
        RECT 34.410 64.550 35.370 64.780 ;
        RECT 31.230 63.390 33.070 64.390 ;
        RECT 31.230 62.820 32.970 63.390 ;
        RECT 33.360 63.230 33.880 64.550 ;
        RECT 34.130 63.390 34.360 64.390 ;
        RECT 34.630 63.230 35.150 64.550 ;
        RECT 35.530 64.390 36.070 65.660 ;
        RECT 35.420 63.390 36.070 64.390 ;
        RECT 33.120 63.000 34.080 63.230 ;
        RECT 34.410 63.000 35.370 63.230 ;
        RECT 35.530 62.860 36.070 63.390 ;
        RECT 31.250 62.800 32.970 62.820 ;
        RECT 28.930 62.385 29.890 62.615 ;
        RECT 30.220 62.385 31.180 62.615 ;
        RECT 31.940 62.390 32.630 62.800 ;
        RECT 35.520 62.740 36.070 62.860 ;
        RECT 31.930 61.770 32.630 62.390 ;
        RECT 28.930 60.965 29.890 61.195 ;
        RECT 30.220 61.170 31.180 61.195 ;
        RECT 31.940 61.170 32.630 61.770 ;
        RECT 35.510 61.600 36.070 62.740 ;
        RECT 30.220 61.000 34.020 61.170 ;
        RECT 30.220 60.965 31.180 61.000 ;
        RECT 26.800 60.760 28.740 60.960 ;
        RECT 26.800 58.960 28.880 60.760 ;
        RECT 26.940 58.760 28.880 58.960 ;
        RECT 23.050 57.910 23.750 58.530 ;
        RECT 24.500 58.525 25.460 58.755 ;
        RECT 25.790 58.525 26.750 58.755 ;
        RECT 26.940 58.160 28.740 58.760 ;
        RECT 29.100 58.555 29.620 60.965 ;
        RECT 29.940 58.760 30.170 60.760 ;
        RECT 30.430 58.555 30.950 60.965 ;
        RECT 31.250 60.760 32.970 60.780 ;
        RECT 31.230 60.330 32.970 60.760 ;
        RECT 33.180 60.720 34.020 61.000 ;
        RECT 33.120 60.490 34.080 60.720 ;
        RECT 34.410 60.490 35.370 60.720 ;
        RECT 31.230 59.330 33.070 60.330 ;
        RECT 31.230 58.760 32.970 59.330 ;
        RECT 33.360 59.170 33.880 60.490 ;
        RECT 34.130 59.330 34.360 60.330 ;
        RECT 34.630 59.170 35.150 60.490 ;
        RECT 35.530 60.330 36.070 61.600 ;
        RECT 35.420 59.330 36.070 60.330 ;
        RECT 33.120 58.940 34.080 59.170 ;
        RECT 34.410 58.940 35.370 59.170 ;
        RECT 35.530 58.800 36.070 59.330 ;
        RECT 31.250 58.740 32.970 58.760 ;
        RECT 28.930 58.325 29.890 58.555 ;
        RECT 30.220 58.325 31.180 58.555 ;
        RECT 31.940 58.330 32.630 58.740 ;
        RECT 35.520 58.680 36.070 58.800 ;
        RECT 19.610 56.480 20.150 57.740 ;
        RECT 23.050 57.320 23.740 57.910 ;
        RECT 24.500 57.320 25.460 57.345 ;
        RECT 21.660 57.150 25.460 57.320 ;
        RECT 21.660 56.870 22.500 57.150 ;
        RECT 24.500 57.115 25.460 57.150 ;
        RECT 25.790 57.115 26.750 57.345 ;
        RECT 22.710 56.910 24.430 56.930 ;
        RECT 20.310 56.640 21.270 56.870 ;
        RECT 21.600 56.640 22.560 56.870 ;
        RECT 19.610 55.480 20.260 56.480 ;
        RECT 19.610 54.950 20.150 55.480 ;
        RECT 20.530 55.320 21.050 56.640 ;
        RECT 21.320 55.480 21.550 56.480 ;
        RECT 21.800 55.320 22.320 56.640 ;
        RECT 22.710 56.480 24.450 56.910 ;
        RECT 22.610 55.480 24.450 56.480 ;
        RECT 20.310 55.090 21.270 55.320 ;
        RECT 21.600 55.090 22.560 55.320 ;
        RECT 19.610 54.830 20.160 54.950 ;
        RECT 22.710 54.910 24.450 55.480 ;
        RECT 22.710 54.890 24.430 54.910 ;
        RECT 19.610 53.690 20.170 54.830 ;
        RECT 23.050 54.480 23.740 54.890 ;
        RECT 24.730 54.705 25.250 57.115 ;
        RECT 25.510 54.910 25.740 56.910 ;
        RECT 26.060 54.705 26.580 57.115 ;
        RECT 26.940 56.910 28.745 58.160 ;
        RECT 31.930 57.710 32.630 58.330 ;
        RECT 26.800 56.220 28.745 56.910 ;
        RECT 31.935 57.410 32.625 57.710 ;
        RECT 35.510 57.540 36.070 58.680 ;
        RECT 28.930 56.425 29.890 56.655 ;
        RECT 30.220 56.630 31.180 56.655 ;
        RECT 31.935 56.630 32.630 57.410 ;
        RECT 30.220 56.460 34.020 56.630 ;
        RECT 30.220 56.425 31.180 56.460 ;
        RECT 26.800 54.910 28.880 56.220 ;
        RECT 23.050 53.860 23.750 54.480 ;
        RECT 24.500 54.475 25.460 54.705 ;
        RECT 25.790 54.475 26.750 54.705 ;
        RECT 26.940 54.220 28.880 54.910 ;
        RECT 19.610 52.430 20.150 53.690 ;
        RECT 23.050 53.270 23.740 53.860 ;
        RECT 24.500 53.270 25.460 53.295 ;
        RECT 21.660 53.100 25.460 53.270 ;
        RECT 21.660 52.820 22.500 53.100 ;
        RECT 24.500 53.065 25.460 53.100 ;
        RECT 25.790 53.065 26.750 53.295 ;
        RECT 26.940 53.130 28.745 54.220 ;
        RECT 29.100 54.015 29.620 56.425 ;
        RECT 29.940 54.220 30.170 56.220 ;
        RECT 30.430 54.015 30.950 56.425 ;
        RECT 31.250 56.220 32.970 56.240 ;
        RECT 31.230 55.790 32.970 56.220 ;
        RECT 33.180 56.180 34.020 56.460 ;
        RECT 33.120 55.950 34.080 56.180 ;
        RECT 34.410 55.950 35.370 56.180 ;
        RECT 31.230 54.790 33.070 55.790 ;
        RECT 31.230 54.220 32.970 54.790 ;
        RECT 33.360 54.630 33.880 55.950 ;
        RECT 34.130 54.790 34.360 55.790 ;
        RECT 34.630 54.630 35.150 55.950 ;
        RECT 35.530 55.790 36.070 57.540 ;
        RECT 35.420 54.790 36.070 55.790 ;
        RECT 33.120 54.400 34.080 54.630 ;
        RECT 34.410 54.400 35.370 54.630 ;
        RECT 35.530 54.260 36.070 54.790 ;
        RECT 31.250 54.200 32.970 54.220 ;
        RECT 28.930 53.785 29.890 54.015 ;
        RECT 30.220 53.785 31.180 54.015 ;
        RECT 31.655 53.180 32.750 54.200 ;
        RECT 35.520 54.140 36.070 54.260 ;
        RECT 22.710 52.860 24.430 52.880 ;
        RECT 20.310 52.590 21.270 52.820 ;
        RECT 21.600 52.590 22.560 52.820 ;
        RECT 19.610 51.430 20.260 52.430 ;
        RECT 19.610 50.900 20.150 51.430 ;
        RECT 20.530 51.270 21.050 52.590 ;
        RECT 21.320 51.430 21.550 52.430 ;
        RECT 21.800 51.270 22.320 52.590 ;
        RECT 22.710 52.430 24.450 52.860 ;
        RECT 22.610 51.430 24.450 52.430 ;
        RECT 20.310 51.040 21.270 51.270 ;
        RECT 21.600 51.040 22.560 51.270 ;
        RECT 19.610 50.780 20.160 50.900 ;
        RECT 22.710 50.860 24.450 51.430 ;
        RECT 22.710 50.840 24.430 50.860 ;
        RECT 19.610 49.640 20.170 50.780 ;
        RECT 23.050 50.430 23.740 50.840 ;
        RECT 24.730 50.655 25.250 53.065 ;
        RECT 25.510 50.860 25.740 52.860 ;
        RECT 26.060 50.655 26.580 53.065 ;
        RECT 26.940 53.000 28.740 53.130 ;
        RECT 26.940 52.860 27.840 53.000 ;
        RECT 26.800 50.860 27.840 52.860 ;
        RECT 31.690 51.665 32.750 53.180 ;
        RECT 35.510 53.000 36.070 54.140 ;
        RECT 23.050 49.810 23.750 50.430 ;
        RECT 24.500 50.425 25.460 50.655 ;
        RECT 25.790 50.425 26.750 50.655 ;
        RECT 19.610 48.380 20.150 49.640 ;
        RECT 23.050 49.220 23.740 49.810 ;
        RECT 24.500 49.220 25.460 49.245 ;
        RECT 21.660 49.050 25.460 49.220 ;
        RECT 21.660 48.770 22.500 49.050 ;
        RECT 24.500 49.015 25.460 49.050 ;
        RECT 25.790 49.015 26.750 49.245 ;
        RECT 22.710 48.810 24.430 48.830 ;
        RECT 20.310 48.540 21.270 48.770 ;
        RECT 21.600 48.540 22.560 48.770 ;
        RECT 19.610 47.380 20.260 48.380 ;
        RECT 19.610 46.850 20.150 47.380 ;
        RECT 20.530 47.220 21.050 48.540 ;
        RECT 21.320 47.380 21.550 48.380 ;
        RECT 21.800 47.220 22.320 48.540 ;
        RECT 22.710 48.380 24.450 48.810 ;
        RECT 22.610 47.380 24.450 48.380 ;
        RECT 20.310 46.990 21.270 47.220 ;
        RECT 21.600 46.990 22.560 47.220 ;
        RECT 19.610 46.730 20.160 46.850 ;
        RECT 22.710 46.810 24.450 47.380 ;
        RECT 22.710 46.790 24.430 46.810 ;
        RECT 19.610 45.590 20.170 46.730 ;
        RECT 23.050 46.380 23.740 46.790 ;
        RECT 24.730 46.605 25.250 49.015 ;
        RECT 25.510 46.810 25.740 48.810 ;
        RECT 26.060 46.605 26.580 49.015 ;
        RECT 26.940 48.810 27.840 50.860 ;
        RECT 26.800 46.810 27.840 48.810 ;
        RECT 23.050 45.760 23.750 46.380 ;
        RECT 24.500 46.375 25.460 46.605 ;
        RECT 25.790 46.375 26.750 46.605 ;
        RECT 19.610 44.330 20.150 45.590 ;
        RECT 23.050 45.170 23.740 45.760 ;
        RECT 24.500 45.170 25.460 45.195 ;
        RECT 21.660 45.000 25.460 45.170 ;
        RECT 21.660 44.720 22.500 45.000 ;
        RECT 24.500 44.965 25.460 45.000 ;
        RECT 25.790 44.965 26.750 45.195 ;
        RECT 22.710 44.760 24.430 44.780 ;
        RECT 20.310 44.490 21.270 44.720 ;
        RECT 21.600 44.490 22.560 44.720 ;
        RECT 19.610 43.330 20.260 44.330 ;
        RECT 19.610 42.800 20.150 43.330 ;
        RECT 20.530 43.170 21.050 44.490 ;
        RECT 21.320 43.330 21.550 44.330 ;
        RECT 21.800 43.170 22.320 44.490 ;
        RECT 22.710 44.330 24.450 44.760 ;
        RECT 22.610 43.330 24.450 44.330 ;
        RECT 20.310 42.940 21.270 43.170 ;
        RECT 21.600 42.940 22.560 43.170 ;
        RECT 19.610 42.680 20.160 42.800 ;
        RECT 22.710 42.760 24.450 43.330 ;
        RECT 22.710 42.740 24.430 42.760 ;
        RECT 19.610 41.540 20.170 42.680 ;
        RECT 23.050 42.330 23.740 42.740 ;
        RECT 24.730 42.555 25.250 44.965 ;
        RECT 25.510 42.760 25.740 44.760 ;
        RECT 26.060 42.555 26.580 44.965 ;
        RECT 26.940 44.760 27.840 46.810 ;
        RECT 26.800 42.760 27.840 44.760 ;
        RECT 31.655 51.580 32.750 51.665 ;
        RECT 31.655 44.375 32.655 51.580 ;
        RECT 23.050 41.710 23.750 42.330 ;
        RECT 24.500 42.325 25.460 42.555 ;
        RECT 25.790 42.325 26.750 42.555 ;
        RECT 19.610 40.280 20.150 41.540 ;
        RECT 23.050 41.120 23.740 41.710 ;
        RECT 24.500 41.120 25.460 41.145 ;
        RECT 21.660 40.950 25.460 41.120 ;
        RECT 21.660 40.670 22.500 40.950 ;
        RECT 24.500 40.915 25.460 40.950 ;
        RECT 25.790 40.915 26.750 41.145 ;
        RECT 22.710 40.710 24.430 40.730 ;
        RECT 20.310 40.440 21.270 40.670 ;
        RECT 21.600 40.440 22.560 40.670 ;
        RECT 19.610 39.280 20.260 40.280 ;
        RECT 19.610 38.750 20.150 39.280 ;
        RECT 20.530 39.120 21.050 40.440 ;
        RECT 21.320 39.280 21.550 40.280 ;
        RECT 21.800 39.120 22.320 40.440 ;
        RECT 22.710 40.280 24.450 40.710 ;
        RECT 22.610 39.280 24.450 40.280 ;
        RECT 20.310 38.890 21.270 39.120 ;
        RECT 21.600 38.890 22.560 39.120 ;
        RECT 19.610 38.630 20.160 38.750 ;
        RECT 22.710 38.710 24.450 39.280 ;
        RECT 22.710 38.690 24.430 38.710 ;
        RECT 19.610 37.490 20.170 38.630 ;
        RECT 23.050 38.280 23.740 38.690 ;
        RECT 24.730 38.505 25.250 40.915 ;
        RECT 25.510 38.710 25.740 40.710 ;
        RECT 26.060 38.505 26.580 40.915 ;
        RECT 26.940 40.710 27.840 42.760 ;
        RECT 26.800 38.710 27.840 40.710 ;
        RECT 23.050 37.660 23.750 38.280 ;
        RECT 24.500 38.275 25.460 38.505 ;
        RECT 25.790 38.275 26.750 38.505 ;
        RECT 19.610 36.230 20.150 37.490 ;
        RECT 23.050 37.070 23.740 37.660 ;
        RECT 24.500 37.070 25.460 37.095 ;
        RECT 21.660 36.900 25.460 37.070 ;
        RECT 21.660 36.620 22.500 36.900 ;
        RECT 24.500 36.865 25.460 36.900 ;
        RECT 25.790 36.865 26.750 37.095 ;
        RECT 22.710 36.660 24.430 36.680 ;
        RECT 20.310 36.390 21.270 36.620 ;
        RECT 21.600 36.390 22.560 36.620 ;
        RECT 19.610 35.230 20.260 36.230 ;
        RECT 19.610 34.700 20.150 35.230 ;
        RECT 20.530 35.070 21.050 36.390 ;
        RECT 21.320 35.230 21.550 36.230 ;
        RECT 21.800 35.070 22.320 36.390 ;
        RECT 22.710 36.230 24.450 36.660 ;
        RECT 22.610 35.230 24.450 36.230 ;
        RECT 20.310 34.840 21.270 35.070 ;
        RECT 21.600 34.840 22.560 35.070 ;
        RECT 19.610 34.580 20.160 34.700 ;
        RECT 22.710 34.660 24.450 35.230 ;
        RECT 22.710 34.640 24.430 34.660 ;
        RECT 19.610 33.440 20.170 34.580 ;
        RECT 23.050 34.230 23.740 34.640 ;
        RECT 24.730 34.455 25.250 36.865 ;
        RECT 25.510 34.660 25.740 36.660 ;
        RECT 26.060 34.455 26.580 36.865 ;
        RECT 26.940 36.660 27.840 38.710 ;
        RECT 26.800 34.660 27.840 36.660 ;
        RECT 23.050 33.610 23.750 34.230 ;
        RECT 24.500 34.225 25.460 34.455 ;
        RECT 25.790 34.225 26.750 34.455 ;
        RECT 19.610 32.180 20.150 33.440 ;
        RECT 23.050 33.020 23.740 33.610 ;
        RECT 24.500 33.020 25.460 33.045 ;
        RECT 21.660 32.850 25.460 33.020 ;
        RECT 21.660 32.570 22.500 32.850 ;
        RECT 24.500 32.815 25.460 32.850 ;
        RECT 25.790 32.815 26.750 33.045 ;
        RECT 22.710 32.610 24.430 32.630 ;
        RECT 20.310 32.340 21.270 32.570 ;
        RECT 21.600 32.340 22.560 32.570 ;
        RECT 19.610 31.180 20.260 32.180 ;
        RECT 19.610 30.650 20.150 31.180 ;
        RECT 20.530 31.020 21.050 32.340 ;
        RECT 21.320 31.180 21.550 32.180 ;
        RECT 21.800 31.020 22.320 32.340 ;
        RECT 22.710 32.180 24.450 32.610 ;
        RECT 22.610 31.180 24.450 32.180 ;
        RECT 20.310 30.790 21.270 31.020 ;
        RECT 21.600 30.790 22.560 31.020 ;
        RECT 19.610 30.530 20.160 30.650 ;
        RECT 22.710 30.610 24.450 31.180 ;
        RECT 22.710 30.590 24.430 30.610 ;
        RECT 19.610 29.390 20.170 30.530 ;
        RECT 23.050 30.180 23.740 30.590 ;
        RECT 24.730 30.405 25.250 32.815 ;
        RECT 25.510 30.610 25.740 32.610 ;
        RECT 26.060 30.405 26.580 32.815 ;
        RECT 26.940 32.610 27.840 34.660 ;
        RECT 26.800 30.610 27.840 32.610 ;
        RECT 23.050 29.560 23.750 30.180 ;
        RECT 24.500 30.175 25.460 30.405 ;
        RECT 25.790 30.175 26.750 30.405 ;
        RECT 19.610 28.130 20.150 29.390 ;
        RECT 23.050 28.970 23.740 29.560 ;
        RECT 24.500 28.970 25.460 28.995 ;
        RECT 21.660 28.800 25.460 28.970 ;
        RECT 21.660 28.520 22.500 28.800 ;
        RECT 24.500 28.765 25.460 28.800 ;
        RECT 25.790 28.765 26.750 28.995 ;
        RECT 22.710 28.560 24.430 28.580 ;
        RECT 20.310 28.290 21.270 28.520 ;
        RECT 21.600 28.290 22.560 28.520 ;
        RECT 19.610 27.130 20.260 28.130 ;
        RECT 19.610 26.600 20.150 27.130 ;
        RECT 20.530 26.970 21.050 28.290 ;
        RECT 21.320 27.130 21.550 28.130 ;
        RECT 21.800 26.970 22.320 28.290 ;
        RECT 22.710 28.130 24.450 28.560 ;
        RECT 22.610 27.130 24.450 28.130 ;
        RECT 20.310 26.740 21.270 26.970 ;
        RECT 21.600 26.740 22.560 26.970 ;
        RECT 19.610 26.480 20.160 26.600 ;
        RECT 22.710 26.560 24.450 27.130 ;
        RECT 22.710 26.540 24.430 26.560 ;
        RECT 19.610 25.340 20.170 26.480 ;
        RECT 23.050 26.130 23.740 26.540 ;
        RECT 24.730 26.355 25.250 28.765 ;
        RECT 25.510 26.560 25.740 28.560 ;
        RECT 26.060 26.355 26.580 28.765 ;
        RECT 26.940 28.560 27.840 30.610 ;
        RECT 26.800 26.560 27.840 28.560 ;
        RECT 23.050 25.510 23.750 26.130 ;
        RECT 24.500 26.125 25.460 26.355 ;
        RECT 25.790 26.125 26.750 26.355 ;
        RECT 19.610 24.045 20.150 25.340 ;
        RECT 23.050 24.885 23.740 25.510 ;
        RECT 24.500 24.885 25.460 24.910 ;
        RECT 21.660 24.715 25.460 24.885 ;
        RECT 21.660 24.435 22.500 24.715 ;
        RECT 24.500 24.680 25.460 24.715 ;
        RECT 25.790 24.680 26.750 24.910 ;
        RECT 22.710 24.475 24.430 24.495 ;
        RECT 20.310 24.205 21.270 24.435 ;
        RECT 21.600 24.205 22.560 24.435 ;
        RECT 19.610 23.045 20.260 24.045 ;
        RECT 19.610 22.515 20.150 23.045 ;
        RECT 20.530 22.885 21.050 24.205 ;
        RECT 21.320 23.045 21.550 24.045 ;
        RECT 21.800 22.885 22.320 24.205 ;
        RECT 22.710 24.045 24.450 24.475 ;
        RECT 22.610 23.045 24.450 24.045 ;
        RECT 20.310 22.655 21.270 22.885 ;
        RECT 21.600 22.655 22.560 22.885 ;
        RECT 19.610 22.395 20.160 22.515 ;
        RECT 22.710 22.475 24.450 23.045 ;
        RECT 22.710 22.455 24.430 22.475 ;
        RECT 19.610 21.255 20.170 22.395 ;
        RECT 23.050 22.045 23.740 22.455 ;
        RECT 24.730 22.270 25.250 24.680 ;
        RECT 25.510 22.475 25.740 24.475 ;
        RECT 26.060 22.270 26.580 24.680 ;
        RECT 26.940 24.475 27.840 26.560 ;
        RECT 26.800 22.475 27.840 24.475 ;
        RECT 23.050 21.425 23.750 22.045 ;
        RECT 24.500 22.040 25.460 22.270 ;
        RECT 25.790 22.040 26.750 22.270 ;
        RECT 19.610 19.920 20.150 21.255 ;
        RECT 23.050 20.760 23.740 21.425 ;
        RECT 24.500 20.760 25.460 20.785 ;
        RECT 21.660 20.590 25.460 20.760 ;
        RECT 21.660 20.310 22.500 20.590 ;
        RECT 24.500 20.555 25.460 20.590 ;
        RECT 25.790 20.555 26.750 20.785 ;
        RECT 22.710 20.350 24.430 20.370 ;
        RECT 20.310 20.080 21.270 20.310 ;
        RECT 21.600 20.080 22.560 20.310 ;
        RECT 19.610 18.920 20.260 19.920 ;
        RECT 19.610 18.390 20.150 18.920 ;
        RECT 20.530 18.760 21.050 20.080 ;
        RECT 21.320 18.920 21.550 19.920 ;
        RECT 21.800 18.760 22.320 20.080 ;
        RECT 22.710 19.920 24.450 20.350 ;
        RECT 22.610 18.920 24.450 19.920 ;
        RECT 20.310 18.530 21.270 18.760 ;
        RECT 21.600 18.530 22.560 18.760 ;
        RECT 19.610 18.270 20.160 18.390 ;
        RECT 22.710 18.350 24.450 18.920 ;
        RECT 22.710 18.330 24.430 18.350 ;
        RECT 19.610 17.130 20.170 18.270 ;
        RECT 23.050 17.920 23.740 18.330 ;
        RECT 24.730 18.145 25.250 20.555 ;
        RECT 25.510 18.350 25.740 20.350 ;
        RECT 26.060 18.145 26.580 20.555 ;
        RECT 26.940 20.350 27.840 22.475 ;
        RECT 26.800 18.350 27.840 20.350 ;
        RECT 23.050 17.300 23.750 17.920 ;
        RECT 24.500 17.915 25.460 18.145 ;
        RECT 25.790 17.915 26.750 18.145 ;
        RECT 19.610 15.365 20.150 17.130 ;
        RECT 23.055 16.985 23.745 17.300 ;
        RECT 23.050 16.495 23.745 16.985 ;
        RECT 23.050 16.205 23.740 16.495 ;
        RECT 24.500 16.205 25.460 16.230 ;
        RECT 21.660 16.035 25.460 16.205 ;
        RECT 21.660 15.755 22.500 16.035 ;
        RECT 24.500 16.000 25.460 16.035 ;
        RECT 25.790 16.000 26.750 16.230 ;
        RECT 22.710 15.795 24.430 15.815 ;
        RECT 20.310 15.525 21.270 15.755 ;
        RECT 21.600 15.525 22.560 15.755 ;
        RECT 19.610 14.365 20.260 15.365 ;
        RECT 19.610 13.835 20.150 14.365 ;
        RECT 20.530 14.205 21.050 15.525 ;
        RECT 21.320 14.365 21.550 15.365 ;
        RECT 21.800 14.205 22.320 15.525 ;
        RECT 22.710 15.365 24.450 15.795 ;
        RECT 22.610 14.365 24.450 15.365 ;
        RECT 20.310 13.975 21.270 14.205 ;
        RECT 21.600 13.975 22.560 14.205 ;
        RECT 19.610 13.715 20.160 13.835 ;
        RECT 22.710 13.795 24.450 14.365 ;
        RECT 22.710 13.775 24.430 13.795 ;
        RECT 19.610 12.575 20.170 13.715 ;
        RECT 22.905 13.275 23.910 13.775 ;
        RECT 24.730 13.590 25.250 16.000 ;
        RECT 25.510 13.795 25.740 15.795 ;
        RECT 26.060 13.590 26.580 16.000 ;
        RECT 26.940 15.795 27.840 18.350 ;
        RECT 26.800 13.795 27.840 15.795 ;
        RECT 24.500 13.360 25.460 13.590 ;
        RECT 25.790 13.360 26.750 13.590 ;
        RECT 22.885 5.970 23.910 13.275 ;
        RECT 26.940 12.965 27.840 13.795 ;
        RECT 26.945 12.785 27.840 12.965 ;
        RECT 26.940 12.575 27.840 12.785 ;
        RECT 31.660 9.285 32.650 44.375 ;
        RECT 31.660 8.295 138.840 9.285 ;
        RECT 134.355 6.625 135.205 8.295 ;
        RECT 22.885 4.945 131.895 5.970 ;
        RECT 134.325 5.775 135.235 6.625 ;
        RECT 156.320 5.965 157.345 5.995 ;
        RECT 130.870 4.020 131.895 4.945 ;
        RECT 137.340 4.940 157.345 5.965 ;
        RECT 137.340 4.020 138.365 4.940 ;
        RECT 156.320 4.910 157.345 4.940 ;
        RECT 130.870 2.995 138.365 4.020 ;
      LAYER via ;
        RECT 23.135 142.325 23.685 143.090 ;
        RECT 27.030 142.310 28.600 143.310 ;
        RECT 32.005 142.470 32.565 143.060 ;
        RECT 19.660 141.360 20.110 141.830 ;
        RECT 20.530 140.530 21.050 141.010 ;
        RECT 19.720 138.910 20.100 139.570 ;
        RECT 26.060 141.330 26.580 141.830 ;
        RECT 26.860 140.540 27.130 140.990 ;
        RECT 28.550 140.540 28.820 140.990 ;
        RECT 29.100 141.330 29.620 141.830 ;
        RECT 19.660 137.360 20.110 137.830 ;
        RECT 20.530 136.530 21.050 137.010 ;
        RECT 34.630 140.530 35.150 141.010 ;
        RECT 35.570 141.360 36.020 141.830 ;
        RECT 36.420 141.695 38.070 143.365 ;
        RECT 35.580 138.930 35.930 139.570 ;
        RECT 26.060 137.330 26.580 137.830 ;
        RECT 26.860 136.540 27.130 136.990 ;
        RECT 28.550 136.480 28.820 136.930 ;
        RECT 29.100 137.270 29.620 137.770 ;
        RECT 19.660 133.260 20.110 133.730 ;
        RECT 20.530 132.430 21.050 132.910 ;
        RECT 34.630 136.470 35.150 136.950 ;
        RECT 35.570 137.300 36.020 137.770 ;
        RECT 26.060 133.230 26.580 133.730 ;
        RECT 26.860 132.440 27.130 132.890 ;
        RECT 28.550 132.420 28.820 132.870 ;
        RECT 29.100 133.210 29.620 133.710 ;
        RECT 19.660 129.210 20.110 129.680 ;
        RECT 20.530 128.380 21.050 128.860 ;
        RECT 34.630 132.410 35.150 132.890 ;
        RECT 35.570 133.240 36.020 133.710 ;
        RECT 26.060 129.180 26.580 129.680 ;
        RECT 26.860 128.390 27.130 128.840 ;
        RECT 28.550 128.360 28.820 128.810 ;
        RECT 29.100 129.150 29.620 129.650 ;
        RECT 19.660 125.160 20.110 125.630 ;
        RECT 20.530 124.330 21.050 124.810 ;
        RECT 34.630 128.350 35.150 128.830 ;
        RECT 35.570 129.180 36.020 129.650 ;
        RECT 26.060 125.130 26.580 125.630 ;
        RECT 26.860 124.340 27.130 124.790 ;
        RECT 28.550 124.300 28.820 124.750 ;
        RECT 29.100 125.090 29.620 125.590 ;
        RECT 19.660 121.110 20.110 121.580 ;
        RECT 20.530 120.280 21.050 120.760 ;
        RECT 34.630 124.290 35.150 124.770 ;
        RECT 35.570 125.120 36.020 125.590 ;
        RECT 26.060 121.080 26.580 121.580 ;
        RECT 26.860 120.290 27.130 120.740 ;
        RECT 28.550 120.240 28.820 120.690 ;
        RECT 29.100 121.030 29.620 121.530 ;
        RECT 19.660 117.060 20.110 117.530 ;
        RECT 20.530 116.230 21.050 116.710 ;
        RECT 34.630 120.230 35.150 120.710 ;
        RECT 35.570 121.060 36.020 121.530 ;
        RECT 26.060 117.030 26.580 117.530 ;
        RECT 26.860 116.240 27.130 116.690 ;
        RECT 28.550 116.180 28.820 116.630 ;
        RECT 29.100 116.970 29.620 117.470 ;
        RECT 19.660 113.010 20.110 113.480 ;
        RECT 20.530 112.180 21.050 112.660 ;
        RECT 34.630 116.170 35.150 116.650 ;
        RECT 35.570 117.000 36.020 117.470 ;
        RECT 26.060 112.980 26.580 113.480 ;
        RECT 26.860 112.190 27.130 112.640 ;
        RECT 28.550 112.120 28.820 112.570 ;
        RECT 29.100 112.910 29.620 113.410 ;
        RECT 19.660 108.960 20.110 109.430 ;
        RECT 20.530 108.130 21.050 108.610 ;
        RECT 34.630 112.110 35.150 112.590 ;
        RECT 35.570 112.940 36.020 113.410 ;
        RECT 26.060 108.930 26.580 109.430 ;
        RECT 26.860 108.140 27.130 108.590 ;
        RECT 28.550 108.060 28.820 108.510 ;
        RECT 29.100 108.850 29.620 109.350 ;
        RECT 19.660 104.910 20.110 105.380 ;
        RECT 20.530 104.080 21.050 104.560 ;
        RECT 34.630 108.050 35.150 108.530 ;
        RECT 35.570 108.880 36.020 109.350 ;
        RECT 26.060 104.880 26.580 105.380 ;
        RECT 26.860 104.090 27.130 104.540 ;
        RECT 28.550 104.000 28.820 104.450 ;
        RECT 29.100 104.790 29.620 105.290 ;
        RECT 19.660 100.860 20.110 101.330 ;
        RECT 20.530 100.030 21.050 100.510 ;
        RECT 34.630 103.990 35.150 104.470 ;
        RECT 35.570 104.820 36.020 105.290 ;
        RECT 26.060 100.830 26.580 101.330 ;
        RECT 26.860 100.040 27.130 100.490 ;
        RECT 28.550 99.940 28.820 100.390 ;
        RECT 29.100 100.730 29.620 101.230 ;
        RECT 19.660 96.810 20.110 97.280 ;
        RECT 20.530 95.980 21.050 96.460 ;
        RECT 34.630 99.930 35.150 100.410 ;
        RECT 35.570 100.760 36.020 101.230 ;
        RECT 26.060 96.780 26.580 97.280 ;
        RECT 26.860 95.990 27.130 96.440 ;
        RECT 28.550 95.880 28.820 96.330 ;
        RECT 29.100 96.670 29.620 97.170 ;
        RECT 19.660 92.760 20.110 93.230 ;
        RECT 20.530 91.930 21.050 92.410 ;
        RECT 34.630 95.870 35.150 96.350 ;
        RECT 35.570 96.700 36.020 97.170 ;
        RECT 26.060 92.730 26.580 93.230 ;
        RECT 26.860 91.940 27.130 92.390 ;
        RECT 28.550 91.820 28.820 92.270 ;
        RECT 29.100 92.610 29.620 93.110 ;
        RECT 19.660 88.710 20.110 89.180 ;
        RECT 20.530 87.880 21.050 88.360 ;
        RECT 34.630 91.810 35.150 92.290 ;
        RECT 35.570 92.640 36.020 93.110 ;
        RECT 26.060 88.680 26.580 89.180 ;
        RECT 26.860 87.890 27.130 88.340 ;
        RECT 28.550 87.760 28.820 88.210 ;
        RECT 29.100 88.550 29.620 89.050 ;
        RECT 19.660 84.660 20.110 85.130 ;
        RECT 20.530 83.830 21.050 84.310 ;
        RECT 34.630 87.750 35.150 88.230 ;
        RECT 35.570 88.580 36.020 89.050 ;
        RECT 26.060 84.630 26.580 85.130 ;
        RECT 26.860 83.840 27.130 84.290 ;
        RECT 28.550 83.700 28.820 84.150 ;
        RECT 29.100 84.490 29.620 84.990 ;
        RECT 19.660 80.610 20.110 81.080 ;
        RECT 20.530 79.780 21.050 80.260 ;
        RECT 34.630 83.690 35.150 84.170 ;
        RECT 35.570 84.520 36.020 84.990 ;
        RECT 26.060 80.580 26.580 81.080 ;
        RECT 26.860 79.790 27.130 80.240 ;
        RECT 28.550 79.640 28.820 80.090 ;
        RECT 29.100 80.430 29.620 80.930 ;
        RECT 19.660 76.560 20.110 77.030 ;
        RECT 20.530 75.730 21.050 76.210 ;
        RECT 34.630 79.630 35.150 80.110 ;
        RECT 35.570 80.460 36.020 80.930 ;
        RECT 26.060 76.530 26.580 77.030 ;
        RECT 26.860 75.740 27.130 76.190 ;
        RECT 28.550 75.580 28.820 76.030 ;
        RECT 29.100 76.370 29.620 76.870 ;
        RECT 19.660 72.510 20.110 72.980 ;
        RECT 20.530 71.680 21.050 72.160 ;
        RECT 34.630 75.570 35.150 76.050 ;
        RECT 35.570 76.400 36.020 76.870 ;
        RECT 26.060 72.480 26.580 72.980 ;
        RECT 26.860 71.690 27.130 72.140 ;
        RECT 28.550 71.520 28.820 71.970 ;
        RECT 29.100 72.310 29.620 72.810 ;
        RECT 19.660 68.460 20.110 68.930 ;
        RECT 20.530 67.630 21.050 68.110 ;
        RECT 34.630 71.510 35.150 71.990 ;
        RECT 35.570 72.340 36.020 72.810 ;
        RECT 26.060 68.430 26.580 68.930 ;
        RECT 26.860 67.640 27.130 68.090 ;
        RECT 28.550 67.460 28.820 67.910 ;
        RECT 29.100 68.250 29.620 68.750 ;
        RECT 19.660 64.410 20.110 64.880 ;
        RECT 20.530 63.580 21.050 64.060 ;
        RECT 34.630 67.450 35.150 67.930 ;
        RECT 35.570 68.280 36.020 68.750 ;
        RECT 26.060 64.380 26.580 64.880 ;
        RECT 26.860 63.590 27.130 64.040 ;
        RECT 28.550 63.400 28.820 63.850 ;
        RECT 29.100 64.190 29.620 64.690 ;
        RECT 19.660 60.360 20.110 60.830 ;
        RECT 20.530 59.530 21.050 60.010 ;
        RECT 34.630 63.390 35.150 63.870 ;
        RECT 35.570 64.220 36.020 64.690 ;
        RECT 26.060 60.330 26.580 60.830 ;
        RECT 26.860 59.540 27.130 59.990 ;
        RECT 28.550 59.340 28.820 59.790 ;
        RECT 29.100 60.130 29.620 60.630 ;
        RECT 34.630 59.330 35.150 59.810 ;
        RECT 35.570 60.160 36.020 60.630 ;
        RECT 19.660 56.310 20.110 56.780 ;
        RECT 20.530 55.480 21.050 55.960 ;
        RECT 31.995 57.760 32.565 58.530 ;
        RECT 26.060 56.280 26.580 56.780 ;
        RECT 26.860 55.490 27.130 55.940 ;
        RECT 28.550 54.800 28.820 55.250 ;
        RECT 29.100 55.590 29.620 56.090 ;
        RECT 34.630 54.790 35.150 55.270 ;
        RECT 35.570 55.620 36.020 56.090 ;
        RECT 19.660 52.260 20.110 52.730 ;
        RECT 20.530 51.430 21.050 51.910 ;
        RECT 26.060 52.230 26.580 52.730 ;
        RECT 26.860 51.440 27.130 51.890 ;
        RECT 19.660 48.210 20.110 48.680 ;
        RECT 20.530 47.380 21.050 47.860 ;
        RECT 26.060 48.180 26.580 48.680 ;
        RECT 26.860 47.390 27.130 47.840 ;
        RECT 19.660 44.160 20.110 44.630 ;
        RECT 20.530 43.330 21.050 43.810 ;
        RECT 26.060 44.130 26.580 44.630 ;
        RECT 26.860 43.340 27.130 43.790 ;
        RECT 19.660 40.110 20.110 40.580 ;
        RECT 20.530 39.280 21.050 39.760 ;
        RECT 26.060 40.080 26.580 40.580 ;
        RECT 26.860 39.290 27.130 39.740 ;
        RECT 19.660 36.060 20.110 36.530 ;
        RECT 20.530 35.230 21.050 35.710 ;
        RECT 26.060 36.030 26.580 36.530 ;
        RECT 26.860 35.240 27.130 35.690 ;
        RECT 19.660 32.010 20.110 32.480 ;
        RECT 20.530 31.180 21.050 31.660 ;
        RECT 26.060 31.980 26.580 32.480 ;
        RECT 26.860 31.190 27.130 31.640 ;
        RECT 19.660 27.960 20.110 28.430 ;
        RECT 20.530 27.130 21.050 27.610 ;
        RECT 26.060 27.930 26.580 28.430 ;
        RECT 26.860 27.140 27.130 27.590 ;
        RECT 19.660 23.875 20.110 24.345 ;
        RECT 20.530 23.045 21.050 23.525 ;
        RECT 26.060 23.845 26.580 24.345 ;
        RECT 26.860 23.055 27.130 23.505 ;
        RECT 19.660 19.750 20.110 20.220 ;
        RECT 20.530 18.920 21.050 19.400 ;
        RECT 23.110 17.420 23.695 18.190 ;
        RECT 26.060 19.720 26.580 20.220 ;
        RECT 26.860 18.930 27.130 19.380 ;
        RECT 19.660 15.195 20.110 15.665 ;
        RECT 20.530 14.365 21.050 14.845 ;
        RECT 26.060 15.165 26.580 15.665 ;
        RECT 26.860 14.375 27.130 14.825 ;
        RECT 134.355 5.775 135.205 6.625 ;
        RECT 156.320 4.940 157.345 5.965 ;
      LAYER met2 ;
        RECT 6.070 145.620 28.725 147.415 ;
        RECT 23.055 142.225 23.755 143.145 ;
        RECT 26.930 142.230 28.725 145.620 ;
        RECT 36.420 143.355 38.070 143.395 ;
        RECT 31.925 142.380 32.625 143.150 ;
        RECT 19.630 141.300 26.620 141.870 ;
        RECT 29.060 141.300 36.050 141.870 ;
        RECT 36.420 141.705 41.840 143.355 ;
        RECT 36.420 141.665 38.070 141.705 ;
        RECT 20.470 140.490 27.170 141.060 ;
        RECT 28.510 140.490 35.210 141.060 ;
        RECT 19.690 138.850 35.990 139.670 ;
        RECT 19.630 137.300 26.620 137.870 ;
        RECT 29.060 137.240 36.050 137.810 ;
        RECT 20.470 136.490 27.170 137.060 ;
        RECT 28.510 136.430 35.210 137.000 ;
        RECT 19.630 133.200 26.620 133.770 ;
        RECT 29.060 133.180 36.050 133.750 ;
        RECT 20.470 132.390 27.170 132.960 ;
        RECT 28.510 132.370 35.210 132.940 ;
        RECT 19.630 129.150 26.620 129.720 ;
        RECT 29.060 129.120 36.050 129.690 ;
        RECT 20.470 128.340 27.170 128.910 ;
        RECT 28.510 128.310 35.210 128.880 ;
        RECT 19.630 125.100 26.620 125.670 ;
        RECT 29.060 125.060 36.050 125.630 ;
        RECT 20.470 124.290 27.170 124.860 ;
        RECT 28.510 124.250 35.210 124.820 ;
        RECT 19.630 121.050 26.620 121.620 ;
        RECT 29.060 121.000 36.050 121.570 ;
        RECT 20.470 120.240 27.170 120.810 ;
        RECT 28.510 120.190 35.210 120.760 ;
        RECT 19.630 117.000 26.620 117.570 ;
        RECT 29.060 116.940 36.050 117.510 ;
        RECT 20.470 116.190 27.170 116.760 ;
        RECT 28.510 116.130 35.210 116.700 ;
        RECT 19.630 112.950 26.620 113.520 ;
        RECT 29.060 112.880 36.050 113.450 ;
        RECT 20.470 112.140 27.170 112.710 ;
        RECT 28.510 112.070 35.210 112.640 ;
        RECT 19.630 108.900 26.620 109.470 ;
        RECT 29.060 108.820 36.050 109.390 ;
        RECT 20.470 108.090 27.170 108.660 ;
        RECT 28.510 108.010 35.210 108.580 ;
        RECT 19.630 104.850 26.620 105.420 ;
        RECT 29.060 104.760 36.050 105.330 ;
        RECT 20.470 104.040 27.170 104.610 ;
        RECT 28.510 103.950 35.210 104.520 ;
        RECT 19.630 100.800 26.620 101.370 ;
        RECT 29.060 100.700 36.050 101.270 ;
        RECT 20.470 99.990 27.170 100.560 ;
        RECT 28.510 99.890 35.210 100.460 ;
        RECT 19.630 96.750 26.620 97.320 ;
        RECT 29.060 96.640 36.050 97.210 ;
        RECT 20.470 95.940 27.170 96.510 ;
        RECT 28.510 95.830 35.210 96.400 ;
        RECT 19.630 92.700 26.620 93.270 ;
        RECT 29.060 92.580 36.050 93.150 ;
        RECT 20.470 91.890 27.170 92.460 ;
        RECT 28.510 91.770 35.210 92.340 ;
        RECT 19.630 88.650 26.620 89.220 ;
        RECT 29.060 88.520 36.050 89.090 ;
        RECT 20.470 87.840 27.170 88.410 ;
        RECT 28.510 87.710 35.210 88.280 ;
        RECT 19.630 84.600 26.620 85.170 ;
        RECT 29.060 84.460 36.050 85.030 ;
        RECT 20.470 83.790 27.170 84.360 ;
        RECT 28.510 83.650 35.210 84.220 ;
        RECT 19.630 80.550 26.620 81.120 ;
        RECT 29.060 80.400 36.050 80.970 ;
        RECT 20.470 79.740 27.170 80.310 ;
        RECT 28.510 79.590 35.210 80.160 ;
        RECT 19.630 76.500 26.620 77.070 ;
        RECT 29.060 76.340 36.050 76.910 ;
        RECT 20.470 75.690 27.170 76.260 ;
        RECT 28.510 75.530 35.210 76.100 ;
        RECT 19.630 72.450 26.620 73.020 ;
        RECT 29.060 72.280 36.050 72.850 ;
        RECT 20.470 71.640 27.170 72.210 ;
        RECT 28.510 71.470 35.210 72.040 ;
        RECT 19.630 68.400 26.620 68.970 ;
        RECT 29.060 68.220 36.050 68.790 ;
        RECT 20.470 67.590 27.170 68.160 ;
        RECT 28.510 67.410 35.210 67.980 ;
        RECT 19.630 64.350 26.620 64.920 ;
        RECT 29.060 64.160 36.050 64.730 ;
        RECT 20.470 63.540 27.170 64.110 ;
        RECT 28.510 63.350 35.210 63.920 ;
        RECT 19.630 60.300 26.620 60.870 ;
        RECT 29.060 60.100 36.050 60.670 ;
        RECT 20.470 59.490 27.170 60.060 ;
        RECT 28.510 59.290 35.210 59.860 ;
        RECT 31.925 57.710 32.625 58.580 ;
        RECT 19.630 56.250 26.620 56.820 ;
        RECT 20.470 55.440 27.170 56.010 ;
        RECT 29.060 55.560 36.050 56.130 ;
        RECT 28.510 54.750 35.210 55.320 ;
        RECT 19.630 52.200 26.620 52.770 ;
        RECT 20.470 51.390 27.170 51.960 ;
        RECT 19.630 48.150 26.620 48.720 ;
        RECT 20.470 47.340 27.170 47.910 ;
        RECT 19.630 44.100 26.620 44.670 ;
        RECT 20.470 43.290 27.170 43.860 ;
        RECT 19.630 40.050 26.620 40.620 ;
        RECT 20.470 39.240 27.170 39.810 ;
        RECT 19.630 36.000 26.620 36.570 ;
        RECT 20.470 35.190 27.170 35.760 ;
        RECT 19.630 31.950 26.620 32.520 ;
        RECT 20.470 31.140 27.170 31.710 ;
        RECT 19.630 27.900 26.620 28.470 ;
        RECT 20.470 27.090 27.170 27.660 ;
        RECT 19.630 23.815 26.620 24.385 ;
        RECT 20.470 23.005 27.170 23.575 ;
        RECT 19.630 19.690 26.620 20.260 ;
        RECT 20.470 18.880 27.170 19.450 ;
        RECT 23.055 17.340 23.755 18.300 ;
        RECT 19.630 15.135 26.620 15.705 ;
        RECT 20.470 14.325 27.170 14.895 ;
        RECT 134.355 5.630 135.205 6.655 ;
        RECT 156.320 5.965 157.345 6.010 ;
        RECT 134.335 4.830 135.225 5.630 ;
        RECT 156.290 4.940 157.375 5.965 ;
        RECT 156.320 4.895 157.345 4.940 ;
        RECT 134.355 4.805 135.205 4.830 ;
      LAYER via2 ;
        RECT 6.115 145.620 7.910 147.415 ;
        RECT 23.135 142.325 23.685 143.090 ;
        RECT 32.005 142.470 32.565 143.060 ;
        RECT 40.145 141.705 41.795 143.355 ;
        RECT 31.995 57.760 32.565 58.530 ;
        RECT 23.110 17.420 23.695 18.190 ;
        RECT 134.380 4.830 135.180 5.630 ;
        RECT 156.320 4.940 157.345 5.965 ;
      LAYER met3 ;
        RECT 6.060 145.595 7.935 147.440 ;
        RECT 40.120 143.355 41.820 143.380 ;
        RECT 23.055 17.305 23.750 143.145 ;
        RECT 31.925 57.710 32.625 143.150 ;
        RECT 40.120 141.705 45.705 143.355 ;
        RECT 40.120 141.680 41.820 141.705 ;
        RECT 134.355 2.610 135.205 5.655 ;
        RECT 156.295 4.915 157.370 5.990 ;
        RECT 156.320 3.350 157.345 4.915 ;
        RECT 134.330 1.770 135.230 2.610 ;
        RECT 134.355 1.765 135.205 1.770 ;
        RECT 156.465 0.325 157.200 3.350 ;
      LAYER via3 ;
        RECT 6.090 145.595 7.885 147.440 ;
        RECT 44.025 141.705 45.675 143.355 ;
        RECT 156.320 3.380 157.345 4.405 ;
        RECT 134.360 1.770 135.200 2.610 ;
      LAYER met4 ;
        RECT 3.990 223.220 4.290 224.760 ;
        RECT 7.670 223.220 7.970 224.760 ;
        RECT 11.350 223.220 11.650 224.760 ;
        RECT 15.030 223.220 15.330 224.760 ;
        RECT 18.710 223.220 19.010 224.760 ;
        RECT 22.390 223.220 22.690 224.760 ;
        RECT 26.070 223.220 26.370 224.760 ;
        RECT 29.750 223.220 30.050 224.760 ;
        RECT 33.430 223.220 33.730 224.760 ;
        RECT 37.110 223.220 37.410 224.760 ;
        RECT 40.790 223.220 41.090 224.760 ;
        RECT 44.470 223.220 44.770 224.760 ;
        RECT 48.150 223.220 48.450 224.760 ;
        RECT 51.830 223.220 52.130 224.760 ;
        RECT 55.510 223.220 55.810 224.760 ;
        RECT 59.190 223.220 59.490 224.760 ;
        RECT 62.870 223.220 63.170 224.760 ;
        RECT 66.550 223.220 66.850 224.760 ;
        RECT 70.230 223.220 70.530 224.760 ;
        RECT 73.910 223.220 74.210 224.760 ;
        RECT 77.590 223.220 77.890 224.760 ;
        RECT 81.270 223.220 81.570 224.760 ;
        RECT 84.950 223.220 85.250 224.760 ;
        RECT 88.630 223.220 88.930 224.760 ;
        RECT 2.970 221.620 89.590 223.220 ;
        RECT 49.000 220.760 50.500 221.620 ;
        RECT 6.085 147.415 7.890 147.445 ;
        RECT 2.500 145.620 7.890 147.415 ;
        RECT 6.085 145.590 7.890 145.620 ;
        RECT 44.020 143.355 45.680 143.360 ;
        RECT 44.020 141.705 49.000 143.355 ;
        RECT 44.020 141.700 45.680 141.705 ;
        RECT 156.315 3.375 157.350 4.410 ;
        RECT 134.355 1.000 135.205 2.615 ;
        RECT 156.535 1.000 157.130 3.375 ;
  END
END tt_um_devinatkin_dual_oscillator
END LIBRARY

