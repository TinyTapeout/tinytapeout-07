VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_devinatkin_dual_oscillator
  CLASS BLOCK ;
  FOREIGN tt_um_devinatkin_dual_oscillator ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 20.000000 ;
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 20.000000 ;
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 84.000000 ;
    ANTENNADIFFAREA 410.998810 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.390 4.940 147.890 220.700 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  OBS
      LAYER pwell ;
        RECT 29.930 192.440 94.510 195.400 ;
        RECT 29.920 190.450 47.880 192.440 ;
        RECT 14.160 121.620 17.950 183.010 ;
        RECT 19.900 152.050 26.950 183.010 ;
      LAYER nwell ;
        RECT 28.440 170.140 45.540 184.010 ;
      LAYER pwell ;
        RECT 61.720 183.760 70.940 184.010 ;
        RECT 45.550 170.140 70.940 183.760 ;
        RECT 71.450 173.830 94.510 192.440 ;
      LAYER nwell ;
        RECT 94.510 178.140 105.760 195.410 ;
      LAYER pwell ;
        RECT 105.760 178.140 113.960 195.410 ;
      LAYER nwell ;
        RECT 122.725 184.375 127.175 189.005 ;
      LAYER pwell ;
        RECT 127.175 184.375 130.955 189.005 ;
      LAYER nwell ;
        RECT 94.510 173.830 106.850 178.140 ;
      LAYER pwell ;
        RECT 71.450 171.370 94.500 173.830 ;
      LAYER nwell ;
        RECT 94.500 171.370 106.850 173.830 ;
      LAYER pwell ;
        RECT 106.850 171.370 113.950 178.140 ;
      LAYER nwell ;
        RECT 122.725 176.275 127.175 180.905 ;
      LAYER pwell ;
        RECT 127.175 176.275 130.955 180.905 ;
        RECT 71.450 171.360 104.730 171.370 ;
        RECT 28.440 170.130 61.720 170.140 ;
        RECT 28.440 167.670 51.490 170.130 ;
      LAYER nwell ;
        RECT 51.490 167.670 63.840 170.130 ;
      LAYER pwell ;
        RECT 28.440 146.100 51.500 167.670 ;
      LAYER nwell ;
        RECT 51.500 163.360 63.840 167.670 ;
      LAYER pwell ;
        RECT 63.840 163.360 70.940 170.130 ;
      LAYER nwell ;
        RECT 51.500 146.090 62.750 163.360 ;
      LAYER pwell ;
        RECT 62.750 146.090 70.950 163.360 ;
      LAYER nwell ;
        RECT 71.450 142.860 88.550 171.360 ;
      LAYER pwell ;
        RECT 88.560 157.740 113.950 171.360 ;
      LAYER nwell ;
        RECT 122.725 168.175 127.175 172.805 ;
      LAYER pwell ;
        RECT 127.175 168.175 130.955 172.805 ;
      LAYER nwell ;
        RECT 122.725 163.580 127.175 164.705 ;
      LAYER pwell ;
        RECT 104.730 157.490 113.950 157.740 ;
        RECT 104.730 156.480 113.950 156.730 ;
        RECT 88.560 142.860 113.950 156.480 ;
        RECT 71.450 142.850 104.730 142.860 ;
        RECT 71.450 140.390 94.500 142.850 ;
      LAYER nwell ;
        RECT 94.500 140.390 106.850 142.850 ;
      LAYER pwell ;
        RECT 14.170 44.220 17.960 105.610 ;
        RECT 71.450 96.920 94.510 140.390 ;
      LAYER nwell ;
        RECT 94.510 136.080 106.850 140.390 ;
      LAYER pwell ;
        RECT 106.850 136.080 113.950 142.850 ;
        RECT 114.545 138.170 118.325 163.580 ;
      LAYER nwell ;
        RECT 118.325 160.075 127.175 163.580 ;
      LAYER pwell ;
        RECT 127.175 160.075 130.955 164.705 ;
      LAYER nwell ;
        RECT 118.325 156.605 122.775 160.075 ;
        RECT 118.325 151.975 127.175 156.605 ;
      LAYER pwell ;
        RECT 127.175 151.975 130.955 156.605 ;
      LAYER nwell ;
        RECT 118.325 148.505 122.775 151.975 ;
        RECT 118.325 143.875 127.175 148.505 ;
      LAYER pwell ;
        RECT 127.175 143.875 130.955 148.505 ;
      LAYER nwell ;
        RECT 118.325 140.405 122.775 143.875 ;
        RECT 118.325 138.170 127.175 140.405 ;
        RECT 94.510 101.230 105.760 136.080 ;
      LAYER pwell ;
        RECT 105.760 118.810 113.960 136.080 ;
      LAYER nwell ;
        RECT 121.380 135.775 127.175 138.170 ;
      LAYER pwell ;
        RECT 127.175 135.775 130.955 140.405 ;
      LAYER nwell ;
        RECT 121.380 134.680 122.780 135.775 ;
      LAYER pwell ;
        RECT 105.760 101.230 113.960 118.500 ;
      LAYER nwell ;
        RECT 94.510 96.920 106.850 101.230 ;
      LAYER pwell ;
        RECT 71.450 94.460 94.500 96.920 ;
      LAYER nwell ;
        RECT 94.500 94.460 106.850 96.920 ;
      LAYER pwell ;
        RECT 106.850 94.460 113.950 101.230 ;
        RECT 114.545 97.570 118.325 134.680 ;
      LAYER nwell ;
        RECT 118.325 134.590 122.780 134.680 ;
        RECT 118.325 132.305 122.775 134.590 ;
        RECT 118.325 127.675 127.175 132.305 ;
      LAYER pwell ;
        RECT 127.175 127.675 130.955 132.305 ;
      LAYER nwell ;
        RECT 118.325 124.205 122.775 127.675 ;
        RECT 118.325 119.575 127.175 124.205 ;
      LAYER pwell ;
        RECT 127.175 119.575 130.955 124.205 ;
      LAYER nwell ;
        RECT 118.325 116.105 122.775 119.575 ;
        RECT 118.325 111.475 127.175 116.105 ;
      LAYER pwell ;
        RECT 127.175 111.475 130.955 116.105 ;
      LAYER nwell ;
        RECT 118.325 108.005 122.775 111.475 ;
        RECT 118.325 97.570 127.175 108.005 ;
      LAYER pwell ;
        RECT 71.450 94.450 104.730 94.460 ;
        RECT 19.910 44.220 26.960 75.180 ;
        RECT 28.450 59.560 51.510 81.130 ;
      LAYER nwell ;
        RECT 51.510 63.870 62.760 81.140 ;
      LAYER pwell ;
        RECT 62.760 63.870 70.960 81.140 ;
      LAYER nwell ;
        RECT 71.450 67.260 88.550 94.450 ;
      LAYER pwell ;
        RECT 88.560 67.260 113.950 94.450 ;
      LAYER nwell ;
        RECT 122.725 94.080 127.175 97.570 ;
      LAYER pwell ;
        RECT 114.545 73.210 118.325 94.080 ;
      LAYER nwell ;
        RECT 118.325 73.210 127.175 94.080 ;
      LAYER pwell ;
        RECT 71.450 67.250 104.730 67.260 ;
        RECT 71.450 64.790 94.500 67.250 ;
      LAYER nwell ;
        RECT 94.500 64.790 106.850 67.250 ;
        RECT 51.510 59.560 63.850 63.870 ;
      LAYER pwell ;
        RECT 28.450 57.100 51.500 59.560 ;
      LAYER nwell ;
        RECT 51.500 57.100 63.850 59.560 ;
      LAYER pwell ;
        RECT 63.850 57.100 70.950 63.870 ;
        RECT 28.450 57.090 61.730 57.100 ;
      LAYER nwell ;
        RECT 28.450 43.220 45.550 57.090 ;
      LAYER pwell ;
        RECT 45.560 43.470 70.950 57.090 ;
        RECT 61.730 43.220 70.950 43.470 ;
        RECT 71.450 43.220 94.510 64.790 ;
      LAYER nwell ;
        RECT 94.510 60.480 106.850 64.790 ;
      LAYER pwell ;
        RECT 106.850 60.480 113.950 67.250 ;
      LAYER nwell ;
        RECT 94.510 43.210 105.760 60.480 ;
      LAYER pwell ;
        RECT 105.760 43.210 113.960 60.480 ;
      LAYER nwell ;
        RECT 122.725 58.210 127.175 73.210 ;
      LAYER pwell ;
        RECT 127.175 58.210 130.955 108.005 ;
      LAYER li1 ;
        RECT 30.110 195.050 71.850 195.220 ;
        RECT 30.110 192.790 30.280 195.050 ;
        RECT 30.960 194.480 71.000 194.650 ;
        RECT 30.620 193.420 30.790 194.420 ;
        RECT 71.170 193.420 71.340 194.420 ;
        RECT 30.960 193.190 71.000 193.360 ;
        RECT 71.680 192.790 71.850 195.050 ;
        RECT 30.110 192.620 71.850 192.790 ;
        RECT 106.350 194.910 113.660 195.090 ;
        RECT 30.100 192.090 47.700 192.260 ;
        RECT 30.100 191.870 30.270 192.090 ;
        RECT 30.100 191.180 30.280 191.870 ;
        RECT 30.830 191.530 31.000 191.610 ;
        RECT 46.800 191.530 46.970 191.610 ;
        RECT 30.830 191.360 32.815 191.530 ;
        RECT 44.985 191.360 46.970 191.530 ;
        RECT 30.830 191.280 31.000 191.360 ;
        RECT 46.800 191.280 46.970 191.360 ;
        RECT 30.100 190.800 30.270 191.180 ;
        RECT 47.530 190.800 47.700 192.090 ;
        RECT 30.100 190.630 47.700 190.800 ;
        RECT 98.770 191.530 105.540 191.700 ;
        RECT 29.090 183.410 45.200 183.590 ;
        RECT 14.340 182.660 17.770 182.830 ;
        RECT 14.340 152.400 14.510 182.660 ;
        RECT 14.990 181.930 15.490 182.100 ;
        RECT 15.070 180.115 15.410 181.930 ;
        RECT 15.070 153.130 15.410 154.945 ;
        RECT 14.990 152.960 15.490 153.130 ;
        RECT 15.970 152.400 16.140 182.660 ;
        RECT 16.620 181.930 17.120 182.100 ;
        RECT 16.700 180.115 17.040 181.930 ;
        RECT 16.700 153.130 17.040 154.945 ;
        RECT 16.620 152.960 17.120 153.130 ;
        RECT 17.600 152.400 17.770 182.660 ;
        RECT 14.340 152.230 17.770 152.400 ;
        RECT 20.080 182.660 26.770 182.830 ;
        RECT 20.080 152.400 20.250 182.660 ;
        RECT 20.730 181.930 21.230 182.100 ;
        RECT 20.810 180.115 21.150 181.930 ;
        RECT 20.810 153.130 21.150 154.945 ;
        RECT 20.730 152.960 21.230 153.130 ;
        RECT 21.710 152.400 21.880 182.660 ;
        RECT 22.360 181.930 22.860 182.100 ;
        RECT 22.440 180.115 22.780 181.930 ;
        RECT 22.440 153.130 22.780 154.945 ;
        RECT 22.360 152.960 22.860 153.130 ;
        RECT 23.340 152.400 23.510 182.660 ;
        RECT 23.990 181.930 24.490 182.100 ;
        RECT 24.070 180.115 24.410 181.930 ;
        RECT 24.070 153.130 24.410 154.945 ;
        RECT 23.990 152.960 24.490 153.130 ;
        RECT 24.970 152.400 25.140 182.660 ;
        RECT 25.620 181.930 26.120 182.100 ;
        RECT 25.700 180.115 26.040 181.930 ;
        RECT 25.700 153.130 26.040 154.945 ;
        RECT 25.620 152.960 26.120 153.130 ;
        RECT 26.600 152.400 26.770 182.660 ;
        RECT 29.090 170.750 29.270 183.410 ;
        RECT 30.020 182.600 35.060 182.770 ;
        RECT 39.020 182.600 44.060 182.770 ;
        RECT 29.635 182.040 29.805 182.540 ;
        RECT 35.275 182.040 35.445 182.540 ;
        RECT 38.635 182.040 38.805 182.540 ;
        RECT 44.275 182.040 44.445 182.540 ;
        RECT 30.020 181.810 35.060 181.980 ;
        RECT 39.020 181.810 44.060 181.980 ;
        RECT 30.020 178.100 35.060 178.270 ;
        RECT 39.020 178.100 44.060 178.270 ;
        RECT 29.635 177.540 29.805 178.040 ;
        RECT 35.275 177.540 35.445 178.040 ;
        RECT 38.635 177.540 38.805 178.040 ;
        RECT 44.275 177.540 44.445 178.040 ;
        RECT 30.020 177.310 35.060 177.480 ;
        RECT 39.020 177.310 44.060 177.480 ;
        RECT 30.020 173.600 35.060 173.770 ;
        RECT 39.020 173.600 44.060 173.770 ;
        RECT 29.635 173.040 29.805 173.540 ;
        RECT 35.275 173.040 35.445 173.540 ;
        RECT 38.635 173.040 38.805 173.540 ;
        RECT 44.275 173.040 44.445 173.540 ;
        RECT 30.020 172.810 35.060 172.980 ;
        RECT 39.020 172.810 44.060 172.980 ;
        RECT 45.020 170.750 45.200 183.410 ;
        RECT 29.090 170.570 45.200 170.750 ;
        RECT 45.860 183.240 61.420 183.410 ;
        RECT 45.860 170.720 46.030 183.240 ;
        RECT 47.740 181.620 52.780 181.790 ;
        RECT 54.740 181.620 59.780 181.790 ;
        RECT 47.400 180.560 47.570 181.560 ;
        RECT 52.950 180.560 53.120 181.560 ;
        RECT 54.400 180.560 54.570 181.560 ;
        RECT 59.950 180.560 60.120 181.560 ;
        RECT 47.740 180.330 52.780 180.500 ;
        RECT 54.740 180.330 59.780 180.500 ;
        RECT 47.740 179.620 52.780 179.790 ;
        RECT 54.740 179.620 59.780 179.790 ;
        RECT 47.400 178.560 47.570 179.560 ;
        RECT 52.950 178.560 53.120 179.560 ;
        RECT 54.400 178.560 54.570 179.560 ;
        RECT 59.950 178.560 60.120 179.560 ;
        RECT 47.740 178.330 52.780 178.500 ;
        RECT 54.740 178.330 59.780 178.500 ;
        RECT 47.740 175.620 52.780 175.790 ;
        RECT 54.740 175.620 59.780 175.790 ;
        RECT 47.400 174.560 47.570 175.560 ;
        RECT 52.950 174.560 53.120 175.560 ;
        RECT 54.400 174.560 54.570 175.560 ;
        RECT 59.950 174.560 60.120 175.560 ;
        RECT 47.740 174.330 52.780 174.500 ;
        RECT 54.740 174.330 59.780 174.500 ;
        RECT 47.740 173.620 52.780 173.790 ;
        RECT 54.740 173.620 59.780 173.790 ;
        RECT 47.400 172.560 47.570 173.560 ;
        RECT 52.950 172.560 53.120 173.560 ;
        RECT 54.400 172.560 54.570 173.560 ;
        RECT 59.950 172.560 60.120 173.560 ;
        RECT 47.740 172.330 52.780 172.500 ;
        RECT 54.740 172.330 59.780 172.500 ;
        RECT 61.250 170.720 61.420 183.240 ;
        RECT 45.860 170.550 61.420 170.720 ;
        RECT 62.280 183.380 70.680 183.550 ;
        RECT 62.280 170.580 62.450 183.380 ;
        RECT 63.200 181.340 68.240 181.510 ;
        RECT 62.860 180.280 63.030 181.280 ;
        RECT 68.410 180.280 68.580 181.280 ;
        RECT 63.200 180.050 68.240 180.220 ;
        RECT 62.860 178.990 63.030 179.990 ;
        RECT 68.410 178.990 68.580 179.990 ;
        RECT 63.200 178.760 68.240 178.930 ;
        RECT 62.860 177.700 63.030 178.700 ;
        RECT 68.410 177.700 68.580 178.700 ;
        RECT 63.200 177.470 68.240 177.640 ;
        RECT 62.860 176.410 63.030 177.410 ;
        RECT 68.410 176.410 68.580 177.410 ;
        RECT 63.200 176.180 68.240 176.350 ;
        RECT 62.860 175.120 63.030 176.120 ;
        RECT 68.410 175.120 68.580 176.120 ;
        RECT 63.200 174.890 68.240 175.060 ;
        RECT 62.860 173.830 63.030 174.830 ;
        RECT 68.410 173.830 68.580 174.830 ;
        RECT 63.200 173.600 68.240 173.770 ;
        RECT 62.860 172.540 63.030 173.540 ;
        RECT 68.410 172.540 68.580 173.540 ;
        RECT 63.200 172.310 68.240 172.480 ;
        RECT 62.860 171.250 63.030 172.250 ;
        RECT 68.410 171.250 68.580 172.250 ;
        RECT 63.200 171.020 68.240 171.190 ;
        RECT 70.510 170.580 70.680 183.380 ;
        RECT 98.770 178.770 98.940 191.530 ;
        RECT 99.620 190.580 104.660 190.750 ;
        RECT 99.235 190.020 99.405 190.520 ;
        RECT 104.875 190.020 105.045 190.520 ;
        RECT 99.620 189.790 104.660 189.960 ;
        RECT 99.235 189.230 99.405 189.730 ;
        RECT 104.875 189.230 105.045 189.730 ;
        RECT 99.620 189.000 104.660 189.170 ;
        RECT 99.235 188.440 99.405 188.940 ;
        RECT 104.875 188.440 105.045 188.940 ;
        RECT 99.620 188.210 104.660 188.380 ;
        RECT 99.235 187.650 99.405 188.150 ;
        RECT 104.875 187.650 105.045 188.150 ;
        RECT 99.620 187.420 104.660 187.590 ;
        RECT 99.235 186.860 99.405 187.360 ;
        RECT 104.875 186.860 105.045 187.360 ;
        RECT 99.620 186.630 104.660 186.800 ;
        RECT 99.235 186.070 99.405 186.570 ;
        RECT 104.875 186.070 105.045 186.570 ;
        RECT 99.620 185.840 104.660 186.010 ;
        RECT 99.235 185.280 99.405 185.780 ;
        RECT 104.875 185.280 105.045 185.780 ;
        RECT 99.620 185.050 104.660 185.220 ;
        RECT 99.235 184.490 99.405 184.990 ;
        RECT 104.875 184.490 105.045 184.990 ;
        RECT 99.620 184.260 104.660 184.430 ;
        RECT 99.235 183.700 99.405 184.200 ;
        RECT 104.875 183.700 105.045 184.200 ;
        RECT 99.620 183.470 104.660 183.640 ;
        RECT 99.235 182.910 99.405 183.410 ;
        RECT 104.875 182.910 105.045 183.410 ;
        RECT 99.620 182.680 104.660 182.850 ;
        RECT 99.235 182.120 99.405 182.620 ;
        RECT 104.875 182.120 105.045 182.620 ;
        RECT 99.620 181.890 104.660 182.060 ;
        RECT 99.235 181.330 99.405 181.830 ;
        RECT 104.875 181.330 105.045 181.830 ;
        RECT 99.620 181.100 104.660 181.270 ;
        RECT 99.235 180.540 99.405 181.040 ;
        RECT 104.875 180.540 105.045 181.040 ;
        RECT 99.620 180.310 104.660 180.480 ;
        RECT 99.235 179.750 99.405 180.250 ;
        RECT 104.875 179.750 105.045 180.250 ;
        RECT 99.620 179.520 104.660 179.690 ;
        RECT 105.370 178.770 105.540 191.530 ;
        RECT 98.770 178.600 105.540 178.770 ;
        RECT 106.350 178.780 106.520 194.910 ;
        RECT 107.680 194.350 112.720 194.520 ;
        RECT 107.340 193.790 107.510 194.290 ;
        RECT 112.890 193.790 113.060 194.290 ;
        RECT 107.680 193.560 112.720 193.730 ;
        RECT 107.340 193.000 107.510 193.500 ;
        RECT 112.890 193.000 113.060 193.500 ;
        RECT 107.680 192.770 112.720 192.940 ;
        RECT 107.340 192.210 107.510 192.710 ;
        RECT 112.890 192.210 113.060 192.710 ;
        RECT 107.680 191.980 112.720 192.150 ;
        RECT 107.340 191.420 107.510 191.920 ;
        RECT 112.890 191.420 113.060 191.920 ;
        RECT 107.680 191.190 112.720 191.360 ;
        RECT 107.340 190.630 107.510 191.130 ;
        RECT 112.890 190.630 113.060 191.130 ;
        RECT 107.680 190.400 112.720 190.570 ;
        RECT 107.340 189.840 107.510 190.340 ;
        RECT 112.890 189.840 113.060 190.340 ;
        RECT 107.680 189.610 112.720 189.780 ;
        RECT 107.340 189.050 107.510 189.550 ;
        RECT 112.890 189.050 113.060 189.550 ;
        RECT 107.680 188.820 112.720 188.990 ;
        RECT 107.340 188.260 107.510 188.760 ;
        RECT 112.890 188.260 113.060 188.760 ;
        RECT 107.680 188.030 112.720 188.200 ;
        RECT 107.340 187.470 107.510 187.970 ;
        RECT 112.890 187.470 113.060 187.970 ;
        RECT 107.680 187.240 112.720 187.410 ;
        RECT 107.340 186.680 107.510 187.180 ;
        RECT 112.890 186.680 113.060 187.180 ;
        RECT 107.680 186.450 112.720 186.620 ;
        RECT 107.340 185.890 107.510 186.390 ;
        RECT 112.890 185.890 113.060 186.390 ;
        RECT 107.680 185.660 112.720 185.830 ;
        RECT 107.340 185.100 107.510 185.600 ;
        RECT 112.890 185.100 113.060 185.600 ;
        RECT 107.680 184.870 112.720 185.040 ;
        RECT 107.340 184.310 107.510 184.810 ;
        RECT 112.890 184.310 113.060 184.810 ;
        RECT 107.680 184.080 112.720 184.250 ;
        RECT 107.340 183.520 107.510 184.020 ;
        RECT 112.890 183.520 113.060 184.020 ;
        RECT 107.680 183.290 112.720 183.460 ;
        RECT 107.340 182.730 107.510 183.230 ;
        RECT 112.890 182.730 113.060 183.230 ;
        RECT 107.680 182.500 112.720 182.670 ;
        RECT 107.340 181.940 107.510 182.440 ;
        RECT 112.890 181.940 113.060 182.440 ;
        RECT 107.680 181.710 112.720 181.880 ;
        RECT 107.340 181.150 107.510 181.650 ;
        RECT 112.890 181.150 113.060 181.650 ;
        RECT 107.680 180.920 112.720 181.090 ;
        RECT 107.340 180.360 107.510 180.860 ;
        RECT 112.890 180.360 113.060 180.860 ;
        RECT 107.680 180.130 112.720 180.300 ;
        RECT 107.340 179.570 107.510 180.070 ;
        RECT 112.890 179.570 113.060 180.070 ;
        RECT 107.680 179.340 112.720 179.510 ;
        RECT 113.490 178.780 113.660 194.910 ;
        RECT 126.085 188.825 126.885 188.835 ;
        RECT 122.895 188.655 126.995 188.825 ;
        RECT 122.895 184.765 123.075 188.655 ;
        RECT 123.795 187.830 124.795 188.000 ;
        RECT 125.085 187.830 126.085 188.000 ;
        RECT 123.565 185.575 123.735 187.615 ;
        RECT 124.855 185.575 125.025 187.615 ;
        RECT 126.145 185.575 126.315 187.615 ;
        RECT 123.795 185.190 124.795 185.360 ;
        RECT 125.085 185.190 126.085 185.360 ;
        RECT 126.825 184.765 126.995 188.655 ;
        RECT 122.895 184.555 126.995 184.765 ;
        RECT 127.345 188.655 130.845 188.825 ;
        RECT 127.345 188.645 130.855 188.655 ;
        RECT 127.345 184.765 127.515 188.645 ;
        RECT 130.675 187.545 130.855 188.645 ;
        RECT 127.985 187.355 128.985 187.525 ;
        RECT 129.275 187.355 130.275 187.525 ;
        RECT 127.755 186.145 127.925 187.185 ;
        RECT 129.045 186.145 129.215 187.185 ;
        RECT 130.335 186.145 130.505 187.185 ;
        RECT 127.985 185.805 128.985 185.975 ;
        RECT 129.275 185.805 130.275 185.975 ;
        RECT 130.675 184.765 130.845 187.545 ;
        RECT 127.345 184.555 130.845 184.765 ;
        RECT 126.085 180.725 126.885 180.735 ;
        RECT 106.350 178.600 113.660 178.780 ;
        RECT 122.895 180.555 126.995 180.725 ;
        RECT 95.175 177.785 104.005 177.955 ;
        RECT 95.175 177.470 95.345 177.785 ;
        RECT 95.175 176.330 95.350 177.470 ;
        RECT 96.070 177.215 103.110 177.385 ;
        RECT 95.685 176.655 95.855 177.155 ;
        RECT 103.325 176.655 103.495 177.155 ;
        RECT 96.070 176.425 103.110 176.595 ;
        RECT 95.175 176.025 95.345 176.330 ;
        RECT 103.835 176.025 104.005 177.785 ;
        RECT 122.895 176.665 123.075 180.555 ;
        RECT 123.795 179.730 124.795 179.900 ;
        RECT 125.085 179.730 126.085 179.900 ;
        RECT 123.565 177.475 123.735 179.515 ;
        RECT 124.855 177.475 125.025 179.515 ;
        RECT 126.145 177.475 126.315 179.515 ;
        RECT 123.795 177.090 124.795 177.260 ;
        RECT 125.085 177.090 126.085 177.260 ;
        RECT 126.825 176.665 126.995 180.555 ;
        RECT 122.895 176.455 126.995 176.665 ;
        RECT 127.345 180.555 130.845 180.725 ;
        RECT 127.345 180.545 130.855 180.555 ;
        RECT 127.345 176.665 127.515 180.545 ;
        RECT 130.675 179.445 130.855 180.545 ;
        RECT 127.985 179.255 128.985 179.425 ;
        RECT 129.275 179.255 130.275 179.425 ;
        RECT 127.755 178.045 127.925 179.085 ;
        RECT 129.045 178.045 129.215 179.085 ;
        RECT 130.335 178.045 130.505 179.085 ;
        RECT 127.985 177.705 128.985 177.875 ;
        RECT 129.275 177.705 130.275 177.875 ;
        RECT 130.675 176.665 130.845 179.445 ;
        RECT 127.345 176.455 130.845 176.665 ;
        RECT 95.175 175.855 104.005 176.025 ;
        RECT 95.175 175.540 95.345 175.855 ;
        RECT 95.175 174.400 95.350 175.540 ;
        RECT 96.070 175.285 103.110 175.455 ;
        RECT 95.685 174.725 95.855 175.225 ;
        RECT 103.325 174.725 103.495 175.225 ;
        RECT 96.070 174.495 103.110 174.665 ;
        RECT 95.175 174.095 95.345 174.400 ;
        RECT 103.835 174.095 104.005 175.855 ;
        RECT 95.175 173.925 104.005 174.095 ;
        RECT 107.030 173.985 113.770 174.155 ;
        RECT 97.830 173.920 102.780 173.925 ;
        RECT 94.680 173.480 106.670 173.650 ;
        RECT 94.680 171.720 94.850 173.480 ;
        RECT 95.575 172.910 103.115 173.080 ;
        RECT 95.190 172.350 95.360 172.850 ;
        RECT 103.330 172.350 103.500 172.850 ;
        RECT 95.575 172.120 103.115 172.290 ;
        RECT 103.840 171.720 104.010 173.480 ;
        RECT 104.735 172.910 105.775 173.080 ;
        RECT 104.350 172.350 104.520 172.850 ;
        RECT 105.990 172.350 106.160 172.850 ;
        RECT 104.735 172.120 105.775 172.290 ;
        RECT 106.500 171.720 106.670 173.480 ;
        RECT 94.680 171.550 106.670 171.720 ;
        RECT 107.030 171.725 107.200 173.985 ;
        RECT 107.880 173.415 112.920 173.585 ;
        RECT 107.540 172.355 107.710 173.355 ;
        RECT 113.090 172.355 113.260 173.355 ;
        RECT 107.880 172.125 112.920 172.295 ;
        RECT 113.600 171.725 113.770 173.985 ;
        RECT 126.085 172.625 126.885 172.635 ;
        RECT 107.030 171.555 113.770 171.725 ;
        RECT 122.895 172.455 126.995 172.625 ;
        RECT 108.420 171.550 109.060 171.555 ;
        RECT 109.600 171.550 110.240 171.555 ;
        RECT 111.000 171.550 111.640 171.555 ;
        RECT 112.650 171.550 113.290 171.555 ;
        RECT 62.280 170.410 70.680 170.580 ;
        RECT 72.100 170.750 88.210 170.930 ;
        RECT 51.670 169.780 63.660 169.950 ;
        RECT 65.410 169.945 66.050 169.950 ;
        RECT 66.590 169.945 67.230 169.950 ;
        RECT 67.990 169.945 68.630 169.950 ;
        RECT 69.640 169.945 70.280 169.950 ;
        RECT 51.670 168.020 51.840 169.780 ;
        RECT 52.565 169.210 60.105 169.380 ;
        RECT 52.180 168.650 52.350 169.150 ;
        RECT 60.320 168.650 60.490 169.150 ;
        RECT 52.565 168.420 60.105 168.590 ;
        RECT 60.830 168.020 61.000 169.780 ;
        RECT 61.725 169.210 62.765 169.380 ;
        RECT 61.340 168.650 61.510 169.150 ;
        RECT 62.980 168.650 63.150 169.150 ;
        RECT 61.725 168.420 62.765 168.590 ;
        RECT 63.490 168.020 63.660 169.780 ;
        RECT 51.670 167.850 63.660 168.020 ;
        RECT 64.020 169.775 70.760 169.945 ;
        RECT 54.820 167.575 59.770 167.580 ;
        RECT 52.165 167.405 60.995 167.575 ;
        RECT 52.165 167.100 52.335 167.405 ;
        RECT 52.165 165.960 52.340 167.100 ;
        RECT 53.060 166.835 60.100 167.005 ;
        RECT 52.675 166.275 52.845 166.775 ;
        RECT 60.315 166.275 60.485 166.775 ;
        RECT 53.060 166.045 60.100 166.215 ;
        RECT 52.165 165.645 52.335 165.960 ;
        RECT 60.825 165.645 60.995 167.405 ;
        RECT 64.020 167.515 64.190 169.775 ;
        RECT 64.870 169.205 69.910 169.375 ;
        RECT 64.530 168.145 64.700 169.145 ;
        RECT 70.080 168.145 70.250 169.145 ;
        RECT 64.870 167.915 69.910 168.085 ;
        RECT 70.590 167.515 70.760 169.775 ;
        RECT 64.020 167.345 70.760 167.515 ;
        RECT 52.165 165.475 60.995 165.645 ;
        RECT 52.165 165.170 52.335 165.475 ;
        RECT 52.165 164.030 52.340 165.170 ;
        RECT 53.060 164.905 60.100 165.075 ;
        RECT 52.675 164.345 52.845 164.845 ;
        RECT 60.315 164.345 60.485 164.845 ;
        RECT 53.060 164.115 60.100 164.285 ;
        RECT 52.165 163.715 52.335 164.030 ;
        RECT 60.825 163.715 60.995 165.475 ;
        RECT 52.165 163.545 60.995 163.715 ;
        RECT 20.080 152.230 26.770 152.400 ;
        RECT 55.760 162.730 62.530 162.900 ;
        RECT 14.340 121.970 14.510 152.230 ;
        RECT 14.990 151.500 15.490 151.670 ;
        RECT 15.070 149.685 15.410 151.500 ;
        RECT 15.070 122.700 15.410 124.515 ;
        RECT 14.990 122.530 15.490 122.700 ;
        RECT 15.970 121.970 16.140 152.230 ;
        RECT 16.620 151.500 17.120 151.670 ;
        RECT 16.700 149.685 17.040 151.500 ;
        RECT 16.700 122.700 17.040 124.515 ;
        RECT 16.620 122.530 17.120 122.700 ;
        RECT 17.600 121.970 17.770 152.230 ;
        RECT 55.760 149.970 55.930 162.730 ;
        RECT 56.610 161.810 61.650 161.980 ;
        RECT 56.225 161.250 56.395 161.750 ;
        RECT 61.865 161.250 62.035 161.750 ;
        RECT 56.610 161.020 61.650 161.190 ;
        RECT 56.225 160.460 56.395 160.960 ;
        RECT 61.865 160.460 62.035 160.960 ;
        RECT 56.610 160.230 61.650 160.400 ;
        RECT 56.225 159.670 56.395 160.170 ;
        RECT 61.865 159.670 62.035 160.170 ;
        RECT 56.610 159.440 61.650 159.610 ;
        RECT 56.225 158.880 56.395 159.380 ;
        RECT 61.865 158.880 62.035 159.380 ;
        RECT 56.610 158.650 61.650 158.820 ;
        RECT 56.225 158.090 56.395 158.590 ;
        RECT 61.865 158.090 62.035 158.590 ;
        RECT 56.610 157.860 61.650 158.030 ;
        RECT 56.225 157.300 56.395 157.800 ;
        RECT 61.865 157.300 62.035 157.800 ;
        RECT 56.610 157.070 61.650 157.240 ;
        RECT 56.225 156.510 56.395 157.010 ;
        RECT 61.865 156.510 62.035 157.010 ;
        RECT 56.610 156.280 61.650 156.450 ;
        RECT 56.225 155.720 56.395 156.220 ;
        RECT 61.865 155.720 62.035 156.220 ;
        RECT 56.610 155.490 61.650 155.660 ;
        RECT 56.225 154.930 56.395 155.430 ;
        RECT 61.865 154.930 62.035 155.430 ;
        RECT 56.610 154.700 61.650 154.870 ;
        RECT 56.225 154.140 56.395 154.640 ;
        RECT 61.865 154.140 62.035 154.640 ;
        RECT 56.610 153.910 61.650 154.080 ;
        RECT 56.225 153.350 56.395 153.850 ;
        RECT 61.865 153.350 62.035 153.850 ;
        RECT 56.610 153.120 61.650 153.290 ;
        RECT 56.225 152.560 56.395 153.060 ;
        RECT 61.865 152.560 62.035 153.060 ;
        RECT 56.610 152.330 61.650 152.500 ;
        RECT 56.225 151.770 56.395 152.270 ;
        RECT 61.865 151.770 62.035 152.270 ;
        RECT 56.610 151.540 61.650 151.710 ;
        RECT 56.225 150.980 56.395 151.480 ;
        RECT 61.865 150.980 62.035 151.480 ;
        RECT 56.610 150.750 61.650 150.920 ;
        RECT 62.360 149.970 62.530 162.730 ;
        RECT 55.760 149.800 62.530 149.970 ;
        RECT 63.340 162.720 70.650 162.900 ;
        RECT 63.340 146.590 63.510 162.720 ;
        RECT 64.670 161.990 69.710 162.160 ;
        RECT 64.330 161.430 64.500 161.930 ;
        RECT 69.880 161.430 70.050 161.930 ;
        RECT 64.670 161.200 69.710 161.370 ;
        RECT 64.330 160.640 64.500 161.140 ;
        RECT 69.880 160.640 70.050 161.140 ;
        RECT 64.670 160.410 69.710 160.580 ;
        RECT 64.330 159.850 64.500 160.350 ;
        RECT 69.880 159.850 70.050 160.350 ;
        RECT 64.670 159.620 69.710 159.790 ;
        RECT 64.330 159.060 64.500 159.560 ;
        RECT 69.880 159.060 70.050 159.560 ;
        RECT 64.670 158.830 69.710 159.000 ;
        RECT 64.330 158.270 64.500 158.770 ;
        RECT 69.880 158.270 70.050 158.770 ;
        RECT 64.670 158.040 69.710 158.210 ;
        RECT 64.330 157.480 64.500 157.980 ;
        RECT 69.880 157.480 70.050 157.980 ;
        RECT 64.670 157.250 69.710 157.420 ;
        RECT 64.330 156.690 64.500 157.190 ;
        RECT 69.880 156.690 70.050 157.190 ;
        RECT 64.670 156.460 69.710 156.630 ;
        RECT 64.330 155.900 64.500 156.400 ;
        RECT 69.880 155.900 70.050 156.400 ;
        RECT 64.670 155.670 69.710 155.840 ;
        RECT 64.330 155.110 64.500 155.610 ;
        RECT 69.880 155.110 70.050 155.610 ;
        RECT 64.670 154.880 69.710 155.050 ;
        RECT 64.330 154.320 64.500 154.820 ;
        RECT 69.880 154.320 70.050 154.820 ;
        RECT 64.670 154.090 69.710 154.260 ;
        RECT 64.330 153.530 64.500 154.030 ;
        RECT 69.880 153.530 70.050 154.030 ;
        RECT 64.670 153.300 69.710 153.470 ;
        RECT 64.330 152.740 64.500 153.240 ;
        RECT 69.880 152.740 70.050 153.240 ;
        RECT 64.670 152.510 69.710 152.680 ;
        RECT 64.330 151.950 64.500 152.450 ;
        RECT 69.880 151.950 70.050 152.450 ;
        RECT 64.670 151.720 69.710 151.890 ;
        RECT 64.330 151.160 64.500 151.660 ;
        RECT 69.880 151.160 70.050 151.660 ;
        RECT 64.670 150.930 69.710 151.100 ;
        RECT 64.330 150.370 64.500 150.870 ;
        RECT 69.880 150.370 70.050 150.870 ;
        RECT 64.670 150.140 69.710 150.310 ;
        RECT 64.330 149.580 64.500 150.080 ;
        RECT 69.880 149.580 70.050 150.080 ;
        RECT 64.670 149.350 69.710 149.520 ;
        RECT 64.330 148.790 64.500 149.290 ;
        RECT 69.880 148.790 70.050 149.290 ;
        RECT 64.670 148.560 69.710 148.730 ;
        RECT 64.330 148.000 64.500 148.500 ;
        RECT 69.880 148.000 70.050 148.500 ;
        RECT 64.670 147.770 69.710 147.940 ;
        RECT 64.330 147.210 64.500 147.710 ;
        RECT 69.880 147.210 70.050 147.710 ;
        RECT 64.670 146.980 69.710 147.150 ;
        RECT 70.480 146.590 70.650 162.720 ;
        RECT 72.100 158.090 72.280 170.750 ;
        RECT 73.030 168.520 78.070 168.690 ;
        RECT 82.030 168.520 87.070 168.690 ;
        RECT 72.645 167.960 72.815 168.460 ;
        RECT 78.285 167.960 78.455 168.460 ;
        RECT 81.645 167.960 81.815 168.460 ;
        RECT 87.285 167.960 87.455 168.460 ;
        RECT 73.030 167.730 78.070 167.900 ;
        RECT 82.030 167.730 87.070 167.900 ;
        RECT 73.030 164.020 78.070 164.190 ;
        RECT 82.030 164.020 87.070 164.190 ;
        RECT 72.645 163.460 72.815 163.960 ;
        RECT 78.285 163.460 78.455 163.960 ;
        RECT 81.645 163.460 81.815 163.960 ;
        RECT 87.285 163.460 87.455 163.960 ;
        RECT 73.030 163.230 78.070 163.400 ;
        RECT 82.030 163.230 87.070 163.400 ;
        RECT 73.030 159.520 78.070 159.690 ;
        RECT 82.030 159.520 87.070 159.690 ;
        RECT 72.645 158.960 72.815 159.460 ;
        RECT 78.285 158.960 78.455 159.460 ;
        RECT 81.645 158.960 81.815 159.460 ;
        RECT 87.285 158.960 87.455 159.460 ;
        RECT 73.030 158.730 78.070 158.900 ;
        RECT 82.030 158.730 87.070 158.900 ;
        RECT 88.030 158.090 88.210 170.750 ;
        RECT 88.870 170.780 104.430 170.950 ;
        RECT 88.870 158.260 89.040 170.780 ;
        RECT 90.750 169.000 95.790 169.170 ;
        RECT 97.750 169.000 102.790 169.170 ;
        RECT 90.410 167.940 90.580 168.940 ;
        RECT 95.960 167.940 96.130 168.940 ;
        RECT 97.410 167.940 97.580 168.940 ;
        RECT 102.960 167.940 103.130 168.940 ;
        RECT 90.750 167.710 95.790 167.880 ;
        RECT 97.750 167.710 102.790 167.880 ;
        RECT 90.750 167.000 95.790 167.170 ;
        RECT 97.750 167.000 102.790 167.170 ;
        RECT 90.410 165.940 90.580 166.940 ;
        RECT 95.960 165.940 96.130 166.940 ;
        RECT 97.410 165.940 97.580 166.940 ;
        RECT 102.960 165.940 103.130 166.940 ;
        RECT 90.750 165.710 95.790 165.880 ;
        RECT 97.750 165.710 102.790 165.880 ;
        RECT 90.750 163.000 95.790 163.170 ;
        RECT 97.750 163.000 102.790 163.170 ;
        RECT 90.410 161.940 90.580 162.940 ;
        RECT 95.960 161.940 96.130 162.940 ;
        RECT 97.410 161.940 97.580 162.940 ;
        RECT 102.960 161.940 103.130 162.940 ;
        RECT 90.750 161.710 95.790 161.880 ;
        RECT 97.750 161.710 102.790 161.880 ;
        RECT 90.750 161.000 95.790 161.170 ;
        RECT 97.750 161.000 102.790 161.170 ;
        RECT 90.410 159.940 90.580 160.940 ;
        RECT 95.960 159.940 96.130 160.940 ;
        RECT 97.410 159.940 97.580 160.940 ;
        RECT 102.960 159.940 103.130 160.940 ;
        RECT 90.750 159.710 95.790 159.880 ;
        RECT 97.750 159.710 102.790 159.880 ;
        RECT 104.260 158.260 104.430 170.780 ;
        RECT 88.870 158.090 104.430 158.260 ;
        RECT 105.290 170.920 113.690 171.090 ;
        RECT 105.290 158.120 105.460 170.920 ;
        RECT 106.210 170.310 111.250 170.480 ;
        RECT 105.870 169.250 106.040 170.250 ;
        RECT 111.420 169.250 111.590 170.250 ;
        RECT 106.210 169.020 111.250 169.190 ;
        RECT 105.870 167.960 106.040 168.960 ;
        RECT 111.420 167.960 111.590 168.960 ;
        RECT 106.210 167.730 111.250 167.900 ;
        RECT 105.870 166.670 106.040 167.670 ;
        RECT 111.420 166.670 111.590 167.670 ;
        RECT 106.210 166.440 111.250 166.610 ;
        RECT 105.870 165.380 106.040 166.380 ;
        RECT 111.420 165.380 111.590 166.380 ;
        RECT 106.210 165.150 111.250 165.320 ;
        RECT 105.870 164.090 106.040 165.090 ;
        RECT 111.420 164.090 111.590 165.090 ;
        RECT 106.210 163.860 111.250 164.030 ;
        RECT 105.870 162.800 106.040 163.800 ;
        RECT 111.420 162.800 111.590 163.800 ;
        RECT 106.210 162.570 111.250 162.740 ;
        RECT 105.870 161.510 106.040 162.510 ;
        RECT 111.420 161.510 111.590 162.510 ;
        RECT 106.210 161.280 111.250 161.450 ;
        RECT 105.870 160.220 106.040 161.220 ;
        RECT 111.420 160.220 111.590 161.220 ;
        RECT 106.210 159.990 111.250 160.160 ;
        RECT 113.520 158.120 113.690 170.920 ;
        RECT 122.895 168.565 123.075 172.455 ;
        RECT 123.795 171.630 124.795 171.800 ;
        RECT 125.085 171.630 126.085 171.800 ;
        RECT 123.565 169.375 123.735 171.415 ;
        RECT 124.855 169.375 125.025 171.415 ;
        RECT 126.145 169.375 126.315 171.415 ;
        RECT 123.795 168.990 124.795 169.160 ;
        RECT 125.085 168.990 126.085 169.160 ;
        RECT 126.825 168.565 126.995 172.455 ;
        RECT 122.895 168.355 126.995 168.565 ;
        RECT 127.345 172.455 130.845 172.625 ;
        RECT 127.345 172.445 130.855 172.455 ;
        RECT 127.345 168.565 127.515 172.445 ;
        RECT 130.675 171.345 130.855 172.445 ;
        RECT 127.985 171.155 128.985 171.325 ;
        RECT 129.275 171.155 130.275 171.325 ;
        RECT 127.755 169.945 127.925 170.985 ;
        RECT 129.045 169.945 129.215 170.985 ;
        RECT 130.335 169.945 130.505 170.985 ;
        RECT 127.985 169.605 128.985 169.775 ;
        RECT 129.275 169.605 130.275 169.775 ;
        RECT 130.675 168.565 130.845 171.345 ;
        RECT 127.345 168.355 130.845 168.565 ;
        RECT 126.085 164.525 126.885 164.535 ;
        RECT 122.895 164.355 126.995 164.525 ;
        RECT 114.655 163.190 118.155 163.400 ;
        RECT 114.655 160.410 114.825 163.190 ;
        RECT 115.225 161.980 116.225 162.150 ;
        RECT 116.515 161.980 117.515 162.150 ;
        RECT 114.995 160.770 115.165 161.810 ;
        RECT 116.285 160.770 116.455 161.810 ;
        RECT 117.575 160.770 117.745 161.810 ;
        RECT 115.225 160.430 116.225 160.600 ;
        RECT 116.515 160.430 117.515 160.600 ;
        RECT 114.645 159.310 114.825 160.410 ;
        RECT 117.985 159.310 118.155 163.190 ;
        RECT 114.645 159.300 118.155 159.310 ;
        RECT 114.655 159.130 118.155 159.300 ;
        RECT 118.505 163.190 122.605 163.400 ;
        RECT 118.505 159.300 118.675 163.190 ;
        RECT 119.415 162.595 120.415 162.765 ;
        RECT 120.705 162.595 121.705 162.765 ;
        RECT 119.185 160.340 119.355 162.380 ;
        RECT 120.475 160.340 120.645 162.380 ;
        RECT 121.765 160.340 121.935 162.380 ;
        RECT 119.415 159.955 120.415 160.125 ;
        RECT 120.705 159.955 121.705 160.125 ;
        RECT 122.425 159.300 122.605 163.190 ;
        RECT 122.895 160.465 123.075 164.355 ;
        RECT 123.795 163.530 124.795 163.700 ;
        RECT 125.085 163.530 126.085 163.700 ;
        RECT 123.565 161.275 123.735 163.315 ;
        RECT 124.855 161.275 125.025 163.315 ;
        RECT 126.145 161.275 126.315 163.315 ;
        RECT 123.795 160.890 124.795 161.060 ;
        RECT 125.085 160.890 126.085 161.060 ;
        RECT 126.825 160.465 126.995 164.355 ;
        RECT 122.895 160.255 126.995 160.465 ;
        RECT 127.345 164.355 130.845 164.525 ;
        RECT 127.345 164.345 130.855 164.355 ;
        RECT 127.345 160.465 127.515 164.345 ;
        RECT 130.675 163.245 130.855 164.345 ;
        RECT 127.985 163.055 128.985 163.225 ;
        RECT 129.275 163.055 130.275 163.225 ;
        RECT 127.755 161.845 127.925 162.885 ;
        RECT 129.045 161.845 129.215 162.885 ;
        RECT 130.335 161.845 130.505 162.885 ;
        RECT 127.985 161.505 128.985 161.675 ;
        RECT 129.275 161.505 130.275 161.675 ;
        RECT 130.675 160.465 130.845 163.245 ;
        RECT 127.345 160.255 130.845 160.465 ;
        RECT 118.505 159.130 122.605 159.300 ;
        RECT 118.615 159.120 119.415 159.130 ;
        RECT 72.100 157.910 88.210 158.090 ;
        RECT 105.290 157.950 113.690 158.120 ;
        RECT 114.655 158.650 118.155 158.860 ;
        RECT 63.340 146.410 70.650 146.590 ;
        RECT 72.100 156.130 88.210 156.310 ;
        RECT 72.100 143.470 72.280 156.130 ;
        RECT 73.030 155.320 78.070 155.490 ;
        RECT 82.030 155.320 87.070 155.490 ;
        RECT 72.645 154.760 72.815 155.260 ;
        RECT 78.285 154.760 78.455 155.260 ;
        RECT 81.645 154.760 81.815 155.260 ;
        RECT 87.285 154.760 87.455 155.260 ;
        RECT 73.030 154.530 78.070 154.700 ;
        RECT 82.030 154.530 87.070 154.700 ;
        RECT 73.030 150.820 78.070 150.990 ;
        RECT 82.030 150.820 87.070 150.990 ;
        RECT 72.645 150.260 72.815 150.760 ;
        RECT 78.285 150.260 78.455 150.760 ;
        RECT 81.645 150.260 81.815 150.760 ;
        RECT 87.285 150.260 87.455 150.760 ;
        RECT 73.030 150.030 78.070 150.200 ;
        RECT 82.030 150.030 87.070 150.200 ;
        RECT 73.030 146.320 78.070 146.490 ;
        RECT 82.030 146.320 87.070 146.490 ;
        RECT 72.645 145.760 72.815 146.260 ;
        RECT 78.285 145.760 78.455 146.260 ;
        RECT 81.645 145.760 81.815 146.260 ;
        RECT 87.285 145.760 87.455 146.260 ;
        RECT 73.030 145.530 78.070 145.700 ;
        RECT 82.030 145.530 87.070 145.700 ;
        RECT 88.030 143.470 88.210 156.130 ;
        RECT 72.100 143.290 88.210 143.470 ;
        RECT 88.870 155.960 104.430 156.130 ;
        RECT 88.870 143.440 89.040 155.960 ;
        RECT 90.750 154.340 95.790 154.510 ;
        RECT 97.750 154.340 102.790 154.510 ;
        RECT 90.410 153.280 90.580 154.280 ;
        RECT 95.960 153.280 96.130 154.280 ;
        RECT 97.410 153.280 97.580 154.280 ;
        RECT 102.960 153.280 103.130 154.280 ;
        RECT 90.750 153.050 95.790 153.220 ;
        RECT 97.750 153.050 102.790 153.220 ;
        RECT 90.750 152.340 95.790 152.510 ;
        RECT 97.750 152.340 102.790 152.510 ;
        RECT 90.410 151.280 90.580 152.280 ;
        RECT 95.960 151.280 96.130 152.280 ;
        RECT 97.410 151.280 97.580 152.280 ;
        RECT 102.960 151.280 103.130 152.280 ;
        RECT 90.750 151.050 95.790 151.220 ;
        RECT 97.750 151.050 102.790 151.220 ;
        RECT 90.750 148.340 95.790 148.510 ;
        RECT 97.750 148.340 102.790 148.510 ;
        RECT 90.410 147.280 90.580 148.280 ;
        RECT 95.960 147.280 96.130 148.280 ;
        RECT 97.410 147.280 97.580 148.280 ;
        RECT 102.960 147.280 103.130 148.280 ;
        RECT 90.750 147.050 95.790 147.220 ;
        RECT 97.750 147.050 102.790 147.220 ;
        RECT 90.750 146.340 95.790 146.510 ;
        RECT 97.750 146.340 102.790 146.510 ;
        RECT 90.410 145.280 90.580 146.280 ;
        RECT 95.960 145.280 96.130 146.280 ;
        RECT 97.410 145.280 97.580 146.280 ;
        RECT 102.960 145.280 103.130 146.280 ;
        RECT 90.750 145.050 95.790 145.220 ;
        RECT 97.750 145.050 102.790 145.220 ;
        RECT 104.260 143.440 104.430 155.960 ;
        RECT 88.870 143.270 104.430 143.440 ;
        RECT 105.290 156.100 113.690 156.270 ;
        RECT 105.290 143.300 105.460 156.100 ;
        RECT 106.210 154.060 111.250 154.230 ;
        RECT 105.870 153.000 106.040 154.000 ;
        RECT 111.420 153.000 111.590 154.000 ;
        RECT 106.210 152.770 111.250 152.940 ;
        RECT 105.870 151.710 106.040 152.710 ;
        RECT 111.420 151.710 111.590 152.710 ;
        RECT 106.210 151.480 111.250 151.650 ;
        RECT 105.870 150.420 106.040 151.420 ;
        RECT 111.420 150.420 111.590 151.420 ;
        RECT 106.210 150.190 111.250 150.360 ;
        RECT 105.870 149.130 106.040 150.130 ;
        RECT 111.420 149.130 111.590 150.130 ;
        RECT 106.210 148.900 111.250 149.070 ;
        RECT 105.870 147.840 106.040 148.840 ;
        RECT 111.420 147.840 111.590 148.840 ;
        RECT 106.210 147.610 111.250 147.780 ;
        RECT 105.870 146.550 106.040 147.550 ;
        RECT 111.420 146.550 111.590 147.550 ;
        RECT 106.210 146.320 111.250 146.490 ;
        RECT 105.870 145.260 106.040 146.260 ;
        RECT 111.420 145.260 111.590 146.260 ;
        RECT 106.210 145.030 111.250 145.200 ;
        RECT 105.870 143.970 106.040 144.970 ;
        RECT 111.420 143.970 111.590 144.970 ;
        RECT 106.210 143.740 111.250 143.910 ;
        RECT 113.520 143.300 113.690 156.100 ;
        RECT 114.655 155.870 114.825 158.650 ;
        RECT 115.225 157.440 116.225 157.610 ;
        RECT 116.515 157.440 117.515 157.610 ;
        RECT 114.995 156.230 115.165 157.270 ;
        RECT 116.285 156.230 116.455 157.270 ;
        RECT 117.575 156.230 117.745 157.270 ;
        RECT 115.225 155.890 116.225 156.060 ;
        RECT 116.515 155.890 117.515 156.060 ;
        RECT 114.645 154.800 114.825 155.870 ;
        RECT 117.985 154.800 118.155 158.650 ;
        RECT 114.645 154.760 118.155 154.800 ;
        RECT 114.655 154.590 118.155 154.760 ;
        RECT 114.655 151.810 114.825 154.590 ;
        RECT 115.225 153.380 116.225 153.550 ;
        RECT 116.515 153.380 117.515 153.550 ;
        RECT 114.995 152.170 115.165 153.210 ;
        RECT 116.285 152.170 116.455 153.210 ;
        RECT 117.575 152.170 117.745 153.210 ;
        RECT 115.225 151.830 116.225 152.000 ;
        RECT 116.515 151.830 117.515 152.000 ;
        RECT 114.645 150.740 114.825 151.810 ;
        RECT 117.985 150.740 118.155 154.590 ;
        RECT 114.645 150.700 118.155 150.740 ;
        RECT 114.655 150.530 118.155 150.700 ;
        RECT 114.655 147.750 114.825 150.530 ;
        RECT 115.225 149.320 116.225 149.490 ;
        RECT 116.515 149.320 117.515 149.490 ;
        RECT 114.995 148.110 115.165 149.150 ;
        RECT 116.285 148.110 116.455 149.150 ;
        RECT 117.575 148.110 117.745 149.150 ;
        RECT 115.225 147.770 116.225 147.940 ;
        RECT 116.515 147.770 117.515 147.940 ;
        RECT 114.645 146.680 114.825 147.750 ;
        RECT 117.985 146.680 118.155 150.530 ;
        RECT 114.645 146.640 118.155 146.680 ;
        RECT 114.655 146.470 118.155 146.640 ;
        RECT 114.655 143.690 114.825 146.470 ;
        RECT 115.225 145.260 116.225 145.430 ;
        RECT 116.515 145.260 117.515 145.430 ;
        RECT 114.995 144.050 115.165 145.090 ;
        RECT 116.285 144.050 116.455 145.090 ;
        RECT 117.575 144.050 117.745 145.090 ;
        RECT 115.225 143.710 116.225 143.880 ;
        RECT 116.515 143.710 117.515 143.880 ;
        RECT 105.290 143.130 113.690 143.300 ;
        RECT 94.680 142.500 106.670 142.670 ;
        RECT 108.420 142.665 109.060 142.670 ;
        RECT 109.600 142.665 110.240 142.670 ;
        RECT 111.000 142.665 111.640 142.670 ;
        RECT 112.650 142.665 113.290 142.670 ;
        RECT 94.680 140.740 94.850 142.500 ;
        RECT 95.575 141.930 103.115 142.100 ;
        RECT 95.190 141.370 95.360 141.870 ;
        RECT 103.330 141.370 103.500 141.870 ;
        RECT 95.575 141.140 103.115 141.310 ;
        RECT 103.840 140.740 104.010 142.500 ;
        RECT 104.735 141.930 105.775 142.100 ;
        RECT 104.350 141.370 104.520 141.870 ;
        RECT 105.990 141.370 106.160 141.870 ;
        RECT 104.735 141.140 105.775 141.310 ;
        RECT 106.500 140.740 106.670 142.500 ;
        RECT 94.680 140.570 106.670 140.740 ;
        RECT 107.030 142.495 113.770 142.665 ;
        RECT 114.645 142.620 114.825 143.690 ;
        RECT 117.985 142.620 118.155 146.470 ;
        RECT 114.645 142.580 118.155 142.620 ;
        RECT 97.830 140.295 102.780 140.300 ;
        RECT 95.175 140.125 104.005 140.295 ;
        RECT 95.175 139.820 95.345 140.125 ;
        RECT 95.175 138.680 95.350 139.820 ;
        RECT 96.070 139.555 103.110 139.725 ;
        RECT 95.685 138.995 95.855 139.495 ;
        RECT 103.325 138.995 103.495 139.495 ;
        RECT 96.070 138.765 103.110 138.935 ;
        RECT 95.175 138.365 95.345 138.680 ;
        RECT 103.835 138.365 104.005 140.125 ;
        RECT 107.030 140.235 107.200 142.495 ;
        RECT 107.880 141.925 112.920 142.095 ;
        RECT 107.540 140.865 107.710 141.865 ;
        RECT 113.090 140.865 113.260 141.865 ;
        RECT 107.880 140.635 112.920 140.805 ;
        RECT 113.600 140.235 113.770 142.495 ;
        RECT 107.030 140.065 113.770 140.235 ;
        RECT 114.655 142.410 118.155 142.580 ;
        RECT 114.655 139.630 114.825 142.410 ;
        RECT 115.225 141.200 116.225 141.370 ;
        RECT 116.515 141.200 117.515 141.370 ;
        RECT 114.995 139.990 115.165 141.030 ;
        RECT 116.285 139.990 116.455 141.030 ;
        RECT 117.575 139.990 117.745 141.030 ;
        RECT 115.225 139.650 116.225 139.820 ;
        RECT 116.515 139.650 117.515 139.820 ;
        RECT 114.645 138.530 114.825 139.630 ;
        RECT 117.985 138.530 118.155 142.410 ;
        RECT 114.645 138.520 118.155 138.530 ;
        RECT 95.175 138.195 104.005 138.365 ;
        RECT 114.655 138.350 118.155 138.520 ;
        RECT 118.505 158.650 122.605 158.860 ;
        RECT 118.505 154.800 118.675 158.650 ;
        RECT 119.415 158.055 120.415 158.225 ;
        RECT 120.705 158.055 121.705 158.225 ;
        RECT 119.185 155.800 119.355 157.840 ;
        RECT 120.475 155.800 120.645 157.840 ;
        RECT 121.765 155.800 121.935 157.840 ;
        RECT 119.415 155.415 120.415 155.585 ;
        RECT 120.705 155.415 121.705 155.585 ;
        RECT 122.425 154.800 122.605 158.650 ;
        RECT 126.085 156.425 126.885 156.435 ;
        RECT 118.505 154.590 122.605 154.800 ;
        RECT 118.505 154.580 119.415 154.590 ;
        RECT 118.505 150.740 118.675 154.580 ;
        RECT 119.415 153.995 120.415 154.165 ;
        RECT 120.705 153.995 121.705 154.165 ;
        RECT 119.185 151.740 119.355 153.780 ;
        RECT 120.475 151.740 120.645 153.780 ;
        RECT 121.765 151.740 121.935 153.780 ;
        RECT 119.415 151.355 120.415 151.525 ;
        RECT 120.705 151.355 121.705 151.525 ;
        RECT 122.425 150.740 122.605 154.590 ;
        RECT 122.895 156.255 126.995 156.425 ;
        RECT 122.895 152.365 123.075 156.255 ;
        RECT 123.795 155.430 124.795 155.600 ;
        RECT 125.085 155.430 126.085 155.600 ;
        RECT 123.565 153.175 123.735 155.215 ;
        RECT 124.855 153.175 125.025 155.215 ;
        RECT 126.145 153.175 126.315 155.215 ;
        RECT 123.795 152.790 124.795 152.960 ;
        RECT 125.085 152.790 126.085 152.960 ;
        RECT 126.825 152.365 126.995 156.255 ;
        RECT 122.895 152.155 126.995 152.365 ;
        RECT 127.345 156.255 130.845 156.425 ;
        RECT 127.345 156.245 130.855 156.255 ;
        RECT 127.345 152.365 127.515 156.245 ;
        RECT 130.675 155.145 130.855 156.245 ;
        RECT 127.985 154.955 128.985 155.125 ;
        RECT 129.275 154.955 130.275 155.125 ;
        RECT 127.755 153.745 127.925 154.785 ;
        RECT 129.045 153.745 129.215 154.785 ;
        RECT 130.335 153.745 130.505 154.785 ;
        RECT 127.985 153.405 128.985 153.575 ;
        RECT 129.275 153.405 130.275 153.575 ;
        RECT 130.675 152.365 130.845 155.145 ;
        RECT 127.345 152.155 130.845 152.365 ;
        RECT 118.505 150.530 122.605 150.740 ;
        RECT 118.505 150.520 119.415 150.530 ;
        RECT 118.505 146.680 118.675 150.520 ;
        RECT 119.415 149.935 120.415 150.105 ;
        RECT 120.705 149.935 121.705 150.105 ;
        RECT 119.185 147.680 119.355 149.720 ;
        RECT 120.475 147.680 120.645 149.720 ;
        RECT 121.765 147.680 121.935 149.720 ;
        RECT 119.415 147.295 120.415 147.465 ;
        RECT 120.705 147.295 121.705 147.465 ;
        RECT 122.425 146.680 122.605 150.530 ;
        RECT 126.085 148.325 126.885 148.335 ;
        RECT 118.505 146.470 122.605 146.680 ;
        RECT 118.505 146.460 119.415 146.470 ;
        RECT 118.505 142.620 118.675 146.460 ;
        RECT 119.415 145.875 120.415 146.045 ;
        RECT 120.705 145.875 121.705 146.045 ;
        RECT 119.185 143.620 119.355 145.660 ;
        RECT 120.475 143.620 120.645 145.660 ;
        RECT 121.765 143.620 121.935 145.660 ;
        RECT 119.415 143.235 120.415 143.405 ;
        RECT 120.705 143.235 121.705 143.405 ;
        RECT 122.425 142.620 122.605 146.470 ;
        RECT 122.895 148.155 126.995 148.325 ;
        RECT 122.895 144.265 123.075 148.155 ;
        RECT 123.795 147.330 124.795 147.500 ;
        RECT 125.085 147.330 126.085 147.500 ;
        RECT 123.565 145.075 123.735 147.115 ;
        RECT 124.855 145.075 125.025 147.115 ;
        RECT 126.145 145.075 126.315 147.115 ;
        RECT 123.795 144.690 124.795 144.860 ;
        RECT 125.085 144.690 126.085 144.860 ;
        RECT 126.825 144.265 126.995 148.155 ;
        RECT 122.895 144.055 126.995 144.265 ;
        RECT 127.345 148.155 130.845 148.325 ;
        RECT 127.345 148.145 130.855 148.155 ;
        RECT 127.345 144.265 127.515 148.145 ;
        RECT 130.675 147.045 130.855 148.145 ;
        RECT 127.985 146.855 128.985 147.025 ;
        RECT 129.275 146.855 130.275 147.025 ;
        RECT 127.755 145.645 127.925 146.685 ;
        RECT 129.045 145.645 129.215 146.685 ;
        RECT 130.335 145.645 130.505 146.685 ;
        RECT 127.985 145.305 128.985 145.475 ;
        RECT 129.275 145.305 130.275 145.475 ;
        RECT 130.675 144.265 130.845 147.045 ;
        RECT 127.345 144.055 130.845 144.265 ;
        RECT 118.505 142.410 122.605 142.620 ;
        RECT 118.505 142.400 119.415 142.410 ;
        RECT 118.505 138.520 118.675 142.400 ;
        RECT 119.415 141.815 120.415 141.985 ;
        RECT 120.705 141.815 121.705 141.985 ;
        RECT 119.185 139.560 119.355 141.600 ;
        RECT 120.475 139.560 120.645 141.600 ;
        RECT 121.765 139.560 121.935 141.600 ;
        RECT 119.415 139.175 120.415 139.345 ;
        RECT 120.705 139.175 121.705 139.345 ;
        RECT 122.425 138.520 122.605 142.410 ;
        RECT 126.085 140.225 126.885 140.235 ;
        RECT 118.505 138.350 122.605 138.520 ;
        RECT 122.895 140.055 126.995 140.225 ;
        RECT 118.615 138.340 119.415 138.350 ;
        RECT 95.175 137.890 95.345 138.195 ;
        RECT 95.175 136.750 95.350 137.890 ;
        RECT 96.070 137.625 103.110 137.795 ;
        RECT 95.685 137.065 95.855 137.565 ;
        RECT 103.325 137.065 103.495 137.565 ;
        RECT 96.070 136.835 103.110 137.005 ;
        RECT 95.175 136.435 95.345 136.750 ;
        RECT 103.835 136.435 104.005 138.195 ;
        RECT 95.175 136.265 104.005 136.435 ;
        RECT 122.895 136.165 123.075 140.055 ;
        RECT 123.795 139.230 124.795 139.400 ;
        RECT 125.085 139.230 126.085 139.400 ;
        RECT 123.565 136.975 123.735 139.015 ;
        RECT 124.855 136.975 125.025 139.015 ;
        RECT 126.145 136.975 126.315 139.015 ;
        RECT 123.795 136.590 124.795 136.760 ;
        RECT 125.085 136.590 126.085 136.760 ;
        RECT 126.825 136.165 126.995 140.055 ;
        RECT 122.895 135.955 126.995 136.165 ;
        RECT 127.345 140.055 130.845 140.225 ;
        RECT 127.345 140.045 130.855 140.055 ;
        RECT 127.345 136.165 127.515 140.045 ;
        RECT 130.675 138.945 130.855 140.045 ;
        RECT 127.985 138.755 128.985 138.925 ;
        RECT 129.275 138.755 130.275 138.925 ;
        RECT 127.755 137.545 127.925 138.585 ;
        RECT 129.045 137.545 129.215 138.585 ;
        RECT 130.335 137.545 130.505 138.585 ;
        RECT 127.985 137.205 128.985 137.375 ;
        RECT 129.275 137.205 130.275 137.375 ;
        RECT 130.675 136.165 130.845 138.945 ;
        RECT 127.345 135.955 130.845 136.165 ;
        RECT 98.770 135.450 105.540 135.620 ;
        RECT 98.770 122.690 98.940 135.450 ;
        RECT 99.620 134.530 104.660 134.700 ;
        RECT 99.235 133.970 99.405 134.470 ;
        RECT 104.875 133.970 105.045 134.470 ;
        RECT 99.620 133.740 104.660 133.910 ;
        RECT 99.235 133.180 99.405 133.680 ;
        RECT 104.875 133.180 105.045 133.680 ;
        RECT 99.620 132.950 104.660 133.120 ;
        RECT 99.235 132.390 99.405 132.890 ;
        RECT 104.875 132.390 105.045 132.890 ;
        RECT 99.620 132.160 104.660 132.330 ;
        RECT 99.235 131.600 99.405 132.100 ;
        RECT 104.875 131.600 105.045 132.100 ;
        RECT 99.620 131.370 104.660 131.540 ;
        RECT 99.235 130.810 99.405 131.310 ;
        RECT 104.875 130.810 105.045 131.310 ;
        RECT 99.620 130.580 104.660 130.750 ;
        RECT 99.235 130.020 99.405 130.520 ;
        RECT 104.875 130.020 105.045 130.520 ;
        RECT 99.620 129.790 104.660 129.960 ;
        RECT 99.235 129.230 99.405 129.730 ;
        RECT 104.875 129.230 105.045 129.730 ;
        RECT 99.620 129.000 104.660 129.170 ;
        RECT 99.235 128.440 99.405 128.940 ;
        RECT 104.875 128.440 105.045 128.940 ;
        RECT 99.620 128.210 104.660 128.380 ;
        RECT 99.235 127.650 99.405 128.150 ;
        RECT 104.875 127.650 105.045 128.150 ;
        RECT 99.620 127.420 104.660 127.590 ;
        RECT 99.235 126.860 99.405 127.360 ;
        RECT 104.875 126.860 105.045 127.360 ;
        RECT 99.620 126.630 104.660 126.800 ;
        RECT 99.235 126.070 99.405 126.570 ;
        RECT 104.875 126.070 105.045 126.570 ;
        RECT 99.620 125.840 104.660 126.010 ;
        RECT 99.235 125.280 99.405 125.780 ;
        RECT 104.875 125.280 105.045 125.780 ;
        RECT 99.620 125.050 104.660 125.220 ;
        RECT 99.235 124.490 99.405 124.990 ;
        RECT 104.875 124.490 105.045 124.990 ;
        RECT 99.620 124.260 104.660 124.430 ;
        RECT 99.235 123.700 99.405 124.200 ;
        RECT 104.875 123.700 105.045 124.200 ;
        RECT 99.620 123.470 104.660 123.640 ;
        RECT 105.370 122.690 105.540 135.450 ;
        RECT 98.770 122.520 105.540 122.690 ;
        RECT 106.350 135.440 113.660 135.620 ;
        RECT 14.340 121.800 17.770 121.970 ;
        RECT 106.350 119.310 106.520 135.440 ;
        RECT 107.680 134.710 112.720 134.880 ;
        RECT 107.340 134.150 107.510 134.650 ;
        RECT 112.890 134.150 113.060 134.650 ;
        RECT 107.680 133.920 112.720 134.090 ;
        RECT 107.340 133.360 107.510 133.860 ;
        RECT 112.890 133.360 113.060 133.860 ;
        RECT 107.680 133.130 112.720 133.300 ;
        RECT 107.340 132.570 107.510 133.070 ;
        RECT 112.890 132.570 113.060 133.070 ;
        RECT 107.680 132.340 112.720 132.510 ;
        RECT 107.340 131.780 107.510 132.280 ;
        RECT 112.890 131.780 113.060 132.280 ;
        RECT 107.680 131.550 112.720 131.720 ;
        RECT 107.340 130.990 107.510 131.490 ;
        RECT 112.890 130.990 113.060 131.490 ;
        RECT 107.680 130.760 112.720 130.930 ;
        RECT 107.340 130.200 107.510 130.700 ;
        RECT 112.890 130.200 113.060 130.700 ;
        RECT 107.680 129.970 112.720 130.140 ;
        RECT 107.340 129.410 107.510 129.910 ;
        RECT 112.890 129.410 113.060 129.910 ;
        RECT 107.680 129.180 112.720 129.350 ;
        RECT 107.340 128.620 107.510 129.120 ;
        RECT 112.890 128.620 113.060 129.120 ;
        RECT 107.680 128.390 112.720 128.560 ;
        RECT 107.340 127.830 107.510 128.330 ;
        RECT 112.890 127.830 113.060 128.330 ;
        RECT 107.680 127.600 112.720 127.770 ;
        RECT 107.340 127.040 107.510 127.540 ;
        RECT 112.890 127.040 113.060 127.540 ;
        RECT 107.680 126.810 112.720 126.980 ;
        RECT 107.340 126.250 107.510 126.750 ;
        RECT 112.890 126.250 113.060 126.750 ;
        RECT 107.680 126.020 112.720 126.190 ;
        RECT 107.340 125.460 107.510 125.960 ;
        RECT 112.890 125.460 113.060 125.960 ;
        RECT 107.680 125.230 112.720 125.400 ;
        RECT 107.340 124.670 107.510 125.170 ;
        RECT 112.890 124.670 113.060 125.170 ;
        RECT 107.680 124.440 112.720 124.610 ;
        RECT 107.340 123.880 107.510 124.380 ;
        RECT 112.890 123.880 113.060 124.380 ;
        RECT 107.680 123.650 112.720 123.820 ;
        RECT 107.340 123.090 107.510 123.590 ;
        RECT 112.890 123.090 113.060 123.590 ;
        RECT 107.680 122.860 112.720 123.030 ;
        RECT 107.340 122.300 107.510 122.800 ;
        RECT 112.890 122.300 113.060 122.800 ;
        RECT 107.680 122.070 112.720 122.240 ;
        RECT 107.340 121.510 107.510 122.010 ;
        RECT 112.890 121.510 113.060 122.010 ;
        RECT 107.680 121.280 112.720 121.450 ;
        RECT 107.340 120.720 107.510 121.220 ;
        RECT 112.890 120.720 113.060 121.220 ;
        RECT 107.680 120.490 112.720 120.660 ;
        RECT 107.340 119.930 107.510 120.430 ;
        RECT 112.890 119.930 113.060 120.430 ;
        RECT 107.680 119.700 112.720 119.870 ;
        RECT 113.490 119.310 113.660 135.440 ;
        RECT 114.655 134.290 118.155 134.500 ;
        RECT 114.655 131.510 114.825 134.290 ;
        RECT 115.225 133.080 116.225 133.250 ;
        RECT 116.515 133.080 117.515 133.250 ;
        RECT 114.995 131.870 115.165 132.910 ;
        RECT 116.285 131.870 116.455 132.910 ;
        RECT 117.575 131.870 117.745 132.910 ;
        RECT 115.225 131.530 116.225 131.700 ;
        RECT 116.515 131.530 117.515 131.700 ;
        RECT 114.645 130.440 114.825 131.510 ;
        RECT 117.985 130.440 118.155 134.290 ;
        RECT 114.645 130.400 118.155 130.440 ;
        RECT 114.655 130.230 118.155 130.400 ;
        RECT 114.655 127.450 114.825 130.230 ;
        RECT 115.225 129.020 116.225 129.190 ;
        RECT 116.515 129.020 117.515 129.190 ;
        RECT 114.995 127.810 115.165 128.850 ;
        RECT 116.285 127.810 116.455 128.850 ;
        RECT 117.575 127.810 117.745 128.850 ;
        RECT 115.225 127.470 116.225 127.640 ;
        RECT 116.515 127.470 117.515 127.640 ;
        RECT 114.645 126.380 114.825 127.450 ;
        RECT 117.985 126.380 118.155 130.230 ;
        RECT 114.645 126.340 118.155 126.380 ;
        RECT 114.655 126.170 118.155 126.340 ;
        RECT 114.655 123.390 114.825 126.170 ;
        RECT 115.225 124.960 116.225 125.130 ;
        RECT 116.515 124.960 117.515 125.130 ;
        RECT 114.995 123.750 115.165 124.790 ;
        RECT 116.285 123.750 116.455 124.790 ;
        RECT 117.575 123.750 117.745 124.790 ;
        RECT 115.225 123.410 116.225 123.580 ;
        RECT 116.515 123.410 117.515 123.580 ;
        RECT 114.645 122.320 114.825 123.390 ;
        RECT 117.985 122.320 118.155 126.170 ;
        RECT 114.645 122.280 118.155 122.320 ;
        RECT 114.655 122.110 118.155 122.280 ;
        RECT 114.655 119.330 114.825 122.110 ;
        RECT 115.225 120.900 116.225 121.070 ;
        RECT 116.515 120.900 117.515 121.070 ;
        RECT 114.995 119.690 115.165 120.730 ;
        RECT 116.285 119.690 116.455 120.730 ;
        RECT 117.575 119.690 117.745 120.730 ;
        RECT 115.225 119.350 116.225 119.520 ;
        RECT 116.515 119.350 117.515 119.520 ;
        RECT 106.350 119.130 113.660 119.310 ;
        RECT 114.645 118.260 114.825 119.330 ;
        RECT 117.985 118.260 118.155 122.110 ;
        RECT 114.645 118.220 118.155 118.260 ;
        RECT 106.350 118.000 113.660 118.180 ;
        RECT 98.770 114.620 105.540 114.790 ;
        RECT 14.350 105.260 17.780 105.430 ;
        RECT 14.350 75.000 14.520 105.260 ;
        RECT 15.000 104.530 15.500 104.700 ;
        RECT 15.080 102.715 15.420 104.530 ;
        RECT 15.080 75.730 15.420 77.545 ;
        RECT 15.000 75.560 15.500 75.730 ;
        RECT 15.980 75.000 16.150 105.260 ;
        RECT 16.630 104.530 17.130 104.700 ;
        RECT 16.710 102.715 17.050 104.530 ;
        RECT 16.710 75.730 17.050 77.545 ;
        RECT 16.630 75.560 17.130 75.730 ;
        RECT 17.610 75.000 17.780 105.260 ;
        RECT 98.770 101.860 98.940 114.620 ;
        RECT 99.620 113.670 104.660 113.840 ;
        RECT 99.235 113.110 99.405 113.610 ;
        RECT 104.875 113.110 105.045 113.610 ;
        RECT 99.620 112.880 104.660 113.050 ;
        RECT 99.235 112.320 99.405 112.820 ;
        RECT 104.875 112.320 105.045 112.820 ;
        RECT 99.620 112.090 104.660 112.260 ;
        RECT 99.235 111.530 99.405 112.030 ;
        RECT 104.875 111.530 105.045 112.030 ;
        RECT 99.620 111.300 104.660 111.470 ;
        RECT 99.235 110.740 99.405 111.240 ;
        RECT 104.875 110.740 105.045 111.240 ;
        RECT 99.620 110.510 104.660 110.680 ;
        RECT 99.235 109.950 99.405 110.450 ;
        RECT 104.875 109.950 105.045 110.450 ;
        RECT 99.620 109.720 104.660 109.890 ;
        RECT 99.235 109.160 99.405 109.660 ;
        RECT 104.875 109.160 105.045 109.660 ;
        RECT 99.620 108.930 104.660 109.100 ;
        RECT 99.235 108.370 99.405 108.870 ;
        RECT 104.875 108.370 105.045 108.870 ;
        RECT 99.620 108.140 104.660 108.310 ;
        RECT 99.235 107.580 99.405 108.080 ;
        RECT 104.875 107.580 105.045 108.080 ;
        RECT 99.620 107.350 104.660 107.520 ;
        RECT 99.235 106.790 99.405 107.290 ;
        RECT 104.875 106.790 105.045 107.290 ;
        RECT 99.620 106.560 104.660 106.730 ;
        RECT 99.235 106.000 99.405 106.500 ;
        RECT 104.875 106.000 105.045 106.500 ;
        RECT 99.620 105.770 104.660 105.940 ;
        RECT 99.235 105.210 99.405 105.710 ;
        RECT 104.875 105.210 105.045 105.710 ;
        RECT 99.620 104.980 104.660 105.150 ;
        RECT 99.235 104.420 99.405 104.920 ;
        RECT 104.875 104.420 105.045 104.920 ;
        RECT 99.620 104.190 104.660 104.360 ;
        RECT 99.235 103.630 99.405 104.130 ;
        RECT 104.875 103.630 105.045 104.130 ;
        RECT 99.620 103.400 104.660 103.570 ;
        RECT 99.235 102.840 99.405 103.340 ;
        RECT 104.875 102.840 105.045 103.340 ;
        RECT 99.620 102.610 104.660 102.780 ;
        RECT 105.370 101.860 105.540 114.620 ;
        RECT 98.770 101.690 105.540 101.860 ;
        RECT 106.350 101.870 106.520 118.000 ;
        RECT 107.680 117.440 112.720 117.610 ;
        RECT 107.340 116.880 107.510 117.380 ;
        RECT 112.890 116.880 113.060 117.380 ;
        RECT 107.680 116.650 112.720 116.820 ;
        RECT 107.340 116.090 107.510 116.590 ;
        RECT 112.890 116.090 113.060 116.590 ;
        RECT 107.680 115.860 112.720 116.030 ;
        RECT 107.340 115.300 107.510 115.800 ;
        RECT 112.890 115.300 113.060 115.800 ;
        RECT 107.680 115.070 112.720 115.240 ;
        RECT 107.340 114.510 107.510 115.010 ;
        RECT 112.890 114.510 113.060 115.010 ;
        RECT 107.680 114.280 112.720 114.450 ;
        RECT 107.340 113.720 107.510 114.220 ;
        RECT 112.890 113.720 113.060 114.220 ;
        RECT 107.680 113.490 112.720 113.660 ;
        RECT 107.340 112.930 107.510 113.430 ;
        RECT 112.890 112.930 113.060 113.430 ;
        RECT 107.680 112.700 112.720 112.870 ;
        RECT 107.340 112.140 107.510 112.640 ;
        RECT 112.890 112.140 113.060 112.640 ;
        RECT 107.680 111.910 112.720 112.080 ;
        RECT 107.340 111.350 107.510 111.850 ;
        RECT 112.890 111.350 113.060 111.850 ;
        RECT 107.680 111.120 112.720 111.290 ;
        RECT 107.340 110.560 107.510 111.060 ;
        RECT 112.890 110.560 113.060 111.060 ;
        RECT 107.680 110.330 112.720 110.500 ;
        RECT 107.340 109.770 107.510 110.270 ;
        RECT 112.890 109.770 113.060 110.270 ;
        RECT 107.680 109.540 112.720 109.710 ;
        RECT 107.340 108.980 107.510 109.480 ;
        RECT 112.890 108.980 113.060 109.480 ;
        RECT 107.680 108.750 112.720 108.920 ;
        RECT 107.340 108.190 107.510 108.690 ;
        RECT 112.890 108.190 113.060 108.690 ;
        RECT 107.680 107.960 112.720 108.130 ;
        RECT 107.340 107.400 107.510 107.900 ;
        RECT 112.890 107.400 113.060 107.900 ;
        RECT 107.680 107.170 112.720 107.340 ;
        RECT 107.340 106.610 107.510 107.110 ;
        RECT 112.890 106.610 113.060 107.110 ;
        RECT 107.680 106.380 112.720 106.550 ;
        RECT 107.340 105.820 107.510 106.320 ;
        RECT 112.890 105.820 113.060 106.320 ;
        RECT 107.680 105.590 112.720 105.760 ;
        RECT 107.340 105.030 107.510 105.530 ;
        RECT 112.890 105.030 113.060 105.530 ;
        RECT 107.680 104.800 112.720 104.970 ;
        RECT 107.340 104.240 107.510 104.740 ;
        RECT 112.890 104.240 113.060 104.740 ;
        RECT 107.680 104.010 112.720 104.180 ;
        RECT 107.340 103.450 107.510 103.950 ;
        RECT 112.890 103.450 113.060 103.950 ;
        RECT 107.680 103.220 112.720 103.390 ;
        RECT 107.340 102.660 107.510 103.160 ;
        RECT 112.890 102.660 113.060 103.160 ;
        RECT 107.680 102.430 112.720 102.600 ;
        RECT 113.490 101.870 113.660 118.000 ;
        RECT 114.655 118.050 118.155 118.220 ;
        RECT 114.655 115.270 114.825 118.050 ;
        RECT 115.225 116.840 116.225 117.010 ;
        RECT 116.515 116.840 117.515 117.010 ;
        RECT 114.995 115.630 115.165 116.670 ;
        RECT 116.285 115.630 116.455 116.670 ;
        RECT 117.575 115.630 117.745 116.670 ;
        RECT 115.225 115.290 116.225 115.460 ;
        RECT 116.515 115.290 117.515 115.460 ;
        RECT 114.645 114.200 114.825 115.270 ;
        RECT 117.985 114.200 118.155 118.050 ;
        RECT 114.645 114.160 118.155 114.200 ;
        RECT 114.655 113.990 118.155 114.160 ;
        RECT 114.655 111.210 114.825 113.990 ;
        RECT 115.225 112.780 116.225 112.950 ;
        RECT 116.515 112.780 117.515 112.950 ;
        RECT 114.995 111.570 115.165 112.610 ;
        RECT 116.285 111.570 116.455 112.610 ;
        RECT 117.575 111.570 117.745 112.610 ;
        RECT 115.225 111.230 116.225 111.400 ;
        RECT 116.515 111.230 117.515 111.400 ;
        RECT 114.645 110.140 114.825 111.210 ;
        RECT 117.985 110.140 118.155 113.990 ;
        RECT 114.645 110.100 118.155 110.140 ;
        RECT 114.655 109.930 118.155 110.100 ;
        RECT 114.655 107.150 114.825 109.930 ;
        RECT 115.225 108.720 116.225 108.890 ;
        RECT 116.515 108.720 117.515 108.890 ;
        RECT 114.995 107.510 115.165 108.550 ;
        RECT 116.285 107.510 116.455 108.550 ;
        RECT 117.575 107.510 117.745 108.550 ;
        RECT 115.225 107.170 116.225 107.340 ;
        RECT 116.515 107.170 117.515 107.340 ;
        RECT 114.645 106.080 114.825 107.150 ;
        RECT 117.985 106.080 118.155 109.930 ;
        RECT 114.645 106.040 118.155 106.080 ;
        RECT 114.655 105.870 118.155 106.040 ;
        RECT 114.655 103.090 114.825 105.870 ;
        RECT 115.225 104.660 116.225 104.830 ;
        RECT 116.515 104.660 117.515 104.830 ;
        RECT 114.995 103.450 115.165 104.490 ;
        RECT 116.285 103.450 116.455 104.490 ;
        RECT 117.575 103.450 117.745 104.490 ;
        RECT 115.225 103.110 116.225 103.280 ;
        RECT 116.515 103.110 117.515 103.280 ;
        RECT 114.645 102.020 114.825 103.090 ;
        RECT 117.985 102.020 118.155 105.870 ;
        RECT 114.645 101.980 118.155 102.020 ;
        RECT 106.350 101.690 113.660 101.870 ;
        RECT 114.655 101.810 118.155 101.980 ;
        RECT 95.175 100.875 104.005 101.045 ;
        RECT 95.175 100.560 95.345 100.875 ;
        RECT 95.175 99.420 95.350 100.560 ;
        RECT 96.070 100.305 103.110 100.475 ;
        RECT 95.685 99.745 95.855 100.245 ;
        RECT 103.325 99.745 103.495 100.245 ;
        RECT 96.070 99.515 103.110 99.685 ;
        RECT 95.175 99.115 95.345 99.420 ;
        RECT 103.835 99.115 104.005 100.875 ;
        RECT 95.175 98.945 104.005 99.115 ;
        RECT 114.655 99.030 114.825 101.810 ;
        RECT 115.225 100.600 116.225 100.770 ;
        RECT 116.515 100.600 117.515 100.770 ;
        RECT 114.995 99.390 115.165 100.430 ;
        RECT 116.285 99.390 116.455 100.430 ;
        RECT 117.575 99.390 117.745 100.430 ;
        RECT 115.225 99.050 116.225 99.220 ;
        RECT 116.515 99.050 117.515 99.220 ;
        RECT 95.175 98.630 95.345 98.945 ;
        RECT 95.175 97.490 95.350 98.630 ;
        RECT 96.070 98.375 103.110 98.545 ;
        RECT 95.685 97.815 95.855 98.315 ;
        RECT 103.325 97.815 103.495 98.315 ;
        RECT 96.070 97.585 103.110 97.755 ;
        RECT 95.175 97.185 95.345 97.490 ;
        RECT 103.835 97.185 104.005 98.945 ;
        RECT 114.645 97.930 114.825 99.030 ;
        RECT 117.985 97.930 118.155 101.810 ;
        RECT 114.645 97.920 118.155 97.930 ;
        RECT 114.655 97.750 118.155 97.920 ;
        RECT 118.505 134.290 122.605 134.500 ;
        RECT 118.505 130.440 118.675 134.290 ;
        RECT 119.415 133.695 120.415 133.865 ;
        RECT 120.705 133.695 121.705 133.865 ;
        RECT 119.185 131.440 119.355 133.480 ;
        RECT 120.475 131.440 120.645 133.480 ;
        RECT 121.765 131.440 121.935 133.480 ;
        RECT 119.415 131.055 120.415 131.225 ;
        RECT 120.705 131.055 121.705 131.225 ;
        RECT 122.425 130.440 122.605 134.290 ;
        RECT 126.085 132.125 126.885 132.135 ;
        RECT 118.505 130.230 122.605 130.440 ;
        RECT 118.505 130.220 119.415 130.230 ;
        RECT 118.505 126.380 118.675 130.220 ;
        RECT 119.415 129.635 120.415 129.805 ;
        RECT 120.705 129.635 121.705 129.805 ;
        RECT 119.185 127.380 119.355 129.420 ;
        RECT 120.475 127.380 120.645 129.420 ;
        RECT 121.765 127.380 121.935 129.420 ;
        RECT 119.415 126.995 120.415 127.165 ;
        RECT 120.705 126.995 121.705 127.165 ;
        RECT 122.425 126.380 122.605 130.230 ;
        RECT 122.895 131.955 126.995 132.125 ;
        RECT 122.895 128.065 123.075 131.955 ;
        RECT 123.795 131.130 124.795 131.300 ;
        RECT 125.085 131.130 126.085 131.300 ;
        RECT 123.565 128.875 123.735 130.915 ;
        RECT 124.855 128.875 125.025 130.915 ;
        RECT 126.145 128.875 126.315 130.915 ;
        RECT 123.795 128.490 124.795 128.660 ;
        RECT 125.085 128.490 126.085 128.660 ;
        RECT 126.825 128.065 126.995 131.955 ;
        RECT 122.895 127.855 126.995 128.065 ;
        RECT 127.345 131.955 130.845 132.125 ;
        RECT 127.345 131.945 130.855 131.955 ;
        RECT 127.345 128.065 127.515 131.945 ;
        RECT 130.675 130.845 130.855 131.945 ;
        RECT 127.985 130.655 128.985 130.825 ;
        RECT 129.275 130.655 130.275 130.825 ;
        RECT 127.755 129.445 127.925 130.485 ;
        RECT 129.045 129.445 129.215 130.485 ;
        RECT 130.335 129.445 130.505 130.485 ;
        RECT 127.985 129.105 128.985 129.275 ;
        RECT 129.275 129.105 130.275 129.275 ;
        RECT 130.675 128.065 130.845 130.845 ;
        RECT 127.345 127.855 130.845 128.065 ;
        RECT 118.505 126.170 122.605 126.380 ;
        RECT 118.505 126.160 119.415 126.170 ;
        RECT 118.505 122.320 118.675 126.160 ;
        RECT 119.415 125.575 120.415 125.745 ;
        RECT 120.705 125.575 121.705 125.745 ;
        RECT 119.185 123.320 119.355 125.360 ;
        RECT 120.475 123.320 120.645 125.360 ;
        RECT 121.765 123.320 121.935 125.360 ;
        RECT 119.415 122.935 120.415 123.105 ;
        RECT 120.705 122.935 121.705 123.105 ;
        RECT 122.425 122.320 122.605 126.170 ;
        RECT 126.085 124.025 126.885 124.035 ;
        RECT 118.505 122.110 122.605 122.320 ;
        RECT 118.505 122.100 119.415 122.110 ;
        RECT 118.505 118.260 118.675 122.100 ;
        RECT 119.415 121.515 120.415 121.685 ;
        RECT 120.705 121.515 121.705 121.685 ;
        RECT 119.185 119.260 119.355 121.300 ;
        RECT 120.475 119.260 120.645 121.300 ;
        RECT 121.765 119.260 121.935 121.300 ;
        RECT 119.415 118.875 120.415 119.045 ;
        RECT 120.705 118.875 121.705 119.045 ;
        RECT 122.425 118.260 122.605 122.110 ;
        RECT 122.895 123.855 126.995 124.025 ;
        RECT 122.895 119.965 123.075 123.855 ;
        RECT 123.795 123.030 124.795 123.200 ;
        RECT 125.085 123.030 126.085 123.200 ;
        RECT 123.565 120.775 123.735 122.815 ;
        RECT 124.855 120.775 125.025 122.815 ;
        RECT 126.145 120.775 126.315 122.815 ;
        RECT 123.795 120.390 124.795 120.560 ;
        RECT 125.085 120.390 126.085 120.560 ;
        RECT 126.825 119.965 126.995 123.855 ;
        RECT 122.895 119.755 126.995 119.965 ;
        RECT 127.345 123.855 130.845 124.025 ;
        RECT 127.345 123.845 130.855 123.855 ;
        RECT 127.345 119.965 127.515 123.845 ;
        RECT 130.675 122.745 130.855 123.845 ;
        RECT 127.985 122.555 128.985 122.725 ;
        RECT 129.275 122.555 130.275 122.725 ;
        RECT 127.755 121.345 127.925 122.385 ;
        RECT 129.045 121.345 129.215 122.385 ;
        RECT 130.335 121.345 130.505 122.385 ;
        RECT 127.985 121.005 128.985 121.175 ;
        RECT 129.275 121.005 130.275 121.175 ;
        RECT 130.675 119.965 130.845 122.745 ;
        RECT 127.345 119.755 130.845 119.965 ;
        RECT 118.505 118.050 122.605 118.260 ;
        RECT 118.505 118.040 119.415 118.050 ;
        RECT 118.505 114.200 118.675 118.040 ;
        RECT 119.415 117.455 120.415 117.625 ;
        RECT 120.705 117.455 121.705 117.625 ;
        RECT 119.185 115.200 119.355 117.240 ;
        RECT 120.475 115.200 120.645 117.240 ;
        RECT 121.765 115.200 121.935 117.240 ;
        RECT 119.415 114.815 120.415 114.985 ;
        RECT 120.705 114.815 121.705 114.985 ;
        RECT 122.425 114.200 122.605 118.050 ;
        RECT 126.085 115.925 126.885 115.935 ;
        RECT 118.505 113.990 122.605 114.200 ;
        RECT 118.505 113.980 119.415 113.990 ;
        RECT 118.505 110.140 118.675 113.980 ;
        RECT 119.415 113.395 120.415 113.565 ;
        RECT 120.705 113.395 121.705 113.565 ;
        RECT 119.185 111.140 119.355 113.180 ;
        RECT 120.475 111.140 120.645 113.180 ;
        RECT 121.765 111.140 121.935 113.180 ;
        RECT 119.415 110.755 120.415 110.925 ;
        RECT 120.705 110.755 121.705 110.925 ;
        RECT 122.425 110.140 122.605 113.990 ;
        RECT 122.895 115.755 126.995 115.925 ;
        RECT 122.895 111.865 123.075 115.755 ;
        RECT 123.795 114.930 124.795 115.100 ;
        RECT 125.085 114.930 126.085 115.100 ;
        RECT 123.565 112.675 123.735 114.715 ;
        RECT 124.855 112.675 125.025 114.715 ;
        RECT 126.145 112.675 126.315 114.715 ;
        RECT 123.795 112.290 124.795 112.460 ;
        RECT 125.085 112.290 126.085 112.460 ;
        RECT 126.825 111.865 126.995 115.755 ;
        RECT 122.895 111.655 126.995 111.865 ;
        RECT 127.345 115.755 130.845 115.925 ;
        RECT 127.345 115.745 130.855 115.755 ;
        RECT 127.345 111.865 127.515 115.745 ;
        RECT 130.675 114.645 130.855 115.745 ;
        RECT 127.985 114.455 128.985 114.625 ;
        RECT 129.275 114.455 130.275 114.625 ;
        RECT 127.755 113.245 127.925 114.285 ;
        RECT 129.045 113.245 129.215 114.285 ;
        RECT 130.335 113.245 130.505 114.285 ;
        RECT 127.985 112.905 128.985 113.075 ;
        RECT 129.275 112.905 130.275 113.075 ;
        RECT 130.675 111.865 130.845 114.645 ;
        RECT 127.345 111.655 130.845 111.865 ;
        RECT 118.505 109.930 122.605 110.140 ;
        RECT 118.505 109.920 119.415 109.930 ;
        RECT 118.505 106.080 118.675 109.920 ;
        RECT 119.415 109.335 120.415 109.505 ;
        RECT 120.705 109.335 121.705 109.505 ;
        RECT 119.185 107.080 119.355 109.120 ;
        RECT 120.475 107.080 120.645 109.120 ;
        RECT 121.765 107.080 121.935 109.120 ;
        RECT 119.415 106.695 120.415 106.865 ;
        RECT 120.705 106.695 121.705 106.865 ;
        RECT 122.425 106.080 122.605 109.930 ;
        RECT 126.085 107.825 126.885 107.835 ;
        RECT 118.505 105.870 122.605 106.080 ;
        RECT 118.505 105.860 119.415 105.870 ;
        RECT 118.505 102.020 118.675 105.860 ;
        RECT 119.415 105.275 120.415 105.445 ;
        RECT 120.705 105.275 121.705 105.445 ;
        RECT 119.185 103.020 119.355 105.060 ;
        RECT 120.475 103.020 120.645 105.060 ;
        RECT 121.765 103.020 121.935 105.060 ;
        RECT 119.415 102.635 120.415 102.805 ;
        RECT 120.705 102.635 121.705 102.805 ;
        RECT 122.425 102.020 122.605 105.870 ;
        RECT 118.505 101.810 122.605 102.020 ;
        RECT 118.505 101.800 119.415 101.810 ;
        RECT 118.505 97.920 118.675 101.800 ;
        RECT 119.415 101.215 120.415 101.385 ;
        RECT 120.705 101.215 121.705 101.385 ;
        RECT 119.185 98.960 119.355 101.000 ;
        RECT 120.475 98.960 120.645 101.000 ;
        RECT 121.765 98.960 121.935 101.000 ;
        RECT 119.415 98.575 120.415 98.745 ;
        RECT 120.705 98.575 121.705 98.745 ;
        RECT 122.425 97.920 122.605 101.810 ;
        RECT 118.505 97.750 122.605 97.920 ;
        RECT 122.895 107.655 126.995 107.825 ;
        RECT 122.895 103.775 123.075 107.655 ;
        RECT 123.795 106.830 124.795 107.000 ;
        RECT 125.085 106.830 126.085 107.000 ;
        RECT 123.565 104.575 123.735 106.615 ;
        RECT 124.855 104.575 125.025 106.615 ;
        RECT 126.145 104.575 126.315 106.615 ;
        RECT 123.795 104.190 124.795 104.360 ;
        RECT 125.085 104.190 126.085 104.360 ;
        RECT 126.825 103.785 126.995 107.655 ;
        RECT 126.085 103.775 126.995 103.785 ;
        RECT 122.895 103.555 126.995 103.775 ;
        RECT 122.895 99.725 123.075 103.555 ;
        RECT 123.795 102.780 124.795 102.950 ;
        RECT 125.085 102.780 126.085 102.950 ;
        RECT 123.565 100.525 123.735 102.565 ;
        RECT 124.855 100.525 125.025 102.565 ;
        RECT 126.145 100.525 126.315 102.565 ;
        RECT 123.795 100.140 124.795 100.310 ;
        RECT 125.085 100.140 126.085 100.310 ;
        RECT 126.825 99.735 126.995 103.555 ;
        RECT 126.085 99.725 126.995 99.735 ;
        RECT 122.895 99.505 126.995 99.725 ;
        RECT 118.615 97.740 119.415 97.750 ;
        RECT 95.175 97.015 104.005 97.185 ;
        RECT 107.030 97.075 113.770 97.245 ;
        RECT 97.830 97.010 102.780 97.015 ;
        RECT 94.680 96.570 106.670 96.740 ;
        RECT 94.680 94.810 94.850 96.570 ;
        RECT 95.575 96.000 103.115 96.170 ;
        RECT 95.190 95.440 95.360 95.940 ;
        RECT 103.330 95.440 103.500 95.940 ;
        RECT 95.575 95.210 103.115 95.380 ;
        RECT 103.840 94.810 104.010 96.570 ;
        RECT 104.735 96.000 105.775 96.170 ;
        RECT 104.350 95.440 104.520 95.940 ;
        RECT 105.990 95.440 106.160 95.940 ;
        RECT 104.735 95.210 105.775 95.380 ;
        RECT 106.500 94.810 106.670 96.570 ;
        RECT 94.680 94.640 106.670 94.810 ;
        RECT 107.030 94.815 107.200 97.075 ;
        RECT 107.880 96.505 112.920 96.675 ;
        RECT 107.540 95.445 107.710 96.445 ;
        RECT 113.090 95.445 113.260 96.445 ;
        RECT 107.880 95.215 112.920 95.385 ;
        RECT 113.600 94.815 113.770 97.075 ;
        RECT 107.030 94.645 113.770 94.815 ;
        RECT 122.895 95.675 123.075 99.505 ;
        RECT 123.795 98.730 124.795 98.900 ;
        RECT 125.085 98.730 126.085 98.900 ;
        RECT 123.565 96.475 123.735 98.515 ;
        RECT 124.855 96.475 125.025 98.515 ;
        RECT 126.145 96.475 126.315 98.515 ;
        RECT 123.795 96.090 124.795 96.260 ;
        RECT 125.085 96.090 126.085 96.260 ;
        RECT 126.825 95.685 126.995 99.505 ;
        RECT 126.085 95.675 126.995 95.685 ;
        RECT 122.895 95.455 126.995 95.675 ;
        RECT 108.420 94.640 109.060 94.645 ;
        RECT 109.600 94.640 110.240 94.645 ;
        RECT 111.000 94.640 111.640 94.645 ;
        RECT 112.650 94.640 113.290 94.645 ;
        RECT 72.100 93.840 88.210 94.020 ;
        RECT 72.100 81.180 72.280 93.840 ;
        RECT 73.030 91.610 78.070 91.780 ;
        RECT 82.030 91.610 87.070 91.780 ;
        RECT 72.645 91.050 72.815 91.550 ;
        RECT 78.285 91.050 78.455 91.550 ;
        RECT 81.645 91.050 81.815 91.550 ;
        RECT 87.285 91.050 87.455 91.550 ;
        RECT 73.030 90.820 78.070 90.990 ;
        RECT 82.030 90.820 87.070 90.990 ;
        RECT 73.030 87.110 78.070 87.280 ;
        RECT 82.030 87.110 87.070 87.280 ;
        RECT 72.645 86.550 72.815 87.050 ;
        RECT 78.285 86.550 78.455 87.050 ;
        RECT 81.645 86.550 81.815 87.050 ;
        RECT 87.285 86.550 87.455 87.050 ;
        RECT 73.030 86.320 78.070 86.490 ;
        RECT 82.030 86.320 87.070 86.490 ;
        RECT 73.030 82.610 78.070 82.780 ;
        RECT 82.030 82.610 87.070 82.780 ;
        RECT 72.645 82.050 72.815 82.550 ;
        RECT 78.285 82.050 78.455 82.550 ;
        RECT 81.645 82.050 81.815 82.550 ;
        RECT 87.285 82.050 87.455 82.550 ;
        RECT 73.030 81.820 78.070 81.990 ;
        RECT 82.030 81.820 87.070 81.990 ;
        RECT 88.030 81.180 88.210 93.840 ;
        RECT 88.870 93.870 104.430 94.040 ;
        RECT 88.870 81.350 89.040 93.870 ;
        RECT 90.750 92.090 95.790 92.260 ;
        RECT 97.750 92.090 102.790 92.260 ;
        RECT 90.410 91.030 90.580 92.030 ;
        RECT 95.960 91.030 96.130 92.030 ;
        RECT 97.410 91.030 97.580 92.030 ;
        RECT 102.960 91.030 103.130 92.030 ;
        RECT 90.750 90.800 95.790 90.970 ;
        RECT 97.750 90.800 102.790 90.970 ;
        RECT 90.750 90.090 95.790 90.260 ;
        RECT 97.750 90.090 102.790 90.260 ;
        RECT 90.410 89.030 90.580 90.030 ;
        RECT 95.960 89.030 96.130 90.030 ;
        RECT 97.410 89.030 97.580 90.030 ;
        RECT 102.960 89.030 103.130 90.030 ;
        RECT 90.750 88.800 95.790 88.970 ;
        RECT 97.750 88.800 102.790 88.970 ;
        RECT 90.750 86.090 95.790 86.260 ;
        RECT 97.750 86.090 102.790 86.260 ;
        RECT 90.410 85.030 90.580 86.030 ;
        RECT 95.960 85.030 96.130 86.030 ;
        RECT 97.410 85.030 97.580 86.030 ;
        RECT 102.960 85.030 103.130 86.030 ;
        RECT 90.750 84.800 95.790 84.970 ;
        RECT 97.750 84.800 102.790 84.970 ;
        RECT 90.750 84.090 95.790 84.260 ;
        RECT 97.750 84.090 102.790 84.260 ;
        RECT 90.410 83.030 90.580 84.030 ;
        RECT 95.960 83.030 96.130 84.030 ;
        RECT 97.410 83.030 97.580 84.030 ;
        RECT 102.960 83.030 103.130 84.030 ;
        RECT 90.750 82.800 95.790 82.970 ;
        RECT 97.750 82.800 102.790 82.970 ;
        RECT 104.260 81.350 104.430 93.870 ;
        RECT 88.870 81.180 104.430 81.350 ;
        RECT 105.290 94.010 113.690 94.180 ;
        RECT 105.290 81.210 105.460 94.010 ;
        RECT 106.210 93.400 111.250 93.570 ;
        RECT 105.870 92.340 106.040 93.340 ;
        RECT 111.420 92.340 111.590 93.340 ;
        RECT 106.210 92.110 111.250 92.280 ;
        RECT 105.870 91.050 106.040 92.050 ;
        RECT 111.420 91.050 111.590 92.050 ;
        RECT 106.210 90.820 111.250 90.990 ;
        RECT 105.870 89.760 106.040 90.760 ;
        RECT 111.420 89.760 111.590 90.760 ;
        RECT 106.210 89.530 111.250 89.700 ;
        RECT 105.870 88.470 106.040 89.470 ;
        RECT 111.420 88.470 111.590 89.470 ;
        RECT 106.210 88.240 111.250 88.410 ;
        RECT 105.870 87.180 106.040 88.180 ;
        RECT 111.420 87.180 111.590 88.180 ;
        RECT 106.210 86.950 111.250 87.120 ;
        RECT 105.870 85.890 106.040 86.890 ;
        RECT 111.420 85.890 111.590 86.890 ;
        RECT 106.210 85.660 111.250 85.830 ;
        RECT 105.870 84.600 106.040 85.600 ;
        RECT 111.420 84.600 111.590 85.600 ;
        RECT 106.210 84.370 111.250 84.540 ;
        RECT 105.870 83.310 106.040 84.310 ;
        RECT 111.420 83.310 111.590 84.310 ;
        RECT 106.210 83.080 111.250 83.250 ;
        RECT 113.520 81.210 113.690 94.010 ;
        RECT 114.655 93.690 118.155 93.900 ;
        RECT 114.655 90.910 114.825 93.690 ;
        RECT 115.225 92.480 116.225 92.650 ;
        RECT 116.515 92.480 117.515 92.650 ;
        RECT 114.995 91.270 115.165 92.310 ;
        RECT 116.285 91.270 116.455 92.310 ;
        RECT 117.575 91.270 117.745 92.310 ;
        RECT 115.225 90.930 116.225 91.100 ;
        RECT 116.515 90.930 117.515 91.100 ;
        RECT 114.645 89.840 114.825 90.910 ;
        RECT 117.985 89.840 118.155 93.690 ;
        RECT 114.645 89.800 118.155 89.840 ;
        RECT 114.655 89.630 118.155 89.800 ;
        RECT 114.655 86.850 114.825 89.630 ;
        RECT 115.225 88.420 116.225 88.590 ;
        RECT 116.515 88.420 117.515 88.590 ;
        RECT 114.995 87.210 115.165 88.250 ;
        RECT 116.285 87.210 116.455 88.250 ;
        RECT 117.575 87.210 117.745 88.250 ;
        RECT 115.225 86.870 116.225 87.040 ;
        RECT 116.515 86.870 117.515 87.040 ;
        RECT 114.645 85.780 114.825 86.850 ;
        RECT 117.985 85.780 118.155 89.630 ;
        RECT 114.645 85.740 118.155 85.780 ;
        RECT 114.655 85.570 118.155 85.740 ;
        RECT 114.655 82.790 114.825 85.570 ;
        RECT 115.225 84.360 116.225 84.530 ;
        RECT 116.515 84.360 117.515 84.530 ;
        RECT 114.995 83.150 115.165 84.190 ;
        RECT 116.285 83.150 116.455 84.190 ;
        RECT 117.575 83.150 117.745 84.190 ;
        RECT 115.225 82.810 116.225 82.980 ;
        RECT 116.515 82.810 117.515 82.980 ;
        RECT 114.645 81.720 114.825 82.790 ;
        RECT 117.985 81.720 118.155 85.570 ;
        RECT 114.645 81.680 118.155 81.720 ;
        RECT 72.100 81.000 88.210 81.180 ;
        RECT 105.290 81.040 113.690 81.210 ;
        RECT 114.655 81.510 118.155 81.680 ;
        RECT 63.350 80.640 70.660 80.820 ;
        RECT 55.770 77.260 62.540 77.430 ;
        RECT 14.350 74.830 17.780 75.000 ;
        RECT 14.350 44.570 14.520 74.830 ;
        RECT 15.000 74.100 15.500 74.270 ;
        RECT 15.080 72.285 15.420 74.100 ;
        RECT 15.080 45.300 15.420 47.115 ;
        RECT 15.000 45.130 15.500 45.300 ;
        RECT 15.980 44.570 16.150 74.830 ;
        RECT 16.630 74.100 17.130 74.270 ;
        RECT 16.710 72.285 17.050 74.100 ;
        RECT 16.710 45.300 17.050 47.115 ;
        RECT 16.630 45.130 17.130 45.300 ;
        RECT 17.610 44.570 17.780 74.830 ;
        RECT 14.350 44.400 17.780 44.570 ;
        RECT 20.090 74.830 26.780 75.000 ;
        RECT 20.090 44.570 20.260 74.830 ;
        RECT 20.740 74.100 21.240 74.270 ;
        RECT 20.820 72.285 21.160 74.100 ;
        RECT 20.820 45.300 21.160 47.115 ;
        RECT 20.740 45.130 21.240 45.300 ;
        RECT 21.720 44.570 21.890 74.830 ;
        RECT 22.370 74.100 22.870 74.270 ;
        RECT 22.450 72.285 22.790 74.100 ;
        RECT 22.450 45.300 22.790 47.115 ;
        RECT 22.370 45.130 22.870 45.300 ;
        RECT 23.350 44.570 23.520 74.830 ;
        RECT 24.000 74.100 24.500 74.270 ;
        RECT 24.080 72.285 24.420 74.100 ;
        RECT 24.080 45.300 24.420 47.115 ;
        RECT 24.000 45.130 24.500 45.300 ;
        RECT 24.980 44.570 25.150 74.830 ;
        RECT 25.630 74.100 26.130 74.270 ;
        RECT 25.710 72.285 26.050 74.100 ;
        RECT 25.710 45.300 26.050 47.115 ;
        RECT 25.630 45.130 26.130 45.300 ;
        RECT 26.610 44.570 26.780 74.830 ;
        RECT 55.770 64.500 55.940 77.260 ;
        RECT 56.620 76.310 61.660 76.480 ;
        RECT 56.235 75.750 56.405 76.250 ;
        RECT 61.875 75.750 62.045 76.250 ;
        RECT 56.620 75.520 61.660 75.690 ;
        RECT 56.235 74.960 56.405 75.460 ;
        RECT 61.875 74.960 62.045 75.460 ;
        RECT 56.620 74.730 61.660 74.900 ;
        RECT 56.235 74.170 56.405 74.670 ;
        RECT 61.875 74.170 62.045 74.670 ;
        RECT 56.620 73.940 61.660 74.110 ;
        RECT 56.235 73.380 56.405 73.880 ;
        RECT 61.875 73.380 62.045 73.880 ;
        RECT 56.620 73.150 61.660 73.320 ;
        RECT 56.235 72.590 56.405 73.090 ;
        RECT 61.875 72.590 62.045 73.090 ;
        RECT 56.620 72.360 61.660 72.530 ;
        RECT 56.235 71.800 56.405 72.300 ;
        RECT 61.875 71.800 62.045 72.300 ;
        RECT 56.620 71.570 61.660 71.740 ;
        RECT 56.235 71.010 56.405 71.510 ;
        RECT 61.875 71.010 62.045 71.510 ;
        RECT 56.620 70.780 61.660 70.950 ;
        RECT 56.235 70.220 56.405 70.720 ;
        RECT 61.875 70.220 62.045 70.720 ;
        RECT 56.620 69.990 61.660 70.160 ;
        RECT 56.235 69.430 56.405 69.930 ;
        RECT 61.875 69.430 62.045 69.930 ;
        RECT 56.620 69.200 61.660 69.370 ;
        RECT 56.235 68.640 56.405 69.140 ;
        RECT 61.875 68.640 62.045 69.140 ;
        RECT 56.620 68.410 61.660 68.580 ;
        RECT 56.235 67.850 56.405 68.350 ;
        RECT 61.875 67.850 62.045 68.350 ;
        RECT 56.620 67.620 61.660 67.790 ;
        RECT 56.235 67.060 56.405 67.560 ;
        RECT 61.875 67.060 62.045 67.560 ;
        RECT 56.620 66.830 61.660 67.000 ;
        RECT 56.235 66.270 56.405 66.770 ;
        RECT 61.875 66.270 62.045 66.770 ;
        RECT 56.620 66.040 61.660 66.210 ;
        RECT 56.235 65.480 56.405 65.980 ;
        RECT 61.875 65.480 62.045 65.980 ;
        RECT 56.620 65.250 61.660 65.420 ;
        RECT 62.370 64.500 62.540 77.260 ;
        RECT 55.770 64.330 62.540 64.500 ;
        RECT 63.350 64.510 63.520 80.640 ;
        RECT 64.680 80.080 69.720 80.250 ;
        RECT 64.340 79.520 64.510 80.020 ;
        RECT 69.890 79.520 70.060 80.020 ;
        RECT 64.680 79.290 69.720 79.460 ;
        RECT 64.340 78.730 64.510 79.230 ;
        RECT 69.890 78.730 70.060 79.230 ;
        RECT 64.680 78.500 69.720 78.670 ;
        RECT 64.340 77.940 64.510 78.440 ;
        RECT 69.890 77.940 70.060 78.440 ;
        RECT 64.680 77.710 69.720 77.880 ;
        RECT 64.340 77.150 64.510 77.650 ;
        RECT 69.890 77.150 70.060 77.650 ;
        RECT 64.680 76.920 69.720 77.090 ;
        RECT 64.340 76.360 64.510 76.860 ;
        RECT 69.890 76.360 70.060 76.860 ;
        RECT 64.680 76.130 69.720 76.300 ;
        RECT 64.340 75.570 64.510 76.070 ;
        RECT 69.890 75.570 70.060 76.070 ;
        RECT 64.680 75.340 69.720 75.510 ;
        RECT 64.340 74.780 64.510 75.280 ;
        RECT 69.890 74.780 70.060 75.280 ;
        RECT 64.680 74.550 69.720 74.720 ;
        RECT 64.340 73.990 64.510 74.490 ;
        RECT 69.890 73.990 70.060 74.490 ;
        RECT 64.680 73.760 69.720 73.930 ;
        RECT 64.340 73.200 64.510 73.700 ;
        RECT 69.890 73.200 70.060 73.700 ;
        RECT 64.680 72.970 69.720 73.140 ;
        RECT 64.340 72.410 64.510 72.910 ;
        RECT 69.890 72.410 70.060 72.910 ;
        RECT 64.680 72.180 69.720 72.350 ;
        RECT 64.340 71.620 64.510 72.120 ;
        RECT 69.890 71.620 70.060 72.120 ;
        RECT 64.680 71.390 69.720 71.560 ;
        RECT 64.340 70.830 64.510 71.330 ;
        RECT 69.890 70.830 70.060 71.330 ;
        RECT 64.680 70.600 69.720 70.770 ;
        RECT 64.340 70.040 64.510 70.540 ;
        RECT 69.890 70.040 70.060 70.540 ;
        RECT 64.680 69.810 69.720 69.980 ;
        RECT 64.340 69.250 64.510 69.750 ;
        RECT 69.890 69.250 70.060 69.750 ;
        RECT 64.680 69.020 69.720 69.190 ;
        RECT 64.340 68.460 64.510 68.960 ;
        RECT 69.890 68.460 70.060 68.960 ;
        RECT 64.680 68.230 69.720 68.400 ;
        RECT 64.340 67.670 64.510 68.170 ;
        RECT 69.890 67.670 70.060 68.170 ;
        RECT 64.680 67.440 69.720 67.610 ;
        RECT 64.340 66.880 64.510 67.380 ;
        RECT 69.890 66.880 70.060 67.380 ;
        RECT 64.680 66.650 69.720 66.820 ;
        RECT 64.340 66.090 64.510 66.590 ;
        RECT 69.890 66.090 70.060 66.590 ;
        RECT 64.680 65.860 69.720 66.030 ;
        RECT 64.340 65.300 64.510 65.800 ;
        RECT 69.890 65.300 70.060 65.800 ;
        RECT 64.680 65.070 69.720 65.240 ;
        RECT 70.490 64.510 70.660 80.640 ;
        RECT 72.100 80.530 88.210 80.710 ;
        RECT 72.100 67.870 72.280 80.530 ;
        RECT 73.030 79.720 78.070 79.890 ;
        RECT 82.030 79.720 87.070 79.890 ;
        RECT 72.645 79.160 72.815 79.660 ;
        RECT 78.285 79.160 78.455 79.660 ;
        RECT 81.645 79.160 81.815 79.660 ;
        RECT 87.285 79.160 87.455 79.660 ;
        RECT 73.030 78.930 78.070 79.100 ;
        RECT 82.030 78.930 87.070 79.100 ;
        RECT 73.030 75.220 78.070 75.390 ;
        RECT 82.030 75.220 87.070 75.390 ;
        RECT 72.645 74.660 72.815 75.160 ;
        RECT 78.285 74.660 78.455 75.160 ;
        RECT 81.645 74.660 81.815 75.160 ;
        RECT 87.285 74.660 87.455 75.160 ;
        RECT 73.030 74.430 78.070 74.600 ;
        RECT 82.030 74.430 87.070 74.600 ;
        RECT 73.030 70.720 78.070 70.890 ;
        RECT 82.030 70.720 87.070 70.890 ;
        RECT 72.645 70.160 72.815 70.660 ;
        RECT 78.285 70.160 78.455 70.660 ;
        RECT 81.645 70.160 81.815 70.660 ;
        RECT 87.285 70.160 87.455 70.660 ;
        RECT 73.030 69.930 78.070 70.100 ;
        RECT 82.030 69.930 87.070 70.100 ;
        RECT 88.030 67.870 88.210 80.530 ;
        RECT 72.100 67.690 88.210 67.870 ;
        RECT 88.870 80.360 104.430 80.530 ;
        RECT 88.870 67.840 89.040 80.360 ;
        RECT 90.750 78.740 95.790 78.910 ;
        RECT 97.750 78.740 102.790 78.910 ;
        RECT 90.410 77.680 90.580 78.680 ;
        RECT 95.960 77.680 96.130 78.680 ;
        RECT 97.410 77.680 97.580 78.680 ;
        RECT 102.960 77.680 103.130 78.680 ;
        RECT 90.750 77.450 95.790 77.620 ;
        RECT 97.750 77.450 102.790 77.620 ;
        RECT 90.750 76.740 95.790 76.910 ;
        RECT 97.750 76.740 102.790 76.910 ;
        RECT 90.410 75.680 90.580 76.680 ;
        RECT 95.960 75.680 96.130 76.680 ;
        RECT 97.410 75.680 97.580 76.680 ;
        RECT 102.960 75.680 103.130 76.680 ;
        RECT 90.750 75.450 95.790 75.620 ;
        RECT 97.750 75.450 102.790 75.620 ;
        RECT 90.750 72.740 95.790 72.910 ;
        RECT 97.750 72.740 102.790 72.910 ;
        RECT 90.410 71.680 90.580 72.680 ;
        RECT 95.960 71.680 96.130 72.680 ;
        RECT 97.410 71.680 97.580 72.680 ;
        RECT 102.960 71.680 103.130 72.680 ;
        RECT 90.750 71.450 95.790 71.620 ;
        RECT 97.750 71.450 102.790 71.620 ;
        RECT 90.750 70.740 95.790 70.910 ;
        RECT 97.750 70.740 102.790 70.910 ;
        RECT 90.410 69.680 90.580 70.680 ;
        RECT 95.960 69.680 96.130 70.680 ;
        RECT 97.410 69.680 97.580 70.680 ;
        RECT 102.960 69.680 103.130 70.680 ;
        RECT 90.750 69.450 95.790 69.620 ;
        RECT 97.750 69.450 102.790 69.620 ;
        RECT 104.260 67.840 104.430 80.360 ;
        RECT 88.870 67.670 104.430 67.840 ;
        RECT 105.290 80.500 113.690 80.670 ;
        RECT 105.290 67.700 105.460 80.500 ;
        RECT 106.210 78.460 111.250 78.630 ;
        RECT 105.870 77.400 106.040 78.400 ;
        RECT 111.420 77.400 111.590 78.400 ;
        RECT 106.210 77.170 111.250 77.340 ;
        RECT 105.870 76.110 106.040 77.110 ;
        RECT 111.420 76.110 111.590 77.110 ;
        RECT 106.210 75.880 111.250 76.050 ;
        RECT 105.870 74.820 106.040 75.820 ;
        RECT 111.420 74.820 111.590 75.820 ;
        RECT 106.210 74.590 111.250 74.760 ;
        RECT 105.870 73.530 106.040 74.530 ;
        RECT 111.420 73.530 111.590 74.530 ;
        RECT 106.210 73.300 111.250 73.470 ;
        RECT 105.870 72.240 106.040 73.240 ;
        RECT 111.420 72.240 111.590 73.240 ;
        RECT 106.210 72.010 111.250 72.180 ;
        RECT 105.870 70.950 106.040 71.950 ;
        RECT 111.420 70.950 111.590 71.950 ;
        RECT 106.210 70.720 111.250 70.890 ;
        RECT 105.870 69.660 106.040 70.660 ;
        RECT 111.420 69.660 111.590 70.660 ;
        RECT 106.210 69.430 111.250 69.600 ;
        RECT 105.870 68.370 106.040 69.370 ;
        RECT 111.420 68.370 111.590 69.370 ;
        RECT 106.210 68.140 111.250 68.310 ;
        RECT 113.520 67.700 113.690 80.500 ;
        RECT 114.655 78.730 114.825 81.510 ;
        RECT 115.225 80.300 116.225 80.470 ;
        RECT 116.515 80.300 117.515 80.470 ;
        RECT 114.995 79.090 115.165 80.130 ;
        RECT 116.285 79.090 116.455 80.130 ;
        RECT 117.575 79.090 117.745 80.130 ;
        RECT 115.225 78.750 116.225 78.920 ;
        RECT 116.515 78.750 117.515 78.920 ;
        RECT 114.645 77.660 114.825 78.730 ;
        RECT 117.985 77.660 118.155 81.510 ;
        RECT 114.645 77.620 118.155 77.660 ;
        RECT 114.655 77.450 118.155 77.620 ;
        RECT 114.655 74.670 114.825 77.450 ;
        RECT 115.225 76.240 116.225 76.410 ;
        RECT 116.515 76.240 117.515 76.410 ;
        RECT 114.995 75.030 115.165 76.070 ;
        RECT 116.285 75.030 116.455 76.070 ;
        RECT 117.575 75.030 117.745 76.070 ;
        RECT 115.225 74.690 116.225 74.860 ;
        RECT 116.515 74.690 117.515 74.860 ;
        RECT 114.645 73.570 114.825 74.670 ;
        RECT 117.985 73.570 118.155 77.450 ;
        RECT 114.645 73.560 118.155 73.570 ;
        RECT 114.655 73.390 118.155 73.560 ;
        RECT 118.505 93.690 122.605 93.900 ;
        RECT 118.505 89.840 118.675 93.690 ;
        RECT 119.415 93.095 120.415 93.265 ;
        RECT 120.705 93.095 121.705 93.265 ;
        RECT 119.185 90.840 119.355 92.880 ;
        RECT 120.475 90.840 120.645 92.880 ;
        RECT 121.765 90.840 121.935 92.880 ;
        RECT 119.415 90.455 120.415 90.625 ;
        RECT 120.705 90.455 121.705 90.625 ;
        RECT 122.425 89.840 122.605 93.690 ;
        RECT 118.505 89.630 122.605 89.840 ;
        RECT 118.505 89.620 119.415 89.630 ;
        RECT 118.505 85.780 118.675 89.620 ;
        RECT 119.415 89.035 120.415 89.205 ;
        RECT 120.705 89.035 121.705 89.205 ;
        RECT 119.185 86.780 119.355 88.820 ;
        RECT 120.475 86.780 120.645 88.820 ;
        RECT 121.765 86.780 121.935 88.820 ;
        RECT 119.415 86.395 120.415 86.565 ;
        RECT 120.705 86.395 121.705 86.565 ;
        RECT 122.425 85.780 122.605 89.630 ;
        RECT 118.505 85.570 122.605 85.780 ;
        RECT 118.505 85.560 119.415 85.570 ;
        RECT 118.505 81.720 118.675 85.560 ;
        RECT 119.415 84.975 120.415 85.145 ;
        RECT 120.705 84.975 121.705 85.145 ;
        RECT 119.185 82.720 119.355 84.760 ;
        RECT 120.475 82.720 120.645 84.760 ;
        RECT 121.765 82.720 121.935 84.760 ;
        RECT 119.415 82.335 120.415 82.505 ;
        RECT 120.705 82.335 121.705 82.505 ;
        RECT 122.425 81.720 122.605 85.570 ;
        RECT 118.505 81.510 122.605 81.720 ;
        RECT 118.505 81.500 119.415 81.510 ;
        RECT 118.505 77.660 118.675 81.500 ;
        RECT 119.415 80.915 120.415 81.085 ;
        RECT 120.705 80.915 121.705 81.085 ;
        RECT 119.185 78.660 119.355 80.700 ;
        RECT 120.475 78.660 120.645 80.700 ;
        RECT 121.765 78.660 121.935 80.700 ;
        RECT 119.415 78.275 120.415 78.445 ;
        RECT 120.705 78.275 121.705 78.445 ;
        RECT 122.425 77.660 122.605 81.510 ;
        RECT 118.505 77.450 122.605 77.660 ;
        RECT 118.505 77.440 119.415 77.450 ;
        RECT 118.505 73.560 118.675 77.440 ;
        RECT 119.415 76.855 120.415 77.025 ;
        RECT 120.705 76.855 121.705 77.025 ;
        RECT 119.185 74.600 119.355 76.640 ;
        RECT 120.475 74.600 120.645 76.640 ;
        RECT 121.765 74.600 121.935 76.640 ;
        RECT 119.415 74.215 120.415 74.385 ;
        RECT 120.705 74.215 121.705 74.385 ;
        RECT 122.425 73.560 122.605 77.450 ;
        RECT 118.505 73.390 122.605 73.560 ;
        RECT 122.895 91.625 123.075 95.455 ;
        RECT 123.795 94.680 124.795 94.850 ;
        RECT 125.085 94.680 126.085 94.850 ;
        RECT 123.565 92.425 123.735 94.465 ;
        RECT 124.855 92.425 125.025 94.465 ;
        RECT 126.145 92.425 126.315 94.465 ;
        RECT 123.795 92.040 124.795 92.210 ;
        RECT 125.085 92.040 126.085 92.210 ;
        RECT 126.825 91.635 126.995 95.455 ;
        RECT 126.085 91.625 126.995 91.635 ;
        RECT 122.895 91.405 126.995 91.625 ;
        RECT 122.895 87.575 123.075 91.405 ;
        RECT 123.795 90.630 124.795 90.800 ;
        RECT 125.085 90.630 126.085 90.800 ;
        RECT 123.565 88.375 123.735 90.415 ;
        RECT 124.855 88.375 125.025 90.415 ;
        RECT 126.145 88.375 126.315 90.415 ;
        RECT 123.795 87.990 124.795 88.160 ;
        RECT 125.085 87.990 126.085 88.160 ;
        RECT 126.825 87.585 126.995 91.405 ;
        RECT 126.085 87.575 126.995 87.585 ;
        RECT 122.895 87.355 126.995 87.575 ;
        RECT 122.895 83.525 123.075 87.355 ;
        RECT 123.795 86.580 124.795 86.750 ;
        RECT 125.085 86.580 126.085 86.750 ;
        RECT 123.565 84.325 123.735 86.365 ;
        RECT 124.855 84.325 125.025 86.365 ;
        RECT 126.145 84.325 126.315 86.365 ;
        RECT 123.795 83.940 124.795 84.110 ;
        RECT 125.085 83.940 126.085 84.110 ;
        RECT 126.825 83.535 126.995 87.355 ;
        RECT 126.085 83.525 126.995 83.535 ;
        RECT 122.895 83.305 126.995 83.525 ;
        RECT 122.895 79.475 123.075 83.305 ;
        RECT 123.795 82.530 124.795 82.700 ;
        RECT 125.085 82.530 126.085 82.700 ;
        RECT 123.565 80.275 123.735 82.315 ;
        RECT 124.855 80.275 125.025 82.315 ;
        RECT 126.145 80.275 126.315 82.315 ;
        RECT 123.795 79.890 124.795 80.060 ;
        RECT 125.085 79.890 126.085 80.060 ;
        RECT 126.825 79.485 126.995 83.305 ;
        RECT 126.085 79.475 126.995 79.485 ;
        RECT 122.895 79.255 126.995 79.475 ;
        RECT 122.895 75.425 123.075 79.255 ;
        RECT 123.795 78.480 124.795 78.650 ;
        RECT 125.085 78.480 126.085 78.650 ;
        RECT 123.565 76.225 123.735 78.265 ;
        RECT 124.855 76.225 125.025 78.265 ;
        RECT 126.145 76.225 126.315 78.265 ;
        RECT 123.795 75.840 124.795 76.010 ;
        RECT 125.085 75.840 126.085 76.010 ;
        RECT 126.825 75.435 126.995 79.255 ;
        RECT 126.085 75.425 126.995 75.435 ;
        RECT 122.895 75.205 126.995 75.425 ;
        RECT 118.615 73.380 119.415 73.390 ;
        RECT 105.290 67.530 113.690 67.700 ;
        RECT 122.895 71.365 123.075 75.205 ;
        RECT 123.795 74.430 124.795 74.600 ;
        RECT 125.085 74.430 126.085 74.600 ;
        RECT 123.565 72.175 123.735 74.215 ;
        RECT 124.855 72.175 125.025 74.215 ;
        RECT 126.145 72.175 126.315 74.215 ;
        RECT 123.795 71.790 124.795 71.960 ;
        RECT 125.085 71.790 126.085 71.960 ;
        RECT 126.825 71.365 126.995 75.205 ;
        RECT 122.895 71.155 126.995 71.365 ;
        RECT 122.895 67.280 123.075 71.155 ;
        RECT 123.795 70.345 124.795 70.515 ;
        RECT 125.085 70.345 126.085 70.515 ;
        RECT 123.565 68.090 123.735 70.130 ;
        RECT 124.855 68.090 125.025 70.130 ;
        RECT 126.145 68.090 126.315 70.130 ;
        RECT 123.795 67.705 124.795 67.875 ;
        RECT 125.085 67.705 126.085 67.875 ;
        RECT 126.825 67.280 126.995 71.155 ;
        RECT 94.680 66.900 106.670 67.070 ;
        RECT 108.420 67.065 109.060 67.070 ;
        RECT 109.600 67.065 110.240 67.070 ;
        RECT 111.000 67.065 111.640 67.070 ;
        RECT 112.650 67.065 113.290 67.070 ;
        RECT 94.680 65.140 94.850 66.900 ;
        RECT 95.575 66.330 103.115 66.500 ;
        RECT 95.190 65.770 95.360 66.270 ;
        RECT 103.330 65.770 103.500 66.270 ;
        RECT 95.575 65.540 103.115 65.710 ;
        RECT 103.840 65.140 104.010 66.900 ;
        RECT 104.735 66.330 105.775 66.500 ;
        RECT 104.350 65.770 104.520 66.270 ;
        RECT 105.990 65.770 106.160 66.270 ;
        RECT 104.735 65.540 105.775 65.710 ;
        RECT 106.500 65.140 106.670 66.900 ;
        RECT 94.680 64.970 106.670 65.140 ;
        RECT 107.030 66.895 113.770 67.065 ;
        RECT 97.830 64.695 102.780 64.700 ;
        RECT 63.350 64.330 70.660 64.510 ;
        RECT 95.175 64.525 104.005 64.695 ;
        RECT 95.175 64.220 95.345 64.525 ;
        RECT 52.175 63.515 61.005 63.685 ;
        RECT 52.175 63.200 52.345 63.515 ;
        RECT 52.175 62.060 52.350 63.200 ;
        RECT 53.070 62.945 60.110 63.115 ;
        RECT 52.685 62.385 52.855 62.885 ;
        RECT 60.325 62.385 60.495 62.885 ;
        RECT 53.070 62.155 60.110 62.325 ;
        RECT 52.175 61.755 52.345 62.060 ;
        RECT 60.835 61.755 61.005 63.515 ;
        RECT 52.175 61.585 61.005 61.755 ;
        RECT 52.175 61.270 52.345 61.585 ;
        RECT 52.175 60.130 52.350 61.270 ;
        RECT 53.070 61.015 60.110 61.185 ;
        RECT 52.685 60.455 52.855 60.955 ;
        RECT 60.325 60.455 60.495 60.955 ;
        RECT 53.070 60.225 60.110 60.395 ;
        RECT 52.175 59.825 52.345 60.130 ;
        RECT 60.835 59.825 61.005 61.585 ;
        RECT 95.175 63.080 95.350 64.220 ;
        RECT 96.070 63.955 103.110 64.125 ;
        RECT 95.685 63.395 95.855 63.895 ;
        RECT 103.325 63.395 103.495 63.895 ;
        RECT 96.070 63.165 103.110 63.335 ;
        RECT 95.175 62.765 95.345 63.080 ;
        RECT 103.835 62.765 104.005 64.525 ;
        RECT 107.030 64.635 107.200 66.895 ;
        RECT 107.880 66.325 112.920 66.495 ;
        RECT 107.540 65.265 107.710 66.265 ;
        RECT 113.090 65.265 113.260 66.265 ;
        RECT 107.880 65.035 112.920 65.205 ;
        RECT 113.600 64.635 113.770 66.895 ;
        RECT 107.030 64.465 113.770 64.635 ;
        RECT 122.895 67.045 126.995 67.280 ;
        RECT 122.895 63.155 123.075 67.045 ;
        RECT 123.795 66.220 124.795 66.390 ;
        RECT 125.085 66.220 126.085 66.390 ;
        RECT 123.565 63.965 123.735 66.005 ;
        RECT 124.855 63.965 125.025 66.005 ;
        RECT 126.145 63.965 126.315 66.005 ;
        RECT 123.795 63.580 124.795 63.750 ;
        RECT 125.085 63.580 126.085 63.750 ;
        RECT 126.825 63.155 126.995 67.045 ;
        RECT 122.895 62.945 126.995 63.155 ;
        RECT 127.345 107.655 130.845 107.825 ;
        RECT 127.345 107.645 130.855 107.655 ;
        RECT 127.345 103.775 127.515 107.645 ;
        RECT 130.675 106.545 130.855 107.645 ;
        RECT 127.985 106.355 128.985 106.525 ;
        RECT 129.275 106.355 130.275 106.525 ;
        RECT 127.755 105.145 127.925 106.185 ;
        RECT 129.045 105.145 129.215 106.185 ;
        RECT 130.335 105.145 130.505 106.185 ;
        RECT 127.985 104.805 128.985 104.975 ;
        RECT 129.275 104.805 130.275 104.975 ;
        RECT 130.675 103.775 130.845 106.545 ;
        RECT 127.345 103.605 130.845 103.775 ;
        RECT 127.345 103.555 130.855 103.605 ;
        RECT 127.345 99.725 127.515 103.555 ;
        RECT 130.675 102.495 130.855 103.555 ;
        RECT 127.985 102.305 128.985 102.475 ;
        RECT 129.275 102.305 130.275 102.475 ;
        RECT 127.755 101.095 127.925 102.135 ;
        RECT 129.045 101.095 129.215 102.135 ;
        RECT 130.335 101.095 130.505 102.135 ;
        RECT 127.985 100.755 128.985 100.925 ;
        RECT 129.275 100.755 130.275 100.925 ;
        RECT 130.675 99.725 130.845 102.495 ;
        RECT 127.345 99.555 130.845 99.725 ;
        RECT 127.345 99.505 130.855 99.555 ;
        RECT 127.345 95.675 127.515 99.505 ;
        RECT 130.675 98.445 130.855 99.505 ;
        RECT 127.985 98.255 128.985 98.425 ;
        RECT 129.275 98.255 130.275 98.425 ;
        RECT 127.755 97.045 127.925 98.085 ;
        RECT 129.045 97.045 129.215 98.085 ;
        RECT 130.335 97.045 130.505 98.085 ;
        RECT 127.985 96.705 128.985 96.875 ;
        RECT 129.275 96.705 130.275 96.875 ;
        RECT 130.675 95.675 130.845 98.445 ;
        RECT 127.345 95.505 130.845 95.675 ;
        RECT 127.345 95.455 130.855 95.505 ;
        RECT 127.345 91.625 127.515 95.455 ;
        RECT 130.675 94.395 130.855 95.455 ;
        RECT 127.985 94.205 128.985 94.375 ;
        RECT 129.275 94.205 130.275 94.375 ;
        RECT 127.755 92.995 127.925 94.035 ;
        RECT 129.045 92.995 129.215 94.035 ;
        RECT 130.335 92.995 130.505 94.035 ;
        RECT 127.985 92.655 128.985 92.825 ;
        RECT 129.275 92.655 130.275 92.825 ;
        RECT 130.675 91.625 130.845 94.395 ;
        RECT 127.345 91.455 130.845 91.625 ;
        RECT 127.345 91.405 130.855 91.455 ;
        RECT 127.345 87.575 127.515 91.405 ;
        RECT 130.675 90.345 130.855 91.405 ;
        RECT 127.985 90.155 128.985 90.325 ;
        RECT 129.275 90.155 130.275 90.325 ;
        RECT 127.755 88.945 127.925 89.985 ;
        RECT 129.045 88.945 129.215 89.985 ;
        RECT 130.335 88.945 130.505 89.985 ;
        RECT 127.985 88.605 128.985 88.775 ;
        RECT 129.275 88.605 130.275 88.775 ;
        RECT 130.675 87.575 130.845 90.345 ;
        RECT 127.345 87.405 130.845 87.575 ;
        RECT 127.345 87.355 130.855 87.405 ;
        RECT 127.345 83.525 127.515 87.355 ;
        RECT 130.675 86.295 130.855 87.355 ;
        RECT 127.985 86.105 128.985 86.275 ;
        RECT 129.275 86.105 130.275 86.275 ;
        RECT 127.755 84.895 127.925 85.935 ;
        RECT 129.045 84.895 129.215 85.935 ;
        RECT 130.335 84.895 130.505 85.935 ;
        RECT 127.985 84.555 128.985 84.725 ;
        RECT 129.275 84.555 130.275 84.725 ;
        RECT 130.675 83.525 130.845 86.295 ;
        RECT 127.345 83.355 130.845 83.525 ;
        RECT 127.345 83.305 130.855 83.355 ;
        RECT 127.345 79.475 127.515 83.305 ;
        RECT 130.675 82.245 130.855 83.305 ;
        RECT 127.985 82.055 128.985 82.225 ;
        RECT 129.275 82.055 130.275 82.225 ;
        RECT 127.755 80.845 127.925 81.885 ;
        RECT 129.045 80.845 129.215 81.885 ;
        RECT 130.335 80.845 130.505 81.885 ;
        RECT 127.985 80.505 128.985 80.675 ;
        RECT 129.275 80.505 130.275 80.675 ;
        RECT 130.675 79.475 130.845 82.245 ;
        RECT 127.345 79.305 130.845 79.475 ;
        RECT 127.345 79.255 130.855 79.305 ;
        RECT 127.345 75.425 127.515 79.255 ;
        RECT 130.675 78.195 130.855 79.255 ;
        RECT 127.985 78.005 128.985 78.175 ;
        RECT 129.275 78.005 130.275 78.175 ;
        RECT 127.755 76.795 127.925 77.835 ;
        RECT 129.045 76.795 129.215 77.835 ;
        RECT 130.335 76.795 130.505 77.835 ;
        RECT 127.985 76.455 128.985 76.625 ;
        RECT 129.275 76.455 130.275 76.625 ;
        RECT 130.675 75.425 130.845 78.195 ;
        RECT 127.345 75.255 130.845 75.425 ;
        RECT 127.345 75.205 130.855 75.255 ;
        RECT 127.345 71.365 127.515 75.205 ;
        RECT 130.675 74.145 130.855 75.205 ;
        RECT 127.985 73.955 128.985 74.125 ;
        RECT 129.275 73.955 130.275 74.125 ;
        RECT 127.755 72.745 127.925 73.785 ;
        RECT 129.045 72.745 129.215 73.785 ;
        RECT 130.335 72.745 130.505 73.785 ;
        RECT 127.985 72.405 128.985 72.575 ;
        RECT 129.275 72.405 130.275 72.575 ;
        RECT 130.675 71.365 130.845 74.145 ;
        RECT 127.345 71.170 130.845 71.365 ;
        RECT 127.345 71.155 130.855 71.170 ;
        RECT 127.345 67.280 127.515 71.155 ;
        RECT 130.675 70.060 130.855 71.155 ;
        RECT 127.985 69.870 128.985 70.040 ;
        RECT 129.275 69.870 130.275 70.040 ;
        RECT 127.755 68.660 127.925 69.700 ;
        RECT 129.045 68.660 129.215 69.700 ;
        RECT 130.335 68.660 130.505 69.700 ;
        RECT 127.985 68.320 128.985 68.490 ;
        RECT 129.275 68.320 130.275 68.490 ;
        RECT 130.675 67.280 130.845 70.060 ;
        RECT 127.345 67.045 130.845 67.280 ;
        RECT 127.345 67.035 130.855 67.045 ;
        RECT 127.345 63.155 127.515 67.035 ;
        RECT 130.675 65.935 130.855 67.035 ;
        RECT 127.985 65.745 128.985 65.915 ;
        RECT 129.275 65.745 130.275 65.915 ;
        RECT 127.755 64.535 127.925 65.575 ;
        RECT 129.045 64.535 129.215 65.575 ;
        RECT 130.335 64.535 130.505 65.575 ;
        RECT 127.985 64.195 128.985 64.365 ;
        RECT 129.275 64.195 130.275 64.365 ;
        RECT 130.675 63.155 130.845 65.935 ;
        RECT 127.345 62.945 130.845 63.155 ;
        RECT 95.175 62.595 104.005 62.765 ;
        RECT 126.085 62.660 126.885 62.670 ;
        RECT 95.175 62.290 95.345 62.595 ;
        RECT 95.175 61.150 95.350 62.290 ;
        RECT 96.070 62.025 103.110 62.195 ;
        RECT 95.685 61.465 95.855 61.965 ;
        RECT 103.325 61.465 103.495 61.965 ;
        RECT 96.070 61.235 103.110 61.405 ;
        RECT 95.175 60.835 95.345 61.150 ;
        RECT 103.835 60.835 104.005 62.595 ;
        RECT 95.175 60.665 104.005 60.835 ;
        RECT 122.895 62.490 126.995 62.660 ;
        RECT 52.175 59.655 61.005 59.825 ;
        RECT 64.030 59.715 70.770 59.885 ;
        RECT 54.830 59.650 59.780 59.655 ;
        RECT 51.680 59.210 63.670 59.380 ;
        RECT 51.680 57.450 51.850 59.210 ;
        RECT 52.575 58.640 60.115 58.810 ;
        RECT 52.190 58.080 52.360 58.580 ;
        RECT 60.330 58.080 60.500 58.580 ;
        RECT 52.575 57.850 60.115 58.020 ;
        RECT 60.840 57.450 61.010 59.210 ;
        RECT 61.735 58.640 62.775 58.810 ;
        RECT 61.350 58.080 61.520 58.580 ;
        RECT 62.990 58.080 63.160 58.580 ;
        RECT 61.735 57.850 62.775 58.020 ;
        RECT 63.500 57.450 63.670 59.210 ;
        RECT 51.680 57.280 63.670 57.450 ;
        RECT 64.030 57.455 64.200 59.715 ;
        RECT 64.880 59.145 69.920 59.315 ;
        RECT 64.540 58.085 64.710 59.085 ;
        RECT 70.090 58.085 70.260 59.085 ;
        RECT 64.880 57.855 69.920 58.025 ;
        RECT 70.600 57.455 70.770 59.715 ;
        RECT 64.030 57.285 70.770 57.455 ;
        RECT 98.770 59.850 105.540 60.020 ;
        RECT 65.420 57.280 66.060 57.285 ;
        RECT 66.600 57.280 67.240 57.285 ;
        RECT 68.000 57.280 68.640 57.285 ;
        RECT 69.650 57.280 70.290 57.285 ;
        RECT 20.090 44.400 26.780 44.570 ;
        RECT 29.100 56.480 45.210 56.660 ;
        RECT 29.100 43.820 29.280 56.480 ;
        RECT 30.030 54.250 35.070 54.420 ;
        RECT 39.030 54.250 44.070 54.420 ;
        RECT 29.645 53.690 29.815 54.190 ;
        RECT 35.285 53.690 35.455 54.190 ;
        RECT 38.645 53.690 38.815 54.190 ;
        RECT 44.285 53.690 44.455 54.190 ;
        RECT 30.030 53.460 35.070 53.630 ;
        RECT 39.030 53.460 44.070 53.630 ;
        RECT 30.030 49.750 35.070 49.920 ;
        RECT 39.030 49.750 44.070 49.920 ;
        RECT 29.645 49.190 29.815 49.690 ;
        RECT 35.285 49.190 35.455 49.690 ;
        RECT 38.645 49.190 38.815 49.690 ;
        RECT 44.285 49.190 44.455 49.690 ;
        RECT 30.030 48.960 35.070 49.130 ;
        RECT 39.030 48.960 44.070 49.130 ;
        RECT 30.030 45.250 35.070 45.420 ;
        RECT 39.030 45.250 44.070 45.420 ;
        RECT 29.645 44.690 29.815 45.190 ;
        RECT 35.285 44.690 35.455 45.190 ;
        RECT 38.645 44.690 38.815 45.190 ;
        RECT 44.285 44.690 44.455 45.190 ;
        RECT 30.030 44.460 35.070 44.630 ;
        RECT 39.030 44.460 44.070 44.630 ;
        RECT 45.030 43.820 45.210 56.480 ;
        RECT 45.870 56.510 61.430 56.680 ;
        RECT 45.870 43.990 46.040 56.510 ;
        RECT 47.750 54.730 52.790 54.900 ;
        RECT 54.750 54.730 59.790 54.900 ;
        RECT 47.410 53.670 47.580 54.670 ;
        RECT 52.960 53.670 53.130 54.670 ;
        RECT 54.410 53.670 54.580 54.670 ;
        RECT 59.960 53.670 60.130 54.670 ;
        RECT 47.750 53.440 52.790 53.610 ;
        RECT 54.750 53.440 59.790 53.610 ;
        RECT 47.750 52.730 52.790 52.900 ;
        RECT 54.750 52.730 59.790 52.900 ;
        RECT 47.410 51.670 47.580 52.670 ;
        RECT 52.960 51.670 53.130 52.670 ;
        RECT 54.410 51.670 54.580 52.670 ;
        RECT 59.960 51.670 60.130 52.670 ;
        RECT 47.750 51.440 52.790 51.610 ;
        RECT 54.750 51.440 59.790 51.610 ;
        RECT 47.750 48.730 52.790 48.900 ;
        RECT 54.750 48.730 59.790 48.900 ;
        RECT 47.410 47.670 47.580 48.670 ;
        RECT 52.960 47.670 53.130 48.670 ;
        RECT 54.410 47.670 54.580 48.670 ;
        RECT 59.960 47.670 60.130 48.670 ;
        RECT 47.750 47.440 52.790 47.610 ;
        RECT 54.750 47.440 59.790 47.610 ;
        RECT 47.750 46.730 52.790 46.900 ;
        RECT 54.750 46.730 59.790 46.900 ;
        RECT 47.410 45.670 47.580 46.670 ;
        RECT 52.960 45.670 53.130 46.670 ;
        RECT 54.410 45.670 54.580 46.670 ;
        RECT 59.960 45.670 60.130 46.670 ;
        RECT 47.750 45.440 52.790 45.610 ;
        RECT 54.750 45.440 59.790 45.610 ;
        RECT 61.260 43.990 61.430 56.510 ;
        RECT 45.870 43.820 61.430 43.990 ;
        RECT 62.290 56.650 70.690 56.820 ;
        RECT 62.290 43.850 62.460 56.650 ;
        RECT 63.210 56.040 68.250 56.210 ;
        RECT 62.870 54.980 63.040 55.980 ;
        RECT 68.420 54.980 68.590 55.980 ;
        RECT 63.210 54.750 68.250 54.920 ;
        RECT 62.870 53.690 63.040 54.690 ;
        RECT 68.420 53.690 68.590 54.690 ;
        RECT 63.210 53.460 68.250 53.630 ;
        RECT 62.870 52.400 63.040 53.400 ;
        RECT 68.420 52.400 68.590 53.400 ;
        RECT 63.210 52.170 68.250 52.340 ;
        RECT 62.870 51.110 63.040 52.110 ;
        RECT 68.420 51.110 68.590 52.110 ;
        RECT 63.210 50.880 68.250 51.050 ;
        RECT 62.870 49.820 63.040 50.820 ;
        RECT 68.420 49.820 68.590 50.820 ;
        RECT 63.210 49.590 68.250 49.760 ;
        RECT 62.870 48.530 63.040 49.530 ;
        RECT 68.420 48.530 68.590 49.530 ;
        RECT 63.210 48.300 68.250 48.470 ;
        RECT 62.870 47.240 63.040 48.240 ;
        RECT 68.420 47.240 68.590 48.240 ;
        RECT 63.210 47.010 68.250 47.180 ;
        RECT 62.870 45.950 63.040 46.950 ;
        RECT 68.420 45.950 68.590 46.950 ;
        RECT 63.210 45.720 68.250 45.890 ;
        RECT 70.520 43.850 70.690 56.650 ;
        RECT 98.770 47.090 98.940 59.850 ;
        RECT 99.620 58.930 104.660 59.100 ;
        RECT 99.235 58.370 99.405 58.870 ;
        RECT 104.875 58.370 105.045 58.870 ;
        RECT 99.620 58.140 104.660 58.310 ;
        RECT 99.235 57.580 99.405 58.080 ;
        RECT 104.875 57.580 105.045 58.080 ;
        RECT 99.620 57.350 104.660 57.520 ;
        RECT 99.235 56.790 99.405 57.290 ;
        RECT 104.875 56.790 105.045 57.290 ;
        RECT 99.620 56.560 104.660 56.730 ;
        RECT 99.235 56.000 99.405 56.500 ;
        RECT 104.875 56.000 105.045 56.500 ;
        RECT 99.620 55.770 104.660 55.940 ;
        RECT 99.235 55.210 99.405 55.710 ;
        RECT 104.875 55.210 105.045 55.710 ;
        RECT 99.620 54.980 104.660 55.150 ;
        RECT 99.235 54.420 99.405 54.920 ;
        RECT 104.875 54.420 105.045 54.920 ;
        RECT 99.620 54.190 104.660 54.360 ;
        RECT 99.235 53.630 99.405 54.130 ;
        RECT 104.875 53.630 105.045 54.130 ;
        RECT 99.620 53.400 104.660 53.570 ;
        RECT 99.235 52.840 99.405 53.340 ;
        RECT 104.875 52.840 105.045 53.340 ;
        RECT 99.620 52.610 104.660 52.780 ;
        RECT 99.235 52.050 99.405 52.550 ;
        RECT 104.875 52.050 105.045 52.550 ;
        RECT 99.620 51.820 104.660 51.990 ;
        RECT 99.235 51.260 99.405 51.760 ;
        RECT 104.875 51.260 105.045 51.760 ;
        RECT 99.620 51.030 104.660 51.200 ;
        RECT 99.235 50.470 99.405 50.970 ;
        RECT 104.875 50.470 105.045 50.970 ;
        RECT 99.620 50.240 104.660 50.410 ;
        RECT 99.235 49.680 99.405 50.180 ;
        RECT 104.875 49.680 105.045 50.180 ;
        RECT 99.620 49.450 104.660 49.620 ;
        RECT 99.235 48.890 99.405 49.390 ;
        RECT 104.875 48.890 105.045 49.390 ;
        RECT 99.620 48.660 104.660 48.830 ;
        RECT 99.235 48.100 99.405 48.600 ;
        RECT 104.875 48.100 105.045 48.600 ;
        RECT 99.620 47.870 104.660 48.040 ;
        RECT 105.370 47.090 105.540 59.850 ;
        RECT 98.770 46.920 105.540 47.090 ;
        RECT 106.350 59.840 113.660 60.020 ;
        RECT 29.100 43.640 45.210 43.820 ;
        RECT 62.290 43.680 70.690 43.850 ;
        RECT 106.350 43.710 106.520 59.840 ;
        RECT 107.680 59.110 112.720 59.280 ;
        RECT 107.340 58.550 107.510 59.050 ;
        RECT 112.890 58.550 113.060 59.050 ;
        RECT 107.680 58.320 112.720 58.490 ;
        RECT 107.340 57.760 107.510 58.260 ;
        RECT 112.890 57.760 113.060 58.260 ;
        RECT 107.680 57.530 112.720 57.700 ;
        RECT 107.340 56.970 107.510 57.470 ;
        RECT 112.890 56.970 113.060 57.470 ;
        RECT 107.680 56.740 112.720 56.910 ;
        RECT 107.340 56.180 107.510 56.680 ;
        RECT 112.890 56.180 113.060 56.680 ;
        RECT 107.680 55.950 112.720 56.120 ;
        RECT 107.340 55.390 107.510 55.890 ;
        RECT 112.890 55.390 113.060 55.890 ;
        RECT 107.680 55.160 112.720 55.330 ;
        RECT 107.340 54.600 107.510 55.100 ;
        RECT 112.890 54.600 113.060 55.100 ;
        RECT 107.680 54.370 112.720 54.540 ;
        RECT 107.340 53.810 107.510 54.310 ;
        RECT 112.890 53.810 113.060 54.310 ;
        RECT 107.680 53.580 112.720 53.750 ;
        RECT 107.340 53.020 107.510 53.520 ;
        RECT 112.890 53.020 113.060 53.520 ;
        RECT 107.680 52.790 112.720 52.960 ;
        RECT 107.340 52.230 107.510 52.730 ;
        RECT 112.890 52.230 113.060 52.730 ;
        RECT 107.680 52.000 112.720 52.170 ;
        RECT 107.340 51.440 107.510 51.940 ;
        RECT 112.890 51.440 113.060 51.940 ;
        RECT 107.680 51.210 112.720 51.380 ;
        RECT 107.340 50.650 107.510 51.150 ;
        RECT 112.890 50.650 113.060 51.150 ;
        RECT 107.680 50.420 112.720 50.590 ;
        RECT 107.340 49.860 107.510 50.360 ;
        RECT 112.890 49.860 113.060 50.360 ;
        RECT 107.680 49.630 112.720 49.800 ;
        RECT 107.340 49.070 107.510 49.570 ;
        RECT 112.890 49.070 113.060 49.570 ;
        RECT 107.680 48.840 112.720 49.010 ;
        RECT 107.340 48.280 107.510 48.780 ;
        RECT 112.890 48.280 113.060 48.780 ;
        RECT 107.680 48.050 112.720 48.220 ;
        RECT 107.340 47.490 107.510 47.990 ;
        RECT 112.890 47.490 113.060 47.990 ;
        RECT 107.680 47.260 112.720 47.430 ;
        RECT 107.340 46.700 107.510 47.200 ;
        RECT 112.890 46.700 113.060 47.200 ;
        RECT 107.680 46.470 112.720 46.640 ;
        RECT 107.340 45.910 107.510 46.410 ;
        RECT 112.890 45.910 113.060 46.410 ;
        RECT 107.680 45.680 112.720 45.850 ;
        RECT 107.340 45.120 107.510 45.620 ;
        RECT 112.890 45.120 113.060 45.620 ;
        RECT 107.680 44.890 112.720 45.060 ;
        RECT 107.340 44.330 107.510 44.830 ;
        RECT 112.890 44.330 113.060 44.830 ;
        RECT 107.680 44.100 112.720 44.270 ;
        RECT 113.490 43.710 113.660 59.840 ;
        RECT 122.895 58.600 123.075 62.490 ;
        RECT 123.795 61.665 124.795 61.835 ;
        RECT 125.085 61.665 126.085 61.835 ;
        RECT 123.565 59.410 123.735 61.450 ;
        RECT 124.855 59.410 125.025 61.450 ;
        RECT 126.145 59.410 126.315 61.450 ;
        RECT 123.795 59.025 124.795 59.195 ;
        RECT 125.085 59.025 126.085 59.195 ;
        RECT 126.825 58.600 126.995 62.490 ;
        RECT 122.895 58.390 126.995 58.600 ;
        RECT 127.345 62.490 130.845 62.660 ;
        RECT 127.345 62.480 130.855 62.490 ;
        RECT 127.345 58.600 127.515 62.480 ;
        RECT 130.675 61.380 130.855 62.480 ;
        RECT 127.985 61.190 128.985 61.360 ;
        RECT 129.275 61.190 130.275 61.360 ;
        RECT 127.755 59.980 127.925 61.020 ;
        RECT 129.045 59.980 129.215 61.020 ;
        RECT 130.335 59.980 130.505 61.020 ;
        RECT 127.985 59.640 128.985 59.810 ;
        RECT 129.275 59.640 130.275 59.810 ;
        RECT 130.675 58.600 130.845 61.380 ;
        RECT 127.345 58.390 130.845 58.600 ;
        RECT 106.350 43.530 113.660 43.710 ;
      LAYER mcon ;
        RECT 30.590 195.050 70.470 195.220 ;
        RECT 30.110 193.100 30.280 194.740 ;
        RECT 31.040 194.480 70.920 194.650 ;
        RECT 30.620 193.500 30.790 194.340 ;
        RECT 71.170 193.500 71.340 194.340 ;
        RECT 31.040 193.190 70.920 193.360 ;
        RECT 30.110 191.180 30.280 191.870 ;
        RECT 30.830 191.360 32.815 191.530 ;
        RECT 44.985 191.360 46.970 191.530 ;
        RECT 99.700 190.580 104.580 190.750 ;
        RECT 98.770 189.420 98.940 190.560 ;
        RECT 99.235 190.100 99.405 190.440 ;
        RECT 104.875 190.100 105.045 190.440 ;
        RECT 99.700 189.790 104.580 189.960 ;
        RECT 99.235 189.310 99.405 189.650 ;
        RECT 104.875 189.310 105.045 189.650 ;
        RECT 99.700 189.000 104.580 189.170 ;
        RECT 99.235 188.520 99.405 188.860 ;
        RECT 104.875 188.520 105.045 188.860 ;
        RECT 99.700 188.210 104.580 188.380 ;
        RECT 98.770 187.020 98.940 188.160 ;
        RECT 99.235 187.730 99.405 188.070 ;
        RECT 104.875 187.730 105.045 188.070 ;
        RECT 99.700 187.420 104.580 187.590 ;
        RECT 99.235 186.940 99.405 187.280 ;
        RECT 104.875 186.940 105.045 187.280 ;
        RECT 99.700 186.630 104.580 186.800 ;
        RECT 99.235 186.150 99.405 186.490 ;
        RECT 104.875 186.150 105.045 186.490 ;
        RECT 99.700 185.840 104.580 186.010 ;
        RECT 98.770 184.580 98.940 185.720 ;
        RECT 99.235 185.360 99.405 185.700 ;
        RECT 104.875 185.360 105.045 185.700 ;
        RECT 99.700 185.050 104.580 185.220 ;
        RECT 37.650 183.410 38.270 183.590 ;
        RECT 15.070 152.960 15.410 154.945 ;
        RECT 16.700 152.960 17.040 154.945 ;
        RECT 20.810 152.960 21.150 154.945 ;
        RECT 22.440 152.960 22.780 154.945 ;
        RECT 24.070 152.960 24.410 154.945 ;
        RECT 25.700 152.960 26.040 154.945 ;
        RECT 29.090 171.310 29.270 182.980 ;
        RECT 30.100 182.600 34.980 182.770 ;
        RECT 39.100 182.600 43.980 182.770 ;
        RECT 29.635 182.120 29.805 182.460 ;
        RECT 35.275 182.120 35.445 182.460 ;
        RECT 38.635 182.120 38.805 182.460 ;
        RECT 44.275 182.120 44.445 182.460 ;
        RECT 30.100 181.810 34.980 181.980 ;
        RECT 39.100 181.810 43.980 181.980 ;
        RECT 30.100 178.100 34.980 178.270 ;
        RECT 39.100 178.100 43.980 178.270 ;
        RECT 29.635 177.620 29.805 177.960 ;
        RECT 35.275 177.620 35.445 177.960 ;
        RECT 38.635 177.620 38.805 177.960 ;
        RECT 44.275 177.620 44.445 177.960 ;
        RECT 30.100 177.310 34.980 177.480 ;
        RECT 39.100 177.310 43.980 177.480 ;
        RECT 30.100 173.600 34.980 173.770 ;
        RECT 39.100 173.600 43.980 173.770 ;
        RECT 29.635 173.120 29.805 173.460 ;
        RECT 35.275 173.120 35.445 173.460 ;
        RECT 38.635 173.120 38.805 173.460 ;
        RECT 44.275 173.120 44.445 173.460 ;
        RECT 30.100 172.810 34.980 172.980 ;
        RECT 39.100 172.810 43.980 172.980 ;
        RECT 37.320 170.570 38.380 170.750 ;
        RECT 47.820 181.620 52.700 181.790 ;
        RECT 54.820 181.620 59.700 181.790 ;
        RECT 47.400 180.640 47.570 181.480 ;
        RECT 52.950 180.640 53.120 181.480 ;
        RECT 54.400 180.640 54.570 181.480 ;
        RECT 59.950 180.640 60.120 181.480 ;
        RECT 61.250 180.570 61.420 182.780 ;
        RECT 47.820 180.330 52.700 180.500 ;
        RECT 54.820 180.330 59.700 180.500 ;
        RECT 47.820 179.620 52.700 179.790 ;
        RECT 54.820 179.620 59.700 179.790 ;
        RECT 47.400 178.640 47.570 179.480 ;
        RECT 52.950 178.640 53.120 179.480 ;
        RECT 54.400 178.640 54.570 179.480 ;
        RECT 59.950 178.640 60.120 179.480 ;
        RECT 47.820 178.330 52.700 178.500 ;
        RECT 54.820 178.330 59.700 178.500 ;
        RECT 47.820 175.620 52.700 175.790 ;
        RECT 54.820 175.620 59.700 175.790 ;
        RECT 47.400 174.640 47.570 175.480 ;
        RECT 52.950 174.640 53.120 175.480 ;
        RECT 54.400 174.640 54.570 175.480 ;
        RECT 59.950 174.640 60.120 175.480 ;
        RECT 47.820 174.330 52.700 174.500 ;
        RECT 54.820 174.330 59.700 174.500 ;
        RECT 47.820 173.620 52.700 173.790 ;
        RECT 54.820 173.620 59.700 173.790 ;
        RECT 47.400 172.640 47.570 173.480 ;
        RECT 52.950 172.640 53.120 173.480 ;
        RECT 54.400 172.640 54.570 173.480 ;
        RECT 59.950 172.640 60.120 173.480 ;
        RECT 47.820 172.330 52.700 172.500 ;
        RECT 54.820 172.330 59.700 172.500 ;
        RECT 63.280 181.340 68.160 181.510 ;
        RECT 62.860 180.360 63.030 181.200 ;
        RECT 68.410 180.360 68.580 181.200 ;
        RECT 63.280 180.050 68.160 180.220 ;
        RECT 62.860 179.070 63.030 179.910 ;
        RECT 68.410 179.070 68.580 179.910 ;
        RECT 63.280 178.760 68.160 178.930 ;
        RECT 62.860 177.780 63.030 178.620 ;
        RECT 68.410 177.780 68.580 178.620 ;
        RECT 63.280 177.470 68.160 177.640 ;
        RECT 62.860 176.490 63.030 177.330 ;
        RECT 68.410 176.490 68.580 177.330 ;
        RECT 63.280 176.180 68.160 176.350 ;
        RECT 62.860 175.200 63.030 176.040 ;
        RECT 68.410 175.200 68.580 176.040 ;
        RECT 63.280 174.890 68.160 175.060 ;
        RECT 62.860 173.910 63.030 174.750 ;
        RECT 68.410 173.910 68.580 174.750 ;
        RECT 63.280 173.600 68.160 173.770 ;
        RECT 62.860 172.620 63.030 173.460 ;
        RECT 68.410 172.620 68.580 173.460 ;
        RECT 63.280 172.310 68.160 172.480 ;
        RECT 62.860 171.330 63.030 172.170 ;
        RECT 68.410 171.330 68.580 172.170 ;
        RECT 70.510 171.930 70.680 181.640 ;
        RECT 99.235 184.570 99.405 184.910 ;
        RECT 104.875 184.570 105.045 184.910 ;
        RECT 99.700 184.260 104.580 184.430 ;
        RECT 99.235 183.780 99.405 184.120 ;
        RECT 104.875 183.780 105.045 184.120 ;
        RECT 99.700 183.470 104.580 183.640 ;
        RECT 98.770 182.280 98.940 183.420 ;
        RECT 99.235 182.990 99.405 183.330 ;
        RECT 104.875 182.990 105.045 183.330 ;
        RECT 99.700 182.680 104.580 182.850 ;
        RECT 99.235 182.200 99.405 182.540 ;
        RECT 104.875 182.200 105.045 182.540 ;
        RECT 99.700 181.890 104.580 182.060 ;
        RECT 99.235 181.410 99.405 181.750 ;
        RECT 104.875 181.410 105.045 181.750 ;
        RECT 98.770 180.040 98.940 181.180 ;
        RECT 99.700 181.100 104.580 181.270 ;
        RECT 99.235 180.620 99.405 180.960 ;
        RECT 104.875 180.620 105.045 180.960 ;
        RECT 99.700 180.310 104.580 180.480 ;
        RECT 99.235 179.830 99.405 180.170 ;
        RECT 104.875 179.830 105.045 180.170 ;
        RECT 99.700 179.520 104.580 179.690 ;
        RECT 107.760 194.350 112.640 194.520 ;
        RECT 107.340 193.870 107.510 194.210 ;
        RECT 112.890 193.870 113.060 194.210 ;
        RECT 107.760 193.560 112.640 193.730 ;
        RECT 107.340 193.080 107.510 193.420 ;
        RECT 112.890 193.080 113.060 193.420 ;
        RECT 107.760 192.770 112.640 192.940 ;
        RECT 113.490 192.830 113.660 194.300 ;
        RECT 107.340 192.290 107.510 192.630 ;
        RECT 112.890 192.290 113.060 192.630 ;
        RECT 107.760 191.980 112.640 192.150 ;
        RECT 107.340 191.500 107.510 191.840 ;
        RECT 112.890 191.500 113.060 191.840 ;
        RECT 107.760 191.190 112.640 191.360 ;
        RECT 107.340 190.710 107.510 191.050 ;
        RECT 112.890 190.710 113.060 191.050 ;
        RECT 107.760 190.400 112.640 190.570 ;
        RECT 107.340 189.920 107.510 190.260 ;
        RECT 112.890 189.920 113.060 190.260 ;
        RECT 113.490 190.260 113.660 191.730 ;
        RECT 107.760 189.610 112.640 189.780 ;
        RECT 107.340 189.130 107.510 189.470 ;
        RECT 112.890 189.130 113.060 189.470 ;
        RECT 107.760 188.820 112.640 188.990 ;
        RECT 107.340 188.340 107.510 188.680 ;
        RECT 112.890 188.340 113.060 188.680 ;
        RECT 107.760 188.030 112.640 188.200 ;
        RECT 107.340 187.550 107.510 187.890 ;
        RECT 112.890 187.550 113.060 187.890 ;
        RECT 113.490 187.680 113.660 189.150 ;
        RECT 107.760 187.240 112.640 187.410 ;
        RECT 107.340 186.760 107.510 187.100 ;
        RECT 112.890 186.760 113.060 187.100 ;
        RECT 107.760 186.450 112.640 186.620 ;
        RECT 107.340 185.970 107.510 186.310 ;
        RECT 112.890 185.970 113.060 186.310 ;
        RECT 107.760 185.660 112.640 185.830 ;
        RECT 107.340 185.180 107.510 185.520 ;
        RECT 112.890 185.180 113.060 185.520 ;
        RECT 113.490 185.160 113.660 186.630 ;
        RECT 107.760 184.870 112.640 185.040 ;
        RECT 107.340 184.390 107.510 184.730 ;
        RECT 112.890 184.390 113.060 184.730 ;
        RECT 122.895 184.855 123.075 188.525 ;
        RECT 123.875 187.830 124.715 188.000 ;
        RECT 125.165 187.830 126.005 188.000 ;
        RECT 123.565 185.655 123.735 187.535 ;
        RECT 124.855 185.655 125.025 187.535 ;
        RECT 126.145 185.655 126.315 187.535 ;
        RECT 123.875 185.190 124.715 185.360 ;
        RECT 125.165 185.190 126.005 185.360 ;
        RECT 128.065 187.355 128.905 187.525 ;
        RECT 129.355 187.355 130.195 187.525 ;
        RECT 127.755 186.225 127.925 187.105 ;
        RECT 129.045 186.225 129.215 187.105 ;
        RECT 130.335 186.225 130.505 187.105 ;
        RECT 128.065 185.805 128.905 185.975 ;
        RECT 129.355 185.805 130.195 185.975 ;
        RECT 130.675 184.895 130.845 185.335 ;
        RECT 107.760 184.080 112.640 184.250 ;
        RECT 107.340 183.600 107.510 183.940 ;
        RECT 112.890 183.600 113.060 183.940 ;
        RECT 107.760 183.290 112.640 183.460 ;
        RECT 107.340 182.810 107.510 183.150 ;
        RECT 112.890 182.810 113.060 183.150 ;
        RECT 113.490 182.810 113.660 184.280 ;
        RECT 107.760 182.500 112.640 182.670 ;
        RECT 107.340 182.020 107.510 182.360 ;
        RECT 112.890 182.020 113.060 182.360 ;
        RECT 107.760 181.710 112.640 181.880 ;
        RECT 107.340 181.230 107.510 181.570 ;
        RECT 112.890 181.230 113.060 181.570 ;
        RECT 107.760 180.920 112.640 181.090 ;
        RECT 107.340 180.440 107.510 180.780 ;
        RECT 112.890 180.440 113.060 180.780 ;
        RECT 107.760 180.130 112.640 180.300 ;
        RECT 107.340 179.650 107.510 179.990 ;
        RECT 112.890 179.650 113.060 179.990 ;
        RECT 113.490 179.980 113.660 181.450 ;
        RECT 107.760 179.340 112.640 179.510 ;
        RECT 95.180 176.330 95.350 177.470 ;
        RECT 96.150 177.215 103.030 177.385 ;
        RECT 95.685 176.735 95.855 177.075 ;
        RECT 103.325 176.735 103.495 177.075 ;
        RECT 96.150 176.425 103.030 176.595 ;
        RECT 122.895 176.755 123.075 180.425 ;
        RECT 123.875 179.730 124.715 179.900 ;
        RECT 125.165 179.730 126.005 179.900 ;
        RECT 123.565 177.555 123.735 179.435 ;
        RECT 124.855 177.555 125.025 179.435 ;
        RECT 126.145 177.555 126.315 179.435 ;
        RECT 123.875 177.090 124.715 177.260 ;
        RECT 125.165 177.090 126.005 177.260 ;
        RECT 128.065 179.255 128.905 179.425 ;
        RECT 129.355 179.255 130.195 179.425 ;
        RECT 127.755 178.125 127.925 179.005 ;
        RECT 129.045 178.125 129.215 179.005 ;
        RECT 130.335 178.125 130.505 179.005 ;
        RECT 128.065 177.705 128.905 177.875 ;
        RECT 129.355 177.705 130.195 177.875 ;
        RECT 130.675 176.795 130.845 177.235 ;
        RECT 95.180 174.400 95.350 175.540 ;
        RECT 96.150 175.285 103.030 175.455 ;
        RECT 95.685 174.805 95.855 175.145 ;
        RECT 103.325 174.805 103.495 175.145 ;
        RECT 96.150 174.495 103.030 174.665 ;
        RECT 63.280 171.020 68.160 171.190 ;
        RECT 95.860 173.480 97.000 173.650 ;
        RECT 97.830 173.480 102.780 173.650 ;
        RECT 94.680 172.030 94.850 173.170 ;
        RECT 95.655 172.910 103.035 173.080 ;
        RECT 95.190 172.430 95.360 172.770 ;
        RECT 103.330 172.430 103.500 172.770 ;
        RECT 95.655 172.120 103.035 172.290 ;
        RECT 104.815 172.910 105.695 173.080 ;
        RECT 104.350 172.430 104.520 172.770 ;
        RECT 105.990 172.430 106.160 172.770 ;
        RECT 104.815 172.120 105.695 172.290 ;
        RECT 95.570 171.550 96.140 171.720 ;
        RECT 107.960 173.415 112.840 173.585 ;
        RECT 107.540 172.435 107.710 173.275 ;
        RECT 113.090 172.435 113.260 173.275 ;
        RECT 107.960 172.125 112.840 172.295 ;
        RECT 113.600 172.030 113.770 173.670 ;
        RECT 80.330 170.750 81.390 170.930 ;
        RECT 52.560 169.780 53.130 169.950 ;
        RECT 51.670 168.330 51.840 169.470 ;
        RECT 52.645 169.210 60.025 169.380 ;
        RECT 52.180 168.730 52.350 169.070 ;
        RECT 60.320 168.730 60.490 169.070 ;
        RECT 52.645 168.420 60.025 168.590 ;
        RECT 61.805 169.210 62.685 169.380 ;
        RECT 61.340 168.730 61.510 169.070 ;
        RECT 62.980 168.730 63.150 169.070 ;
        RECT 61.805 168.420 62.685 168.590 ;
        RECT 52.850 167.850 53.990 168.020 ;
        RECT 54.820 167.850 59.770 168.020 ;
        RECT 65.410 169.780 66.050 169.950 ;
        RECT 66.590 169.780 67.230 169.950 ;
        RECT 67.990 169.780 68.630 169.950 ;
        RECT 69.640 169.780 70.280 169.950 ;
        RECT 54.820 167.410 59.770 167.580 ;
        RECT 52.170 165.960 52.340 167.100 ;
        RECT 53.140 166.835 60.020 167.005 ;
        RECT 52.675 166.355 52.845 166.695 ;
        RECT 60.315 166.355 60.485 166.695 ;
        RECT 53.140 166.045 60.020 166.215 ;
        RECT 64.950 169.205 69.830 169.375 ;
        RECT 64.530 168.225 64.700 169.065 ;
        RECT 70.080 168.225 70.250 169.065 ;
        RECT 64.950 167.915 69.830 168.085 ;
        RECT 70.590 167.830 70.760 169.470 ;
        RECT 52.170 164.030 52.340 165.170 ;
        RECT 53.140 164.905 60.020 165.075 ;
        RECT 52.675 164.425 52.845 164.765 ;
        RECT 60.315 164.425 60.485 164.765 ;
        RECT 53.140 164.115 60.020 164.285 ;
        RECT 56.690 161.810 61.570 161.980 ;
        RECT 55.760 160.320 55.930 161.460 ;
        RECT 56.225 161.330 56.395 161.670 ;
        RECT 61.865 161.330 62.035 161.670 ;
        RECT 56.690 161.020 61.570 161.190 ;
        RECT 56.225 160.540 56.395 160.880 ;
        RECT 61.865 160.540 62.035 160.880 ;
        RECT 56.690 160.230 61.570 160.400 ;
        RECT 56.225 159.750 56.395 160.090 ;
        RECT 61.865 159.750 62.035 160.090 ;
        RECT 56.690 159.440 61.570 159.610 ;
        RECT 55.760 158.080 55.930 159.220 ;
        RECT 56.225 158.960 56.395 159.300 ;
        RECT 61.865 158.960 62.035 159.300 ;
        RECT 56.690 158.650 61.570 158.820 ;
        RECT 56.225 158.170 56.395 158.510 ;
        RECT 61.865 158.170 62.035 158.510 ;
        RECT 56.690 157.860 61.570 158.030 ;
        RECT 56.225 157.380 56.395 157.720 ;
        RECT 61.865 157.380 62.035 157.720 ;
        RECT 56.690 157.070 61.570 157.240 ;
        RECT 55.760 155.780 55.930 156.920 ;
        RECT 56.225 156.590 56.395 156.930 ;
        RECT 61.865 156.590 62.035 156.930 ;
        RECT 56.690 156.280 61.570 156.450 ;
        RECT 56.225 155.800 56.395 156.140 ;
        RECT 61.865 155.800 62.035 156.140 ;
        RECT 56.690 155.490 61.570 155.660 ;
        RECT 56.225 155.010 56.395 155.350 ;
        RECT 61.865 155.010 62.035 155.350 ;
        RECT 56.690 154.700 61.570 154.870 ;
        RECT 55.760 153.340 55.930 154.480 ;
        RECT 56.225 154.220 56.395 154.560 ;
        RECT 61.865 154.220 62.035 154.560 ;
        RECT 56.690 153.910 61.570 154.080 ;
        RECT 56.225 153.430 56.395 153.770 ;
        RECT 61.865 153.430 62.035 153.770 ;
        RECT 15.070 122.530 15.410 124.515 ;
        RECT 16.700 122.530 17.040 124.515 ;
        RECT 56.690 153.120 61.570 153.290 ;
        RECT 56.225 152.640 56.395 152.980 ;
        RECT 61.865 152.640 62.035 152.980 ;
        RECT 56.690 152.330 61.570 152.500 ;
        RECT 55.760 150.940 55.930 152.080 ;
        RECT 56.225 151.850 56.395 152.190 ;
        RECT 61.865 151.850 62.035 152.190 ;
        RECT 56.690 151.540 61.570 151.710 ;
        RECT 56.225 151.060 56.395 151.400 ;
        RECT 61.865 151.060 62.035 151.400 ;
        RECT 56.690 150.750 61.570 150.920 ;
        RECT 64.750 161.990 69.630 162.160 ;
        RECT 64.330 161.510 64.500 161.850 ;
        RECT 69.880 161.510 70.050 161.850 ;
        RECT 64.750 161.200 69.630 161.370 ;
        RECT 64.330 160.720 64.500 161.060 ;
        RECT 69.880 160.720 70.050 161.060 ;
        RECT 64.750 160.410 69.630 160.580 ;
        RECT 64.330 159.930 64.500 160.270 ;
        RECT 69.880 159.930 70.050 160.270 ;
        RECT 70.480 160.050 70.650 161.520 ;
        RECT 64.750 159.620 69.630 159.790 ;
        RECT 64.330 159.140 64.500 159.480 ;
        RECT 69.880 159.140 70.050 159.480 ;
        RECT 64.750 158.830 69.630 159.000 ;
        RECT 64.330 158.350 64.500 158.690 ;
        RECT 69.880 158.350 70.050 158.690 ;
        RECT 64.750 158.040 69.630 158.210 ;
        RECT 64.330 157.560 64.500 157.900 ;
        RECT 69.880 157.560 70.050 157.900 ;
        RECT 64.750 157.250 69.630 157.420 ;
        RECT 70.480 157.220 70.650 158.690 ;
        RECT 72.100 158.520 72.280 170.190 ;
        RECT 73.110 168.520 77.990 168.690 ;
        RECT 82.110 168.520 86.990 168.690 ;
        RECT 72.645 168.040 72.815 168.380 ;
        RECT 78.285 168.040 78.455 168.380 ;
        RECT 81.645 168.040 81.815 168.380 ;
        RECT 87.285 168.040 87.455 168.380 ;
        RECT 73.110 167.730 77.990 167.900 ;
        RECT 82.110 167.730 86.990 167.900 ;
        RECT 73.110 164.020 77.990 164.190 ;
        RECT 82.110 164.020 86.990 164.190 ;
        RECT 72.645 163.540 72.815 163.880 ;
        RECT 78.285 163.540 78.455 163.880 ;
        RECT 81.645 163.540 81.815 163.880 ;
        RECT 87.285 163.540 87.455 163.880 ;
        RECT 73.110 163.230 77.990 163.400 ;
        RECT 82.110 163.230 86.990 163.400 ;
        RECT 73.110 159.520 77.990 159.690 ;
        RECT 82.110 159.520 86.990 159.690 ;
        RECT 72.645 159.040 72.815 159.380 ;
        RECT 78.285 159.040 78.455 159.380 ;
        RECT 81.645 159.040 81.815 159.380 ;
        RECT 87.285 159.040 87.455 159.380 ;
        RECT 73.110 158.730 77.990 158.900 ;
        RECT 82.110 158.730 86.990 158.900 ;
        RECT 90.830 169.000 95.710 169.170 ;
        RECT 97.830 169.000 102.710 169.170 ;
        RECT 90.410 168.020 90.580 168.860 ;
        RECT 95.960 168.020 96.130 168.860 ;
        RECT 97.410 168.020 97.580 168.860 ;
        RECT 102.960 168.020 103.130 168.860 ;
        RECT 90.830 167.710 95.710 167.880 ;
        RECT 97.830 167.710 102.710 167.880 ;
        RECT 90.830 167.000 95.710 167.170 ;
        RECT 97.830 167.000 102.710 167.170 ;
        RECT 90.410 166.020 90.580 166.860 ;
        RECT 95.960 166.020 96.130 166.860 ;
        RECT 97.410 166.020 97.580 166.860 ;
        RECT 102.960 166.020 103.130 166.860 ;
        RECT 90.830 165.710 95.710 165.880 ;
        RECT 97.830 165.710 102.710 165.880 ;
        RECT 90.830 163.000 95.710 163.170 ;
        RECT 97.830 163.000 102.710 163.170 ;
        RECT 90.410 162.020 90.580 162.860 ;
        RECT 95.960 162.020 96.130 162.860 ;
        RECT 97.410 162.020 97.580 162.860 ;
        RECT 102.960 162.020 103.130 162.860 ;
        RECT 90.830 161.710 95.710 161.880 ;
        RECT 97.830 161.710 102.710 161.880 ;
        RECT 90.830 161.000 95.710 161.170 ;
        RECT 97.830 161.000 102.710 161.170 ;
        RECT 90.410 160.020 90.580 160.860 ;
        RECT 95.960 160.020 96.130 160.860 ;
        RECT 97.410 160.020 97.580 160.860 ;
        RECT 102.960 160.020 103.130 160.860 ;
        RECT 90.830 159.710 95.710 159.880 ;
        RECT 97.830 159.710 102.710 159.880 ;
        RECT 104.260 158.720 104.430 160.930 ;
        RECT 106.290 170.310 111.170 170.480 ;
        RECT 105.870 169.330 106.040 170.170 ;
        RECT 111.420 169.330 111.590 170.170 ;
        RECT 106.290 169.020 111.170 169.190 ;
        RECT 105.870 168.040 106.040 168.880 ;
        RECT 111.420 168.040 111.590 168.880 ;
        RECT 106.290 167.730 111.170 167.900 ;
        RECT 105.870 166.750 106.040 167.590 ;
        RECT 111.420 166.750 111.590 167.590 ;
        RECT 106.290 166.440 111.170 166.610 ;
        RECT 105.870 165.460 106.040 166.300 ;
        RECT 111.420 165.460 111.590 166.300 ;
        RECT 106.290 165.150 111.170 165.320 ;
        RECT 105.870 164.170 106.040 165.010 ;
        RECT 111.420 164.170 111.590 165.010 ;
        RECT 106.290 163.860 111.170 164.030 ;
        RECT 105.870 162.880 106.040 163.720 ;
        RECT 111.420 162.880 111.590 163.720 ;
        RECT 106.290 162.570 111.170 162.740 ;
        RECT 105.870 161.590 106.040 162.430 ;
        RECT 111.420 161.590 111.590 162.430 ;
        RECT 106.290 161.280 111.170 161.450 ;
        RECT 105.870 160.300 106.040 161.140 ;
        RECT 111.420 160.300 111.590 161.140 ;
        RECT 106.290 159.990 111.170 160.160 ;
        RECT 113.520 159.860 113.690 169.570 ;
        RECT 122.895 168.655 123.075 172.325 ;
        RECT 123.875 171.630 124.715 171.800 ;
        RECT 125.165 171.630 126.005 171.800 ;
        RECT 123.565 169.455 123.735 171.335 ;
        RECT 124.855 169.455 125.025 171.335 ;
        RECT 126.145 169.455 126.315 171.335 ;
        RECT 123.875 168.990 124.715 169.160 ;
        RECT 125.165 168.990 126.005 169.160 ;
        RECT 128.065 171.155 128.905 171.325 ;
        RECT 129.355 171.155 130.195 171.325 ;
        RECT 127.755 170.025 127.925 170.905 ;
        RECT 129.045 170.025 129.215 170.905 ;
        RECT 130.335 170.025 130.505 170.905 ;
        RECT 128.065 169.605 128.905 169.775 ;
        RECT 129.355 169.605 130.195 169.775 ;
        RECT 130.675 168.695 130.845 169.135 ;
        RECT 114.655 162.620 114.825 163.060 ;
        RECT 115.305 161.980 116.145 162.150 ;
        RECT 116.595 161.980 117.435 162.150 ;
        RECT 114.995 160.850 115.165 161.730 ;
        RECT 116.285 160.850 116.455 161.730 ;
        RECT 117.575 160.850 117.745 161.730 ;
        RECT 115.305 160.430 116.145 160.600 ;
        RECT 116.595 160.430 117.435 160.600 ;
        RECT 119.495 162.595 120.335 162.765 ;
        RECT 120.785 162.595 121.625 162.765 ;
        RECT 119.185 160.420 119.355 162.300 ;
        RECT 120.475 160.420 120.645 162.300 ;
        RECT 121.765 160.420 121.935 162.300 ;
        RECT 119.495 159.955 120.335 160.125 ;
        RECT 120.785 159.955 121.625 160.125 ;
        RECT 122.425 159.430 122.605 163.100 ;
        RECT 122.895 160.555 123.075 164.225 ;
        RECT 123.875 163.530 124.715 163.700 ;
        RECT 125.165 163.530 126.005 163.700 ;
        RECT 123.565 161.355 123.735 163.235 ;
        RECT 124.855 161.355 125.025 163.235 ;
        RECT 126.145 161.355 126.315 163.235 ;
        RECT 123.875 160.890 124.715 161.060 ;
        RECT 125.165 160.890 126.005 161.060 ;
        RECT 128.065 163.055 128.905 163.225 ;
        RECT 129.355 163.055 130.195 163.225 ;
        RECT 127.755 161.925 127.925 162.805 ;
        RECT 129.045 161.925 129.215 162.805 ;
        RECT 130.335 161.925 130.505 162.805 ;
        RECT 128.065 161.505 128.905 161.675 ;
        RECT 129.355 161.505 130.195 161.675 ;
        RECT 130.675 160.595 130.845 161.035 ;
        RECT 80.660 157.910 81.280 158.090 ;
        RECT 114.655 158.080 114.825 158.520 ;
        RECT 64.330 156.770 64.500 157.110 ;
        RECT 69.880 156.770 70.050 157.110 ;
        RECT 64.750 156.460 69.630 156.630 ;
        RECT 64.330 155.980 64.500 156.320 ;
        RECT 69.880 155.980 70.050 156.320 ;
        RECT 64.750 155.670 69.630 155.840 ;
        RECT 64.330 155.190 64.500 155.530 ;
        RECT 69.880 155.190 70.050 155.530 ;
        RECT 64.750 154.880 69.630 155.050 ;
        RECT 70.480 154.870 70.650 156.340 ;
        RECT 64.330 154.400 64.500 154.740 ;
        RECT 69.880 154.400 70.050 154.740 ;
        RECT 64.750 154.090 69.630 154.260 ;
        RECT 64.330 153.610 64.500 153.950 ;
        RECT 69.880 153.610 70.050 153.950 ;
        RECT 64.750 153.300 69.630 153.470 ;
        RECT 64.330 152.820 64.500 153.160 ;
        RECT 69.880 152.820 70.050 153.160 ;
        RECT 64.750 152.510 69.630 152.680 ;
        RECT 64.330 152.030 64.500 152.370 ;
        RECT 69.880 152.030 70.050 152.370 ;
        RECT 70.480 152.350 70.650 153.820 ;
        RECT 64.750 151.720 69.630 151.890 ;
        RECT 64.330 151.240 64.500 151.580 ;
        RECT 69.880 151.240 70.050 151.580 ;
        RECT 64.750 150.930 69.630 151.100 ;
        RECT 64.330 150.450 64.500 150.790 ;
        RECT 69.880 150.450 70.050 150.790 ;
        RECT 64.750 150.140 69.630 150.310 ;
        RECT 64.330 149.660 64.500 150.000 ;
        RECT 69.880 149.660 70.050 150.000 ;
        RECT 70.480 149.770 70.650 151.240 ;
        RECT 64.750 149.350 69.630 149.520 ;
        RECT 64.330 148.870 64.500 149.210 ;
        RECT 69.880 148.870 70.050 149.210 ;
        RECT 64.750 148.560 69.630 148.730 ;
        RECT 64.330 148.080 64.500 148.420 ;
        RECT 69.880 148.080 70.050 148.420 ;
        RECT 64.750 147.770 69.630 147.940 ;
        RECT 64.330 147.290 64.500 147.630 ;
        RECT 69.880 147.290 70.050 147.630 ;
        RECT 70.480 147.200 70.650 148.670 ;
        RECT 64.750 146.980 69.630 147.150 ;
        RECT 80.660 156.130 81.280 156.310 ;
        RECT 72.100 144.030 72.280 155.700 ;
        RECT 73.110 155.320 77.990 155.490 ;
        RECT 82.110 155.320 86.990 155.490 ;
        RECT 72.645 154.840 72.815 155.180 ;
        RECT 78.285 154.840 78.455 155.180 ;
        RECT 81.645 154.840 81.815 155.180 ;
        RECT 87.285 154.840 87.455 155.180 ;
        RECT 73.110 154.530 77.990 154.700 ;
        RECT 82.110 154.530 86.990 154.700 ;
        RECT 73.110 150.820 77.990 150.990 ;
        RECT 82.110 150.820 86.990 150.990 ;
        RECT 72.645 150.340 72.815 150.680 ;
        RECT 78.285 150.340 78.455 150.680 ;
        RECT 81.645 150.340 81.815 150.680 ;
        RECT 87.285 150.340 87.455 150.680 ;
        RECT 73.110 150.030 77.990 150.200 ;
        RECT 82.110 150.030 86.990 150.200 ;
        RECT 73.110 146.320 77.990 146.490 ;
        RECT 82.110 146.320 86.990 146.490 ;
        RECT 72.645 145.840 72.815 146.180 ;
        RECT 78.285 145.840 78.455 146.180 ;
        RECT 81.645 145.840 81.815 146.180 ;
        RECT 87.285 145.840 87.455 146.180 ;
        RECT 73.110 145.530 77.990 145.700 ;
        RECT 82.110 145.530 86.990 145.700 ;
        RECT 80.330 143.290 81.390 143.470 ;
        RECT 90.830 154.340 95.710 154.510 ;
        RECT 97.830 154.340 102.710 154.510 ;
        RECT 90.410 153.360 90.580 154.200 ;
        RECT 95.960 153.360 96.130 154.200 ;
        RECT 97.410 153.360 97.580 154.200 ;
        RECT 102.960 153.360 103.130 154.200 ;
        RECT 104.260 153.290 104.430 155.500 ;
        RECT 90.830 153.050 95.710 153.220 ;
        RECT 97.830 153.050 102.710 153.220 ;
        RECT 90.830 152.340 95.710 152.510 ;
        RECT 97.830 152.340 102.710 152.510 ;
        RECT 90.410 151.360 90.580 152.200 ;
        RECT 95.960 151.360 96.130 152.200 ;
        RECT 97.410 151.360 97.580 152.200 ;
        RECT 102.960 151.360 103.130 152.200 ;
        RECT 90.830 151.050 95.710 151.220 ;
        RECT 97.830 151.050 102.710 151.220 ;
        RECT 90.830 148.340 95.710 148.510 ;
        RECT 97.830 148.340 102.710 148.510 ;
        RECT 90.410 147.360 90.580 148.200 ;
        RECT 95.960 147.360 96.130 148.200 ;
        RECT 97.410 147.360 97.580 148.200 ;
        RECT 102.960 147.360 103.130 148.200 ;
        RECT 90.830 147.050 95.710 147.220 ;
        RECT 97.830 147.050 102.710 147.220 ;
        RECT 90.830 146.340 95.710 146.510 ;
        RECT 97.830 146.340 102.710 146.510 ;
        RECT 90.410 145.360 90.580 146.200 ;
        RECT 95.960 145.360 96.130 146.200 ;
        RECT 97.410 145.360 97.580 146.200 ;
        RECT 102.960 145.360 103.130 146.200 ;
        RECT 90.830 145.050 95.710 145.220 ;
        RECT 97.830 145.050 102.710 145.220 ;
        RECT 115.305 157.440 116.145 157.610 ;
        RECT 116.595 157.440 117.435 157.610 ;
        RECT 114.995 156.310 115.165 157.190 ;
        RECT 116.285 156.310 116.455 157.190 ;
        RECT 117.575 156.310 117.745 157.190 ;
        RECT 115.305 155.890 116.145 156.060 ;
        RECT 116.595 155.890 117.435 156.060 ;
        RECT 106.290 154.060 111.170 154.230 ;
        RECT 105.870 153.080 106.040 153.920 ;
        RECT 111.420 153.080 111.590 153.920 ;
        RECT 106.290 152.770 111.170 152.940 ;
        RECT 105.870 151.790 106.040 152.630 ;
        RECT 111.420 151.790 111.590 152.630 ;
        RECT 106.290 151.480 111.170 151.650 ;
        RECT 105.870 150.500 106.040 151.340 ;
        RECT 111.420 150.500 111.590 151.340 ;
        RECT 106.290 150.190 111.170 150.360 ;
        RECT 105.870 149.210 106.040 150.050 ;
        RECT 111.420 149.210 111.590 150.050 ;
        RECT 106.290 148.900 111.170 149.070 ;
        RECT 105.870 147.920 106.040 148.760 ;
        RECT 111.420 147.920 111.590 148.760 ;
        RECT 106.290 147.610 111.170 147.780 ;
        RECT 105.870 146.630 106.040 147.470 ;
        RECT 111.420 146.630 111.590 147.470 ;
        RECT 106.290 146.320 111.170 146.490 ;
        RECT 105.870 145.340 106.040 146.180 ;
        RECT 111.420 145.340 111.590 146.180 ;
        RECT 106.290 145.030 111.170 145.200 ;
        RECT 105.870 144.050 106.040 144.890 ;
        RECT 111.420 144.050 111.590 144.890 ;
        RECT 113.520 144.650 113.690 154.360 ;
        RECT 114.655 154.020 114.825 154.460 ;
        RECT 115.305 153.380 116.145 153.550 ;
        RECT 116.595 153.380 117.435 153.550 ;
        RECT 114.995 152.250 115.165 153.130 ;
        RECT 116.285 152.250 116.455 153.130 ;
        RECT 117.575 152.250 117.745 153.130 ;
        RECT 115.305 151.830 116.145 152.000 ;
        RECT 116.595 151.830 117.435 152.000 ;
        RECT 114.655 149.960 114.825 150.400 ;
        RECT 115.305 149.320 116.145 149.490 ;
        RECT 116.595 149.320 117.435 149.490 ;
        RECT 114.995 148.190 115.165 149.070 ;
        RECT 116.285 148.190 116.455 149.070 ;
        RECT 117.575 148.190 117.745 149.070 ;
        RECT 115.305 147.770 116.145 147.940 ;
        RECT 116.595 147.770 117.435 147.940 ;
        RECT 106.290 143.740 111.170 143.910 ;
        RECT 114.655 145.900 114.825 146.340 ;
        RECT 115.305 145.260 116.145 145.430 ;
        RECT 116.595 145.260 117.435 145.430 ;
        RECT 114.995 144.130 115.165 145.010 ;
        RECT 116.285 144.130 116.455 145.010 ;
        RECT 117.575 144.130 117.745 145.010 ;
        RECT 115.305 143.710 116.145 143.880 ;
        RECT 116.595 143.710 117.435 143.880 ;
        RECT 95.570 142.500 96.140 142.670 ;
        RECT 94.680 141.050 94.850 142.190 ;
        RECT 95.655 141.930 103.035 142.100 ;
        RECT 95.190 141.450 95.360 141.790 ;
        RECT 103.330 141.450 103.500 141.790 ;
        RECT 95.655 141.140 103.035 141.310 ;
        RECT 104.815 141.930 105.695 142.100 ;
        RECT 104.350 141.450 104.520 141.790 ;
        RECT 105.990 141.450 106.160 141.790 ;
        RECT 104.815 141.140 105.695 141.310 ;
        RECT 95.860 140.570 97.000 140.740 ;
        RECT 97.830 140.570 102.780 140.740 ;
        RECT 108.420 142.500 109.060 142.670 ;
        RECT 109.600 142.500 110.240 142.670 ;
        RECT 111.000 142.500 111.640 142.670 ;
        RECT 112.650 142.500 113.290 142.670 ;
        RECT 97.830 140.130 102.780 140.300 ;
        RECT 95.180 138.680 95.350 139.820 ;
        RECT 96.150 139.555 103.030 139.725 ;
        RECT 95.685 139.075 95.855 139.415 ;
        RECT 103.325 139.075 103.495 139.415 ;
        RECT 96.150 138.765 103.030 138.935 ;
        RECT 107.960 141.925 112.840 142.095 ;
        RECT 107.540 140.945 107.710 141.785 ;
        RECT 113.090 140.945 113.260 141.785 ;
        RECT 107.960 140.635 112.840 140.805 ;
        RECT 113.600 140.550 113.770 142.190 ;
        RECT 114.655 141.840 114.825 142.280 ;
        RECT 115.305 141.200 116.145 141.370 ;
        RECT 116.595 141.200 117.435 141.370 ;
        RECT 114.995 140.070 115.165 140.950 ;
        RECT 116.285 140.070 116.455 140.950 ;
        RECT 117.575 140.070 117.745 140.950 ;
        RECT 115.305 139.650 116.145 139.820 ;
        RECT 116.595 139.650 117.435 139.820 ;
        RECT 119.495 158.055 120.335 158.225 ;
        RECT 120.785 158.055 121.625 158.225 ;
        RECT 119.185 155.880 119.355 157.760 ;
        RECT 120.475 155.880 120.645 157.760 ;
        RECT 121.765 155.880 121.935 157.760 ;
        RECT 119.495 155.415 120.335 155.585 ;
        RECT 120.785 155.415 121.625 155.585 ;
        RECT 122.425 154.890 122.605 158.560 ;
        RECT 119.495 153.995 120.335 154.165 ;
        RECT 120.785 153.995 121.625 154.165 ;
        RECT 119.185 151.820 119.355 153.700 ;
        RECT 120.475 151.820 120.645 153.700 ;
        RECT 121.765 151.820 121.935 153.700 ;
        RECT 119.495 151.355 120.335 151.525 ;
        RECT 120.785 151.355 121.625 151.525 ;
        RECT 122.425 150.830 122.605 154.500 ;
        RECT 122.895 152.455 123.075 156.125 ;
        RECT 123.875 155.430 124.715 155.600 ;
        RECT 125.165 155.430 126.005 155.600 ;
        RECT 123.565 153.255 123.735 155.135 ;
        RECT 124.855 153.255 125.025 155.135 ;
        RECT 126.145 153.255 126.315 155.135 ;
        RECT 123.875 152.790 124.715 152.960 ;
        RECT 125.165 152.790 126.005 152.960 ;
        RECT 128.065 154.955 128.905 155.125 ;
        RECT 129.355 154.955 130.195 155.125 ;
        RECT 127.755 153.825 127.925 154.705 ;
        RECT 129.045 153.825 129.215 154.705 ;
        RECT 130.335 153.825 130.505 154.705 ;
        RECT 128.065 153.405 128.905 153.575 ;
        RECT 129.355 153.405 130.195 153.575 ;
        RECT 130.675 152.495 130.845 152.935 ;
        RECT 119.495 149.935 120.335 150.105 ;
        RECT 120.785 149.935 121.625 150.105 ;
        RECT 119.185 147.760 119.355 149.640 ;
        RECT 120.475 147.760 120.645 149.640 ;
        RECT 121.765 147.760 121.935 149.640 ;
        RECT 119.495 147.295 120.335 147.465 ;
        RECT 120.785 147.295 121.625 147.465 ;
        RECT 122.425 146.770 122.605 150.440 ;
        RECT 119.495 145.875 120.335 146.045 ;
        RECT 120.785 145.875 121.625 146.045 ;
        RECT 119.185 143.700 119.355 145.580 ;
        RECT 120.475 143.700 120.645 145.580 ;
        RECT 121.765 143.700 121.935 145.580 ;
        RECT 119.495 143.235 120.335 143.405 ;
        RECT 120.785 143.235 121.625 143.405 ;
        RECT 122.425 142.710 122.605 146.380 ;
        RECT 122.895 144.355 123.075 148.025 ;
        RECT 123.875 147.330 124.715 147.500 ;
        RECT 125.165 147.330 126.005 147.500 ;
        RECT 123.565 145.155 123.735 147.035 ;
        RECT 124.855 145.155 125.025 147.035 ;
        RECT 126.145 145.155 126.315 147.035 ;
        RECT 123.875 144.690 124.715 144.860 ;
        RECT 125.165 144.690 126.005 144.860 ;
        RECT 128.065 146.855 128.905 147.025 ;
        RECT 129.355 146.855 130.195 147.025 ;
        RECT 127.755 145.725 127.925 146.605 ;
        RECT 129.045 145.725 129.215 146.605 ;
        RECT 130.335 145.725 130.505 146.605 ;
        RECT 128.065 145.305 128.905 145.475 ;
        RECT 129.355 145.305 130.195 145.475 ;
        RECT 130.675 144.395 130.845 144.835 ;
        RECT 119.495 141.815 120.335 141.985 ;
        RECT 120.785 141.815 121.625 141.985 ;
        RECT 119.185 139.640 119.355 141.520 ;
        RECT 120.475 139.640 120.645 141.520 ;
        RECT 121.765 139.640 121.935 141.520 ;
        RECT 119.495 139.175 120.335 139.345 ;
        RECT 120.785 139.175 121.625 139.345 ;
        RECT 122.425 138.650 122.605 142.320 ;
        RECT 95.180 136.750 95.350 137.890 ;
        RECT 96.150 137.625 103.030 137.795 ;
        RECT 95.685 137.145 95.855 137.485 ;
        RECT 103.325 137.145 103.495 137.485 ;
        RECT 96.150 136.835 103.030 137.005 ;
        RECT 122.895 136.255 123.075 139.925 ;
        RECT 123.875 139.230 124.715 139.400 ;
        RECT 125.165 139.230 126.005 139.400 ;
        RECT 123.565 137.055 123.735 138.935 ;
        RECT 124.855 137.055 125.025 138.935 ;
        RECT 126.145 137.055 126.315 138.935 ;
        RECT 123.875 136.590 124.715 136.760 ;
        RECT 125.165 136.590 126.005 136.760 ;
        RECT 128.065 138.755 128.905 138.925 ;
        RECT 129.355 138.755 130.195 138.925 ;
        RECT 127.755 137.625 127.925 138.505 ;
        RECT 129.045 137.625 129.215 138.505 ;
        RECT 130.335 137.625 130.505 138.505 ;
        RECT 128.065 137.205 128.905 137.375 ;
        RECT 129.355 137.205 130.195 137.375 ;
        RECT 130.675 136.295 130.845 136.735 ;
        RECT 99.700 134.530 104.580 134.700 ;
        RECT 98.770 133.040 98.940 134.180 ;
        RECT 99.235 134.050 99.405 134.390 ;
        RECT 104.875 134.050 105.045 134.390 ;
        RECT 99.700 133.740 104.580 133.910 ;
        RECT 99.235 133.260 99.405 133.600 ;
        RECT 104.875 133.260 105.045 133.600 ;
        RECT 99.700 132.950 104.580 133.120 ;
        RECT 99.235 132.470 99.405 132.810 ;
        RECT 104.875 132.470 105.045 132.810 ;
        RECT 99.700 132.160 104.580 132.330 ;
        RECT 98.770 130.800 98.940 131.940 ;
        RECT 99.235 131.680 99.405 132.020 ;
        RECT 104.875 131.680 105.045 132.020 ;
        RECT 99.700 131.370 104.580 131.540 ;
        RECT 99.235 130.890 99.405 131.230 ;
        RECT 104.875 130.890 105.045 131.230 ;
        RECT 99.700 130.580 104.580 130.750 ;
        RECT 99.235 130.100 99.405 130.440 ;
        RECT 104.875 130.100 105.045 130.440 ;
        RECT 99.700 129.790 104.580 129.960 ;
        RECT 98.770 128.500 98.940 129.640 ;
        RECT 99.235 129.310 99.405 129.650 ;
        RECT 104.875 129.310 105.045 129.650 ;
        RECT 99.700 129.000 104.580 129.170 ;
        RECT 99.235 128.520 99.405 128.860 ;
        RECT 104.875 128.520 105.045 128.860 ;
        RECT 99.700 128.210 104.580 128.380 ;
        RECT 99.235 127.730 99.405 128.070 ;
        RECT 104.875 127.730 105.045 128.070 ;
        RECT 99.700 127.420 104.580 127.590 ;
        RECT 98.770 126.060 98.940 127.200 ;
        RECT 99.235 126.940 99.405 127.280 ;
        RECT 104.875 126.940 105.045 127.280 ;
        RECT 99.700 126.630 104.580 126.800 ;
        RECT 99.235 126.150 99.405 126.490 ;
        RECT 104.875 126.150 105.045 126.490 ;
        RECT 99.700 125.840 104.580 126.010 ;
        RECT 99.235 125.360 99.405 125.700 ;
        RECT 104.875 125.360 105.045 125.700 ;
        RECT 99.700 125.050 104.580 125.220 ;
        RECT 98.770 123.660 98.940 124.800 ;
        RECT 99.235 124.570 99.405 124.910 ;
        RECT 104.875 124.570 105.045 124.910 ;
        RECT 99.700 124.260 104.580 124.430 ;
        RECT 99.235 123.780 99.405 124.120 ;
        RECT 104.875 123.780 105.045 124.120 ;
        RECT 99.700 123.470 104.580 123.640 ;
        RECT 107.760 134.710 112.640 134.880 ;
        RECT 107.340 134.230 107.510 134.570 ;
        RECT 112.890 134.230 113.060 134.570 ;
        RECT 107.760 133.920 112.640 134.090 ;
        RECT 107.340 133.440 107.510 133.780 ;
        RECT 112.890 133.440 113.060 133.780 ;
        RECT 107.760 133.130 112.640 133.300 ;
        RECT 107.340 132.650 107.510 132.990 ;
        RECT 112.890 132.650 113.060 132.990 ;
        RECT 113.490 132.770 113.660 134.240 ;
        RECT 107.760 132.340 112.640 132.510 ;
        RECT 107.340 131.860 107.510 132.200 ;
        RECT 112.890 131.860 113.060 132.200 ;
        RECT 107.760 131.550 112.640 131.720 ;
        RECT 107.340 131.070 107.510 131.410 ;
        RECT 112.890 131.070 113.060 131.410 ;
        RECT 114.655 133.720 114.825 134.160 ;
        RECT 115.305 133.080 116.145 133.250 ;
        RECT 116.595 133.080 117.435 133.250 ;
        RECT 114.995 131.950 115.165 132.830 ;
        RECT 116.285 131.950 116.455 132.830 ;
        RECT 117.575 131.950 117.745 132.830 ;
        RECT 115.305 131.530 116.145 131.700 ;
        RECT 116.595 131.530 117.435 131.700 ;
        RECT 107.760 130.760 112.640 130.930 ;
        RECT 107.340 130.280 107.510 130.620 ;
        RECT 112.890 130.280 113.060 130.620 ;
        RECT 107.760 129.970 112.640 130.140 ;
        RECT 113.490 129.940 113.660 131.410 ;
        RECT 107.340 129.490 107.510 129.830 ;
        RECT 112.890 129.490 113.060 129.830 ;
        RECT 107.760 129.180 112.640 129.350 ;
        RECT 107.340 128.700 107.510 129.040 ;
        RECT 112.890 128.700 113.060 129.040 ;
        RECT 107.760 128.390 112.640 128.560 ;
        RECT 107.340 127.910 107.510 128.250 ;
        RECT 112.890 127.910 113.060 128.250 ;
        RECT 107.760 127.600 112.640 127.770 ;
        RECT 113.490 127.590 113.660 129.060 ;
        RECT 107.340 127.120 107.510 127.460 ;
        RECT 112.890 127.120 113.060 127.460 ;
        RECT 107.760 126.810 112.640 126.980 ;
        RECT 107.340 126.330 107.510 126.670 ;
        RECT 112.890 126.330 113.060 126.670 ;
        RECT 114.655 129.660 114.825 130.100 ;
        RECT 115.305 129.020 116.145 129.190 ;
        RECT 116.595 129.020 117.435 129.190 ;
        RECT 114.995 127.890 115.165 128.770 ;
        RECT 116.285 127.890 116.455 128.770 ;
        RECT 117.575 127.890 117.745 128.770 ;
        RECT 115.305 127.470 116.145 127.640 ;
        RECT 116.595 127.470 117.435 127.640 ;
        RECT 107.760 126.020 112.640 126.190 ;
        RECT 107.340 125.540 107.510 125.880 ;
        RECT 112.890 125.540 113.060 125.880 ;
        RECT 107.760 125.230 112.640 125.400 ;
        RECT 107.340 124.750 107.510 125.090 ;
        RECT 112.890 124.750 113.060 125.090 ;
        RECT 113.490 125.070 113.660 126.540 ;
        RECT 107.760 124.440 112.640 124.610 ;
        RECT 107.340 123.960 107.510 124.300 ;
        RECT 112.890 123.960 113.060 124.300 ;
        RECT 107.760 123.650 112.640 123.820 ;
        RECT 107.340 123.170 107.510 123.510 ;
        RECT 112.890 123.170 113.060 123.510 ;
        RECT 107.760 122.860 112.640 123.030 ;
        RECT 107.340 122.380 107.510 122.720 ;
        RECT 112.890 122.380 113.060 122.720 ;
        RECT 113.490 122.490 113.660 123.960 ;
        RECT 114.655 125.600 114.825 126.040 ;
        RECT 115.305 124.960 116.145 125.130 ;
        RECT 116.595 124.960 117.435 125.130 ;
        RECT 114.995 123.830 115.165 124.710 ;
        RECT 116.285 123.830 116.455 124.710 ;
        RECT 117.575 123.830 117.745 124.710 ;
        RECT 115.305 123.410 116.145 123.580 ;
        RECT 116.595 123.410 117.435 123.580 ;
        RECT 107.760 122.070 112.640 122.240 ;
        RECT 107.340 121.590 107.510 121.930 ;
        RECT 112.890 121.590 113.060 121.930 ;
        RECT 107.760 121.280 112.640 121.450 ;
        RECT 107.340 120.800 107.510 121.140 ;
        RECT 112.890 120.800 113.060 121.140 ;
        RECT 107.760 120.490 112.640 120.660 ;
        RECT 107.340 120.010 107.510 120.350 ;
        RECT 112.890 120.010 113.060 120.350 ;
        RECT 113.490 119.920 113.660 121.390 ;
        RECT 107.760 119.700 112.640 119.870 ;
        RECT 114.655 121.540 114.825 121.980 ;
        RECT 115.305 120.900 116.145 121.070 ;
        RECT 116.595 120.900 117.435 121.070 ;
        RECT 114.995 119.770 115.165 120.650 ;
        RECT 116.285 119.770 116.455 120.650 ;
        RECT 117.575 119.770 117.745 120.650 ;
        RECT 115.305 119.350 116.145 119.520 ;
        RECT 116.595 119.350 117.435 119.520 ;
        RECT 99.700 113.670 104.580 113.840 ;
        RECT 98.770 112.510 98.940 113.650 ;
        RECT 99.235 113.190 99.405 113.530 ;
        RECT 104.875 113.190 105.045 113.530 ;
        RECT 99.700 112.880 104.580 113.050 ;
        RECT 99.235 112.400 99.405 112.740 ;
        RECT 104.875 112.400 105.045 112.740 ;
        RECT 99.700 112.090 104.580 112.260 ;
        RECT 99.235 111.610 99.405 111.950 ;
        RECT 104.875 111.610 105.045 111.950 ;
        RECT 99.700 111.300 104.580 111.470 ;
        RECT 98.770 110.110 98.940 111.250 ;
        RECT 99.235 110.820 99.405 111.160 ;
        RECT 104.875 110.820 105.045 111.160 ;
        RECT 99.700 110.510 104.580 110.680 ;
        RECT 99.235 110.030 99.405 110.370 ;
        RECT 104.875 110.030 105.045 110.370 ;
        RECT 99.700 109.720 104.580 109.890 ;
        RECT 99.235 109.240 99.405 109.580 ;
        RECT 104.875 109.240 105.045 109.580 ;
        RECT 99.700 108.930 104.580 109.100 ;
        RECT 98.770 107.670 98.940 108.810 ;
        RECT 99.235 108.450 99.405 108.790 ;
        RECT 104.875 108.450 105.045 108.790 ;
        RECT 99.700 108.140 104.580 108.310 ;
        RECT 99.235 107.660 99.405 108.000 ;
        RECT 104.875 107.660 105.045 108.000 ;
        RECT 99.700 107.350 104.580 107.520 ;
        RECT 99.235 106.870 99.405 107.210 ;
        RECT 104.875 106.870 105.045 107.210 ;
        RECT 99.700 106.560 104.580 106.730 ;
        RECT 15.080 75.560 15.420 77.545 ;
        RECT 16.710 75.560 17.050 77.545 ;
        RECT 98.770 105.370 98.940 106.510 ;
        RECT 99.235 106.080 99.405 106.420 ;
        RECT 104.875 106.080 105.045 106.420 ;
        RECT 99.700 105.770 104.580 105.940 ;
        RECT 99.235 105.290 99.405 105.630 ;
        RECT 104.875 105.290 105.045 105.630 ;
        RECT 99.700 104.980 104.580 105.150 ;
        RECT 99.235 104.500 99.405 104.840 ;
        RECT 104.875 104.500 105.045 104.840 ;
        RECT 98.770 103.130 98.940 104.270 ;
        RECT 99.700 104.190 104.580 104.360 ;
        RECT 99.235 103.710 99.405 104.050 ;
        RECT 104.875 103.710 105.045 104.050 ;
        RECT 99.700 103.400 104.580 103.570 ;
        RECT 99.235 102.920 99.405 103.260 ;
        RECT 104.875 102.920 105.045 103.260 ;
        RECT 99.700 102.610 104.580 102.780 ;
        RECT 107.760 117.440 112.640 117.610 ;
        RECT 107.340 116.960 107.510 117.300 ;
        RECT 112.890 116.960 113.060 117.300 ;
        RECT 107.760 116.650 112.640 116.820 ;
        RECT 107.340 116.170 107.510 116.510 ;
        RECT 112.890 116.170 113.060 116.510 ;
        RECT 107.760 115.860 112.640 116.030 ;
        RECT 113.490 115.920 113.660 117.390 ;
        RECT 107.340 115.380 107.510 115.720 ;
        RECT 112.890 115.380 113.060 115.720 ;
        RECT 107.760 115.070 112.640 115.240 ;
        RECT 107.340 114.590 107.510 114.930 ;
        RECT 112.890 114.590 113.060 114.930 ;
        RECT 114.655 117.480 114.825 117.920 ;
        RECT 115.305 116.840 116.145 117.010 ;
        RECT 116.595 116.840 117.435 117.010 ;
        RECT 114.995 115.710 115.165 116.590 ;
        RECT 116.285 115.710 116.455 116.590 ;
        RECT 117.575 115.710 117.745 116.590 ;
        RECT 115.305 115.290 116.145 115.460 ;
        RECT 116.595 115.290 117.435 115.460 ;
        RECT 107.760 114.280 112.640 114.450 ;
        RECT 107.340 113.800 107.510 114.140 ;
        RECT 112.890 113.800 113.060 114.140 ;
        RECT 107.760 113.490 112.640 113.660 ;
        RECT 107.340 113.010 107.510 113.350 ;
        RECT 112.890 113.010 113.060 113.350 ;
        RECT 113.490 113.350 113.660 114.820 ;
        RECT 107.760 112.700 112.640 112.870 ;
        RECT 107.340 112.220 107.510 112.560 ;
        RECT 112.890 112.220 113.060 112.560 ;
        RECT 107.760 111.910 112.640 112.080 ;
        RECT 107.340 111.430 107.510 111.770 ;
        RECT 112.890 111.430 113.060 111.770 ;
        RECT 107.760 111.120 112.640 111.290 ;
        RECT 107.340 110.640 107.510 110.980 ;
        RECT 112.890 110.640 113.060 110.980 ;
        RECT 113.490 110.770 113.660 112.240 ;
        RECT 114.655 113.420 114.825 113.860 ;
        RECT 115.305 112.780 116.145 112.950 ;
        RECT 116.595 112.780 117.435 112.950 ;
        RECT 114.995 111.650 115.165 112.530 ;
        RECT 116.285 111.650 116.455 112.530 ;
        RECT 117.575 111.650 117.745 112.530 ;
        RECT 115.305 111.230 116.145 111.400 ;
        RECT 116.595 111.230 117.435 111.400 ;
        RECT 107.760 110.330 112.640 110.500 ;
        RECT 107.340 109.850 107.510 110.190 ;
        RECT 112.890 109.850 113.060 110.190 ;
        RECT 107.760 109.540 112.640 109.710 ;
        RECT 107.340 109.060 107.510 109.400 ;
        RECT 112.890 109.060 113.060 109.400 ;
        RECT 107.760 108.750 112.640 108.920 ;
        RECT 107.340 108.270 107.510 108.610 ;
        RECT 112.890 108.270 113.060 108.610 ;
        RECT 113.490 108.250 113.660 109.720 ;
        RECT 107.760 107.960 112.640 108.130 ;
        RECT 107.340 107.480 107.510 107.820 ;
        RECT 112.890 107.480 113.060 107.820 ;
        RECT 107.760 107.170 112.640 107.340 ;
        RECT 107.340 106.690 107.510 107.030 ;
        RECT 112.890 106.690 113.060 107.030 ;
        RECT 107.760 106.380 112.640 106.550 ;
        RECT 107.340 105.900 107.510 106.240 ;
        RECT 112.890 105.900 113.060 106.240 ;
        RECT 113.490 105.900 113.660 107.370 ;
        RECT 114.655 109.360 114.825 109.800 ;
        RECT 115.305 108.720 116.145 108.890 ;
        RECT 116.595 108.720 117.435 108.890 ;
        RECT 114.995 107.590 115.165 108.470 ;
        RECT 116.285 107.590 116.455 108.470 ;
        RECT 117.575 107.590 117.745 108.470 ;
        RECT 115.305 107.170 116.145 107.340 ;
        RECT 116.595 107.170 117.435 107.340 ;
        RECT 107.760 105.590 112.640 105.760 ;
        RECT 107.340 105.110 107.510 105.450 ;
        RECT 112.890 105.110 113.060 105.450 ;
        RECT 107.760 104.800 112.640 104.970 ;
        RECT 107.340 104.320 107.510 104.660 ;
        RECT 112.890 104.320 113.060 104.660 ;
        RECT 107.760 104.010 112.640 104.180 ;
        RECT 107.340 103.530 107.510 103.870 ;
        RECT 112.890 103.530 113.060 103.870 ;
        RECT 107.760 103.220 112.640 103.390 ;
        RECT 107.340 102.740 107.510 103.080 ;
        RECT 112.890 102.740 113.060 103.080 ;
        RECT 113.490 103.070 113.660 104.540 ;
        RECT 114.655 105.300 114.825 105.740 ;
        RECT 115.305 104.660 116.145 104.830 ;
        RECT 116.595 104.660 117.435 104.830 ;
        RECT 114.995 103.530 115.165 104.410 ;
        RECT 116.285 103.530 116.455 104.410 ;
        RECT 117.575 103.530 117.745 104.410 ;
        RECT 115.305 103.110 116.145 103.280 ;
        RECT 116.595 103.110 117.435 103.280 ;
        RECT 107.760 102.430 112.640 102.600 ;
        RECT 114.655 101.240 114.825 101.680 ;
        RECT 95.180 99.420 95.350 100.560 ;
        RECT 96.150 100.305 103.030 100.475 ;
        RECT 95.685 99.825 95.855 100.165 ;
        RECT 103.325 99.825 103.495 100.165 ;
        RECT 96.150 99.515 103.030 99.685 ;
        RECT 115.305 100.600 116.145 100.770 ;
        RECT 116.595 100.600 117.435 100.770 ;
        RECT 114.995 99.470 115.165 100.350 ;
        RECT 116.285 99.470 116.455 100.350 ;
        RECT 117.575 99.470 117.745 100.350 ;
        RECT 115.305 99.050 116.145 99.220 ;
        RECT 116.595 99.050 117.435 99.220 ;
        RECT 95.180 97.490 95.350 98.630 ;
        RECT 96.150 98.375 103.030 98.545 ;
        RECT 95.685 97.895 95.855 98.235 ;
        RECT 103.325 97.895 103.495 98.235 ;
        RECT 96.150 97.585 103.030 97.755 ;
        RECT 119.495 133.695 120.335 133.865 ;
        RECT 120.785 133.695 121.625 133.865 ;
        RECT 119.185 131.520 119.355 133.400 ;
        RECT 120.475 131.520 120.645 133.400 ;
        RECT 121.765 131.520 121.935 133.400 ;
        RECT 119.495 131.055 120.335 131.225 ;
        RECT 120.785 131.055 121.625 131.225 ;
        RECT 122.425 130.530 122.605 134.200 ;
        RECT 119.495 129.635 120.335 129.805 ;
        RECT 120.785 129.635 121.625 129.805 ;
        RECT 119.185 127.460 119.355 129.340 ;
        RECT 120.475 127.460 120.645 129.340 ;
        RECT 121.765 127.460 121.935 129.340 ;
        RECT 119.495 126.995 120.335 127.165 ;
        RECT 120.785 126.995 121.625 127.165 ;
        RECT 122.425 126.470 122.605 130.140 ;
        RECT 122.895 128.155 123.075 131.825 ;
        RECT 123.875 131.130 124.715 131.300 ;
        RECT 125.165 131.130 126.005 131.300 ;
        RECT 123.565 128.955 123.735 130.835 ;
        RECT 124.855 128.955 125.025 130.835 ;
        RECT 126.145 128.955 126.315 130.835 ;
        RECT 123.875 128.490 124.715 128.660 ;
        RECT 125.165 128.490 126.005 128.660 ;
        RECT 128.065 130.655 128.905 130.825 ;
        RECT 129.355 130.655 130.195 130.825 ;
        RECT 127.755 129.525 127.925 130.405 ;
        RECT 129.045 129.525 129.215 130.405 ;
        RECT 130.335 129.525 130.505 130.405 ;
        RECT 128.065 129.105 128.905 129.275 ;
        RECT 129.355 129.105 130.195 129.275 ;
        RECT 130.675 128.195 130.845 128.635 ;
        RECT 119.495 125.575 120.335 125.745 ;
        RECT 120.785 125.575 121.625 125.745 ;
        RECT 119.185 123.400 119.355 125.280 ;
        RECT 120.475 123.400 120.645 125.280 ;
        RECT 121.765 123.400 121.935 125.280 ;
        RECT 119.495 122.935 120.335 123.105 ;
        RECT 120.785 122.935 121.625 123.105 ;
        RECT 122.425 122.410 122.605 126.080 ;
        RECT 119.495 121.515 120.335 121.685 ;
        RECT 120.785 121.515 121.625 121.685 ;
        RECT 119.185 119.340 119.355 121.220 ;
        RECT 120.475 119.340 120.645 121.220 ;
        RECT 121.765 119.340 121.935 121.220 ;
        RECT 119.495 118.875 120.335 119.045 ;
        RECT 120.785 118.875 121.625 119.045 ;
        RECT 122.425 118.350 122.605 122.020 ;
        RECT 122.895 120.055 123.075 123.725 ;
        RECT 123.875 123.030 124.715 123.200 ;
        RECT 125.165 123.030 126.005 123.200 ;
        RECT 123.565 120.855 123.735 122.735 ;
        RECT 124.855 120.855 125.025 122.735 ;
        RECT 126.145 120.855 126.315 122.735 ;
        RECT 123.875 120.390 124.715 120.560 ;
        RECT 125.165 120.390 126.005 120.560 ;
        RECT 128.065 122.555 128.905 122.725 ;
        RECT 129.355 122.555 130.195 122.725 ;
        RECT 127.755 121.425 127.925 122.305 ;
        RECT 129.045 121.425 129.215 122.305 ;
        RECT 130.335 121.425 130.505 122.305 ;
        RECT 128.065 121.005 128.905 121.175 ;
        RECT 129.355 121.005 130.195 121.175 ;
        RECT 130.675 120.095 130.845 120.535 ;
        RECT 119.495 117.455 120.335 117.625 ;
        RECT 120.785 117.455 121.625 117.625 ;
        RECT 119.185 115.280 119.355 117.160 ;
        RECT 120.475 115.280 120.645 117.160 ;
        RECT 121.765 115.280 121.935 117.160 ;
        RECT 119.495 114.815 120.335 114.985 ;
        RECT 120.785 114.815 121.625 114.985 ;
        RECT 122.425 114.290 122.605 117.960 ;
        RECT 119.495 113.395 120.335 113.565 ;
        RECT 120.785 113.395 121.625 113.565 ;
        RECT 119.185 111.220 119.355 113.100 ;
        RECT 120.475 111.220 120.645 113.100 ;
        RECT 121.765 111.220 121.935 113.100 ;
        RECT 119.495 110.755 120.335 110.925 ;
        RECT 120.785 110.755 121.625 110.925 ;
        RECT 122.425 110.230 122.605 113.900 ;
        RECT 122.895 111.955 123.075 115.625 ;
        RECT 123.875 114.930 124.715 115.100 ;
        RECT 125.165 114.930 126.005 115.100 ;
        RECT 123.565 112.755 123.735 114.635 ;
        RECT 124.855 112.755 125.025 114.635 ;
        RECT 126.145 112.755 126.315 114.635 ;
        RECT 123.875 112.290 124.715 112.460 ;
        RECT 125.165 112.290 126.005 112.460 ;
        RECT 128.065 114.455 128.905 114.625 ;
        RECT 129.355 114.455 130.195 114.625 ;
        RECT 127.755 113.325 127.925 114.205 ;
        RECT 129.045 113.325 129.215 114.205 ;
        RECT 130.335 113.325 130.505 114.205 ;
        RECT 128.065 112.905 128.905 113.075 ;
        RECT 129.355 112.905 130.195 113.075 ;
        RECT 130.675 111.995 130.845 112.435 ;
        RECT 119.495 109.335 120.335 109.505 ;
        RECT 120.785 109.335 121.625 109.505 ;
        RECT 119.185 107.160 119.355 109.040 ;
        RECT 120.475 107.160 120.645 109.040 ;
        RECT 121.765 107.160 121.935 109.040 ;
        RECT 119.495 106.695 120.335 106.865 ;
        RECT 120.785 106.695 121.625 106.865 ;
        RECT 122.425 106.170 122.605 109.840 ;
        RECT 119.495 105.275 120.335 105.445 ;
        RECT 120.785 105.275 121.625 105.445 ;
        RECT 119.185 103.100 119.355 104.980 ;
        RECT 120.475 103.100 120.645 104.980 ;
        RECT 121.765 103.100 121.935 104.980 ;
        RECT 119.495 102.635 120.335 102.805 ;
        RECT 120.785 102.635 121.625 102.805 ;
        RECT 122.425 102.110 122.605 105.780 ;
        RECT 119.495 101.215 120.335 101.385 ;
        RECT 120.785 101.215 121.625 101.385 ;
        RECT 119.185 99.040 119.355 100.920 ;
        RECT 120.475 99.040 120.645 100.920 ;
        RECT 121.765 99.040 121.935 100.920 ;
        RECT 119.495 98.575 120.335 98.745 ;
        RECT 120.785 98.575 121.625 98.745 ;
        RECT 122.425 98.050 122.605 101.720 ;
        RECT 122.895 103.855 123.075 107.525 ;
        RECT 123.875 106.830 124.715 107.000 ;
        RECT 125.165 106.830 126.005 107.000 ;
        RECT 123.565 104.655 123.735 106.535 ;
        RECT 124.855 104.655 125.025 106.535 ;
        RECT 126.145 104.655 126.315 106.535 ;
        RECT 123.875 104.190 124.715 104.360 ;
        RECT 125.165 104.190 126.005 104.360 ;
        RECT 122.895 99.805 123.075 103.475 ;
        RECT 123.875 102.780 124.715 102.950 ;
        RECT 125.165 102.780 126.005 102.950 ;
        RECT 123.565 100.605 123.735 102.485 ;
        RECT 124.855 100.605 125.025 102.485 ;
        RECT 126.145 100.605 126.315 102.485 ;
        RECT 123.875 100.140 124.715 100.310 ;
        RECT 125.165 100.140 126.005 100.310 ;
        RECT 95.860 96.570 97.000 96.740 ;
        RECT 97.830 96.570 102.780 96.740 ;
        RECT 94.680 95.120 94.850 96.260 ;
        RECT 95.655 96.000 103.035 96.170 ;
        RECT 95.190 95.520 95.360 95.860 ;
        RECT 103.330 95.520 103.500 95.860 ;
        RECT 95.655 95.210 103.035 95.380 ;
        RECT 104.815 96.000 105.695 96.170 ;
        RECT 104.350 95.520 104.520 95.860 ;
        RECT 105.990 95.520 106.160 95.860 ;
        RECT 104.815 95.210 105.695 95.380 ;
        RECT 95.570 94.640 96.140 94.810 ;
        RECT 107.960 96.505 112.840 96.675 ;
        RECT 107.540 95.525 107.710 96.365 ;
        RECT 113.090 95.525 113.260 96.365 ;
        RECT 107.960 95.215 112.840 95.385 ;
        RECT 113.600 95.120 113.770 96.760 ;
        RECT 122.895 95.755 123.075 99.425 ;
        RECT 123.875 98.730 124.715 98.900 ;
        RECT 125.165 98.730 126.005 98.900 ;
        RECT 123.565 96.555 123.735 98.435 ;
        RECT 124.855 96.555 125.025 98.435 ;
        RECT 126.145 96.555 126.315 98.435 ;
        RECT 123.875 96.090 124.715 96.260 ;
        RECT 125.165 96.090 126.005 96.260 ;
        RECT 80.330 93.840 81.390 94.020 ;
        RECT 72.100 81.610 72.280 93.280 ;
        RECT 73.110 91.610 77.990 91.780 ;
        RECT 82.110 91.610 86.990 91.780 ;
        RECT 72.645 91.130 72.815 91.470 ;
        RECT 78.285 91.130 78.455 91.470 ;
        RECT 81.645 91.130 81.815 91.470 ;
        RECT 87.285 91.130 87.455 91.470 ;
        RECT 73.110 90.820 77.990 90.990 ;
        RECT 82.110 90.820 86.990 90.990 ;
        RECT 73.110 87.110 77.990 87.280 ;
        RECT 82.110 87.110 86.990 87.280 ;
        RECT 72.645 86.630 72.815 86.970 ;
        RECT 78.285 86.630 78.455 86.970 ;
        RECT 81.645 86.630 81.815 86.970 ;
        RECT 87.285 86.630 87.455 86.970 ;
        RECT 73.110 86.320 77.990 86.490 ;
        RECT 82.110 86.320 86.990 86.490 ;
        RECT 73.110 82.610 77.990 82.780 ;
        RECT 82.110 82.610 86.990 82.780 ;
        RECT 72.645 82.130 72.815 82.470 ;
        RECT 78.285 82.130 78.455 82.470 ;
        RECT 81.645 82.130 81.815 82.470 ;
        RECT 87.285 82.130 87.455 82.470 ;
        RECT 73.110 81.820 77.990 81.990 ;
        RECT 82.110 81.820 86.990 81.990 ;
        RECT 90.830 92.090 95.710 92.260 ;
        RECT 97.830 92.090 102.710 92.260 ;
        RECT 90.410 91.110 90.580 91.950 ;
        RECT 95.960 91.110 96.130 91.950 ;
        RECT 97.410 91.110 97.580 91.950 ;
        RECT 102.960 91.110 103.130 91.950 ;
        RECT 90.830 90.800 95.710 90.970 ;
        RECT 97.830 90.800 102.710 90.970 ;
        RECT 90.830 90.090 95.710 90.260 ;
        RECT 97.830 90.090 102.710 90.260 ;
        RECT 90.410 89.110 90.580 89.950 ;
        RECT 95.960 89.110 96.130 89.950 ;
        RECT 97.410 89.110 97.580 89.950 ;
        RECT 102.960 89.110 103.130 89.950 ;
        RECT 90.830 88.800 95.710 88.970 ;
        RECT 97.830 88.800 102.710 88.970 ;
        RECT 90.830 86.090 95.710 86.260 ;
        RECT 97.830 86.090 102.710 86.260 ;
        RECT 90.410 85.110 90.580 85.950 ;
        RECT 95.960 85.110 96.130 85.950 ;
        RECT 97.410 85.110 97.580 85.950 ;
        RECT 102.960 85.110 103.130 85.950 ;
        RECT 90.830 84.800 95.710 84.970 ;
        RECT 97.830 84.800 102.710 84.970 ;
        RECT 90.830 84.090 95.710 84.260 ;
        RECT 97.830 84.090 102.710 84.260 ;
        RECT 90.410 83.110 90.580 83.950 ;
        RECT 95.960 83.110 96.130 83.950 ;
        RECT 97.410 83.110 97.580 83.950 ;
        RECT 102.960 83.110 103.130 83.950 ;
        RECT 90.830 82.800 95.710 82.970 ;
        RECT 97.830 82.800 102.710 82.970 ;
        RECT 104.260 81.810 104.430 84.020 ;
        RECT 106.290 93.400 111.170 93.570 ;
        RECT 105.870 92.420 106.040 93.260 ;
        RECT 111.420 92.420 111.590 93.260 ;
        RECT 106.290 92.110 111.170 92.280 ;
        RECT 105.870 91.130 106.040 91.970 ;
        RECT 111.420 91.130 111.590 91.970 ;
        RECT 106.290 90.820 111.170 90.990 ;
        RECT 105.870 89.840 106.040 90.680 ;
        RECT 111.420 89.840 111.590 90.680 ;
        RECT 106.290 89.530 111.170 89.700 ;
        RECT 105.870 88.550 106.040 89.390 ;
        RECT 111.420 88.550 111.590 89.390 ;
        RECT 106.290 88.240 111.170 88.410 ;
        RECT 105.870 87.260 106.040 88.100 ;
        RECT 111.420 87.260 111.590 88.100 ;
        RECT 106.290 86.950 111.170 87.120 ;
        RECT 105.870 85.970 106.040 86.810 ;
        RECT 111.420 85.970 111.590 86.810 ;
        RECT 106.290 85.660 111.170 85.830 ;
        RECT 105.870 84.680 106.040 85.520 ;
        RECT 111.420 84.680 111.590 85.520 ;
        RECT 106.290 84.370 111.170 84.540 ;
        RECT 105.870 83.390 106.040 84.230 ;
        RECT 111.420 83.390 111.590 84.230 ;
        RECT 106.290 83.080 111.170 83.250 ;
        RECT 113.520 82.950 113.690 92.660 ;
        RECT 114.655 93.120 114.825 93.560 ;
        RECT 115.305 92.480 116.145 92.650 ;
        RECT 116.595 92.480 117.435 92.650 ;
        RECT 114.995 91.350 115.165 92.230 ;
        RECT 116.285 91.350 116.455 92.230 ;
        RECT 117.575 91.350 117.745 92.230 ;
        RECT 115.305 90.930 116.145 91.100 ;
        RECT 116.595 90.930 117.435 91.100 ;
        RECT 114.655 89.060 114.825 89.500 ;
        RECT 115.305 88.420 116.145 88.590 ;
        RECT 116.595 88.420 117.435 88.590 ;
        RECT 114.995 87.290 115.165 88.170 ;
        RECT 116.285 87.290 116.455 88.170 ;
        RECT 117.575 87.290 117.745 88.170 ;
        RECT 115.305 86.870 116.145 87.040 ;
        RECT 116.595 86.870 117.435 87.040 ;
        RECT 114.655 85.000 114.825 85.440 ;
        RECT 115.305 84.360 116.145 84.530 ;
        RECT 116.595 84.360 117.435 84.530 ;
        RECT 114.995 83.230 115.165 84.110 ;
        RECT 116.285 83.230 116.455 84.110 ;
        RECT 117.575 83.230 117.745 84.110 ;
        RECT 115.305 82.810 116.145 82.980 ;
        RECT 116.595 82.810 117.435 82.980 ;
        RECT 80.660 81.000 81.280 81.180 ;
        RECT 114.655 80.940 114.825 81.380 ;
        RECT 56.700 76.310 61.580 76.480 ;
        RECT 55.770 75.150 55.940 76.290 ;
        RECT 56.235 75.830 56.405 76.170 ;
        RECT 61.875 75.830 62.045 76.170 ;
        RECT 56.700 75.520 61.580 75.690 ;
        RECT 15.080 45.130 15.420 47.115 ;
        RECT 16.710 45.130 17.050 47.115 ;
        RECT 20.820 45.130 21.160 47.115 ;
        RECT 22.450 45.130 22.790 47.115 ;
        RECT 24.080 45.130 24.420 47.115 ;
        RECT 25.710 45.130 26.050 47.115 ;
        RECT 56.235 75.040 56.405 75.380 ;
        RECT 61.875 75.040 62.045 75.380 ;
        RECT 56.700 74.730 61.580 74.900 ;
        RECT 56.235 74.250 56.405 74.590 ;
        RECT 61.875 74.250 62.045 74.590 ;
        RECT 56.700 73.940 61.580 74.110 ;
        RECT 55.770 72.750 55.940 73.890 ;
        RECT 56.235 73.460 56.405 73.800 ;
        RECT 61.875 73.460 62.045 73.800 ;
        RECT 56.700 73.150 61.580 73.320 ;
        RECT 56.235 72.670 56.405 73.010 ;
        RECT 61.875 72.670 62.045 73.010 ;
        RECT 56.700 72.360 61.580 72.530 ;
        RECT 56.235 71.880 56.405 72.220 ;
        RECT 61.875 71.880 62.045 72.220 ;
        RECT 56.700 71.570 61.580 71.740 ;
        RECT 55.770 70.310 55.940 71.450 ;
        RECT 56.235 71.090 56.405 71.430 ;
        RECT 61.875 71.090 62.045 71.430 ;
        RECT 56.700 70.780 61.580 70.950 ;
        RECT 56.235 70.300 56.405 70.640 ;
        RECT 61.875 70.300 62.045 70.640 ;
        RECT 56.700 69.990 61.580 70.160 ;
        RECT 56.235 69.510 56.405 69.850 ;
        RECT 61.875 69.510 62.045 69.850 ;
        RECT 56.700 69.200 61.580 69.370 ;
        RECT 55.770 68.010 55.940 69.150 ;
        RECT 56.235 68.720 56.405 69.060 ;
        RECT 61.875 68.720 62.045 69.060 ;
        RECT 56.700 68.410 61.580 68.580 ;
        RECT 56.235 67.930 56.405 68.270 ;
        RECT 61.875 67.930 62.045 68.270 ;
        RECT 56.700 67.620 61.580 67.790 ;
        RECT 56.235 67.140 56.405 67.480 ;
        RECT 61.875 67.140 62.045 67.480 ;
        RECT 55.770 65.770 55.940 66.910 ;
        RECT 56.700 66.830 61.580 67.000 ;
        RECT 56.235 66.350 56.405 66.690 ;
        RECT 61.875 66.350 62.045 66.690 ;
        RECT 56.700 66.040 61.580 66.210 ;
        RECT 56.235 65.560 56.405 65.900 ;
        RECT 61.875 65.560 62.045 65.900 ;
        RECT 56.700 65.250 61.580 65.420 ;
        RECT 64.760 80.080 69.640 80.250 ;
        RECT 64.340 79.600 64.510 79.940 ;
        RECT 69.890 79.600 70.060 79.940 ;
        RECT 64.760 79.290 69.640 79.460 ;
        RECT 64.340 78.810 64.510 79.150 ;
        RECT 69.890 78.810 70.060 79.150 ;
        RECT 64.760 78.500 69.640 78.670 ;
        RECT 70.490 78.560 70.660 80.030 ;
        RECT 64.340 78.020 64.510 78.360 ;
        RECT 69.890 78.020 70.060 78.360 ;
        RECT 64.760 77.710 69.640 77.880 ;
        RECT 64.340 77.230 64.510 77.570 ;
        RECT 69.890 77.230 70.060 77.570 ;
        RECT 64.760 76.920 69.640 77.090 ;
        RECT 64.340 76.440 64.510 76.780 ;
        RECT 69.890 76.440 70.060 76.780 ;
        RECT 64.760 76.130 69.640 76.300 ;
        RECT 64.340 75.650 64.510 75.990 ;
        RECT 69.890 75.650 70.060 75.990 ;
        RECT 70.490 75.990 70.660 77.460 ;
        RECT 64.760 75.340 69.640 75.510 ;
        RECT 64.340 74.860 64.510 75.200 ;
        RECT 69.890 74.860 70.060 75.200 ;
        RECT 64.760 74.550 69.640 74.720 ;
        RECT 64.340 74.070 64.510 74.410 ;
        RECT 69.890 74.070 70.060 74.410 ;
        RECT 64.760 73.760 69.640 73.930 ;
        RECT 64.340 73.280 64.510 73.620 ;
        RECT 69.890 73.280 70.060 73.620 ;
        RECT 70.490 73.410 70.660 74.880 ;
        RECT 64.760 72.970 69.640 73.140 ;
        RECT 64.340 72.490 64.510 72.830 ;
        RECT 69.890 72.490 70.060 72.830 ;
        RECT 64.760 72.180 69.640 72.350 ;
        RECT 64.340 71.700 64.510 72.040 ;
        RECT 69.890 71.700 70.060 72.040 ;
        RECT 64.760 71.390 69.640 71.560 ;
        RECT 64.340 70.910 64.510 71.250 ;
        RECT 69.890 70.910 70.060 71.250 ;
        RECT 70.490 70.890 70.660 72.360 ;
        RECT 64.760 70.600 69.640 70.770 ;
        RECT 64.340 70.120 64.510 70.460 ;
        RECT 69.890 70.120 70.060 70.460 ;
        RECT 64.760 69.810 69.640 69.980 ;
        RECT 64.340 69.330 64.510 69.670 ;
        RECT 69.890 69.330 70.060 69.670 ;
        RECT 64.760 69.020 69.640 69.190 ;
        RECT 64.340 68.540 64.510 68.880 ;
        RECT 69.890 68.540 70.060 68.880 ;
        RECT 70.490 68.540 70.660 70.010 ;
        RECT 64.760 68.230 69.640 68.400 ;
        RECT 64.340 67.750 64.510 68.090 ;
        RECT 69.890 67.750 70.060 68.090 ;
        RECT 64.760 67.440 69.640 67.610 ;
        RECT 64.340 66.960 64.510 67.300 ;
        RECT 69.890 66.960 70.060 67.300 ;
        RECT 80.660 80.530 81.280 80.710 ;
        RECT 72.100 68.430 72.280 80.100 ;
        RECT 73.110 79.720 77.990 79.890 ;
        RECT 82.110 79.720 86.990 79.890 ;
        RECT 72.645 79.240 72.815 79.580 ;
        RECT 78.285 79.240 78.455 79.580 ;
        RECT 81.645 79.240 81.815 79.580 ;
        RECT 87.285 79.240 87.455 79.580 ;
        RECT 73.110 78.930 77.990 79.100 ;
        RECT 82.110 78.930 86.990 79.100 ;
        RECT 73.110 75.220 77.990 75.390 ;
        RECT 82.110 75.220 86.990 75.390 ;
        RECT 72.645 74.740 72.815 75.080 ;
        RECT 78.285 74.740 78.455 75.080 ;
        RECT 81.645 74.740 81.815 75.080 ;
        RECT 87.285 74.740 87.455 75.080 ;
        RECT 73.110 74.430 77.990 74.600 ;
        RECT 82.110 74.430 86.990 74.600 ;
        RECT 73.110 70.720 77.990 70.890 ;
        RECT 82.110 70.720 86.990 70.890 ;
        RECT 72.645 70.240 72.815 70.580 ;
        RECT 78.285 70.240 78.455 70.580 ;
        RECT 81.645 70.240 81.815 70.580 ;
        RECT 87.285 70.240 87.455 70.580 ;
        RECT 73.110 69.930 77.990 70.100 ;
        RECT 82.110 69.930 86.990 70.100 ;
        RECT 80.330 67.690 81.390 67.870 ;
        RECT 90.830 78.740 95.710 78.910 ;
        RECT 97.830 78.740 102.710 78.910 ;
        RECT 90.410 77.760 90.580 78.600 ;
        RECT 95.960 77.760 96.130 78.600 ;
        RECT 97.410 77.760 97.580 78.600 ;
        RECT 102.960 77.760 103.130 78.600 ;
        RECT 104.260 77.690 104.430 79.900 ;
        RECT 90.830 77.450 95.710 77.620 ;
        RECT 97.830 77.450 102.710 77.620 ;
        RECT 90.830 76.740 95.710 76.910 ;
        RECT 97.830 76.740 102.710 76.910 ;
        RECT 90.410 75.760 90.580 76.600 ;
        RECT 95.960 75.760 96.130 76.600 ;
        RECT 97.410 75.760 97.580 76.600 ;
        RECT 102.960 75.760 103.130 76.600 ;
        RECT 90.830 75.450 95.710 75.620 ;
        RECT 97.830 75.450 102.710 75.620 ;
        RECT 90.830 72.740 95.710 72.910 ;
        RECT 97.830 72.740 102.710 72.910 ;
        RECT 90.410 71.760 90.580 72.600 ;
        RECT 95.960 71.760 96.130 72.600 ;
        RECT 97.410 71.760 97.580 72.600 ;
        RECT 102.960 71.760 103.130 72.600 ;
        RECT 90.830 71.450 95.710 71.620 ;
        RECT 97.830 71.450 102.710 71.620 ;
        RECT 90.830 70.740 95.710 70.910 ;
        RECT 97.830 70.740 102.710 70.910 ;
        RECT 90.410 69.760 90.580 70.600 ;
        RECT 95.960 69.760 96.130 70.600 ;
        RECT 97.410 69.760 97.580 70.600 ;
        RECT 102.960 69.760 103.130 70.600 ;
        RECT 90.830 69.450 95.710 69.620 ;
        RECT 97.830 69.450 102.710 69.620 ;
        RECT 106.290 78.460 111.170 78.630 ;
        RECT 105.870 77.480 106.040 78.320 ;
        RECT 111.420 77.480 111.590 78.320 ;
        RECT 106.290 77.170 111.170 77.340 ;
        RECT 105.870 76.190 106.040 77.030 ;
        RECT 111.420 76.190 111.590 77.030 ;
        RECT 106.290 75.880 111.170 76.050 ;
        RECT 105.870 74.900 106.040 75.740 ;
        RECT 111.420 74.900 111.590 75.740 ;
        RECT 106.290 74.590 111.170 74.760 ;
        RECT 105.870 73.610 106.040 74.450 ;
        RECT 111.420 73.610 111.590 74.450 ;
        RECT 106.290 73.300 111.170 73.470 ;
        RECT 105.870 72.320 106.040 73.160 ;
        RECT 111.420 72.320 111.590 73.160 ;
        RECT 106.290 72.010 111.170 72.180 ;
        RECT 105.870 71.030 106.040 71.870 ;
        RECT 111.420 71.030 111.590 71.870 ;
        RECT 106.290 70.720 111.170 70.890 ;
        RECT 105.870 69.740 106.040 70.580 ;
        RECT 111.420 69.740 111.590 70.580 ;
        RECT 106.290 69.430 111.170 69.600 ;
        RECT 105.870 68.450 106.040 69.290 ;
        RECT 111.420 68.450 111.590 69.290 ;
        RECT 113.520 69.050 113.690 78.760 ;
        RECT 115.305 80.300 116.145 80.470 ;
        RECT 116.595 80.300 117.435 80.470 ;
        RECT 114.995 79.170 115.165 80.050 ;
        RECT 116.285 79.170 116.455 80.050 ;
        RECT 117.575 79.170 117.745 80.050 ;
        RECT 115.305 78.750 116.145 78.920 ;
        RECT 116.595 78.750 117.435 78.920 ;
        RECT 114.655 76.880 114.825 77.320 ;
        RECT 115.305 76.240 116.145 76.410 ;
        RECT 116.595 76.240 117.435 76.410 ;
        RECT 114.995 75.110 115.165 75.990 ;
        RECT 116.285 75.110 116.455 75.990 ;
        RECT 117.575 75.110 117.745 75.990 ;
        RECT 115.305 74.690 116.145 74.860 ;
        RECT 116.595 74.690 117.435 74.860 ;
        RECT 119.495 93.095 120.335 93.265 ;
        RECT 120.785 93.095 121.625 93.265 ;
        RECT 119.185 90.920 119.355 92.800 ;
        RECT 120.475 90.920 120.645 92.800 ;
        RECT 121.765 90.920 121.935 92.800 ;
        RECT 119.495 90.455 120.335 90.625 ;
        RECT 120.785 90.455 121.625 90.625 ;
        RECT 122.425 89.930 122.605 93.600 ;
        RECT 119.495 89.035 120.335 89.205 ;
        RECT 120.785 89.035 121.625 89.205 ;
        RECT 119.185 86.860 119.355 88.740 ;
        RECT 120.475 86.860 120.645 88.740 ;
        RECT 121.765 86.860 121.935 88.740 ;
        RECT 119.495 86.395 120.335 86.565 ;
        RECT 120.785 86.395 121.625 86.565 ;
        RECT 122.425 85.870 122.605 89.540 ;
        RECT 119.495 84.975 120.335 85.145 ;
        RECT 120.785 84.975 121.625 85.145 ;
        RECT 119.185 82.800 119.355 84.680 ;
        RECT 120.475 82.800 120.645 84.680 ;
        RECT 121.765 82.800 121.935 84.680 ;
        RECT 119.495 82.335 120.335 82.505 ;
        RECT 120.785 82.335 121.625 82.505 ;
        RECT 122.425 81.810 122.605 85.480 ;
        RECT 119.495 80.915 120.335 81.085 ;
        RECT 120.785 80.915 121.625 81.085 ;
        RECT 119.185 78.740 119.355 80.620 ;
        RECT 120.475 78.740 120.645 80.620 ;
        RECT 121.765 78.740 121.935 80.620 ;
        RECT 119.495 78.275 120.335 78.445 ;
        RECT 120.785 78.275 121.625 78.445 ;
        RECT 122.425 77.750 122.605 81.420 ;
        RECT 119.495 76.855 120.335 77.025 ;
        RECT 120.785 76.855 121.625 77.025 ;
        RECT 119.185 74.680 119.355 76.560 ;
        RECT 120.475 74.680 120.645 76.560 ;
        RECT 121.765 74.680 121.935 76.560 ;
        RECT 119.495 74.215 120.335 74.385 ;
        RECT 120.785 74.215 121.625 74.385 ;
        RECT 122.425 73.690 122.605 77.360 ;
        RECT 122.895 91.705 123.075 95.375 ;
        RECT 123.875 94.680 124.715 94.850 ;
        RECT 125.165 94.680 126.005 94.850 ;
        RECT 123.565 92.505 123.735 94.385 ;
        RECT 124.855 92.505 125.025 94.385 ;
        RECT 126.145 92.505 126.315 94.385 ;
        RECT 123.875 92.040 124.715 92.210 ;
        RECT 125.165 92.040 126.005 92.210 ;
        RECT 122.895 87.655 123.075 91.325 ;
        RECT 123.875 90.630 124.715 90.800 ;
        RECT 125.165 90.630 126.005 90.800 ;
        RECT 123.565 88.455 123.735 90.335 ;
        RECT 124.855 88.455 125.025 90.335 ;
        RECT 126.145 88.455 126.315 90.335 ;
        RECT 123.875 87.990 124.715 88.160 ;
        RECT 125.165 87.990 126.005 88.160 ;
        RECT 122.895 83.605 123.075 87.275 ;
        RECT 123.875 86.580 124.715 86.750 ;
        RECT 125.165 86.580 126.005 86.750 ;
        RECT 123.565 84.405 123.735 86.285 ;
        RECT 124.855 84.405 125.025 86.285 ;
        RECT 126.145 84.405 126.315 86.285 ;
        RECT 123.875 83.940 124.715 84.110 ;
        RECT 125.165 83.940 126.005 84.110 ;
        RECT 122.895 79.555 123.075 83.225 ;
        RECT 123.875 82.530 124.715 82.700 ;
        RECT 125.165 82.530 126.005 82.700 ;
        RECT 123.565 80.355 123.735 82.235 ;
        RECT 124.855 80.355 125.025 82.235 ;
        RECT 126.145 80.355 126.315 82.235 ;
        RECT 123.875 79.890 124.715 80.060 ;
        RECT 125.165 79.890 126.005 80.060 ;
        RECT 122.895 75.505 123.075 79.175 ;
        RECT 123.875 78.480 124.715 78.650 ;
        RECT 125.165 78.480 126.005 78.650 ;
        RECT 123.565 76.305 123.735 78.185 ;
        RECT 124.855 76.305 125.025 78.185 ;
        RECT 126.145 76.305 126.315 78.185 ;
        RECT 123.875 75.840 124.715 76.010 ;
        RECT 125.165 75.840 126.005 76.010 ;
        RECT 106.290 68.140 111.170 68.310 ;
        RECT 122.895 71.455 123.075 75.125 ;
        RECT 123.875 74.430 124.715 74.600 ;
        RECT 125.165 74.430 126.005 74.600 ;
        RECT 123.565 72.255 123.735 74.135 ;
        RECT 124.855 72.255 125.025 74.135 ;
        RECT 126.145 72.255 126.315 74.135 ;
        RECT 123.875 71.790 124.715 71.960 ;
        RECT 125.165 71.790 126.005 71.960 ;
        RECT 64.760 66.650 69.640 66.820 ;
        RECT 64.340 66.170 64.510 66.510 ;
        RECT 69.890 66.170 70.060 66.510 ;
        RECT 64.760 65.860 69.640 66.030 ;
        RECT 64.340 65.380 64.510 65.720 ;
        RECT 69.890 65.380 70.060 65.720 ;
        RECT 70.490 65.710 70.660 67.180 ;
        RECT 122.895 67.370 123.075 71.040 ;
        RECT 123.875 70.345 124.715 70.515 ;
        RECT 125.165 70.345 126.005 70.515 ;
        RECT 123.565 68.170 123.735 70.050 ;
        RECT 124.855 68.170 125.025 70.050 ;
        RECT 126.145 68.170 126.315 70.050 ;
        RECT 123.875 67.705 124.715 67.875 ;
        RECT 125.165 67.705 126.005 67.875 ;
        RECT 64.760 65.070 69.640 65.240 ;
        RECT 95.570 66.900 96.140 67.070 ;
        RECT 94.680 65.450 94.850 66.590 ;
        RECT 95.655 66.330 103.035 66.500 ;
        RECT 95.190 65.850 95.360 66.190 ;
        RECT 103.330 65.850 103.500 66.190 ;
        RECT 95.655 65.540 103.035 65.710 ;
        RECT 104.815 66.330 105.695 66.500 ;
        RECT 104.350 65.850 104.520 66.190 ;
        RECT 105.990 65.850 106.160 66.190 ;
        RECT 104.815 65.540 105.695 65.710 ;
        RECT 95.860 64.970 97.000 65.140 ;
        RECT 97.830 64.970 102.780 65.140 ;
        RECT 108.420 66.900 109.060 67.070 ;
        RECT 109.600 66.900 110.240 67.070 ;
        RECT 111.000 66.900 111.640 67.070 ;
        RECT 112.650 66.900 113.290 67.070 ;
        RECT 97.830 64.530 102.780 64.700 ;
        RECT 52.180 62.060 52.350 63.200 ;
        RECT 53.150 62.945 60.030 63.115 ;
        RECT 52.685 62.465 52.855 62.805 ;
        RECT 60.325 62.465 60.495 62.805 ;
        RECT 53.150 62.155 60.030 62.325 ;
        RECT 52.180 60.130 52.350 61.270 ;
        RECT 53.150 61.015 60.030 61.185 ;
        RECT 52.685 60.535 52.855 60.875 ;
        RECT 60.325 60.535 60.495 60.875 ;
        RECT 53.150 60.225 60.030 60.395 ;
        RECT 95.180 63.080 95.350 64.220 ;
        RECT 96.150 63.955 103.030 64.125 ;
        RECT 95.685 63.475 95.855 63.815 ;
        RECT 103.325 63.475 103.495 63.815 ;
        RECT 96.150 63.165 103.030 63.335 ;
        RECT 107.960 66.325 112.840 66.495 ;
        RECT 107.540 65.345 107.710 66.185 ;
        RECT 113.090 65.345 113.260 66.185 ;
        RECT 107.960 65.035 112.840 65.205 ;
        RECT 113.600 64.950 113.770 66.590 ;
        RECT 122.895 63.245 123.075 66.915 ;
        RECT 123.875 66.220 124.715 66.390 ;
        RECT 125.165 66.220 126.005 66.390 ;
        RECT 123.565 64.045 123.735 65.925 ;
        RECT 124.855 64.045 125.025 65.925 ;
        RECT 126.145 64.045 126.315 65.925 ;
        RECT 123.875 63.580 124.715 63.750 ;
        RECT 125.165 63.580 126.005 63.750 ;
        RECT 128.065 106.355 128.905 106.525 ;
        RECT 129.355 106.355 130.195 106.525 ;
        RECT 127.755 105.225 127.925 106.105 ;
        RECT 129.045 105.225 129.215 106.105 ;
        RECT 130.335 105.225 130.505 106.105 ;
        RECT 128.065 104.805 128.905 104.975 ;
        RECT 129.355 104.805 130.195 104.975 ;
        RECT 130.675 103.895 130.845 104.335 ;
        RECT 128.065 102.305 128.905 102.475 ;
        RECT 129.355 102.305 130.195 102.475 ;
        RECT 127.755 101.175 127.925 102.055 ;
        RECT 129.045 101.175 129.215 102.055 ;
        RECT 130.335 101.175 130.505 102.055 ;
        RECT 128.065 100.755 128.905 100.925 ;
        RECT 129.355 100.755 130.195 100.925 ;
        RECT 130.675 99.845 130.845 100.285 ;
        RECT 128.065 98.255 128.905 98.425 ;
        RECT 129.355 98.255 130.195 98.425 ;
        RECT 127.755 97.125 127.925 98.005 ;
        RECT 129.045 97.125 129.215 98.005 ;
        RECT 130.335 97.125 130.505 98.005 ;
        RECT 128.065 96.705 128.905 96.875 ;
        RECT 129.355 96.705 130.195 96.875 ;
        RECT 130.675 95.795 130.845 96.235 ;
        RECT 128.065 94.205 128.905 94.375 ;
        RECT 129.355 94.205 130.195 94.375 ;
        RECT 127.755 93.075 127.925 93.955 ;
        RECT 129.045 93.075 129.215 93.955 ;
        RECT 130.335 93.075 130.505 93.955 ;
        RECT 128.065 92.655 128.905 92.825 ;
        RECT 129.355 92.655 130.195 92.825 ;
        RECT 130.675 91.745 130.845 92.185 ;
        RECT 128.065 90.155 128.905 90.325 ;
        RECT 129.355 90.155 130.195 90.325 ;
        RECT 127.755 89.025 127.925 89.905 ;
        RECT 129.045 89.025 129.215 89.905 ;
        RECT 130.335 89.025 130.505 89.905 ;
        RECT 128.065 88.605 128.905 88.775 ;
        RECT 129.355 88.605 130.195 88.775 ;
        RECT 130.675 87.695 130.845 88.135 ;
        RECT 128.065 86.105 128.905 86.275 ;
        RECT 129.355 86.105 130.195 86.275 ;
        RECT 127.755 84.975 127.925 85.855 ;
        RECT 129.045 84.975 129.215 85.855 ;
        RECT 130.335 84.975 130.505 85.855 ;
        RECT 128.065 84.555 128.905 84.725 ;
        RECT 129.355 84.555 130.195 84.725 ;
        RECT 130.675 83.645 130.845 84.085 ;
        RECT 128.065 82.055 128.905 82.225 ;
        RECT 129.355 82.055 130.195 82.225 ;
        RECT 127.755 80.925 127.925 81.805 ;
        RECT 129.045 80.925 129.215 81.805 ;
        RECT 130.335 80.925 130.505 81.805 ;
        RECT 128.065 80.505 128.905 80.675 ;
        RECT 129.355 80.505 130.195 80.675 ;
        RECT 130.675 79.595 130.845 80.035 ;
        RECT 128.065 78.005 128.905 78.175 ;
        RECT 129.355 78.005 130.195 78.175 ;
        RECT 127.755 76.875 127.925 77.755 ;
        RECT 129.045 76.875 129.215 77.755 ;
        RECT 130.335 76.875 130.505 77.755 ;
        RECT 128.065 76.455 128.905 76.625 ;
        RECT 129.355 76.455 130.195 76.625 ;
        RECT 130.675 75.545 130.845 75.985 ;
        RECT 128.065 73.955 128.905 74.125 ;
        RECT 129.355 73.955 130.195 74.125 ;
        RECT 127.755 72.825 127.925 73.705 ;
        RECT 129.045 72.825 129.215 73.705 ;
        RECT 130.335 72.825 130.505 73.705 ;
        RECT 128.065 72.405 128.905 72.575 ;
        RECT 129.355 72.405 130.195 72.575 ;
        RECT 130.675 71.495 130.845 71.935 ;
        RECT 128.065 69.870 128.905 70.040 ;
        RECT 129.355 69.870 130.195 70.040 ;
        RECT 127.755 68.740 127.925 69.620 ;
        RECT 129.045 68.740 129.215 69.620 ;
        RECT 130.335 68.740 130.505 69.620 ;
        RECT 128.065 68.320 128.905 68.490 ;
        RECT 129.355 68.320 130.195 68.490 ;
        RECT 130.675 67.410 130.845 67.850 ;
        RECT 128.065 65.745 128.905 65.915 ;
        RECT 129.355 65.745 130.195 65.915 ;
        RECT 127.755 64.615 127.925 65.495 ;
        RECT 129.045 64.615 129.215 65.495 ;
        RECT 130.335 64.615 130.505 65.495 ;
        RECT 128.065 64.195 128.905 64.365 ;
        RECT 129.355 64.195 130.195 64.365 ;
        RECT 130.675 63.285 130.845 63.725 ;
        RECT 95.180 61.150 95.350 62.290 ;
        RECT 96.150 62.025 103.030 62.195 ;
        RECT 95.685 61.545 95.855 61.885 ;
        RECT 103.325 61.545 103.495 61.885 ;
        RECT 96.150 61.235 103.030 61.405 ;
        RECT 52.860 59.210 54.000 59.380 ;
        RECT 54.830 59.210 59.780 59.380 ;
        RECT 51.680 57.760 51.850 58.900 ;
        RECT 52.655 58.640 60.035 58.810 ;
        RECT 52.190 58.160 52.360 58.500 ;
        RECT 60.330 58.160 60.500 58.500 ;
        RECT 52.655 57.850 60.035 58.020 ;
        RECT 61.815 58.640 62.695 58.810 ;
        RECT 61.350 58.160 61.520 58.500 ;
        RECT 62.990 58.160 63.160 58.500 ;
        RECT 61.815 57.850 62.695 58.020 ;
        RECT 52.570 57.280 53.140 57.450 ;
        RECT 64.960 59.145 69.840 59.315 ;
        RECT 64.540 58.165 64.710 59.005 ;
        RECT 70.090 58.165 70.260 59.005 ;
        RECT 64.960 57.855 69.840 58.025 ;
        RECT 70.600 57.760 70.770 59.400 ;
        RECT 99.700 58.930 104.580 59.100 ;
        RECT 98.770 57.440 98.940 58.580 ;
        RECT 99.235 58.450 99.405 58.790 ;
        RECT 104.875 58.450 105.045 58.790 ;
        RECT 99.700 58.140 104.580 58.310 ;
        RECT 99.235 57.660 99.405 58.000 ;
        RECT 104.875 57.660 105.045 58.000 ;
        RECT 37.330 56.480 38.390 56.660 ;
        RECT 29.100 44.250 29.280 55.920 ;
        RECT 30.110 54.250 34.990 54.420 ;
        RECT 39.110 54.250 43.990 54.420 ;
        RECT 29.645 53.770 29.815 54.110 ;
        RECT 35.285 53.770 35.455 54.110 ;
        RECT 38.645 53.770 38.815 54.110 ;
        RECT 44.285 53.770 44.455 54.110 ;
        RECT 30.110 53.460 34.990 53.630 ;
        RECT 39.110 53.460 43.990 53.630 ;
        RECT 30.110 49.750 34.990 49.920 ;
        RECT 39.110 49.750 43.990 49.920 ;
        RECT 29.645 49.270 29.815 49.610 ;
        RECT 35.285 49.270 35.455 49.610 ;
        RECT 38.645 49.270 38.815 49.610 ;
        RECT 44.285 49.270 44.455 49.610 ;
        RECT 30.110 48.960 34.990 49.130 ;
        RECT 39.110 48.960 43.990 49.130 ;
        RECT 30.110 45.250 34.990 45.420 ;
        RECT 39.110 45.250 43.990 45.420 ;
        RECT 29.645 44.770 29.815 45.110 ;
        RECT 35.285 44.770 35.455 45.110 ;
        RECT 38.645 44.770 38.815 45.110 ;
        RECT 44.285 44.770 44.455 45.110 ;
        RECT 30.110 44.460 34.990 44.630 ;
        RECT 39.110 44.460 43.990 44.630 ;
        RECT 47.830 54.730 52.710 54.900 ;
        RECT 54.830 54.730 59.710 54.900 ;
        RECT 47.410 53.750 47.580 54.590 ;
        RECT 52.960 53.750 53.130 54.590 ;
        RECT 54.410 53.750 54.580 54.590 ;
        RECT 59.960 53.750 60.130 54.590 ;
        RECT 47.830 53.440 52.710 53.610 ;
        RECT 54.830 53.440 59.710 53.610 ;
        RECT 47.830 52.730 52.710 52.900 ;
        RECT 54.830 52.730 59.710 52.900 ;
        RECT 47.410 51.750 47.580 52.590 ;
        RECT 52.960 51.750 53.130 52.590 ;
        RECT 54.410 51.750 54.580 52.590 ;
        RECT 59.960 51.750 60.130 52.590 ;
        RECT 47.830 51.440 52.710 51.610 ;
        RECT 54.830 51.440 59.710 51.610 ;
        RECT 47.830 48.730 52.710 48.900 ;
        RECT 54.830 48.730 59.710 48.900 ;
        RECT 47.410 47.750 47.580 48.590 ;
        RECT 52.960 47.750 53.130 48.590 ;
        RECT 54.410 47.750 54.580 48.590 ;
        RECT 59.960 47.750 60.130 48.590 ;
        RECT 47.830 47.440 52.710 47.610 ;
        RECT 54.830 47.440 59.710 47.610 ;
        RECT 47.830 46.730 52.710 46.900 ;
        RECT 54.830 46.730 59.710 46.900 ;
        RECT 47.410 45.750 47.580 46.590 ;
        RECT 52.960 45.750 53.130 46.590 ;
        RECT 54.410 45.750 54.580 46.590 ;
        RECT 59.960 45.750 60.130 46.590 ;
        RECT 47.830 45.440 52.710 45.610 ;
        RECT 54.830 45.440 59.710 45.610 ;
        RECT 61.260 44.450 61.430 46.660 ;
        RECT 63.290 56.040 68.170 56.210 ;
        RECT 62.870 55.060 63.040 55.900 ;
        RECT 68.420 55.060 68.590 55.900 ;
        RECT 63.290 54.750 68.170 54.920 ;
        RECT 62.870 53.770 63.040 54.610 ;
        RECT 68.420 53.770 68.590 54.610 ;
        RECT 63.290 53.460 68.170 53.630 ;
        RECT 62.870 52.480 63.040 53.320 ;
        RECT 68.420 52.480 68.590 53.320 ;
        RECT 63.290 52.170 68.170 52.340 ;
        RECT 62.870 51.190 63.040 52.030 ;
        RECT 68.420 51.190 68.590 52.030 ;
        RECT 63.290 50.880 68.170 51.050 ;
        RECT 62.870 49.900 63.040 50.740 ;
        RECT 68.420 49.900 68.590 50.740 ;
        RECT 63.290 49.590 68.170 49.760 ;
        RECT 62.870 48.610 63.040 49.450 ;
        RECT 68.420 48.610 68.590 49.450 ;
        RECT 63.290 48.300 68.170 48.470 ;
        RECT 62.870 47.320 63.040 48.160 ;
        RECT 68.420 47.320 68.590 48.160 ;
        RECT 63.290 47.010 68.170 47.180 ;
        RECT 62.870 46.030 63.040 46.870 ;
        RECT 68.420 46.030 68.590 46.870 ;
        RECT 63.290 45.720 68.170 45.890 ;
        RECT 70.520 45.590 70.690 55.300 ;
        RECT 99.700 57.350 104.580 57.520 ;
        RECT 99.235 56.870 99.405 57.210 ;
        RECT 104.875 56.870 105.045 57.210 ;
        RECT 99.700 56.560 104.580 56.730 ;
        RECT 98.770 55.200 98.940 56.340 ;
        RECT 99.235 56.080 99.405 56.420 ;
        RECT 104.875 56.080 105.045 56.420 ;
        RECT 99.700 55.770 104.580 55.940 ;
        RECT 99.235 55.290 99.405 55.630 ;
        RECT 104.875 55.290 105.045 55.630 ;
        RECT 99.700 54.980 104.580 55.150 ;
        RECT 99.235 54.500 99.405 54.840 ;
        RECT 104.875 54.500 105.045 54.840 ;
        RECT 99.700 54.190 104.580 54.360 ;
        RECT 98.770 52.900 98.940 54.040 ;
        RECT 99.235 53.710 99.405 54.050 ;
        RECT 104.875 53.710 105.045 54.050 ;
        RECT 99.700 53.400 104.580 53.570 ;
        RECT 99.235 52.920 99.405 53.260 ;
        RECT 104.875 52.920 105.045 53.260 ;
        RECT 99.700 52.610 104.580 52.780 ;
        RECT 99.235 52.130 99.405 52.470 ;
        RECT 104.875 52.130 105.045 52.470 ;
        RECT 99.700 51.820 104.580 51.990 ;
        RECT 98.770 50.460 98.940 51.600 ;
        RECT 99.235 51.340 99.405 51.680 ;
        RECT 104.875 51.340 105.045 51.680 ;
        RECT 99.700 51.030 104.580 51.200 ;
        RECT 99.235 50.550 99.405 50.890 ;
        RECT 104.875 50.550 105.045 50.890 ;
        RECT 99.700 50.240 104.580 50.410 ;
        RECT 99.235 49.760 99.405 50.100 ;
        RECT 104.875 49.760 105.045 50.100 ;
        RECT 99.700 49.450 104.580 49.620 ;
        RECT 98.770 48.060 98.940 49.200 ;
        RECT 99.235 48.970 99.405 49.310 ;
        RECT 104.875 48.970 105.045 49.310 ;
        RECT 99.700 48.660 104.580 48.830 ;
        RECT 99.235 48.180 99.405 48.520 ;
        RECT 104.875 48.180 105.045 48.520 ;
        RECT 99.700 47.870 104.580 48.040 ;
        RECT 37.660 43.640 38.280 43.820 ;
        RECT 107.760 59.110 112.640 59.280 ;
        RECT 107.340 58.630 107.510 58.970 ;
        RECT 112.890 58.630 113.060 58.970 ;
        RECT 107.760 58.320 112.640 58.490 ;
        RECT 107.340 57.840 107.510 58.180 ;
        RECT 112.890 57.840 113.060 58.180 ;
        RECT 107.760 57.530 112.640 57.700 ;
        RECT 107.340 57.050 107.510 57.390 ;
        RECT 112.890 57.050 113.060 57.390 ;
        RECT 113.490 57.170 113.660 58.640 ;
        RECT 122.895 58.690 123.075 62.360 ;
        RECT 123.875 61.665 124.715 61.835 ;
        RECT 125.165 61.665 126.005 61.835 ;
        RECT 123.565 59.490 123.735 61.370 ;
        RECT 124.855 59.490 125.025 61.370 ;
        RECT 126.145 59.490 126.315 61.370 ;
        RECT 123.875 59.025 124.715 59.195 ;
        RECT 125.165 59.025 126.005 59.195 ;
        RECT 128.065 61.190 128.905 61.360 ;
        RECT 129.355 61.190 130.195 61.360 ;
        RECT 127.755 60.060 127.925 60.940 ;
        RECT 129.045 60.060 129.215 60.940 ;
        RECT 130.335 60.060 130.505 60.940 ;
        RECT 128.065 59.640 128.905 59.810 ;
        RECT 129.355 59.640 130.195 59.810 ;
        RECT 130.675 58.730 130.845 59.170 ;
        RECT 107.760 56.740 112.640 56.910 ;
        RECT 107.340 56.260 107.510 56.600 ;
        RECT 112.890 56.260 113.060 56.600 ;
        RECT 107.760 55.950 112.640 56.120 ;
        RECT 107.340 55.470 107.510 55.810 ;
        RECT 112.890 55.470 113.060 55.810 ;
        RECT 107.760 55.160 112.640 55.330 ;
        RECT 107.340 54.680 107.510 55.020 ;
        RECT 112.890 54.680 113.060 55.020 ;
        RECT 107.760 54.370 112.640 54.540 ;
        RECT 113.490 54.340 113.660 55.810 ;
        RECT 107.340 53.890 107.510 54.230 ;
        RECT 112.890 53.890 113.060 54.230 ;
        RECT 107.760 53.580 112.640 53.750 ;
        RECT 107.340 53.100 107.510 53.440 ;
        RECT 112.890 53.100 113.060 53.440 ;
        RECT 107.760 52.790 112.640 52.960 ;
        RECT 107.340 52.310 107.510 52.650 ;
        RECT 112.890 52.310 113.060 52.650 ;
        RECT 107.760 52.000 112.640 52.170 ;
        RECT 113.490 51.990 113.660 53.460 ;
        RECT 107.340 51.520 107.510 51.860 ;
        RECT 112.890 51.520 113.060 51.860 ;
        RECT 107.760 51.210 112.640 51.380 ;
        RECT 107.340 50.730 107.510 51.070 ;
        RECT 112.890 50.730 113.060 51.070 ;
        RECT 107.760 50.420 112.640 50.590 ;
        RECT 107.340 49.940 107.510 50.280 ;
        RECT 112.890 49.940 113.060 50.280 ;
        RECT 107.760 49.630 112.640 49.800 ;
        RECT 107.340 49.150 107.510 49.490 ;
        RECT 112.890 49.150 113.060 49.490 ;
        RECT 113.490 49.470 113.660 50.940 ;
        RECT 107.760 48.840 112.640 49.010 ;
        RECT 107.340 48.360 107.510 48.700 ;
        RECT 112.890 48.360 113.060 48.700 ;
        RECT 107.760 48.050 112.640 48.220 ;
        RECT 107.340 47.570 107.510 47.910 ;
        RECT 112.890 47.570 113.060 47.910 ;
        RECT 107.760 47.260 112.640 47.430 ;
        RECT 107.340 46.780 107.510 47.120 ;
        RECT 112.890 46.780 113.060 47.120 ;
        RECT 113.490 46.890 113.660 48.360 ;
        RECT 107.760 46.470 112.640 46.640 ;
        RECT 107.340 45.990 107.510 46.330 ;
        RECT 112.890 45.990 113.060 46.330 ;
        RECT 107.760 45.680 112.640 45.850 ;
        RECT 107.340 45.200 107.510 45.540 ;
        RECT 112.890 45.200 113.060 45.540 ;
        RECT 107.760 44.890 112.640 45.060 ;
        RECT 107.340 44.410 107.510 44.750 ;
        RECT 112.890 44.410 113.060 44.750 ;
        RECT 113.490 44.320 113.660 45.790 ;
        RECT 107.760 44.100 112.640 44.270 ;
      LAYER met1 ;
        RECT 26.470 197.400 28.630 199.050 ;
        RECT 26.960 184.010 28.230 197.400 ;
        RECT 71.670 196.690 73.270 199.800 ;
        RECT 130.110 196.690 131.170 199.800 ;
        RECT 72.240 195.300 72.960 196.690 ;
        RECT 106.270 195.580 107.580 196.490 ;
        RECT 30.040 195.180 72.960 195.300 ;
        RECT 30.040 194.900 72.950 195.180 ;
        RECT 30.040 193.050 30.340 194.900 ;
        RECT 31.040 194.680 70.920 194.900 ;
        RECT 30.980 194.450 70.980 194.680 ;
        RECT 30.590 194.340 30.820 194.400 ;
        RECT 30.590 194.280 30.830 194.340 ;
        RECT 30.590 193.440 31.000 194.280 ;
        RECT 30.610 193.390 31.000 193.440 ;
        RECT 71.140 193.390 71.370 194.400 ;
        RECT 30.610 193.160 71.370 193.390 ;
        RECT 30.110 191.950 30.280 193.050 ;
        RECT 30.020 191.120 30.360 191.950 ;
        RECT 30.610 191.350 32.920 193.160 ;
        RECT 44.900 192.260 47.710 192.270 ;
        RECT 30.770 191.330 32.875 191.350 ;
        RECT 30.110 190.700 30.280 191.120 ;
        RECT 44.890 189.840 47.710 192.260 ;
        RECT 62.050 191.280 69.880 193.160 ;
        RECT 72.240 192.470 72.950 194.900 ;
        RECT 70.320 191.970 72.950 192.470 ;
        RECT 106.640 194.370 107.360 195.580 ;
        RECT 107.810 194.550 109.010 194.650 ;
        RECT 106.640 194.270 107.520 194.370 ;
        RECT 107.700 194.320 112.700 194.550 ;
        RECT 107.810 194.290 109.010 194.320 ;
        RECT 112.870 194.270 113.180 194.380 ;
        RECT 106.640 193.810 107.540 194.270 ;
        RECT 106.640 193.480 107.520 193.810 ;
        RECT 111.220 193.760 112.500 193.860 ;
        RECT 112.860 193.810 113.180 194.270 ;
        RECT 107.700 193.530 112.700 193.760 ;
        RECT 111.220 193.500 112.500 193.530 ;
        RECT 112.870 193.480 113.180 193.810 ;
        RECT 106.640 193.020 107.540 193.480 ;
        RECT 107.810 193.030 108.990 193.060 ;
        RECT 106.640 192.690 107.520 193.020 ;
        RECT 107.810 192.970 109.000 193.030 ;
        RECT 112.860 193.020 113.180 193.480 ;
        RECT 107.700 192.740 112.700 192.970 ;
        RECT 107.810 192.690 109.000 192.740 ;
        RECT 112.870 192.690 113.180 193.020 ;
        RECT 70.320 191.760 72.580 191.970 ;
        RECT 44.890 187.380 66.320 189.840 ;
        RECT 28.690 185.040 66.320 187.380 ;
        RECT 70.320 186.920 70.930 191.760 ;
        RECT 70.320 186.140 70.940 186.920 ;
        RECT 28.690 184.700 47.710 185.040 ;
        RECT 14.990 180.030 17.120 182.180 ;
        RECT 18.360 180.030 21.230 182.180 ;
        RECT 22.360 180.030 24.490 182.180 ;
        RECT 26.950 182.170 28.240 184.010 ;
        RECT 25.620 180.030 28.240 182.170 ;
        RECT 18.360 155.020 19.120 180.030 ;
        RECT 27.350 173.970 28.040 174.600 ;
        RECT 27.340 170.640 28.040 173.970 ;
        RECT 14.990 149.600 15.490 155.020 ;
        RECT 16.590 152.870 19.120 155.020 ;
        RECT 20.730 152.880 22.860 155.030 ;
        RECT 23.990 152.880 26.120 155.030 ;
        RECT 16.600 151.470 19.130 151.750 ;
        RECT 27.350 151.470 28.030 170.640 ;
        RECT 28.750 170.130 29.330 184.700 ;
        RECT 37.620 183.260 38.300 183.740 ;
        RECT 34.060 182.800 35.010 182.880 ;
        RECT 29.520 181.990 29.850 182.600 ;
        RECT 30.040 182.570 35.040 182.800 ;
        RECT 34.060 182.440 35.010 182.570 ;
        RECT 35.220 182.060 35.550 182.550 ;
        RECT 34.260 182.010 35.550 182.060 ;
        RECT 30.040 181.990 35.550 182.010 ;
        RECT 29.520 181.780 35.550 181.990 ;
        RECT 29.520 181.730 30.360 181.780 ;
        RECT 34.260 181.770 35.550 181.780 ;
        RECT 29.520 173.170 29.850 181.730 ;
        RECT 34.080 178.300 35.020 178.490 ;
        RECT 30.040 178.070 35.040 178.300 ;
        RECT 34.080 178.020 35.020 178.070 ;
        RECT 34.080 177.510 35.050 177.610 ;
        RECT 30.040 177.280 35.050 177.510 ;
        RECT 34.080 176.890 35.050 177.280 ;
        RECT 34.080 173.800 35.080 173.950 ;
        RECT 30.040 173.570 35.080 173.800 ;
        RECT 34.080 173.490 35.080 173.570 ;
        RECT 29.520 173.080 30.270 173.170 ;
        RECT 35.220 173.110 35.550 181.770 ;
        RECT 29.550 173.010 30.270 173.080 ;
        RECT 34.250 173.030 35.550 173.110 ;
        RECT 34.250 173.010 35.500 173.030 ;
        RECT 29.550 172.800 35.500 173.010 ;
        RECT 30.040 172.780 35.500 172.800 ;
        RECT 34.250 172.760 35.500 172.780 ;
        RECT 35.740 172.670 36.130 183.130 ;
        RECT 36.670 172.590 37.310 183.080 ;
        RECT 37.790 170.930 38.180 183.260 ;
        RECT 39.180 182.800 39.900 183.000 ;
        RECT 70.330 182.980 70.940 186.140 ;
        RECT 38.500 182.520 38.830 182.580 ;
        RECT 39.040 182.570 44.040 182.800 ;
        RECT 38.500 182.060 38.835 182.520 ;
        RECT 39.180 182.430 39.900 182.570 ;
        RECT 38.500 178.020 38.830 182.060 ;
        RECT 39.000 182.010 39.620 182.070 ;
        RECT 39.000 181.780 44.040 182.010 ;
        RECT 39.000 181.570 39.620 181.780 ;
        RECT 44.200 179.370 44.530 182.570 ;
        RECT 61.030 182.120 70.940 182.980 ;
        RECT 47.790 181.820 49.510 181.960 ;
        RECT 55.190 181.820 56.710 181.920 ;
        RECT 47.760 181.590 52.760 181.820 ;
        RECT 54.760 181.590 59.760 181.820 ;
        RECT 45.920 181.540 47.510 181.570 ;
        RECT 47.790 181.540 49.510 181.590 ;
        RECT 53.710 181.540 54.570 181.550 ;
        RECT 45.920 180.580 47.600 181.540 ;
        RECT 52.920 180.580 53.150 181.540 ;
        RECT 53.700 180.580 54.600 181.540 ;
        RECT 55.190 181.400 56.710 181.590 ;
        RECT 59.920 180.580 60.150 181.540 ;
        RECT 45.920 180.560 47.580 180.580 ;
        RECT 53.700 180.560 54.590 180.580 ;
        RECT 45.920 180.220 47.030 180.560 ;
        RECT 53.700 180.540 54.570 180.560 ;
        RECT 47.760 180.510 52.760 180.530 ;
        RECT 44.200 178.480 44.860 179.370 ;
        RECT 39.130 178.300 39.850 178.420 ;
        RECT 39.040 178.070 44.040 178.300 ;
        RECT 38.500 177.560 38.835 178.020 ;
        RECT 39.130 177.850 39.850 178.070 ;
        RECT 38.500 177.400 38.830 177.560 ;
        RECT 39.040 177.480 44.040 177.510 ;
        RECT 44.200 177.480 44.530 178.480 ;
        RECT 39.040 177.400 44.530 177.480 ;
        RECT 38.500 177.280 44.530 177.400 ;
        RECT 38.500 177.050 39.820 177.280 ;
        RECT 43.870 177.230 44.530 177.280 ;
        RECT 38.500 173.520 38.830 177.050 ;
        RECT 39.070 173.800 39.890 173.970 ;
        RECT 39.040 173.570 44.040 173.800 ;
        RECT 38.500 173.060 38.835 173.520 ;
        RECT 39.070 173.470 39.890 173.570 ;
        RECT 39.010 173.010 39.670 173.030 ;
        RECT 42.020 173.010 43.820 173.160 ;
        RECT 44.200 173.050 44.530 177.230 ;
        RECT 46.710 177.770 47.030 180.220 ;
        RECT 47.740 179.620 52.790 180.510 ;
        RECT 47.760 179.590 52.760 179.620 ;
        RECT 53.700 179.560 54.020 180.540 ;
        RECT 54.760 180.500 59.760 180.530 ;
        RECT 54.730 179.800 59.780 180.500 ;
        RECT 61.030 180.470 61.610 182.120 ;
        RECT 63.220 181.540 64.140 181.610 ;
        RECT 63.220 181.310 68.240 181.540 ;
        RECT 54.740 179.610 59.780 179.800 ;
        RECT 54.760 179.590 59.760 179.610 ;
        RECT 52.960 179.540 54.020 179.560 ;
        RECT 47.370 178.580 47.600 179.540 ;
        RECT 52.920 178.580 54.020 179.540 ;
        RECT 52.960 178.560 54.020 178.580 ;
        RECT 47.760 178.300 52.760 178.530 ;
        RECT 50.070 177.970 51.800 178.300 ;
        RECT 46.710 176.140 47.040 177.770 ;
        RECT 46.710 175.560 47.030 176.140 ;
        RECT 53.700 176.110 54.020 178.560 ;
        RECT 54.320 177.630 54.600 179.570 ;
        RECT 57.280 178.530 58.800 178.620 ;
        RECT 59.920 178.580 60.150 179.540 ;
        RECT 54.760 178.300 59.760 178.530 ;
        RECT 57.280 178.100 58.800 178.300 ;
        RECT 54.210 176.600 54.600 177.630 ;
        RECT 62.780 177.130 63.060 181.280 ;
        RECT 63.220 181.190 64.140 181.310 ;
        RECT 68.410 181.260 68.820 181.280 ;
        RECT 67.140 180.250 68.240 180.450 ;
        RECT 68.380 180.300 68.820 181.260 ;
        RECT 70.330 180.450 70.940 182.120 ;
        RECT 63.220 180.020 68.240 180.250 ;
        RECT 67.140 179.780 68.240 180.020 ;
        RECT 68.410 179.970 68.820 180.300 ;
        RECT 63.220 178.960 64.140 179.030 ;
        RECT 68.380 179.010 68.820 179.970 ;
        RECT 70.160 179.790 70.940 180.450 ;
        RECT 63.220 178.730 68.230 178.960 ;
        RECT 63.220 178.610 64.140 178.730 ;
        RECT 68.410 178.680 68.820 179.010 ;
        RECT 67.220 177.680 68.160 177.750 ;
        RECT 68.380 177.720 68.820 178.680 ;
        RECT 63.270 177.670 68.230 177.680 ;
        RECT 63.220 177.450 68.230 177.670 ;
        RECT 63.220 177.440 68.220 177.450 ;
        RECT 67.220 177.360 68.160 177.440 ;
        RECT 68.410 177.390 68.820 177.720 ;
        RECT 68.380 177.130 68.820 177.390 ;
        RECT 62.780 176.680 63.150 177.130 ;
        RECT 68.330 176.680 68.820 177.130 ;
        RECT 47.750 175.820 49.640 175.940 ;
        RECT 47.750 175.590 52.760 175.820 ;
        RECT 46.710 175.540 47.570 175.560 ;
        RECT 46.710 174.580 47.600 175.540 ;
        RECT 47.750 175.320 49.640 175.590 ;
        RECT 53.690 175.580 54.030 176.110 ;
        RECT 55.180 175.820 56.700 175.950 ;
        RECT 54.760 175.590 59.760 175.820 ;
        RECT 52.920 174.580 53.150 175.540 ;
        RECT 46.710 174.550 47.570 174.580 ;
        RECT 53.690 174.530 54.600 175.580 ;
        RECT 55.180 175.430 56.700 175.590 ;
        RECT 59.920 174.580 60.150 175.540 ;
        RECT 47.760 174.510 52.760 174.530 ;
        RECT 47.730 173.620 52.780 174.510 ;
        RECT 47.760 173.590 52.760 173.620 ;
        RECT 53.690 173.580 54.030 174.530 ;
        RECT 54.760 174.510 59.760 174.530 ;
        RECT 54.760 174.300 59.790 174.510 ;
        RECT 54.970 173.820 59.790 174.300 ;
        RECT 54.760 173.620 59.790 173.820 ;
        RECT 52.950 173.540 54.030 173.580 ;
        RECT 39.010 172.780 44.040 173.010 ;
        RECT 39.010 172.560 39.670 172.780 ;
        RECT 42.020 172.340 43.820 172.780 ;
        RECT 47.370 172.580 47.600 173.540 ;
        RECT 47.760 172.300 52.760 172.530 ;
        RECT 50.070 171.960 51.800 172.300 ;
        RECT 52.920 172.140 54.030 173.540 ;
        RECT 54.260 172.560 54.610 173.600 ;
        RECT 54.760 173.590 59.760 173.620 ;
        RECT 57.250 172.530 58.770 172.630 ;
        RECT 59.920 172.580 60.150 173.540 ;
        RECT 54.760 172.300 59.760 172.530 ;
        RECT 57.250 172.110 58.770 172.300 ;
        RECT 62.780 171.270 63.060 176.680 ;
        RECT 63.220 176.380 64.150 176.440 ;
        RECT 68.380 176.430 68.820 176.680 ;
        RECT 63.220 176.150 68.230 176.380 ;
        RECT 63.220 176.060 64.150 176.150 ;
        RECT 68.410 176.100 68.820 176.430 ;
        RECT 67.220 175.100 68.170 175.190 ;
        RECT 68.380 175.140 68.820 176.100 ;
        RECT 63.270 175.090 68.230 175.100 ;
        RECT 63.220 174.870 68.230 175.090 ;
        RECT 63.220 174.860 68.220 174.870 ;
        RECT 67.220 174.810 68.170 174.860 ;
        RECT 68.410 174.810 68.820 175.140 ;
        RECT 63.220 173.810 64.140 173.880 ;
        RECT 68.380 173.850 68.820 174.810 ;
        RECT 63.220 173.580 68.230 173.810 ;
        RECT 63.220 173.570 68.220 173.580 ;
        RECT 63.220 173.510 64.140 173.570 ;
        RECT 68.410 173.520 68.820 173.850 ;
        RECT 67.220 172.510 68.170 172.590 ;
        RECT 68.380 172.560 68.820 173.520 ;
        RECT 63.220 172.280 68.230 172.510 ;
        RECT 67.220 172.190 68.170 172.280 ;
        RECT 68.410 172.230 68.820 172.560 ;
        RECT 63.210 171.220 64.140 171.270 ;
        RECT 68.370 171.260 69.520 172.230 ;
        RECT 63.210 170.990 68.220 171.220 ;
        RECT 63.210 170.950 64.140 170.990 ;
        RECT 37.230 170.130 38.460 170.930 ;
        RECT 28.750 169.470 53.340 170.130 ;
        RECT 70.330 170.040 70.940 179.790 ;
        RECT 71.670 172.360 72.810 190.300 ;
        RECT 98.590 180.040 99.010 192.240 ;
        RECT 106.640 192.230 107.540 192.690 ;
        RECT 107.810 192.640 108.990 192.690 ;
        RECT 106.640 191.900 107.520 192.230 ;
        RECT 111.230 192.180 112.500 192.310 ;
        RECT 112.860 192.230 113.180 192.690 ;
        RECT 107.700 191.950 112.700 192.180 ;
        RECT 111.230 191.920 112.500 191.950 ;
        RECT 112.870 191.900 113.180 192.230 ;
        RECT 106.640 191.440 107.540 191.900 ;
        RECT 106.640 191.110 107.520 191.440 ;
        RECT 107.850 191.390 109.000 191.480 ;
        RECT 112.860 191.440 113.180 191.900 ;
        RECT 107.700 191.160 112.700 191.390 ;
        RECT 107.850 191.130 109.000 191.160 ;
        RECT 112.870 191.110 113.180 191.440 ;
        RECT 103.220 190.780 104.480 190.870 ;
        RECT 96.550 179.430 99.010 180.040 ;
        RECT 99.150 179.700 99.450 190.650 ;
        RECT 99.640 190.550 104.640 190.780 ;
        RECT 103.220 190.520 104.480 190.550 ;
        RECT 99.800 189.990 100.880 190.100 ;
        RECT 99.640 189.760 104.640 189.990 ;
        RECT 99.800 189.670 100.880 189.760 ;
        RECT 103.220 189.200 104.480 189.280 ;
        RECT 99.640 188.970 104.640 189.200 ;
        RECT 103.220 188.940 104.480 188.970 ;
        RECT 99.780 188.410 100.880 188.520 ;
        RECT 99.640 188.180 104.640 188.410 ;
        RECT 99.780 188.100 100.880 188.180 ;
        RECT 103.220 187.620 104.480 187.650 ;
        RECT 99.640 187.390 104.640 187.620 ;
        RECT 103.220 187.310 104.480 187.390 ;
        RECT 99.730 186.830 100.880 186.960 ;
        RECT 99.640 186.600 104.640 186.830 ;
        RECT 99.730 186.500 100.880 186.600 ;
        RECT 103.220 186.040 104.480 186.120 ;
        RECT 99.640 185.810 104.640 186.040 ;
        RECT 103.220 185.780 104.480 185.810 ;
        RECT 99.720 185.250 100.880 185.370 ;
        RECT 99.640 185.020 104.640 185.250 ;
        RECT 99.720 184.950 100.880 185.020 ;
        RECT 103.220 184.460 104.480 184.540 ;
        RECT 99.640 184.230 104.640 184.460 ;
        RECT 103.220 184.180 104.480 184.230 ;
        RECT 99.790 183.670 100.880 183.770 ;
        RECT 99.640 183.440 104.640 183.670 ;
        RECT 99.790 183.410 100.880 183.440 ;
        RECT 103.220 182.880 104.480 182.940 ;
        RECT 99.640 182.650 104.640 182.880 ;
        RECT 103.220 182.580 104.480 182.650 ;
        RECT 99.760 182.090 100.880 182.170 ;
        RECT 99.640 181.860 104.640 182.090 ;
        RECT 99.760 181.830 100.880 181.860 ;
        RECT 103.230 181.300 104.490 181.350 ;
        RECT 99.640 181.070 104.640 181.300 ;
        RECT 103.230 180.990 104.490 181.070 ;
        RECT 104.800 180.660 105.100 190.670 ;
        RECT 106.640 190.650 107.540 191.110 ;
        RECT 106.640 190.320 107.520 190.650 ;
        RECT 111.230 190.600 112.510 190.690 ;
        RECT 112.860 190.650 113.180 191.110 ;
        RECT 107.700 190.370 112.700 190.600 ;
        RECT 111.230 190.330 112.510 190.370 ;
        RECT 112.870 190.320 113.180 190.650 ;
        RECT 106.640 189.860 107.540 190.320 ;
        RECT 106.640 189.530 107.520 189.860 ;
        RECT 107.810 189.810 109.000 189.900 ;
        RECT 112.860 189.860 113.180 190.320 ;
        RECT 107.700 189.580 112.700 189.810 ;
        RECT 107.810 189.540 109.000 189.580 ;
        RECT 112.870 189.530 113.180 189.860 ;
        RECT 106.640 189.070 107.540 189.530 ;
        RECT 106.640 188.740 107.520 189.070 ;
        RECT 111.230 189.020 112.500 189.090 ;
        RECT 112.860 189.070 113.180 189.530 ;
        RECT 107.700 188.790 112.700 189.020 ;
        RECT 106.640 188.280 107.540 188.740 ;
        RECT 111.230 188.730 112.500 188.790 ;
        RECT 112.870 188.740 113.180 189.070 ;
        RECT 106.640 187.950 107.520 188.280 ;
        RECT 107.850 188.230 109.000 188.320 ;
        RECT 112.860 188.280 113.180 188.740 ;
        RECT 107.700 188.000 112.700 188.230 ;
        RECT 107.850 187.970 109.000 188.000 ;
        RECT 112.870 187.950 113.180 188.280 ;
        RECT 106.640 187.490 107.540 187.950 ;
        RECT 106.640 187.160 107.520 187.490 ;
        RECT 111.230 187.440 112.490 187.520 ;
        RECT 112.860 187.490 113.180 187.950 ;
        RECT 107.700 187.210 112.700 187.440 ;
        RECT 111.230 187.170 112.490 187.210 ;
        RECT 112.870 187.160 113.180 187.490 ;
        RECT 106.640 186.700 107.540 187.160 ;
        RECT 106.640 186.370 107.520 186.700 ;
        RECT 107.880 186.650 109.000 186.720 ;
        RECT 112.860 186.700 113.180 187.160 ;
        RECT 107.700 186.420 112.700 186.650 ;
        RECT 107.880 186.380 109.000 186.420 ;
        RECT 112.870 186.370 113.180 186.700 ;
        RECT 106.640 185.910 107.540 186.370 ;
        RECT 106.640 185.580 107.520 185.910 ;
        RECT 111.240 185.860 112.500 185.970 ;
        RECT 112.860 185.910 113.180 186.370 ;
        RECT 107.700 185.630 112.700 185.860 ;
        RECT 106.640 185.120 107.540 185.580 ;
        RECT 111.240 185.520 112.500 185.630 ;
        RECT 112.870 185.580 113.180 185.910 ;
        RECT 106.640 184.790 107.520 185.120 ;
        RECT 107.860 185.070 109.010 185.180 ;
        RECT 112.860 185.120 113.180 185.580 ;
        RECT 107.700 184.840 112.700 185.070 ;
        RECT 107.860 184.820 109.010 184.840 ;
        RECT 112.870 184.790 113.180 185.120 ;
        RECT 106.640 184.330 107.540 184.790 ;
        RECT 106.640 184.000 107.520 184.330 ;
        RECT 111.220 184.280 112.550 184.390 ;
        RECT 112.860 184.330 113.180 184.790 ;
        RECT 107.700 184.050 112.700 184.280 ;
        RECT 106.640 183.540 107.540 184.000 ;
        RECT 111.220 183.990 112.550 184.050 ;
        RECT 112.870 184.000 113.180 184.330 ;
        RECT 106.640 183.210 107.520 183.540 ;
        RECT 107.760 183.490 109.000 183.560 ;
        RECT 112.860 183.540 113.180 184.000 ;
        RECT 107.700 183.260 112.700 183.490 ;
        RECT 107.760 183.210 109.000 183.260 ;
        RECT 112.870 183.210 113.180 183.540 ;
        RECT 106.640 182.750 107.540 183.210 ;
        RECT 106.640 182.420 107.520 182.750 ;
        RECT 111.230 182.700 112.510 182.800 ;
        RECT 112.860 182.750 113.180 183.210 ;
        RECT 107.700 182.470 112.700 182.700 ;
        RECT 106.640 181.960 107.540 182.420 ;
        RECT 111.230 182.400 112.510 182.470 ;
        RECT 112.870 182.420 113.180 182.750 ;
        RECT 106.640 181.630 107.520 181.960 ;
        RECT 107.780 181.910 109.000 182.000 ;
        RECT 112.860 181.960 113.180 182.420 ;
        RECT 107.700 181.680 112.700 181.910 ;
        RECT 107.780 181.640 109.000 181.680 ;
        RECT 112.870 181.630 113.180 181.960 ;
        RECT 106.640 181.170 107.540 181.630 ;
        RECT 106.640 180.840 107.520 181.170 ;
        RECT 111.230 181.120 112.510 181.200 ;
        RECT 112.860 181.170 113.180 181.630 ;
        RECT 107.700 180.890 112.700 181.120 ;
        RECT 104.800 180.650 105.760 180.660 ;
        RECT 99.770 180.510 100.890 180.610 ;
        RECT 99.640 180.280 104.640 180.510 ;
        RECT 99.770 180.260 100.890 180.280 ;
        RECT 103.220 179.720 104.480 179.780 ;
        RECT 99.640 179.490 104.640 179.720 ;
        RECT 103.220 179.430 104.480 179.490 ;
        RECT 94.510 178.600 99.010 179.430 ;
        RECT 104.800 179.150 105.980 180.650 ;
        RECT 106.640 179.580 107.540 180.840 ;
        RECT 111.230 180.800 112.510 180.890 ;
        RECT 112.870 180.840 113.180 181.170 ;
        RECT 107.780 180.380 108.990 180.410 ;
        RECT 112.860 180.380 113.180 180.840 ;
        RECT 107.780 180.330 109.000 180.380 ;
        RECT 107.700 180.100 112.700 180.330 ;
        RECT 107.780 180.020 109.000 180.100 ;
        RECT 112.870 180.050 113.180 180.380 ;
        RECT 107.780 180.010 108.990 180.020 ;
        RECT 112.860 179.590 113.180 180.050 ;
        RECT 94.510 173.760 95.410 178.600 ;
        RECT 96.550 178.590 98.980 178.600 ;
        RECT 96.150 177.460 97.060 177.660 ;
        RECT 96.130 177.415 103.100 177.460 ;
        RECT 96.090 177.185 103.100 177.415 ;
        RECT 95.610 174.720 95.900 177.150 ;
        RECT 96.130 177.120 103.100 177.185 ;
        RECT 96.150 177.100 97.060 177.120 ;
        RECT 96.090 176.610 103.090 176.625 ;
        RECT 96.080 175.250 103.120 176.610 ;
        RECT 103.290 175.760 103.580 177.150 ;
        RECT 106.670 175.970 107.540 179.580 ;
        RECT 107.840 179.540 112.680 179.590 ;
        RECT 112.870 179.540 113.180 179.590 ;
        RECT 107.700 179.310 112.700 179.540 ;
        RECT 107.840 179.250 112.680 179.310 ;
        RECT 113.350 178.600 113.960 195.090 ;
        RECT 130.420 189.005 130.950 196.690 ;
        RECT 122.725 189.000 123.625 189.005 ;
        RECT 122.720 187.875 123.625 189.000 ;
        RECT 122.725 187.595 123.625 187.875 ;
        RECT 123.815 187.800 124.775 188.030 ;
        RECT 125.105 188.005 126.065 188.030 ;
        RECT 126.825 188.005 127.515 188.785 ;
        RECT 125.105 187.835 128.905 188.005 ;
        RECT 125.105 187.800 126.065 187.835 ;
        RECT 122.725 185.595 123.765 187.595 ;
        RECT 122.725 185.210 123.625 185.595 ;
        RECT 123.985 185.390 124.505 187.800 ;
        RECT 124.825 185.595 125.055 187.595 ;
        RECT 125.315 185.390 125.835 187.800 ;
        RECT 126.135 187.595 127.855 187.615 ;
        RECT 126.115 187.165 127.855 187.595 ;
        RECT 128.065 187.555 128.905 187.835 ;
        RECT 128.005 187.325 128.965 187.555 ;
        RECT 129.295 187.325 130.255 187.555 ;
        RECT 126.115 186.165 127.955 187.165 ;
        RECT 126.115 185.595 127.855 186.165 ;
        RECT 128.245 186.005 128.765 187.325 ;
        RECT 129.015 186.165 129.245 187.165 ;
        RECT 129.515 186.005 130.035 187.325 ;
        RECT 130.415 187.165 130.955 189.005 ;
        RECT 130.305 186.165 130.955 187.165 ;
        RECT 128.005 185.775 128.965 186.005 ;
        RECT 129.295 185.775 130.255 186.005 ;
        RECT 130.415 185.635 130.955 186.165 ;
        RECT 126.135 185.575 127.855 185.595 ;
        RECT 122.725 184.555 123.650 185.210 ;
        RECT 123.815 185.160 124.775 185.390 ;
        RECT 125.105 185.160 126.065 185.390 ;
        RECT 126.825 185.165 127.515 185.575 ;
        RECT 130.405 185.515 130.955 185.635 ;
        RECT 122.720 184.210 123.650 184.555 ;
        RECT 126.815 184.825 127.515 185.165 ;
        RECT 126.815 184.545 127.520 184.825 ;
        RECT 122.720 179.755 123.630 184.210 ;
        RECT 126.820 180.325 127.520 184.545 ;
        RECT 130.395 184.595 130.955 185.515 ;
        RECT 130.395 184.375 130.960 184.595 ;
        RECT 130.410 180.435 130.960 184.375 ;
        RECT 122.725 179.560 123.625 179.755 ;
        RECT 123.815 179.700 124.775 179.930 ;
        RECT 125.105 179.905 126.065 179.930 ;
        RECT 126.825 179.905 127.515 180.325 ;
        RECT 125.105 179.735 128.905 179.905 ;
        RECT 125.105 179.700 126.065 179.735 ;
        RECT 103.290 174.840 103.590 175.760 ;
        RECT 96.130 174.695 103.100 174.790 ;
        RECT 96.090 174.465 103.100 174.695 ;
        RECT 103.290 174.540 104.010 174.840 ;
        RECT 96.130 174.450 103.100 174.465 ;
        RECT 96.150 174.130 97.060 174.450 ;
        RECT 97.420 173.760 103.040 174.160 ;
        RECT 94.510 173.410 103.040 173.760 ;
        RECT 103.840 173.890 104.010 174.540 ;
        RECT 103.840 173.880 106.240 173.890 ;
        RECT 107.410 173.880 108.110 173.940 ;
        RECT 103.840 173.750 112.930 173.880 ;
        RECT 103.840 173.640 107.630 173.750 ;
        RECT 94.510 173.200 95.410 173.410 ;
        RECT 94.510 172.360 95.000 173.200 ;
        RECT 95.595 172.920 103.535 173.110 ;
        RECT 95.190 172.880 103.535 172.920 ;
        RECT 103.840 172.880 106.240 173.640 ;
        RECT 107.895 173.610 112.930 173.750 ;
        RECT 107.900 173.400 112.930 173.610 ;
        RECT 107.900 173.385 112.900 173.400 ;
        RECT 95.190 172.830 96.170 172.880 ;
        RECT 95.160 172.580 96.170 172.830 ;
        RECT 95.160 172.370 95.390 172.580 ;
        RECT 103.300 172.370 103.535 172.880 ;
        RECT 104.165 172.370 104.555 172.880 ;
        RECT 71.670 172.030 95.000 172.360 ;
        RECT 95.595 172.290 103.095 172.320 ;
        RECT 95.570 172.090 103.095 172.290 ;
        RECT 103.305 172.200 103.535 172.370 ;
        RECT 105.950 172.350 106.240 172.880 ;
        RECT 107.510 172.970 107.740 173.335 ;
        RECT 113.060 172.970 113.290 173.335 ;
        RECT 107.510 172.630 113.290 172.970 ;
        RECT 107.510 172.375 107.740 172.630 ;
        RECT 113.060 172.375 113.290 172.630 ;
        RECT 103.710 172.200 104.090 172.230 ;
        RECT 103.305 172.180 104.090 172.200 ;
        RECT 104.755 172.180 105.755 172.320 ;
        RECT 107.900 172.300 112.900 172.325 ;
        RECT 113.470 172.300 113.960 178.600 ;
        RECT 121.570 179.495 123.625 179.560 ;
        RECT 121.570 177.580 123.765 179.495 ;
        RECT 122.725 177.495 123.765 177.580 ;
        RECT 122.725 177.090 123.625 177.495 ;
        RECT 123.985 177.290 124.505 179.700 ;
        RECT 124.825 177.495 125.055 179.495 ;
        RECT 125.315 177.290 125.835 179.700 ;
        RECT 126.135 179.495 127.855 179.515 ;
        RECT 126.115 179.065 127.855 179.495 ;
        RECT 128.065 179.455 128.905 179.735 ;
        RECT 128.005 179.225 128.965 179.455 ;
        RECT 129.295 179.225 130.255 179.455 ;
        RECT 126.115 178.065 127.955 179.065 ;
        RECT 126.115 177.495 127.855 178.065 ;
        RECT 128.245 177.905 128.765 179.225 ;
        RECT 129.015 178.065 129.245 179.065 ;
        RECT 129.515 177.905 130.035 179.225 ;
        RECT 130.415 179.065 130.955 180.435 ;
        RECT 130.305 178.065 130.955 179.065 ;
        RECT 128.005 177.675 128.965 177.905 ;
        RECT 129.295 177.675 130.255 177.905 ;
        RECT 130.415 177.535 130.955 178.065 ;
        RECT 126.135 177.475 127.855 177.495 ;
        RECT 122.725 176.355 123.640 177.090 ;
        RECT 123.815 177.060 124.775 177.290 ;
        RECT 125.105 177.060 126.065 177.290 ;
        RECT 126.825 177.065 127.515 177.475 ;
        RECT 130.405 177.415 130.955 177.535 ;
        RECT 126.815 176.615 127.515 177.065 ;
        RECT 126.815 176.445 127.520 176.615 ;
        RECT 103.305 172.090 105.755 172.180 ;
        RECT 107.880 172.150 112.900 172.300 ;
        RECT 113.450 172.150 113.960 172.300 ;
        RECT 122.720 176.090 123.640 176.355 ;
        RECT 122.720 172.195 123.630 176.090 ;
        RECT 126.820 172.345 127.520 176.445 ;
        RECT 130.395 176.275 130.955 177.415 ;
        RECT 130.410 172.805 130.950 176.275 ;
        RECT 95.570 172.030 96.350 172.090 ;
        RECT 71.670 171.690 96.350 172.030 ;
        RECT 103.305 171.970 105.730 172.090 ;
        RECT 28.750 169.140 51.990 169.470 ;
        RECT 52.560 169.410 53.340 169.470 ;
        RECT 60.295 169.410 62.720 169.530 ;
        RECT 52.560 169.210 60.085 169.410 ;
        RECT 52.585 169.180 60.085 169.210 ;
        RECT 60.295 169.320 62.745 169.410 ;
        RECT 60.295 169.300 61.080 169.320 ;
        RECT 51.500 168.300 51.990 169.140 ;
        RECT 60.295 169.130 60.525 169.300 ;
        RECT 60.700 169.270 61.080 169.300 ;
        RECT 61.745 169.180 62.745 169.320 ;
        RECT 64.870 169.350 70.940 170.040 ;
        RECT 64.870 169.200 69.890 169.350 ;
        RECT 70.440 169.200 70.940 169.350 ;
        RECT 64.890 169.175 69.890 169.200 ;
        RECT 52.150 168.920 52.380 169.130 ;
        RECT 52.150 168.670 53.160 168.920 ;
        RECT 52.180 168.620 53.160 168.670 ;
        RECT 60.290 168.620 60.525 169.130 ;
        RECT 61.155 168.620 61.545 169.130 ;
        RECT 62.940 168.620 63.230 169.150 ;
        RECT 52.180 168.580 60.525 168.620 ;
        RECT 52.585 168.390 60.525 168.580 ;
        RECT 51.500 168.090 52.400 168.300 ;
        RECT 51.500 167.740 60.030 168.090 ;
        RECT 51.500 162.900 52.400 167.740 ;
        RECT 53.140 167.050 54.050 167.370 ;
        RECT 54.410 167.340 60.030 167.740 ;
        RECT 60.830 167.860 63.230 168.620 ;
        RECT 64.500 168.870 64.730 169.125 ;
        RECT 70.050 168.870 70.280 169.125 ;
        RECT 64.500 168.530 70.280 168.870 ;
        RECT 64.500 168.165 64.730 168.530 ;
        RECT 70.050 168.165 70.280 168.530 ;
        RECT 64.890 168.100 69.890 168.115 ;
        RECT 64.890 167.890 69.920 168.100 ;
        RECT 60.830 167.750 64.620 167.860 ;
        RECT 64.885 167.750 69.920 167.890 ;
        RECT 60.830 167.620 69.920 167.750 ;
        RECT 60.830 167.610 63.230 167.620 ;
        RECT 53.120 167.035 60.090 167.050 ;
        RECT 53.080 166.805 60.090 167.035 ;
        RECT 60.830 166.960 61.000 167.610 ;
        RECT 64.400 167.560 65.100 167.620 ;
        RECT 52.600 164.350 52.890 166.780 ;
        RECT 53.120 166.710 60.090 166.805 ;
        RECT 60.280 166.660 61.000 166.960 ;
        RECT 53.070 164.890 60.110 166.250 ;
        RECT 60.280 165.740 60.580 166.660 ;
        RECT 53.080 164.875 60.080 164.890 ;
        RECT 53.140 164.380 54.050 164.400 ;
        RECT 53.120 164.315 60.090 164.380 ;
        RECT 60.280 164.350 60.570 165.740 ;
        RECT 53.080 164.085 60.090 164.315 ;
        RECT 53.120 164.040 60.090 164.085 ;
        RECT 53.140 163.840 54.050 164.040 ;
        RECT 51.500 162.070 56.000 162.900 ;
        RECT 16.600 150.790 28.030 151.470 ;
        RECT 16.600 149.600 19.700 150.790 ;
        RECT 19.090 131.340 19.700 149.600 ;
        RECT 55.580 149.260 56.000 162.070 ;
        RECT 60.210 162.010 61.470 162.070 ;
        RECT 56.140 150.850 56.440 161.800 ;
        RECT 56.630 161.780 61.630 162.010 ;
        RECT 60.210 161.720 61.470 161.780 ;
        RECT 56.760 161.220 57.880 161.240 ;
        RECT 56.630 160.990 61.630 161.220 ;
        RECT 56.760 160.890 57.880 160.990 ;
        RECT 61.790 160.850 62.970 162.350 ;
        RECT 63.660 161.070 64.530 165.530 ;
        RECT 70.460 162.900 70.940 169.200 ;
        RECT 64.830 162.190 69.670 162.250 ;
        RECT 64.690 161.960 69.690 162.190 ;
        RECT 64.830 161.910 69.670 161.960 ;
        RECT 69.860 161.910 70.170 161.960 ;
        RECT 64.770 161.480 65.980 161.490 ;
        RECT 64.770 161.400 65.990 161.480 ;
        RECT 69.850 161.450 70.170 161.910 ;
        RECT 64.690 161.170 69.690 161.400 ;
        RECT 64.770 161.120 65.990 161.170 ;
        RECT 69.860 161.120 70.170 161.450 ;
        RECT 64.770 161.090 65.980 161.120 ;
        RECT 63.680 161.020 64.530 161.070 ;
        RECT 61.790 160.840 62.750 160.850 ;
        RECT 60.220 160.430 61.480 160.510 ;
        RECT 56.630 160.200 61.630 160.430 ;
        RECT 60.220 160.150 61.480 160.200 ;
        RECT 56.750 159.640 57.870 159.670 ;
        RECT 56.630 159.410 61.630 159.640 ;
        RECT 56.750 159.330 57.870 159.410 ;
        RECT 60.210 158.850 61.470 158.920 ;
        RECT 56.630 158.620 61.630 158.850 ;
        RECT 60.210 158.560 61.470 158.620 ;
        RECT 56.780 158.060 57.870 158.090 ;
        RECT 56.630 157.830 61.630 158.060 ;
        RECT 56.780 157.730 57.870 157.830 ;
        RECT 60.210 157.270 61.470 157.320 ;
        RECT 56.630 157.040 61.630 157.270 ;
        RECT 60.210 156.960 61.470 157.040 ;
        RECT 56.710 156.480 57.870 156.550 ;
        RECT 56.630 156.250 61.630 156.480 ;
        RECT 56.710 156.130 57.870 156.250 ;
        RECT 60.210 155.690 61.470 155.720 ;
        RECT 56.630 155.460 61.630 155.690 ;
        RECT 60.210 155.380 61.470 155.460 ;
        RECT 56.720 154.900 57.870 155.000 ;
        RECT 56.630 154.670 61.630 154.900 ;
        RECT 56.720 154.540 57.870 154.670 ;
        RECT 60.210 154.110 61.470 154.190 ;
        RECT 56.630 153.880 61.630 154.110 ;
        RECT 60.210 153.850 61.470 153.880 ;
        RECT 56.770 153.320 57.870 153.400 ;
        RECT 56.630 153.090 61.630 153.320 ;
        RECT 56.770 152.980 57.870 153.090 ;
        RECT 60.210 152.530 61.470 152.560 ;
        RECT 56.630 152.300 61.630 152.530 ;
        RECT 60.210 152.220 61.470 152.300 ;
        RECT 56.790 151.740 57.870 151.830 ;
        RECT 56.630 151.510 61.630 151.740 ;
        RECT 56.790 151.400 57.870 151.510 ;
        RECT 60.210 150.950 61.470 150.980 ;
        RECT 56.630 150.720 61.630 150.950 ;
        RECT 61.790 150.830 62.090 160.840 ;
        RECT 64.200 160.660 64.530 161.020 ;
        RECT 64.200 160.330 64.510 160.660 ;
        RECT 68.220 160.610 69.500 160.700 ;
        RECT 69.850 160.660 70.170 161.120 ;
        RECT 64.690 160.380 69.690 160.610 ;
        RECT 64.200 159.870 64.530 160.330 ;
        RECT 68.220 160.300 69.500 160.380 ;
        RECT 69.860 160.330 70.170 160.660 ;
        RECT 69.850 159.870 70.170 160.330 ;
        RECT 64.200 159.540 64.510 159.870 ;
        RECT 64.770 159.820 65.990 159.860 ;
        RECT 64.690 159.590 69.690 159.820 ;
        RECT 64.200 159.080 64.530 159.540 ;
        RECT 64.770 159.500 65.990 159.590 ;
        RECT 69.860 159.540 70.170 159.870 ;
        RECT 64.200 158.750 64.510 159.080 ;
        RECT 68.220 159.030 69.500 159.100 ;
        RECT 69.850 159.080 70.170 159.540 ;
        RECT 64.690 158.800 69.690 159.030 ;
        RECT 64.200 158.290 64.530 158.750 ;
        RECT 68.220 158.700 69.500 158.800 ;
        RECT 69.860 158.750 70.170 159.080 ;
        RECT 69.850 158.290 70.170 158.750 ;
        RECT 64.200 157.960 64.510 158.290 ;
        RECT 64.750 158.240 65.990 158.290 ;
        RECT 64.690 158.010 69.690 158.240 ;
        RECT 64.200 157.500 64.530 157.960 ;
        RECT 64.750 157.940 65.990 158.010 ;
        RECT 69.860 157.960 70.170 158.290 ;
        RECT 64.200 157.170 64.510 157.500 ;
        RECT 68.210 157.450 69.540 157.510 ;
        RECT 69.850 157.500 70.170 157.960 ;
        RECT 64.690 157.220 69.690 157.450 ;
        RECT 64.200 156.710 64.530 157.170 ;
        RECT 68.210 157.110 69.540 157.220 ;
        RECT 69.860 157.170 70.170 157.500 ;
        RECT 69.850 156.710 70.170 157.170 ;
        RECT 64.200 156.380 64.510 156.710 ;
        RECT 64.850 156.660 66.000 156.680 ;
        RECT 64.690 156.430 69.690 156.660 ;
        RECT 64.200 155.920 64.530 156.380 ;
        RECT 64.850 156.320 66.000 156.430 ;
        RECT 69.860 156.380 70.170 156.710 ;
        RECT 64.200 155.590 64.510 155.920 ;
        RECT 68.230 155.870 69.490 155.980 ;
        RECT 69.850 155.920 70.170 156.380 ;
        RECT 64.690 155.640 69.690 155.870 ;
        RECT 64.200 155.130 64.530 155.590 ;
        RECT 68.230 155.530 69.490 155.640 ;
        RECT 69.860 155.590 70.170 155.920 ;
        RECT 69.850 155.130 70.170 155.590 ;
        RECT 64.200 154.800 64.510 155.130 ;
        RECT 64.870 155.080 65.990 155.120 ;
        RECT 64.690 154.850 69.690 155.080 ;
        RECT 64.200 154.340 64.530 154.800 ;
        RECT 64.870 154.780 65.990 154.850 ;
        RECT 69.860 154.800 70.170 155.130 ;
        RECT 69.850 154.340 70.170 154.800 ;
        RECT 64.200 154.010 64.510 154.340 ;
        RECT 68.220 154.290 69.480 154.330 ;
        RECT 64.690 154.060 69.690 154.290 ;
        RECT 64.200 153.550 64.530 154.010 ;
        RECT 68.220 153.980 69.480 154.060 ;
        RECT 69.860 154.010 70.170 154.340 ;
        RECT 69.850 153.550 70.170 154.010 ;
        RECT 64.200 153.220 64.510 153.550 ;
        RECT 64.840 153.500 65.990 153.530 ;
        RECT 64.690 153.270 69.690 153.500 ;
        RECT 64.200 152.760 64.530 153.220 ;
        RECT 64.840 153.180 65.990 153.270 ;
        RECT 69.860 153.220 70.170 153.550 ;
        RECT 64.200 152.430 64.510 152.760 ;
        RECT 68.220 152.710 69.490 152.770 ;
        RECT 69.850 152.760 70.170 153.220 ;
        RECT 64.690 152.480 69.690 152.710 ;
        RECT 64.200 151.970 64.530 152.430 ;
        RECT 68.220 152.410 69.490 152.480 ;
        RECT 69.860 152.430 70.170 152.760 ;
        RECT 69.850 151.970 70.170 152.430 ;
        RECT 64.200 151.640 64.510 151.970 ;
        RECT 64.800 151.920 65.990 151.960 ;
        RECT 64.690 151.690 69.690 151.920 ;
        RECT 64.200 151.180 64.530 151.640 ;
        RECT 64.800 151.600 65.990 151.690 ;
        RECT 69.860 151.640 70.170 151.970 ;
        RECT 69.850 151.180 70.170 151.640 ;
        RECT 64.200 150.850 64.510 151.180 ;
        RECT 68.220 151.130 69.500 151.170 ;
        RECT 64.690 150.900 69.690 151.130 ;
        RECT 60.210 150.630 61.470 150.720 ;
        RECT 64.200 150.390 64.530 150.850 ;
        RECT 68.220 150.810 69.500 150.900 ;
        RECT 69.860 150.850 70.170 151.180 ;
        RECT 69.850 150.390 70.170 150.850 ;
        RECT 64.200 150.060 64.510 150.390 ;
        RECT 64.840 150.340 65.990 150.370 ;
        RECT 64.690 150.110 69.690 150.340 ;
        RECT 64.200 149.600 64.530 150.060 ;
        RECT 64.840 150.020 65.990 150.110 ;
        RECT 69.860 150.060 70.170 150.390 ;
        RECT 69.850 149.600 70.170 150.060 ;
        RECT 60.200 147.820 61.460 149.320 ;
        RECT 64.200 149.270 64.510 149.600 ;
        RECT 68.220 149.550 69.490 149.580 ;
        RECT 64.690 149.320 69.690 149.550 ;
        RECT 64.200 148.810 64.530 149.270 ;
        RECT 68.220 149.190 69.490 149.320 ;
        RECT 69.860 149.270 70.170 149.600 ;
        RECT 64.800 148.810 65.980 148.860 ;
        RECT 69.850 148.810 70.170 149.270 ;
        RECT 64.200 148.480 64.510 148.810 ;
        RECT 64.800 148.760 65.990 148.810 ;
        RECT 64.690 148.530 69.690 148.760 ;
        RECT 64.200 148.020 64.530 148.480 ;
        RECT 64.800 148.470 65.990 148.530 ;
        RECT 69.860 148.480 70.170 148.810 ;
        RECT 64.800 148.440 65.980 148.470 ;
        RECT 69.850 148.020 70.170 148.480 ;
        RECT 60.200 147.480 60.820 147.820 ;
        RECT 60.190 146.490 60.820 147.480 ;
        RECT 64.200 147.760 64.510 148.020 ;
        RECT 68.210 147.970 69.490 148.000 ;
        RECT 64.200 147.130 64.540 147.760 ;
        RECT 64.690 147.740 69.690 147.970 ;
        RECT 68.210 147.640 69.490 147.740 ;
        RECT 69.860 147.690 70.170 148.020 ;
        RECT 69.850 147.230 70.170 147.690 ;
        RECT 70.340 147.340 70.940 162.900 ;
        RECT 64.800 147.180 66.000 147.210 ;
        RECT 64.210 146.820 64.540 147.130 ;
        RECT 64.690 146.950 69.690 147.180 ;
        RECT 69.860 147.120 70.170 147.230 ;
        RECT 64.800 146.850 66.000 146.950 ;
        RECT 60.190 145.060 60.810 146.490 ;
        RECT 63.700 145.960 64.540 146.820 ;
        RECT 20.760 144.440 60.810 145.060 ;
        RECT 20.760 141.780 21.380 144.440 ;
        RECT 19.260 130.280 19.810 130.820 ;
        RECT 14.990 122.450 17.120 124.600 ;
        RECT 19.450 121.600 19.700 130.280 ;
        RECT 70.330 130.270 70.940 147.340 ;
        RECT 59.800 129.900 70.940 130.270 ;
        RECT 18.560 120.230 19.840 121.600 ;
        RECT 70.330 115.870 70.940 129.900 ;
        RECT 71.770 171.370 96.350 171.690 ;
        RECT 107.880 171.460 113.960 172.150 ;
        RECT 71.770 142.850 72.340 171.370 ;
        RECT 80.240 170.570 81.470 171.370 ;
        RECT 77.260 168.720 78.510 168.740 ;
        RECT 73.050 168.700 78.510 168.720 ;
        RECT 72.560 168.490 78.510 168.700 ;
        RECT 72.560 168.420 73.280 168.490 ;
        RECT 72.530 168.330 73.280 168.420 ;
        RECT 77.260 168.470 78.510 168.490 ;
        RECT 77.260 168.390 78.560 168.470 ;
        RECT 72.530 159.770 72.860 168.330 ;
        RECT 77.090 167.930 78.090 168.010 ;
        RECT 73.050 167.700 78.090 167.930 ;
        RECT 77.090 167.550 78.090 167.700 ;
        RECT 77.090 164.220 78.060 164.610 ;
        RECT 73.050 163.990 78.060 164.220 ;
        RECT 77.090 163.890 78.060 163.990 ;
        RECT 77.090 163.430 78.030 163.480 ;
        RECT 73.050 163.200 78.050 163.430 ;
        RECT 77.090 163.010 78.030 163.200 ;
        RECT 72.530 159.720 73.370 159.770 ;
        RECT 78.230 159.730 78.560 168.390 ;
        RECT 77.270 159.720 78.560 159.730 ;
        RECT 72.530 159.510 78.560 159.720 ;
        RECT 72.530 158.900 72.860 159.510 ;
        RECT 73.050 159.490 78.560 159.510 ;
        RECT 77.270 159.440 78.560 159.490 ;
        RECT 77.070 158.930 78.020 159.060 ;
        RECT 78.230 158.950 78.560 159.440 ;
        RECT 73.050 158.700 78.050 158.930 ;
        RECT 77.070 158.620 78.020 158.700 ;
        RECT 78.750 158.370 79.140 168.830 ;
        RECT 79.680 158.420 80.320 168.910 ;
        RECT 80.800 158.240 81.190 170.570 ;
        RECT 106.220 170.510 107.150 170.550 ;
        RECT 106.220 170.280 111.230 170.510 ;
        RECT 106.220 170.230 107.150 170.280 ;
        RECT 93.080 169.200 94.810 169.540 ;
        RECT 82.020 168.720 82.680 168.940 ;
        RECT 85.030 168.720 86.830 169.160 ;
        RECT 90.770 168.970 95.770 169.200 ;
        RECT 82.020 168.490 87.050 168.720 ;
        RECT 82.020 168.470 82.680 168.490 ;
        RECT 81.510 167.980 81.845 168.440 ;
        RECT 85.030 168.340 86.830 168.490 ;
        RECT 81.510 164.450 81.840 167.980 ;
        RECT 82.080 167.930 82.900 168.030 ;
        RECT 82.050 167.700 87.050 167.930 ;
        RECT 82.080 167.530 82.900 167.700 ;
        RECT 81.510 164.220 82.830 164.450 ;
        RECT 87.210 164.270 87.540 168.450 ;
        RECT 90.380 167.960 90.610 168.920 ;
        RECT 95.930 167.960 97.040 169.360 ;
        RECT 100.260 169.200 101.780 169.390 ;
        RECT 97.770 168.970 102.770 169.200 ;
        RECT 95.960 167.920 97.040 167.960 ;
        RECT 90.770 167.880 95.770 167.910 ;
        RECT 90.740 166.990 95.790 167.880 ;
        RECT 90.770 166.970 95.770 166.990 ;
        RECT 96.700 166.970 97.040 167.920 ;
        RECT 97.270 167.900 97.620 168.940 ;
        RECT 100.260 168.870 101.780 168.970 ;
        RECT 102.930 167.960 103.160 168.920 ;
        RECT 97.770 167.880 102.770 167.910 ;
        RECT 97.770 167.680 102.800 167.880 ;
        RECT 97.980 167.200 102.800 167.680 ;
        RECT 97.770 166.990 102.800 167.200 ;
        RECT 97.770 166.970 102.770 166.990 ;
        RECT 86.880 164.220 87.540 164.270 ;
        RECT 81.510 164.100 87.540 164.220 ;
        RECT 81.510 163.940 81.840 164.100 ;
        RECT 82.050 164.020 87.540 164.100 ;
        RECT 82.050 163.990 87.050 164.020 ;
        RECT 81.510 163.480 81.845 163.940 ;
        RECT 81.510 159.440 81.840 163.480 ;
        RECT 82.140 163.430 82.860 163.650 ;
        RECT 82.050 163.200 87.050 163.430 ;
        RECT 82.140 163.080 82.860 163.200 ;
        RECT 87.210 163.020 87.540 164.020 ;
        RECT 89.720 166.920 90.580 166.950 ;
        RECT 89.720 165.960 90.610 166.920 ;
        RECT 89.720 165.940 90.580 165.960 ;
        RECT 89.720 165.360 90.040 165.940 ;
        RECT 90.760 165.910 92.650 166.180 ;
        RECT 95.930 165.960 96.160 166.920 ;
        RECT 96.700 165.920 97.610 166.970 ;
        RECT 90.760 165.680 95.770 165.910 ;
        RECT 90.760 165.560 92.650 165.680 ;
        RECT 96.700 165.390 97.040 165.920 ;
        RECT 98.190 165.910 99.710 166.070 ;
        RECT 102.930 165.960 103.160 166.920 ;
        RECT 97.770 165.680 102.770 165.910 ;
        RECT 98.190 165.550 99.710 165.680 ;
        RECT 89.720 163.730 90.050 165.360 ;
        RECT 87.210 162.130 87.870 163.020 ;
        RECT 82.010 159.720 82.630 159.930 ;
        RECT 82.010 159.490 87.050 159.720 ;
        RECT 81.510 158.980 81.845 159.440 ;
        RECT 82.010 159.430 82.630 159.490 ;
        RECT 81.510 158.920 81.840 158.980 ;
        RECT 82.190 158.930 82.910 159.070 ;
        RECT 87.210 158.930 87.540 162.130 ;
        RECT 89.720 161.280 90.040 163.730 ;
        RECT 93.080 163.200 94.810 163.530 ;
        RECT 90.770 162.970 95.770 163.200 ;
        RECT 96.710 162.940 97.030 165.390 ;
        RECT 97.220 163.870 97.610 164.900 ;
        RECT 95.970 162.920 97.030 162.940 ;
        RECT 90.380 161.960 90.610 162.920 ;
        RECT 95.930 161.960 97.030 162.920 ;
        RECT 95.970 161.940 97.030 161.960 ;
        RECT 90.770 161.880 95.770 161.910 ;
        RECT 88.930 160.940 90.040 161.280 ;
        RECT 90.750 160.990 95.800 161.880 ;
        RECT 90.770 160.970 95.770 160.990 ;
        RECT 96.710 160.960 97.030 161.940 ;
        RECT 97.330 161.930 97.610 163.870 ;
        RECT 105.790 164.820 106.070 170.230 ;
        RECT 110.230 169.220 111.180 169.310 ;
        RECT 111.380 169.270 112.530 170.240 ;
        RECT 106.230 168.990 111.240 169.220 ;
        RECT 110.230 168.910 111.180 168.990 ;
        RECT 111.420 168.940 111.810 169.270 ;
        RECT 106.230 167.930 107.150 167.990 ;
        RECT 111.390 167.980 111.810 168.940 ;
        RECT 106.230 167.920 111.230 167.930 ;
        RECT 106.230 167.690 111.240 167.920 ;
        RECT 106.230 167.620 107.150 167.690 ;
        RECT 111.420 167.650 111.810 167.980 ;
        RECT 111.390 166.690 111.810 167.650 ;
        RECT 110.230 166.640 111.180 166.690 ;
        RECT 106.230 166.630 111.230 166.640 ;
        RECT 106.230 166.410 111.240 166.630 ;
        RECT 106.280 166.400 111.240 166.410 ;
        RECT 110.230 166.310 111.180 166.400 ;
        RECT 111.420 166.360 111.810 166.690 ;
        RECT 106.230 165.350 107.160 165.440 ;
        RECT 111.390 165.400 111.810 166.360 ;
        RECT 106.230 165.120 111.240 165.350 ;
        RECT 106.230 165.060 107.160 165.120 ;
        RECT 111.420 165.070 111.810 165.400 ;
        RECT 111.390 164.820 111.810 165.070 ;
        RECT 105.790 164.370 106.160 164.820 ;
        RECT 111.340 164.370 111.810 164.820 ;
        RECT 100.290 163.200 101.810 163.400 ;
        RECT 97.770 162.970 102.770 163.200 ;
        RECT 100.290 162.880 101.810 162.970 ;
        RECT 102.930 161.960 103.160 162.920 ;
        RECT 97.770 161.890 102.770 161.910 ;
        RECT 97.750 161.700 102.790 161.890 ;
        RECT 97.740 161.000 102.790 161.700 ;
        RECT 97.770 160.970 102.770 161.000 ;
        RECT 96.710 160.940 97.580 160.960 ;
        RECT 88.930 160.920 90.590 160.940 ;
        RECT 96.710 160.920 97.600 160.940 ;
        RECT 88.930 159.960 90.610 160.920 ;
        RECT 95.930 159.960 96.160 160.920 ;
        RECT 96.710 159.960 97.610 160.920 ;
        RECT 88.930 159.930 90.520 159.960 ;
        RECT 90.800 159.910 92.520 159.960 ;
        RECT 96.720 159.950 97.580 159.960 ;
        RECT 98.200 159.910 99.720 160.100 ;
        RECT 102.930 159.960 103.160 160.920 ;
        RECT 90.770 159.680 95.770 159.910 ;
        RECT 97.770 159.680 102.770 159.910 ;
        RECT 90.800 159.540 92.520 159.680 ;
        RECT 98.200 159.580 99.720 159.680 ;
        RECT 104.040 159.380 104.620 161.030 ;
        RECT 105.790 160.220 106.070 164.370 ;
        RECT 110.230 164.060 111.170 164.140 ;
        RECT 111.390 164.110 111.810 164.370 ;
        RECT 106.230 164.050 111.230 164.060 ;
        RECT 106.230 163.830 111.240 164.050 ;
        RECT 106.280 163.820 111.240 163.830 ;
        RECT 110.230 163.750 111.170 163.820 ;
        RECT 111.420 163.780 111.810 164.110 ;
        RECT 106.230 162.770 107.150 162.890 ;
        RECT 111.390 162.820 111.810 163.780 ;
        RECT 106.230 162.540 111.240 162.770 ;
        RECT 106.230 162.470 107.150 162.540 ;
        RECT 111.420 162.490 111.810 162.820 ;
        RECT 110.150 161.480 111.250 161.720 ;
        RECT 111.390 161.530 111.810 162.490 ;
        RECT 113.340 163.580 113.960 171.460 ;
        RECT 122.725 171.395 123.625 172.195 ;
        RECT 123.815 171.600 124.775 171.830 ;
        RECT 125.105 171.805 126.065 171.830 ;
        RECT 126.825 171.805 127.515 172.345 ;
        RECT 130.410 172.285 130.955 172.805 ;
        RECT 125.105 171.635 128.905 171.805 ;
        RECT 125.105 171.600 126.065 171.635 ;
        RECT 122.725 169.395 123.765 171.395 ;
        RECT 122.725 168.565 123.625 169.395 ;
        RECT 123.985 169.190 124.505 171.600 ;
        RECT 124.825 169.395 125.055 171.395 ;
        RECT 125.315 169.190 125.835 171.600 ;
        RECT 126.135 171.395 127.855 171.415 ;
        RECT 126.115 170.965 127.855 171.395 ;
        RECT 128.065 171.355 128.905 171.635 ;
        RECT 128.005 171.125 128.965 171.355 ;
        RECT 129.295 171.125 130.255 171.355 ;
        RECT 126.115 169.965 127.955 170.965 ;
        RECT 126.115 169.395 127.855 169.965 ;
        RECT 128.245 169.805 128.765 171.125 ;
        RECT 129.015 169.965 129.245 170.965 ;
        RECT 129.515 169.805 130.035 171.125 ;
        RECT 130.415 170.965 130.955 172.285 ;
        RECT 130.305 169.965 130.955 170.965 ;
        RECT 128.005 169.575 128.965 169.805 ;
        RECT 129.295 169.575 130.255 169.805 ;
        RECT 130.415 169.435 130.955 169.965 ;
        RECT 126.135 169.375 127.855 169.395 ;
        RECT 123.815 168.960 124.775 169.190 ;
        RECT 125.105 168.960 126.065 169.190 ;
        RECT 126.825 168.965 127.515 169.375 ;
        RECT 130.405 169.315 130.955 169.435 ;
        RECT 122.725 168.385 123.205 168.565 ;
        RECT 116.950 164.850 119.550 167.100 ;
        RECT 113.340 162.440 115.105 163.580 ;
        RECT 117.990 163.410 118.960 164.850 ;
        RECT 122.720 164.435 123.640 168.385 ;
        RECT 126.815 168.345 127.515 168.965 ;
        RECT 130.395 168.795 130.955 169.315 ;
        RECT 126.830 164.485 127.500 168.345 ;
        RECT 130.395 168.175 130.960 168.795 ;
        RECT 130.420 164.705 130.960 168.175 ;
        RECT 122.725 163.580 123.625 164.435 ;
        RECT 121.875 163.450 123.625 163.580 ;
        RECT 123.815 163.500 124.775 163.730 ;
        RECT 125.105 163.705 126.065 163.730 ;
        RECT 126.825 163.705 127.515 164.485 ;
        RECT 130.415 163.895 130.960 164.705 ;
        RECT 125.105 163.535 128.905 163.705 ;
        RECT 125.105 163.500 126.065 163.535 ;
        RECT 113.340 162.320 115.095 162.440 ;
        RECT 117.985 162.380 118.960 163.410 ;
        RECT 121.870 163.295 123.625 163.450 ;
        RECT 119.435 162.565 120.395 162.795 ;
        RECT 120.725 162.565 121.685 162.795 ;
        RECT 117.645 162.360 119.365 162.380 ;
        RECT 113.340 161.790 115.085 162.320 ;
        RECT 115.245 161.950 116.205 162.180 ;
        RECT 116.535 161.950 117.495 162.180 ;
        RECT 113.340 161.710 115.195 161.790 ;
        RECT 106.230 161.250 111.250 161.480 ;
        RECT 110.150 161.050 111.250 161.250 ;
        RECT 111.420 161.200 111.810 161.530 ;
        RECT 106.230 160.190 107.150 160.310 ;
        RECT 111.390 160.240 111.810 161.200 ;
        RECT 113.170 161.050 115.195 161.710 ;
        RECT 111.420 160.220 111.810 160.240 ;
        RECT 113.340 160.790 115.195 161.050 ;
        RECT 106.230 159.960 111.250 160.190 ;
        RECT 106.230 159.890 107.150 159.960 ;
        RECT 113.340 159.380 115.085 160.790 ;
        RECT 115.465 160.630 115.985 161.950 ;
        RECT 116.255 160.790 116.485 161.790 ;
        RECT 116.735 160.630 117.255 161.950 ;
        RECT 117.645 161.790 119.385 162.360 ;
        RECT 117.545 160.790 119.385 161.790 ;
        RECT 115.245 160.400 116.205 160.630 ;
        RECT 116.535 160.400 117.495 160.630 ;
        RECT 116.595 160.120 117.435 160.400 ;
        RECT 117.645 160.360 119.385 160.790 ;
        RECT 117.645 160.340 119.365 160.360 ;
        RECT 119.665 160.155 120.185 162.565 ;
        RECT 120.445 160.360 120.675 162.360 ;
        RECT 120.995 160.155 121.515 162.565 ;
        RECT 121.870 162.360 123.765 163.295 ;
        RECT 121.735 161.295 123.765 162.360 ;
        RECT 121.735 160.605 123.625 161.295 ;
        RECT 123.985 161.090 124.505 163.500 ;
        RECT 124.825 161.295 125.055 163.295 ;
        RECT 125.315 161.090 125.835 163.500 ;
        RECT 126.135 163.295 127.855 163.315 ;
        RECT 126.115 162.865 127.855 163.295 ;
        RECT 128.065 163.255 128.905 163.535 ;
        RECT 128.005 163.025 128.965 163.255 ;
        RECT 129.295 163.025 130.255 163.255 ;
        RECT 126.115 161.865 127.955 162.865 ;
        RECT 126.115 161.295 127.855 161.865 ;
        RECT 128.245 161.705 128.765 163.025 ;
        RECT 129.015 161.865 129.245 162.865 ;
        RECT 129.515 161.705 130.035 163.025 ;
        RECT 130.415 162.865 130.955 163.895 ;
        RECT 130.305 161.865 130.955 162.865 ;
        RECT 128.005 161.475 128.965 161.705 ;
        RECT 129.295 161.475 130.255 161.705 ;
        RECT 130.415 161.335 130.955 161.865 ;
        RECT 126.135 161.275 127.855 161.295 ;
        RECT 123.815 160.860 124.775 161.090 ;
        RECT 125.105 160.860 126.065 161.090 ;
        RECT 126.825 160.865 127.515 161.275 ;
        RECT 130.405 161.215 130.955 161.335 ;
        RECT 121.735 160.360 123.630 160.605 ;
        RECT 119.435 160.120 120.395 160.155 ;
        RECT 116.595 159.950 120.395 160.120 ;
        RECT 104.040 159.040 115.085 159.380 ;
        RECT 117.985 159.170 118.680 159.950 ;
        RECT 119.435 159.925 120.395 159.950 ;
        RECT 120.725 159.925 121.685 160.155 ;
        RECT 121.870 159.955 123.630 160.360 ;
        RECT 126.815 160.245 127.515 160.865 ;
        RECT 130.395 160.605 130.955 161.215 ;
        RECT 82.050 158.700 87.050 158.930 ;
        RECT 82.190 158.500 82.910 158.700 ;
        RECT 104.040 158.520 115.105 159.040 ;
        RECT 117.990 158.870 118.680 159.170 ;
        RECT 80.630 157.760 81.310 158.240 ;
        RECT 113.340 157.900 115.105 158.520 ;
        RECT 117.985 158.250 118.685 158.870 ;
        RECT 121.870 158.420 123.620 159.955 ;
        RECT 113.340 157.780 115.095 157.900 ;
        RECT 117.985 157.840 118.675 158.250 ;
        RECT 119.435 158.025 120.395 158.255 ;
        RECT 120.725 158.025 121.685 158.255 ;
        RECT 117.645 157.820 119.365 157.840 ;
        RECT 113.340 157.250 115.085 157.780 ;
        RECT 115.245 157.410 116.205 157.640 ;
        RECT 116.535 157.410 117.495 157.640 ;
        RECT 80.630 155.980 81.310 156.460 ;
        RECT 113.340 156.250 115.195 157.250 ;
        RECT 77.070 155.520 78.020 155.600 ;
        RECT 72.530 154.710 72.860 155.320 ;
        RECT 73.050 155.290 78.050 155.520 ;
        RECT 77.070 155.160 78.020 155.290 ;
        RECT 78.230 154.780 78.560 155.270 ;
        RECT 77.270 154.730 78.560 154.780 ;
        RECT 73.050 154.710 78.560 154.730 ;
        RECT 72.530 154.500 78.560 154.710 ;
        RECT 72.530 154.450 73.370 154.500 ;
        RECT 77.270 154.490 78.560 154.500 ;
        RECT 72.530 145.890 72.860 154.450 ;
        RECT 77.090 151.020 78.030 151.210 ;
        RECT 73.050 150.790 78.050 151.020 ;
        RECT 77.090 150.740 78.030 150.790 ;
        RECT 77.090 150.230 78.060 150.330 ;
        RECT 73.050 150.000 78.060 150.230 ;
        RECT 77.090 149.610 78.060 150.000 ;
        RECT 77.090 146.520 78.090 146.670 ;
        RECT 73.050 146.290 78.090 146.520 ;
        RECT 77.090 146.210 78.090 146.290 ;
        RECT 72.530 145.800 73.280 145.890 ;
        RECT 78.230 145.830 78.560 154.490 ;
        RECT 72.560 145.730 73.280 145.800 ;
        RECT 77.260 145.750 78.560 145.830 ;
        RECT 77.260 145.730 78.510 145.750 ;
        RECT 72.560 145.520 78.510 145.730 ;
        RECT 73.050 145.500 78.510 145.520 ;
        RECT 77.260 145.480 78.510 145.500 ;
        RECT 78.750 145.390 79.140 155.850 ;
        RECT 79.680 145.310 80.320 155.800 ;
        RECT 80.800 143.650 81.190 155.980 ;
        RECT 82.190 155.520 82.910 155.720 ;
        RECT 113.340 155.700 115.085 156.250 ;
        RECT 115.465 156.090 115.985 157.410 ;
        RECT 116.255 156.250 116.485 157.250 ;
        RECT 116.735 156.090 117.255 157.410 ;
        RECT 117.645 157.250 119.385 157.820 ;
        RECT 117.545 156.250 119.385 157.250 ;
        RECT 115.245 155.860 116.205 156.090 ;
        RECT 116.535 155.860 117.495 156.090 ;
        RECT 81.510 155.240 81.840 155.300 ;
        RECT 82.050 155.290 87.050 155.520 ;
        RECT 81.510 154.780 81.845 155.240 ;
        RECT 82.190 155.150 82.910 155.290 ;
        RECT 81.510 150.740 81.840 154.780 ;
        RECT 82.010 154.730 82.630 154.790 ;
        RECT 82.010 154.500 87.050 154.730 ;
        RECT 82.010 154.290 82.630 154.500 ;
        RECT 87.210 152.090 87.540 155.290 ;
        RECT 104.040 154.980 115.085 155.700 ;
        RECT 116.595 155.580 117.435 155.860 ;
        RECT 117.645 155.820 119.385 156.250 ;
        RECT 117.645 155.800 119.365 155.820 ;
        RECT 119.665 155.615 120.185 158.025 ;
        RECT 120.445 155.820 120.675 157.820 ;
        RECT 120.995 155.615 121.515 158.025 ;
        RECT 121.875 157.820 123.620 158.420 ;
        RECT 121.735 156.605 123.620 157.820 ;
        RECT 121.735 155.820 123.625 156.605 ;
        RECT 126.820 156.385 127.510 160.245 ;
        RECT 130.395 160.075 130.960 160.605 ;
        RECT 126.820 155.945 127.515 156.385 ;
        RECT 119.435 155.580 120.395 155.615 ;
        RECT 116.595 155.410 120.395 155.580 ;
        RECT 104.040 154.840 115.105 154.980 ;
        RECT 90.800 154.540 92.520 154.680 ;
        RECT 98.200 154.540 99.720 154.640 ;
        RECT 90.770 154.310 95.770 154.540 ;
        RECT 97.770 154.310 102.770 154.540 ;
        RECT 88.930 154.260 90.520 154.290 ;
        RECT 90.800 154.260 92.520 154.310 ;
        RECT 96.720 154.260 97.580 154.270 ;
        RECT 88.930 153.300 90.610 154.260 ;
        RECT 95.930 153.300 96.160 154.260 ;
        RECT 96.710 153.300 97.610 154.260 ;
        RECT 98.200 154.120 99.720 154.310 ;
        RECT 102.930 153.300 103.160 154.260 ;
        RECT 88.930 153.280 90.590 153.300 ;
        RECT 96.710 153.280 97.600 153.300 ;
        RECT 88.930 152.940 90.040 153.280 ;
        RECT 96.710 153.260 97.580 153.280 ;
        RECT 90.770 153.230 95.770 153.250 ;
        RECT 87.210 151.200 87.870 152.090 ;
        RECT 82.140 151.020 82.860 151.140 ;
        RECT 82.050 150.790 87.050 151.020 ;
        RECT 81.510 150.280 81.845 150.740 ;
        RECT 82.140 150.570 82.860 150.790 ;
        RECT 81.510 150.120 81.840 150.280 ;
        RECT 82.050 150.200 87.050 150.230 ;
        RECT 87.210 150.200 87.540 151.200 ;
        RECT 82.050 150.120 87.540 150.200 ;
        RECT 81.510 150.000 87.540 150.120 ;
        RECT 81.510 149.770 82.830 150.000 ;
        RECT 86.880 149.950 87.540 150.000 ;
        RECT 81.510 146.240 81.840 149.770 ;
        RECT 82.080 146.520 82.900 146.690 ;
        RECT 82.050 146.290 87.050 146.520 ;
        RECT 81.510 145.780 81.845 146.240 ;
        RECT 82.080 146.190 82.900 146.290 ;
        RECT 82.020 145.730 82.680 145.750 ;
        RECT 85.030 145.730 86.830 145.880 ;
        RECT 87.210 145.770 87.540 149.950 ;
        RECT 89.720 150.490 90.040 152.940 ;
        RECT 90.750 152.340 95.800 153.230 ;
        RECT 90.770 152.310 95.770 152.340 ;
        RECT 96.710 152.280 97.030 153.260 ;
        RECT 97.770 153.220 102.770 153.250 ;
        RECT 97.740 152.520 102.790 153.220 ;
        RECT 104.040 153.190 104.620 154.840 ;
        RECT 106.230 154.260 107.150 154.330 ;
        RECT 106.230 154.030 111.250 154.260 ;
        RECT 97.750 152.330 102.790 152.520 ;
        RECT 97.770 152.310 102.770 152.330 ;
        RECT 95.970 152.260 97.030 152.280 ;
        RECT 90.380 151.300 90.610 152.260 ;
        RECT 95.930 151.300 97.030 152.260 ;
        RECT 95.970 151.280 97.030 151.300 ;
        RECT 90.770 151.020 95.770 151.250 ;
        RECT 93.080 150.690 94.810 151.020 ;
        RECT 89.720 148.860 90.050 150.490 ;
        RECT 89.720 148.280 90.040 148.860 ;
        RECT 96.710 148.830 97.030 151.280 ;
        RECT 97.330 150.350 97.610 152.290 ;
        RECT 100.290 151.250 101.810 151.340 ;
        RECT 102.930 151.300 103.160 152.260 ;
        RECT 97.770 151.020 102.770 151.250 ;
        RECT 100.290 150.820 101.810 151.020 ;
        RECT 97.220 149.320 97.610 150.350 ;
        RECT 105.790 149.850 106.070 154.000 ;
        RECT 106.230 153.910 107.150 154.030 ;
        RECT 111.420 153.980 111.810 154.000 ;
        RECT 110.150 152.970 111.250 153.170 ;
        RECT 111.390 153.020 111.810 153.980 ;
        RECT 113.340 153.840 115.105 154.840 ;
        RECT 117.985 154.810 118.675 155.410 ;
        RECT 119.435 155.385 120.395 155.410 ;
        RECT 120.725 155.385 121.685 155.615 ;
        RECT 121.875 155.195 123.625 155.820 ;
        RECT 123.815 155.400 124.775 155.630 ;
        RECT 125.105 155.605 126.065 155.630 ;
        RECT 126.825 155.605 127.515 155.945 ;
        RECT 125.105 155.435 128.905 155.605 ;
        RECT 125.105 155.400 126.065 155.435 ;
        RECT 117.985 154.190 118.685 154.810 ;
        RECT 113.340 153.720 115.095 153.840 ;
        RECT 117.985 153.780 118.675 154.190 ;
        RECT 119.435 153.965 120.395 154.195 ;
        RECT 120.725 153.965 121.685 154.195 ;
        RECT 117.645 153.760 119.365 153.780 ;
        RECT 113.340 153.190 115.085 153.720 ;
        RECT 115.245 153.350 116.205 153.580 ;
        RECT 116.535 153.350 117.495 153.580 ;
        RECT 113.340 153.170 115.195 153.190 ;
        RECT 106.230 152.740 111.250 152.970 ;
        RECT 110.150 152.500 111.250 152.740 ;
        RECT 111.420 152.690 111.810 153.020 ;
        RECT 106.230 151.680 107.150 151.750 ;
        RECT 111.390 151.730 111.810 152.690 ;
        RECT 113.170 152.510 115.195 153.170 ;
        RECT 106.230 151.450 111.240 151.680 ;
        RECT 106.230 151.330 107.150 151.450 ;
        RECT 111.420 151.400 111.810 151.730 ;
        RECT 110.230 150.400 111.170 150.470 ;
        RECT 111.390 150.440 111.810 151.400 ;
        RECT 106.280 150.390 111.240 150.400 ;
        RECT 106.230 150.170 111.240 150.390 ;
        RECT 106.230 150.160 111.230 150.170 ;
        RECT 110.230 150.080 111.170 150.160 ;
        RECT 111.420 150.110 111.810 150.440 ;
        RECT 111.390 149.850 111.810 150.110 ;
        RECT 105.790 149.400 106.160 149.850 ;
        RECT 111.340 149.400 111.810 149.850 ;
        RECT 90.760 148.540 92.650 148.660 ;
        RECT 90.760 148.310 95.770 148.540 ;
        RECT 89.720 148.260 90.580 148.280 ;
        RECT 89.720 147.300 90.610 148.260 ;
        RECT 90.760 148.040 92.650 148.310 ;
        RECT 96.700 148.300 97.040 148.830 ;
        RECT 98.190 148.540 99.710 148.670 ;
        RECT 97.770 148.310 102.770 148.540 ;
        RECT 95.930 147.300 96.160 148.260 ;
        RECT 89.720 147.270 90.580 147.300 ;
        RECT 96.700 147.250 97.610 148.300 ;
        RECT 98.190 148.150 99.710 148.310 ;
        RECT 102.930 147.300 103.160 148.260 ;
        RECT 90.770 147.230 95.770 147.250 ;
        RECT 90.740 146.340 95.790 147.230 ;
        RECT 90.770 146.310 95.770 146.340 ;
        RECT 96.700 146.300 97.040 147.250 ;
        RECT 97.770 147.230 102.770 147.250 ;
        RECT 97.770 147.020 102.800 147.230 ;
        RECT 97.980 146.540 102.800 147.020 ;
        RECT 97.770 146.340 102.800 146.540 ;
        RECT 95.960 146.260 97.040 146.300 ;
        RECT 82.020 145.500 87.050 145.730 ;
        RECT 82.020 145.280 82.680 145.500 ;
        RECT 85.030 145.060 86.830 145.500 ;
        RECT 90.380 145.300 90.610 146.260 ;
        RECT 90.770 145.020 95.770 145.250 ;
        RECT 93.080 144.680 94.810 145.020 ;
        RECT 95.930 144.860 97.040 146.260 ;
        RECT 97.270 145.280 97.620 146.320 ;
        RECT 97.770 146.310 102.770 146.340 ;
        RECT 100.260 145.250 101.780 145.350 ;
        RECT 102.930 145.300 103.160 146.260 ;
        RECT 97.770 145.020 102.770 145.250 ;
        RECT 100.260 144.830 101.780 145.020 ;
        RECT 105.790 143.990 106.070 149.400 ;
        RECT 106.230 149.100 107.160 149.160 ;
        RECT 111.390 149.150 111.810 149.400 ;
        RECT 106.230 148.870 111.240 149.100 ;
        RECT 106.230 148.780 107.160 148.870 ;
        RECT 111.420 148.820 111.810 149.150 ;
        RECT 110.230 147.820 111.180 147.910 ;
        RECT 111.390 147.860 111.810 148.820 ;
        RECT 106.280 147.810 111.240 147.820 ;
        RECT 106.230 147.590 111.240 147.810 ;
        RECT 106.230 147.580 111.230 147.590 ;
        RECT 110.230 147.530 111.180 147.580 ;
        RECT 111.420 147.530 111.810 147.860 ;
        RECT 106.230 146.530 107.150 146.600 ;
        RECT 111.390 146.570 111.810 147.530 ;
        RECT 106.230 146.300 111.240 146.530 ;
        RECT 106.230 146.290 111.230 146.300 ;
        RECT 106.230 146.230 107.150 146.290 ;
        RECT 111.420 146.240 111.810 146.570 ;
        RECT 110.230 145.230 111.180 145.310 ;
        RECT 111.390 145.280 111.810 146.240 ;
        RECT 106.230 145.000 111.240 145.230 ;
        RECT 110.230 144.910 111.180 145.000 ;
        RECT 111.420 144.950 111.810 145.280 ;
        RECT 113.340 152.190 115.195 152.510 ;
        RECT 113.340 150.920 115.085 152.190 ;
        RECT 115.465 152.030 115.985 153.350 ;
        RECT 116.255 152.190 116.485 153.190 ;
        RECT 116.735 152.030 117.255 153.350 ;
        RECT 117.645 153.190 119.385 153.760 ;
        RECT 117.545 152.190 119.385 153.190 ;
        RECT 115.245 151.800 116.205 152.030 ;
        RECT 116.535 151.800 117.495 152.030 ;
        RECT 116.595 151.520 117.435 151.800 ;
        RECT 117.645 151.760 119.385 152.190 ;
        RECT 117.645 151.740 119.365 151.760 ;
        RECT 119.665 151.555 120.185 153.965 ;
        RECT 120.445 151.760 120.675 153.760 ;
        RECT 120.995 151.555 121.515 153.965 ;
        RECT 121.875 153.760 123.765 155.195 ;
        RECT 121.735 153.195 123.765 153.760 ;
        RECT 121.735 152.365 123.625 153.195 ;
        RECT 123.985 152.990 124.505 155.400 ;
        RECT 124.825 153.195 125.055 155.195 ;
        RECT 125.315 152.990 125.835 155.400 ;
        RECT 126.135 155.195 127.855 155.215 ;
        RECT 126.115 154.765 127.855 155.195 ;
        RECT 128.065 155.155 128.905 155.435 ;
        RECT 128.005 154.925 128.965 155.155 ;
        RECT 129.295 154.925 130.255 155.155 ;
        RECT 126.115 153.765 127.955 154.765 ;
        RECT 126.115 153.195 127.855 153.765 ;
        RECT 128.245 153.605 128.765 154.925 ;
        RECT 129.015 153.765 129.245 154.765 ;
        RECT 129.515 153.605 130.035 154.925 ;
        RECT 130.410 154.765 130.960 160.075 ;
        RECT 130.305 153.765 130.960 154.765 ;
        RECT 128.005 153.375 128.965 153.605 ;
        RECT 129.295 153.375 130.255 153.605 ;
        RECT 130.410 153.235 130.960 153.765 ;
        RECT 126.135 153.175 127.855 153.195 ;
        RECT 123.815 152.760 124.775 152.990 ;
        RECT 125.105 152.760 126.065 152.990 ;
        RECT 126.825 152.765 127.515 153.175 ;
        RECT 130.405 153.115 130.960 153.235 ;
        RECT 126.815 152.495 127.515 152.765 ;
        RECT 121.735 152.185 123.205 152.365 ;
        RECT 121.735 152.105 123.625 152.185 ;
        RECT 126.815 152.145 127.520 152.495 ;
        RECT 121.735 151.760 123.630 152.105 ;
        RECT 119.435 151.520 120.395 151.555 ;
        RECT 116.595 151.350 120.395 151.520 ;
        RECT 113.340 149.780 115.105 150.920 ;
        RECT 117.985 150.750 118.675 151.350 ;
        RECT 119.435 151.325 120.395 151.350 ;
        RECT 120.725 151.325 121.685 151.555 ;
        RECT 117.985 150.130 118.685 150.750 ;
        RECT 113.340 149.660 115.095 149.780 ;
        RECT 117.985 149.720 118.675 150.130 ;
        RECT 119.435 149.905 120.395 150.135 ;
        RECT 120.725 149.905 121.685 150.135 ;
        RECT 117.645 149.700 119.365 149.720 ;
        RECT 113.340 149.130 115.085 149.660 ;
        RECT 115.245 149.290 116.205 149.520 ;
        RECT 116.535 149.290 117.495 149.520 ;
        RECT 113.340 148.130 115.195 149.130 ;
        RECT 113.340 146.860 115.085 148.130 ;
        RECT 115.465 147.970 115.985 149.290 ;
        RECT 116.255 148.130 116.485 149.130 ;
        RECT 116.735 147.970 117.255 149.290 ;
        RECT 117.645 149.130 119.385 149.700 ;
        RECT 117.545 148.130 119.385 149.130 ;
        RECT 115.245 147.740 116.205 147.970 ;
        RECT 116.535 147.740 117.495 147.970 ;
        RECT 116.595 147.460 117.435 147.740 ;
        RECT 117.645 147.700 119.385 148.130 ;
        RECT 117.645 147.680 119.365 147.700 ;
        RECT 119.665 147.495 120.185 149.905 ;
        RECT 120.445 147.700 120.675 149.700 ;
        RECT 120.995 147.495 121.515 149.905 ;
        RECT 121.875 149.700 123.630 151.760 ;
        RECT 121.735 148.145 123.630 149.700 ;
        RECT 121.735 147.700 123.625 148.145 ;
        RECT 126.820 147.995 127.520 152.145 ;
        RECT 130.395 151.975 130.960 153.115 ;
        RECT 130.410 148.405 130.960 151.975 ;
        RECT 119.435 147.460 120.395 147.495 ;
        RECT 116.595 147.290 120.395 147.460 ;
        RECT 113.340 145.720 115.105 146.860 ;
        RECT 117.985 146.690 118.675 147.290 ;
        RECT 119.435 147.265 120.395 147.290 ;
        RECT 120.725 147.265 121.685 147.495 ;
        RECT 121.875 147.095 123.625 147.700 ;
        RECT 123.815 147.300 124.775 147.530 ;
        RECT 125.105 147.505 126.065 147.530 ;
        RECT 126.825 147.505 127.515 147.995 ;
        RECT 125.105 147.335 128.905 147.505 ;
        RECT 125.105 147.300 126.065 147.335 ;
        RECT 117.985 146.070 118.685 146.690 ;
        RECT 113.340 145.600 115.095 145.720 ;
        RECT 117.985 145.660 118.675 146.070 ;
        RECT 119.435 145.845 120.395 146.075 ;
        RECT 120.725 145.845 121.685 146.075 ;
        RECT 117.645 145.640 119.365 145.660 ;
        RECT 113.340 145.070 115.085 145.600 ;
        RECT 115.245 145.230 116.205 145.460 ;
        RECT 116.535 145.230 117.495 145.460 ;
        RECT 106.220 143.940 107.150 143.990 ;
        RECT 111.380 143.980 112.530 144.950 ;
        RECT 113.340 144.070 115.195 145.070 ;
        RECT 106.220 143.710 111.230 143.940 ;
        RECT 106.220 143.670 107.150 143.710 ;
        RECT 80.240 142.850 81.470 143.650 ;
        RECT 71.770 142.190 96.350 142.850 ;
        RECT 113.340 142.800 115.085 144.070 ;
        RECT 115.465 143.910 115.985 145.230 ;
        RECT 116.255 144.070 116.485 145.070 ;
        RECT 116.735 143.910 117.255 145.230 ;
        RECT 117.645 145.070 119.385 145.640 ;
        RECT 117.545 144.070 119.385 145.070 ;
        RECT 115.245 143.680 116.205 143.910 ;
        RECT 116.535 143.680 117.495 143.910 ;
        RECT 116.595 143.400 117.435 143.680 ;
        RECT 117.645 143.640 119.385 144.070 ;
        RECT 117.645 143.620 119.365 143.640 ;
        RECT 119.665 143.435 120.185 145.845 ;
        RECT 120.445 143.640 120.675 145.640 ;
        RECT 120.995 143.435 121.515 145.845 ;
        RECT 121.875 145.640 123.765 147.095 ;
        RECT 121.735 145.095 123.765 145.640 ;
        RECT 121.735 144.405 123.625 145.095 ;
        RECT 123.985 144.890 124.505 147.300 ;
        RECT 124.825 145.095 125.055 147.095 ;
        RECT 125.315 144.890 125.835 147.300 ;
        RECT 126.135 147.095 127.855 147.115 ;
        RECT 126.115 146.665 127.855 147.095 ;
        RECT 128.065 147.055 128.905 147.335 ;
        RECT 128.005 146.825 128.965 147.055 ;
        RECT 129.295 146.825 130.255 147.055 ;
        RECT 126.115 145.665 127.955 146.665 ;
        RECT 126.115 145.095 127.855 145.665 ;
        RECT 128.245 145.505 128.765 146.825 ;
        RECT 129.015 145.665 129.245 146.665 ;
        RECT 129.515 145.505 130.035 146.825 ;
        RECT 130.415 146.665 130.955 148.405 ;
        RECT 130.305 145.665 130.955 146.665 ;
        RECT 128.005 145.275 128.965 145.505 ;
        RECT 129.295 145.275 130.255 145.505 ;
        RECT 130.415 145.135 130.955 145.665 ;
        RECT 126.135 145.075 127.855 145.095 ;
        RECT 123.815 144.660 124.775 144.890 ;
        RECT 125.105 144.660 126.065 144.890 ;
        RECT 126.825 144.665 127.515 145.075 ;
        RECT 130.405 145.015 130.955 145.135 ;
        RECT 121.735 143.640 123.630 144.405 ;
        RECT 126.815 144.385 127.515 144.665 ;
        RECT 126.815 144.045 127.520 144.385 ;
        RECT 119.435 143.400 120.395 143.435 ;
        RECT 116.595 143.230 120.395 143.400 ;
        RECT 113.340 142.760 115.105 142.800 ;
        RECT 71.770 141.860 95.000 142.190 ;
        RECT 95.570 142.130 96.350 142.190 ;
        RECT 103.305 142.130 105.730 142.250 ;
        RECT 95.570 141.930 103.095 142.130 ;
        RECT 95.595 141.900 103.095 141.930 ;
        RECT 103.305 142.040 105.755 142.130 ;
        RECT 103.305 142.020 104.090 142.040 ;
        RECT 71.770 124.610 72.690 141.860 ;
        RECT 94.510 141.020 95.000 141.860 ;
        RECT 103.305 141.850 103.535 142.020 ;
        RECT 103.710 141.990 104.090 142.020 ;
        RECT 104.755 141.900 105.755 142.040 ;
        RECT 107.880 142.070 115.105 142.760 ;
        RECT 107.880 141.920 112.900 142.070 ;
        RECT 113.450 141.920 115.105 142.070 ;
        RECT 107.900 141.895 112.900 141.920 ;
        RECT 95.160 141.640 95.390 141.850 ;
        RECT 95.160 141.390 96.170 141.640 ;
        RECT 95.190 141.340 96.170 141.390 ;
        RECT 103.300 141.340 103.535 141.850 ;
        RECT 104.165 141.340 104.555 141.850 ;
        RECT 105.950 141.340 106.240 141.870 ;
        RECT 95.190 141.300 103.535 141.340 ;
        RECT 95.595 141.110 103.535 141.300 ;
        RECT 94.510 140.810 95.410 141.020 ;
        RECT 94.510 140.460 103.040 140.810 ;
        RECT 94.510 135.620 95.410 140.460 ;
        RECT 96.150 139.770 97.060 140.090 ;
        RECT 97.420 140.060 103.040 140.460 ;
        RECT 103.840 140.580 106.240 141.340 ;
        RECT 107.510 141.590 107.740 141.845 ;
        RECT 113.060 141.590 113.290 141.845 ;
        RECT 107.510 141.250 113.290 141.590 ;
        RECT 107.510 140.885 107.740 141.250 ;
        RECT 113.060 140.885 113.290 141.250 ;
        RECT 113.470 141.660 115.105 141.920 ;
        RECT 117.985 142.630 118.675 143.230 ;
        RECT 119.435 143.205 120.395 143.230 ;
        RECT 120.725 143.205 121.685 143.435 ;
        RECT 117.985 142.010 118.685 142.630 ;
        RECT 113.470 141.540 115.095 141.660 ;
        RECT 117.985 141.600 118.675 142.010 ;
        RECT 119.435 141.785 120.395 142.015 ;
        RECT 120.725 141.785 121.685 142.015 ;
        RECT 117.645 141.580 119.365 141.600 ;
        RECT 113.470 141.010 115.085 141.540 ;
        RECT 115.245 141.170 116.205 141.400 ;
        RECT 116.535 141.170 117.495 141.400 ;
        RECT 107.900 140.820 112.900 140.835 ;
        RECT 107.900 140.610 112.930 140.820 ;
        RECT 103.840 140.470 107.630 140.580 ;
        RECT 107.895 140.470 112.930 140.610 ;
        RECT 103.840 140.340 112.930 140.470 ;
        RECT 103.840 140.330 106.240 140.340 ;
        RECT 96.130 139.755 103.100 139.770 ;
        RECT 96.090 139.525 103.100 139.755 ;
        RECT 103.840 139.680 104.010 140.330 ;
        RECT 107.410 140.280 108.110 140.340 ;
        RECT 95.610 137.070 95.900 139.500 ;
        RECT 96.130 139.430 103.100 139.525 ;
        RECT 103.290 139.380 104.010 139.680 ;
        RECT 113.470 140.010 115.195 141.010 ;
        RECT 96.080 137.610 103.120 138.970 ;
        RECT 103.290 138.460 103.590 139.380 ;
        RECT 96.090 137.595 103.090 137.610 ;
        RECT 96.150 137.100 97.060 137.120 ;
        RECT 96.130 137.035 103.100 137.100 ;
        RECT 103.290 137.070 103.580 138.460 ;
        RECT 96.090 136.805 103.100 137.035 ;
        RECT 96.130 136.760 103.100 136.805 ;
        RECT 96.150 136.560 97.060 136.760 ;
        RECT 94.510 134.790 99.010 135.620 ;
        RECT 70.330 111.400 70.950 115.870 ;
        RECT 18.560 105.450 19.960 106.670 ;
        RECT 15.000 102.630 17.130 104.780 ;
        RECT 19.460 96.950 19.710 105.450 ;
        RECT 70.340 97.330 70.950 111.400 ;
        RECT 59.810 96.960 70.950 97.330 ;
        RECT 19.270 96.410 19.820 96.950 ;
        RECT 19.100 77.630 19.710 95.890 ;
        RECT 20.770 82.790 21.390 85.450 ;
        RECT 20.770 82.170 60.820 82.790 ;
        RECT 60.200 80.740 60.820 82.170 ;
        RECT 60.200 79.750 60.830 80.740 ;
        RECT 63.890 80.000 64.520 81.150 ;
        RECT 64.810 80.280 66.010 80.380 ;
        RECT 64.700 80.050 69.700 80.280 ;
        RECT 64.810 80.020 66.010 80.050 ;
        RECT 69.870 80.000 70.180 80.110 ;
        RECT 63.890 79.930 64.540 80.000 ;
        RECT 60.210 79.410 60.830 79.750 ;
        RECT 64.210 79.540 64.540 79.930 ;
        RECT 15.000 72.210 15.500 77.630 ;
        RECT 16.610 76.440 19.710 77.630 ;
        RECT 16.610 75.760 28.040 76.440 ;
        RECT 16.610 75.480 19.140 75.760 ;
        RECT 16.600 72.210 19.130 74.360 ;
        RECT 18.370 47.200 19.130 72.210 ;
        RECT 20.740 72.200 22.870 74.350 ;
        RECT 24.000 72.200 26.130 74.350 ;
        RECT 27.360 56.590 28.040 75.760 ;
        RECT 55.590 65.160 56.010 77.970 ;
        RECT 60.210 77.910 61.470 79.410 ;
        RECT 64.210 79.210 64.520 79.540 ;
        RECT 68.220 79.490 69.500 79.590 ;
        RECT 69.860 79.540 70.180 80.000 ;
        RECT 70.340 79.890 70.950 96.960 ;
        RECT 64.700 79.260 69.700 79.490 ;
        RECT 68.220 79.230 69.500 79.260 ;
        RECT 69.870 79.210 70.180 79.540 ;
        RECT 64.210 78.750 64.540 79.210 ;
        RECT 64.810 78.760 65.990 78.790 ;
        RECT 64.210 78.420 64.520 78.750 ;
        RECT 64.810 78.700 66.000 78.760 ;
        RECT 69.860 78.750 70.180 79.210 ;
        RECT 64.700 78.470 69.700 78.700 ;
        RECT 64.810 78.420 66.000 78.470 ;
        RECT 69.870 78.420 70.180 78.750 ;
        RECT 64.210 77.960 64.540 78.420 ;
        RECT 64.810 78.370 65.990 78.420 ;
        RECT 64.210 77.630 64.520 77.960 ;
        RECT 68.230 77.910 69.500 78.040 ;
        RECT 69.860 77.960 70.180 78.420 ;
        RECT 64.700 77.680 69.700 77.910 ;
        RECT 68.230 77.650 69.500 77.680 ;
        RECT 69.870 77.630 70.180 77.960 ;
        RECT 64.210 77.170 64.540 77.630 ;
        RECT 64.210 76.840 64.520 77.170 ;
        RECT 64.850 77.120 66.000 77.210 ;
        RECT 69.860 77.170 70.180 77.630 ;
        RECT 64.700 76.890 69.700 77.120 ;
        RECT 64.850 76.860 66.000 76.890 ;
        RECT 69.870 76.840 70.180 77.170 ;
        RECT 60.220 76.510 61.480 76.600 ;
        RECT 56.150 65.430 56.450 76.380 ;
        RECT 56.640 76.280 61.640 76.510 ;
        RECT 60.220 76.250 61.480 76.280 ;
        RECT 56.800 75.720 57.880 75.830 ;
        RECT 56.640 75.490 61.640 75.720 ;
        RECT 56.800 75.400 57.880 75.490 ;
        RECT 60.220 74.930 61.480 75.010 ;
        RECT 56.640 74.700 61.640 74.930 ;
        RECT 60.220 74.670 61.480 74.700 ;
        RECT 56.780 74.140 57.880 74.250 ;
        RECT 56.640 73.910 61.640 74.140 ;
        RECT 56.780 73.830 57.880 73.910 ;
        RECT 60.220 73.350 61.480 73.380 ;
        RECT 56.640 73.120 61.640 73.350 ;
        RECT 60.220 73.040 61.480 73.120 ;
        RECT 56.730 72.560 57.880 72.690 ;
        RECT 56.640 72.330 61.640 72.560 ;
        RECT 56.730 72.230 57.880 72.330 ;
        RECT 60.220 71.770 61.480 71.850 ;
        RECT 56.640 71.540 61.640 71.770 ;
        RECT 60.220 71.510 61.480 71.540 ;
        RECT 56.720 70.980 57.880 71.100 ;
        RECT 56.640 70.750 61.640 70.980 ;
        RECT 56.720 70.680 57.880 70.750 ;
        RECT 60.220 70.190 61.480 70.270 ;
        RECT 56.640 69.960 61.640 70.190 ;
        RECT 60.220 69.910 61.480 69.960 ;
        RECT 56.790 69.400 57.880 69.500 ;
        RECT 56.640 69.170 61.640 69.400 ;
        RECT 56.790 69.140 57.880 69.170 ;
        RECT 60.220 68.610 61.480 68.670 ;
        RECT 56.640 68.380 61.640 68.610 ;
        RECT 60.220 68.310 61.480 68.380 ;
        RECT 56.760 67.820 57.880 67.900 ;
        RECT 56.640 67.590 61.640 67.820 ;
        RECT 56.760 67.560 57.880 67.590 ;
        RECT 60.230 67.030 61.490 67.080 ;
        RECT 56.640 66.800 61.640 67.030 ;
        RECT 60.230 66.720 61.490 66.800 ;
        RECT 61.800 66.390 62.100 76.400 ;
        RECT 64.210 76.380 64.540 76.840 ;
        RECT 64.210 76.050 64.520 76.380 ;
        RECT 68.230 76.330 69.510 76.420 ;
        RECT 69.860 76.380 70.180 76.840 ;
        RECT 64.700 76.100 69.700 76.330 ;
        RECT 68.230 76.060 69.510 76.100 ;
        RECT 69.870 76.050 70.180 76.380 ;
        RECT 64.210 75.590 64.540 76.050 ;
        RECT 64.210 75.260 64.520 75.590 ;
        RECT 64.810 75.540 66.000 75.630 ;
        RECT 69.860 75.590 70.180 76.050 ;
        RECT 64.700 75.310 69.700 75.540 ;
        RECT 64.810 75.270 66.000 75.310 ;
        RECT 69.870 75.260 70.180 75.590 ;
        RECT 64.210 74.800 64.540 75.260 ;
        RECT 64.210 74.470 64.520 74.800 ;
        RECT 68.230 74.750 69.500 74.820 ;
        RECT 69.860 74.800 70.180 75.260 ;
        RECT 64.700 74.520 69.700 74.750 ;
        RECT 64.210 74.010 64.540 74.470 ;
        RECT 68.230 74.460 69.500 74.520 ;
        RECT 69.870 74.470 70.180 74.800 ;
        RECT 64.210 73.680 64.520 74.010 ;
        RECT 64.850 73.960 66.000 74.050 ;
        RECT 69.860 74.010 70.180 74.470 ;
        RECT 64.700 73.730 69.700 73.960 ;
        RECT 64.850 73.700 66.000 73.730 ;
        RECT 69.870 73.680 70.180 74.010 ;
        RECT 64.210 73.220 64.540 73.680 ;
        RECT 64.210 72.890 64.520 73.220 ;
        RECT 68.230 73.170 69.490 73.250 ;
        RECT 69.860 73.220 70.180 73.680 ;
        RECT 64.700 72.940 69.700 73.170 ;
        RECT 68.230 72.900 69.490 72.940 ;
        RECT 69.870 72.890 70.180 73.220 ;
        RECT 64.210 72.430 64.540 72.890 ;
        RECT 64.210 72.100 64.520 72.430 ;
        RECT 64.880 72.380 66.000 72.450 ;
        RECT 69.860 72.430 70.180 72.890 ;
        RECT 64.700 72.150 69.700 72.380 ;
        RECT 64.880 72.110 66.000 72.150 ;
        RECT 69.870 72.100 70.180 72.430 ;
        RECT 64.210 71.640 64.540 72.100 ;
        RECT 64.210 71.310 64.520 71.640 ;
        RECT 68.240 71.590 69.500 71.700 ;
        RECT 69.860 71.640 70.180 72.100 ;
        RECT 64.700 71.360 69.700 71.590 ;
        RECT 64.210 70.850 64.540 71.310 ;
        RECT 68.240 71.250 69.500 71.360 ;
        RECT 69.870 71.310 70.180 71.640 ;
        RECT 64.210 70.520 64.520 70.850 ;
        RECT 64.860 70.800 66.010 70.910 ;
        RECT 69.860 70.850 70.180 71.310 ;
        RECT 64.700 70.570 69.700 70.800 ;
        RECT 64.860 70.550 66.010 70.570 ;
        RECT 69.870 70.520 70.180 70.850 ;
        RECT 64.210 70.060 64.540 70.520 ;
        RECT 64.210 69.730 64.520 70.060 ;
        RECT 68.220 70.010 69.550 70.120 ;
        RECT 69.860 70.060 70.180 70.520 ;
        RECT 64.700 69.780 69.700 70.010 ;
        RECT 64.210 69.270 64.540 69.730 ;
        RECT 68.220 69.720 69.550 69.780 ;
        RECT 69.870 69.730 70.180 70.060 ;
        RECT 64.210 68.940 64.520 69.270 ;
        RECT 64.760 69.220 66.000 69.290 ;
        RECT 69.860 69.270 70.180 69.730 ;
        RECT 64.700 68.990 69.700 69.220 ;
        RECT 64.760 68.940 66.000 68.990 ;
        RECT 69.870 68.940 70.180 69.270 ;
        RECT 64.210 68.480 64.540 68.940 ;
        RECT 64.210 68.150 64.520 68.480 ;
        RECT 68.230 68.430 69.510 68.530 ;
        RECT 69.860 68.480 70.180 68.940 ;
        RECT 64.700 68.200 69.700 68.430 ;
        RECT 64.210 67.690 64.540 68.150 ;
        RECT 68.230 68.130 69.510 68.200 ;
        RECT 69.870 68.150 70.180 68.480 ;
        RECT 64.210 67.360 64.520 67.690 ;
        RECT 64.780 67.640 66.000 67.730 ;
        RECT 69.860 67.690 70.180 68.150 ;
        RECT 64.700 67.410 69.700 67.640 ;
        RECT 64.780 67.370 66.000 67.410 ;
        RECT 69.870 67.360 70.180 67.690 ;
        RECT 64.210 66.900 64.540 67.360 ;
        RECT 64.210 66.570 64.520 66.900 ;
        RECT 68.230 66.850 69.510 66.930 ;
        RECT 69.860 66.900 70.180 67.360 ;
        RECT 64.700 66.620 69.700 66.850 ;
        RECT 61.800 66.380 62.760 66.390 ;
        RECT 56.770 66.240 57.890 66.340 ;
        RECT 56.640 66.010 61.640 66.240 ;
        RECT 56.770 65.990 57.890 66.010 ;
        RECT 60.220 65.450 61.480 65.510 ;
        RECT 56.640 65.220 61.640 65.450 ;
        RECT 60.220 65.160 61.480 65.220 ;
        RECT 51.510 64.330 56.010 65.160 ;
        RECT 61.800 64.880 62.980 66.380 ;
        RECT 64.210 66.210 64.540 66.570 ;
        RECT 68.230 66.530 69.510 66.620 ;
        RECT 69.870 66.570 70.180 66.900 ;
        RECT 63.690 66.160 64.540 66.210 ;
        RECT 51.510 59.490 52.410 64.330 ;
        RECT 53.150 63.190 54.060 63.390 ;
        RECT 53.130 63.145 60.100 63.190 ;
        RECT 53.090 62.915 60.100 63.145 ;
        RECT 52.610 60.450 52.900 62.880 ;
        RECT 53.130 62.850 60.100 62.915 ;
        RECT 53.150 62.830 54.060 62.850 ;
        RECT 53.090 62.340 60.090 62.355 ;
        RECT 53.080 60.980 60.120 62.340 ;
        RECT 60.290 61.490 60.580 62.880 ;
        RECT 63.670 61.700 64.540 66.160 ;
        RECT 64.780 66.110 65.990 66.140 ;
        RECT 69.860 66.110 70.180 66.570 ;
        RECT 64.780 66.060 66.000 66.110 ;
        RECT 64.700 65.830 69.700 66.060 ;
        RECT 64.780 65.750 66.000 65.830 ;
        RECT 69.870 65.780 70.180 66.110 ;
        RECT 64.780 65.740 65.990 65.750 ;
        RECT 69.860 65.320 70.180 65.780 ;
        RECT 64.840 65.270 69.680 65.320 ;
        RECT 69.870 65.270 70.180 65.320 ;
        RECT 64.700 65.040 69.700 65.270 ;
        RECT 64.840 64.980 69.680 65.040 ;
        RECT 70.350 64.330 70.950 79.890 ;
        RECT 60.290 60.570 60.590 61.490 ;
        RECT 53.130 60.425 60.100 60.520 ;
        RECT 53.090 60.195 60.100 60.425 ;
        RECT 60.290 60.270 61.010 60.570 ;
        RECT 53.130 60.180 60.100 60.195 ;
        RECT 53.150 59.860 54.060 60.180 ;
        RECT 54.420 59.490 60.040 59.890 ;
        RECT 51.510 59.140 60.040 59.490 ;
        RECT 60.840 59.620 61.010 60.270 ;
        RECT 60.840 59.610 63.240 59.620 ;
        RECT 64.410 59.610 65.110 59.670 ;
        RECT 60.840 59.480 69.930 59.610 ;
        RECT 60.840 59.370 64.630 59.480 ;
        RECT 51.510 58.930 52.410 59.140 ;
        RECT 51.510 58.090 52.000 58.930 ;
        RECT 52.595 58.650 60.535 58.840 ;
        RECT 52.190 58.610 60.535 58.650 ;
        RECT 60.840 58.610 63.240 59.370 ;
        RECT 64.895 59.340 69.930 59.480 ;
        RECT 64.900 59.130 69.930 59.340 ;
        RECT 64.900 59.115 69.900 59.130 ;
        RECT 52.190 58.560 53.170 58.610 ;
        RECT 52.160 58.310 53.170 58.560 ;
        RECT 52.160 58.100 52.390 58.310 ;
        RECT 60.300 58.100 60.535 58.610 ;
        RECT 61.165 58.100 61.555 58.610 ;
        RECT 28.760 57.760 52.000 58.090 ;
        RECT 52.595 58.020 60.095 58.050 ;
        RECT 52.570 57.820 60.095 58.020 ;
        RECT 60.305 57.930 60.535 58.100 ;
        RECT 62.950 58.080 63.240 58.610 ;
        RECT 64.510 58.700 64.740 59.065 ;
        RECT 70.060 58.700 70.290 59.065 ;
        RECT 64.510 58.360 70.290 58.700 ;
        RECT 64.510 58.105 64.740 58.360 ;
        RECT 70.060 58.105 70.290 58.360 ;
        RECT 60.710 57.930 61.090 57.960 ;
        RECT 60.305 57.910 61.090 57.930 ;
        RECT 61.755 57.910 62.755 58.050 ;
        RECT 64.900 58.030 69.900 58.055 ;
        RECT 70.470 58.030 70.950 64.330 ;
        RECT 60.305 57.820 62.755 57.910 ;
        RECT 64.880 57.880 69.900 58.030 ;
        RECT 70.450 57.880 70.950 58.030 ;
        RECT 52.570 57.760 53.350 57.820 ;
        RECT 28.760 57.100 53.350 57.760 ;
        RECT 60.305 57.700 62.730 57.820 ;
        RECT 64.880 57.190 70.950 57.880 ;
        RECT 27.350 53.260 28.050 56.590 ;
        RECT 27.360 52.630 28.050 53.260 ;
        RECT 15.000 45.050 17.130 47.200 ;
        RECT 18.370 45.050 21.240 47.200 ;
        RECT 22.370 45.050 24.500 47.200 ;
        RECT 25.630 45.060 28.250 47.200 ;
        RECT 26.960 44.090 28.250 45.060 ;
        RECT 26.950 43.220 28.250 44.090 ;
        RECT 26.950 40.800 28.190 43.220 ;
        RECT 28.760 38.880 29.340 57.100 ;
        RECT 37.240 56.300 38.470 57.100 ;
        RECT 34.260 54.450 35.510 54.470 ;
        RECT 30.050 54.430 35.510 54.450 ;
        RECT 29.560 54.220 35.510 54.430 ;
        RECT 29.560 54.150 30.280 54.220 ;
        RECT 29.530 54.060 30.280 54.150 ;
        RECT 34.260 54.200 35.510 54.220 ;
        RECT 34.260 54.120 35.560 54.200 ;
        RECT 29.530 45.500 29.860 54.060 ;
        RECT 34.090 53.660 35.090 53.740 ;
        RECT 30.050 53.430 35.090 53.660 ;
        RECT 34.090 53.280 35.090 53.430 ;
        RECT 34.090 49.950 35.060 50.340 ;
        RECT 30.050 49.720 35.060 49.950 ;
        RECT 34.090 49.620 35.060 49.720 ;
        RECT 34.090 49.160 35.030 49.210 ;
        RECT 30.050 48.930 35.050 49.160 ;
        RECT 34.090 48.740 35.030 48.930 ;
        RECT 29.530 45.450 30.370 45.500 ;
        RECT 35.230 45.460 35.560 54.120 ;
        RECT 34.270 45.450 35.560 45.460 ;
        RECT 29.530 45.240 35.560 45.450 ;
        RECT 29.530 44.630 29.860 45.240 ;
        RECT 30.050 45.220 35.560 45.240 ;
        RECT 34.270 45.170 35.560 45.220 ;
        RECT 34.070 44.660 35.020 44.790 ;
        RECT 35.230 44.680 35.560 45.170 ;
        RECT 30.050 44.430 35.050 44.660 ;
        RECT 34.070 44.350 35.020 44.430 ;
        RECT 35.750 44.100 36.140 54.560 ;
        RECT 36.680 44.150 37.320 54.640 ;
        RECT 37.800 43.970 38.190 56.300 ;
        RECT 63.220 56.240 64.150 56.280 ;
        RECT 63.220 56.010 68.230 56.240 ;
        RECT 63.220 55.960 64.150 56.010 ;
        RECT 50.080 54.930 51.810 55.270 ;
        RECT 39.020 54.450 39.680 54.670 ;
        RECT 42.030 54.450 43.830 54.890 ;
        RECT 47.770 54.700 52.770 54.930 ;
        RECT 39.020 54.220 44.050 54.450 ;
        RECT 39.020 54.200 39.680 54.220 ;
        RECT 38.510 53.710 38.845 54.170 ;
        RECT 42.030 54.070 43.830 54.220 ;
        RECT 38.510 50.180 38.840 53.710 ;
        RECT 39.080 53.660 39.900 53.760 ;
        RECT 39.050 53.430 44.050 53.660 ;
        RECT 39.080 53.260 39.900 53.430 ;
        RECT 38.510 49.950 39.830 50.180 ;
        RECT 44.210 50.000 44.540 54.180 ;
        RECT 47.380 53.690 47.610 54.650 ;
        RECT 52.930 53.690 54.040 55.090 ;
        RECT 57.260 54.930 58.780 55.120 ;
        RECT 54.770 54.700 59.770 54.930 ;
        RECT 52.960 53.650 54.040 53.690 ;
        RECT 47.770 53.610 52.770 53.640 ;
        RECT 47.740 52.720 52.790 53.610 ;
        RECT 47.770 52.700 52.770 52.720 ;
        RECT 53.700 52.700 54.040 53.650 ;
        RECT 54.270 53.630 54.620 54.670 ;
        RECT 57.260 54.600 58.780 54.700 ;
        RECT 59.930 53.690 60.160 54.650 ;
        RECT 54.770 53.610 59.770 53.640 ;
        RECT 54.770 53.410 59.800 53.610 ;
        RECT 54.980 52.930 59.800 53.410 ;
        RECT 54.770 52.720 59.800 52.930 ;
        RECT 54.770 52.700 59.770 52.720 ;
        RECT 43.880 49.950 44.540 50.000 ;
        RECT 38.510 49.830 44.540 49.950 ;
        RECT 38.510 49.670 38.840 49.830 ;
        RECT 39.050 49.750 44.540 49.830 ;
        RECT 39.050 49.720 44.050 49.750 ;
        RECT 38.510 49.210 38.845 49.670 ;
        RECT 38.510 45.170 38.840 49.210 ;
        RECT 39.140 49.160 39.860 49.380 ;
        RECT 39.050 48.930 44.050 49.160 ;
        RECT 39.140 48.810 39.860 48.930 ;
        RECT 44.210 48.750 44.540 49.750 ;
        RECT 46.720 52.650 47.580 52.680 ;
        RECT 46.720 51.690 47.610 52.650 ;
        RECT 46.720 51.670 47.580 51.690 ;
        RECT 46.720 51.090 47.040 51.670 ;
        RECT 47.760 51.640 49.650 51.910 ;
        RECT 52.930 51.690 53.160 52.650 ;
        RECT 53.700 51.650 54.610 52.700 ;
        RECT 47.760 51.410 52.770 51.640 ;
        RECT 47.760 51.290 49.650 51.410 ;
        RECT 53.700 51.120 54.040 51.650 ;
        RECT 55.190 51.640 56.710 51.800 ;
        RECT 59.930 51.690 60.160 52.650 ;
        RECT 54.770 51.410 59.770 51.640 ;
        RECT 55.190 51.280 56.710 51.410 ;
        RECT 46.720 49.460 47.050 51.090 ;
        RECT 44.210 47.860 44.870 48.750 ;
        RECT 39.010 45.450 39.630 45.660 ;
        RECT 39.010 45.220 44.050 45.450 ;
        RECT 38.510 44.710 38.845 45.170 ;
        RECT 39.010 45.160 39.630 45.220 ;
        RECT 38.510 44.650 38.840 44.710 ;
        RECT 39.190 44.660 39.910 44.800 ;
        RECT 44.210 44.660 44.540 47.860 ;
        RECT 46.720 47.010 47.040 49.460 ;
        RECT 50.080 48.930 51.810 49.260 ;
        RECT 47.770 48.700 52.770 48.930 ;
        RECT 53.710 48.670 54.030 51.120 ;
        RECT 54.220 49.600 54.610 50.630 ;
        RECT 52.970 48.650 54.030 48.670 ;
        RECT 47.380 47.690 47.610 48.650 ;
        RECT 52.930 47.690 54.030 48.650 ;
        RECT 52.970 47.670 54.030 47.690 ;
        RECT 47.770 47.610 52.770 47.640 ;
        RECT 45.930 46.670 47.040 47.010 ;
        RECT 47.750 46.720 52.800 47.610 ;
        RECT 47.770 46.700 52.770 46.720 ;
        RECT 53.710 46.690 54.030 47.670 ;
        RECT 54.330 47.660 54.610 49.600 ;
        RECT 62.790 50.550 63.070 55.960 ;
        RECT 67.230 54.950 68.180 55.040 ;
        RECT 68.380 55.000 69.530 55.970 ;
        RECT 63.230 54.720 68.240 54.950 ;
        RECT 67.230 54.640 68.180 54.720 ;
        RECT 68.420 54.670 68.830 55.000 ;
        RECT 63.230 53.660 64.150 53.720 ;
        RECT 68.390 53.710 68.830 54.670 ;
        RECT 63.230 53.650 68.230 53.660 ;
        RECT 63.230 53.420 68.240 53.650 ;
        RECT 63.230 53.350 64.150 53.420 ;
        RECT 68.420 53.380 68.830 53.710 ;
        RECT 68.390 52.420 68.830 53.380 ;
        RECT 67.230 52.370 68.180 52.420 ;
        RECT 63.230 52.360 68.230 52.370 ;
        RECT 63.230 52.140 68.240 52.360 ;
        RECT 63.280 52.130 68.240 52.140 ;
        RECT 67.230 52.040 68.180 52.130 ;
        RECT 68.420 52.090 68.830 52.420 ;
        RECT 63.230 51.080 64.160 51.170 ;
        RECT 68.390 51.130 68.830 52.090 ;
        RECT 63.230 50.850 68.240 51.080 ;
        RECT 63.230 50.790 64.160 50.850 ;
        RECT 68.420 50.800 68.830 51.130 ;
        RECT 68.390 50.550 68.830 50.800 ;
        RECT 62.790 50.100 63.160 50.550 ;
        RECT 68.340 50.100 68.830 50.550 ;
        RECT 57.290 48.930 58.810 49.130 ;
        RECT 54.770 48.700 59.770 48.930 ;
        RECT 57.290 48.610 58.810 48.700 ;
        RECT 59.930 47.690 60.160 48.650 ;
        RECT 54.770 47.620 59.770 47.640 ;
        RECT 54.750 47.430 59.790 47.620 ;
        RECT 54.740 46.730 59.790 47.430 ;
        RECT 54.770 46.700 59.770 46.730 ;
        RECT 53.710 46.670 54.580 46.690 ;
        RECT 45.930 46.650 47.590 46.670 ;
        RECT 53.710 46.650 54.600 46.670 ;
        RECT 45.930 45.690 47.610 46.650 ;
        RECT 52.930 45.690 53.160 46.650 ;
        RECT 53.710 45.690 54.610 46.650 ;
        RECT 45.930 45.660 47.520 45.690 ;
        RECT 47.800 45.640 49.520 45.690 ;
        RECT 53.720 45.680 54.580 45.690 ;
        RECT 55.200 45.640 56.720 45.830 ;
        RECT 59.930 45.690 60.160 46.650 ;
        RECT 47.770 45.410 52.770 45.640 ;
        RECT 54.770 45.410 59.770 45.640 ;
        RECT 47.800 45.270 49.520 45.410 ;
        RECT 55.200 45.310 56.720 45.410 ;
        RECT 61.040 45.110 61.620 46.760 ;
        RECT 62.790 45.950 63.070 50.100 ;
        RECT 67.230 49.790 68.170 49.870 ;
        RECT 68.390 49.840 68.830 50.100 ;
        RECT 63.230 49.780 68.230 49.790 ;
        RECT 63.230 49.560 68.240 49.780 ;
        RECT 63.280 49.550 68.240 49.560 ;
        RECT 67.230 49.480 68.170 49.550 ;
        RECT 68.420 49.510 68.830 49.840 ;
        RECT 63.230 48.500 64.150 48.620 ;
        RECT 68.390 48.550 68.830 49.510 ;
        RECT 63.230 48.270 68.240 48.500 ;
        RECT 63.230 48.200 64.150 48.270 ;
        RECT 68.420 48.220 68.830 48.550 ;
        RECT 67.150 47.210 68.250 47.450 ;
        RECT 68.390 47.260 68.830 48.220 ;
        RECT 70.340 47.440 70.950 57.190 ;
        RECT 63.230 46.980 68.250 47.210 ;
        RECT 67.150 46.780 68.250 46.980 ;
        RECT 68.420 46.930 68.830 47.260 ;
        RECT 63.230 45.920 64.150 46.040 ;
        RECT 68.390 45.970 68.830 46.930 ;
        RECT 70.170 46.780 70.950 47.440 ;
        RECT 68.420 45.950 68.830 45.970 ;
        RECT 63.230 45.690 68.250 45.920 ;
        RECT 63.230 45.620 64.150 45.690 ;
        RECT 70.340 45.110 70.950 46.780 ;
        RECT 39.050 44.430 44.050 44.660 ;
        RECT 39.190 44.230 39.910 44.430 ;
        RECT 61.040 44.250 70.950 45.110 ;
        RECT 37.630 43.490 38.310 43.970 ;
        RECT 70.340 43.680 70.950 44.250 ;
        RECT 71.770 112.980 72.340 124.610 ;
        RECT 98.590 119.310 99.010 134.790 ;
        RECT 103.220 134.730 104.480 134.790 ;
        RECT 99.150 123.570 99.450 134.520 ;
        RECT 99.640 134.500 104.640 134.730 ;
        RECT 103.220 134.440 104.480 134.500 ;
        RECT 99.770 133.940 100.890 133.960 ;
        RECT 99.640 133.710 104.640 133.940 ;
        RECT 99.770 133.610 100.890 133.710 ;
        RECT 104.800 133.570 105.980 135.070 ;
        RECT 104.800 133.560 105.760 133.570 ;
        RECT 103.230 133.150 104.490 133.230 ;
        RECT 99.640 132.920 104.640 133.150 ;
        RECT 103.230 132.870 104.490 132.920 ;
        RECT 99.760 132.360 100.880 132.390 ;
        RECT 99.640 132.130 104.640 132.360 ;
        RECT 99.760 132.050 100.880 132.130 ;
        RECT 103.220 131.570 104.480 131.640 ;
        RECT 99.640 131.340 104.640 131.570 ;
        RECT 103.220 131.280 104.480 131.340 ;
        RECT 99.790 130.780 100.880 130.810 ;
        RECT 99.640 130.550 104.640 130.780 ;
        RECT 99.790 130.450 100.880 130.550 ;
        RECT 103.220 129.990 104.480 130.040 ;
        RECT 99.640 129.760 104.640 129.990 ;
        RECT 103.220 129.680 104.480 129.760 ;
        RECT 99.720 129.200 100.880 129.270 ;
        RECT 99.640 128.970 104.640 129.200 ;
        RECT 99.720 128.850 100.880 128.970 ;
        RECT 103.220 128.410 104.480 128.440 ;
        RECT 99.640 128.180 104.640 128.410 ;
        RECT 103.220 128.100 104.480 128.180 ;
        RECT 99.730 127.620 100.880 127.720 ;
        RECT 99.640 127.390 104.640 127.620 ;
        RECT 99.730 127.260 100.880 127.390 ;
        RECT 103.220 126.830 104.480 126.910 ;
        RECT 99.640 126.600 104.640 126.830 ;
        RECT 103.220 126.570 104.480 126.600 ;
        RECT 99.780 126.040 100.880 126.120 ;
        RECT 99.640 125.810 104.640 126.040 ;
        RECT 99.780 125.700 100.880 125.810 ;
        RECT 103.220 125.250 104.480 125.280 ;
        RECT 99.640 125.020 104.640 125.250 ;
        RECT 103.220 124.940 104.480 125.020 ;
        RECT 99.800 124.460 100.880 124.550 ;
        RECT 99.640 124.230 104.640 124.460 ;
        RECT 99.800 124.120 100.880 124.230 ;
        RECT 103.220 123.670 104.480 123.700 ;
        RECT 99.640 123.440 104.640 123.670 ;
        RECT 104.800 123.550 105.100 133.560 ;
        RECT 106.670 133.380 107.540 138.250 ;
        RECT 113.470 138.170 115.085 140.010 ;
        RECT 115.465 139.850 115.985 141.170 ;
        RECT 116.255 140.010 116.485 141.010 ;
        RECT 116.735 139.850 117.255 141.170 ;
        RECT 117.645 141.010 119.385 141.580 ;
        RECT 117.545 140.010 119.385 141.010 ;
        RECT 115.245 139.620 116.205 139.850 ;
        RECT 116.535 139.620 117.495 139.850 ;
        RECT 116.595 139.340 117.435 139.620 ;
        RECT 117.645 139.580 119.385 140.010 ;
        RECT 117.645 139.560 119.365 139.580 ;
        RECT 119.665 139.375 120.185 141.785 ;
        RECT 120.445 139.580 120.675 141.580 ;
        RECT 120.995 139.375 121.515 141.785 ;
        RECT 121.875 141.580 123.630 143.640 ;
        RECT 121.735 140.185 123.630 141.580 ;
        RECT 121.735 139.580 123.625 140.185 ;
        RECT 126.820 139.965 127.520 144.045 ;
        RECT 130.395 143.875 130.955 145.015 ;
        RECT 130.410 140.195 130.955 143.875 ;
        RECT 119.435 139.340 120.395 139.375 ;
        RECT 116.595 139.170 120.395 139.340 ;
        RECT 117.985 138.750 118.675 139.170 ;
        RECT 119.435 139.145 120.395 139.170 ;
        RECT 120.725 139.145 121.685 139.375 ;
        RECT 121.875 138.995 123.625 139.580 ;
        RECT 123.815 139.200 124.775 139.430 ;
        RECT 125.105 139.405 126.065 139.430 ;
        RECT 126.825 139.405 127.515 139.965 ;
        RECT 125.105 139.235 128.905 139.405 ;
        RECT 125.105 139.200 126.065 139.235 ;
        RECT 121.875 138.770 123.765 138.995 ;
        RECT 117.985 138.390 118.680 138.750 ;
        RECT 113.470 136.110 115.080 138.170 ;
        RECT 113.470 135.620 115.450 136.110 ;
        RECT 107.840 134.910 112.680 134.970 ;
        RECT 107.700 134.680 112.700 134.910 ;
        RECT 107.840 134.630 112.680 134.680 ;
        RECT 112.870 134.630 113.180 134.680 ;
        RECT 107.780 134.200 108.990 134.210 ;
        RECT 107.780 134.120 109.000 134.200 ;
        RECT 112.860 134.170 113.180 134.630 ;
        RECT 107.700 133.890 112.700 134.120 ;
        RECT 107.780 133.840 109.000 133.890 ;
        RECT 112.870 133.840 113.180 134.170 ;
        RECT 107.780 133.810 108.990 133.840 ;
        RECT 106.670 133.050 107.520 133.380 ;
        RECT 111.230 133.330 112.510 133.420 ;
        RECT 112.860 133.380 113.180 133.840 ;
        RECT 107.700 133.100 112.700 133.330 ;
        RECT 106.670 132.590 107.540 133.050 ;
        RECT 111.230 133.020 112.510 133.100 ;
        RECT 112.870 133.050 113.180 133.380 ;
        RECT 112.860 132.590 113.180 133.050 ;
        RECT 106.670 132.260 107.520 132.590 ;
        RECT 107.780 132.540 109.000 132.580 ;
        RECT 107.700 132.310 112.700 132.540 ;
        RECT 106.670 131.800 107.540 132.260 ;
        RECT 107.780 132.220 109.000 132.310 ;
        RECT 112.870 132.260 113.180 132.590 ;
        RECT 106.670 131.470 107.520 131.800 ;
        RECT 111.230 131.750 112.510 131.820 ;
        RECT 112.860 131.800 113.180 132.260 ;
        RECT 107.700 131.520 112.700 131.750 ;
        RECT 106.670 131.010 107.540 131.470 ;
        RECT 111.230 131.420 112.510 131.520 ;
        RECT 112.870 131.470 113.180 131.800 ;
        RECT 112.860 131.010 113.180 131.470 ;
        RECT 106.670 130.680 107.520 131.010 ;
        RECT 107.760 130.960 109.000 131.010 ;
        RECT 107.700 130.730 112.700 130.960 ;
        RECT 106.670 130.220 107.540 130.680 ;
        RECT 107.760 130.660 109.000 130.730 ;
        RECT 112.870 130.680 113.180 131.010 ;
        RECT 106.670 129.890 107.520 130.220 ;
        RECT 111.220 130.170 112.550 130.230 ;
        RECT 112.860 130.220 113.180 130.680 ;
        RECT 107.700 129.940 112.700 130.170 ;
        RECT 106.670 129.430 107.540 129.890 ;
        RECT 111.220 129.830 112.550 129.940 ;
        RECT 112.870 129.890 113.180 130.220 ;
        RECT 112.860 129.430 113.180 129.890 ;
        RECT 106.670 129.100 107.520 129.430 ;
        RECT 107.860 129.380 109.010 129.400 ;
        RECT 107.700 129.150 112.700 129.380 ;
        RECT 106.670 128.640 107.540 129.100 ;
        RECT 107.860 129.040 109.010 129.150 ;
        RECT 112.870 129.100 113.180 129.430 ;
        RECT 106.670 128.310 107.520 128.640 ;
        RECT 111.240 128.590 112.500 128.700 ;
        RECT 112.860 128.640 113.180 129.100 ;
        RECT 107.700 128.360 112.700 128.590 ;
        RECT 106.670 127.850 107.540 128.310 ;
        RECT 111.240 128.250 112.500 128.360 ;
        RECT 112.870 128.310 113.180 128.640 ;
        RECT 112.860 127.850 113.180 128.310 ;
        RECT 106.670 127.520 107.520 127.850 ;
        RECT 107.880 127.800 109.000 127.840 ;
        RECT 107.700 127.570 112.700 127.800 ;
        RECT 106.670 127.060 107.540 127.520 ;
        RECT 107.880 127.500 109.000 127.570 ;
        RECT 112.870 127.520 113.180 127.850 ;
        RECT 112.860 127.060 113.180 127.520 ;
        RECT 106.670 126.730 107.520 127.060 ;
        RECT 111.230 127.010 112.490 127.050 ;
        RECT 107.700 126.780 112.700 127.010 ;
        RECT 106.670 126.270 107.540 126.730 ;
        RECT 111.230 126.700 112.490 126.780 ;
        RECT 112.870 126.730 113.180 127.060 ;
        RECT 112.860 126.270 113.180 126.730 ;
        RECT 106.670 125.940 107.520 126.270 ;
        RECT 107.850 126.220 109.000 126.250 ;
        RECT 107.700 125.990 112.700 126.220 ;
        RECT 106.670 125.480 107.540 125.940 ;
        RECT 107.850 125.900 109.000 125.990 ;
        RECT 112.870 125.940 113.180 126.270 ;
        RECT 106.670 125.150 107.520 125.480 ;
        RECT 111.230 125.430 112.500 125.490 ;
        RECT 112.860 125.480 113.180 125.940 ;
        RECT 107.700 125.200 112.700 125.430 ;
        RECT 106.670 124.690 107.540 125.150 ;
        RECT 111.230 125.130 112.500 125.200 ;
        RECT 112.870 125.150 113.180 125.480 ;
        RECT 112.860 124.690 113.180 125.150 ;
        RECT 106.670 124.360 107.520 124.690 ;
        RECT 107.810 124.640 109.000 124.680 ;
        RECT 107.700 124.410 112.700 124.640 ;
        RECT 106.670 123.900 107.540 124.360 ;
        RECT 107.810 124.320 109.000 124.410 ;
        RECT 112.870 124.360 113.180 124.690 ;
        RECT 112.860 123.900 113.180 124.360 ;
        RECT 106.670 123.570 107.520 123.900 ;
        RECT 111.230 123.850 112.510 123.890 ;
        RECT 107.700 123.620 112.700 123.850 ;
        RECT 103.220 123.350 104.480 123.440 ;
        RECT 106.670 123.110 107.540 123.570 ;
        RECT 111.230 123.530 112.510 123.620 ;
        RECT 112.870 123.570 113.180 123.900 ;
        RECT 112.860 123.110 113.180 123.570 ;
        RECT 113.350 134.210 115.450 135.620 ;
        RECT 117.990 134.510 118.680 138.390 ;
        RECT 121.870 136.995 123.765 138.770 ;
        RECT 121.870 136.305 123.625 136.995 ;
        RECT 123.985 136.790 124.505 139.200 ;
        RECT 124.825 136.995 125.055 138.995 ;
        RECT 125.315 136.790 125.835 139.200 ;
        RECT 126.135 138.995 127.855 139.015 ;
        RECT 126.115 138.565 127.855 138.995 ;
        RECT 128.065 138.955 128.905 139.235 ;
        RECT 128.005 138.725 128.965 138.955 ;
        RECT 129.295 138.725 130.255 138.955 ;
        RECT 126.115 137.565 127.955 138.565 ;
        RECT 126.115 136.995 127.855 137.565 ;
        RECT 128.245 137.405 128.765 138.725 ;
        RECT 129.015 137.565 129.245 138.565 ;
        RECT 129.515 137.405 130.035 138.725 ;
        RECT 130.415 138.565 130.955 140.195 ;
        RECT 130.305 137.565 130.955 138.565 ;
        RECT 128.005 137.175 128.965 137.405 ;
        RECT 129.295 137.175 130.255 137.405 ;
        RECT 130.415 137.035 130.955 137.565 ;
        RECT 126.135 136.975 127.855 136.995 ;
        RECT 123.815 136.560 124.775 136.790 ;
        RECT 125.105 136.560 126.065 136.790 ;
        RECT 126.825 136.565 127.515 136.975 ;
        RECT 130.405 136.915 130.955 137.035 ;
        RECT 113.350 133.540 115.105 134.210 ;
        RECT 117.985 133.890 118.685 134.510 ;
        RECT 121.870 134.260 123.630 136.305 ;
        RECT 126.815 135.945 127.515 136.565 ;
        RECT 130.395 136.120 130.955 136.915 ;
        RECT 113.350 133.420 115.095 133.540 ;
        RECT 117.985 133.480 118.675 133.890 ;
        RECT 119.435 133.665 120.395 133.895 ;
        RECT 120.725 133.665 121.685 133.895 ;
        RECT 117.645 133.460 119.365 133.480 ;
        RECT 113.350 132.890 115.085 133.420 ;
        RECT 115.245 133.050 116.205 133.280 ;
        RECT 116.535 133.050 117.495 133.280 ;
        RECT 113.350 131.890 115.195 132.890 ;
        RECT 113.350 130.620 115.085 131.890 ;
        RECT 115.465 131.730 115.985 133.050 ;
        RECT 116.255 131.890 116.485 132.890 ;
        RECT 116.735 131.730 117.255 133.050 ;
        RECT 117.645 132.890 119.385 133.460 ;
        RECT 117.545 131.890 119.385 132.890 ;
        RECT 115.245 131.500 116.205 131.730 ;
        RECT 116.535 131.500 117.495 131.730 ;
        RECT 116.595 131.220 117.435 131.500 ;
        RECT 117.645 131.460 119.385 131.890 ;
        RECT 117.645 131.440 119.365 131.460 ;
        RECT 119.665 131.255 120.185 133.665 ;
        RECT 120.445 131.460 120.675 133.460 ;
        RECT 120.995 131.255 121.515 133.665 ;
        RECT 121.875 133.460 123.630 134.260 ;
        RECT 121.735 131.715 123.630 133.460 ;
        RECT 126.820 132.085 127.510 135.945 ;
        RECT 129.770 134.200 130.960 136.120 ;
        RECT 130.420 132.305 130.960 134.200 ;
        RECT 126.820 131.825 127.515 132.085 ;
        RECT 121.735 131.460 123.625 131.715 ;
        RECT 119.435 131.220 120.395 131.255 ;
        RECT 116.595 131.050 120.395 131.220 ;
        RECT 113.350 129.480 115.105 130.620 ;
        RECT 117.985 130.450 118.675 131.050 ;
        RECT 119.435 131.025 120.395 131.050 ;
        RECT 120.725 131.025 121.685 131.255 ;
        RECT 121.875 130.895 123.625 131.460 ;
        RECT 123.815 131.100 124.775 131.330 ;
        RECT 125.105 131.305 126.065 131.330 ;
        RECT 126.825 131.305 127.515 131.825 ;
        RECT 130.415 132.075 130.960 132.305 ;
        RECT 125.105 131.135 128.905 131.305 ;
        RECT 125.105 131.100 126.065 131.135 ;
        RECT 117.985 129.830 118.685 130.450 ;
        RECT 113.350 129.360 115.095 129.480 ;
        RECT 117.985 129.420 118.675 129.830 ;
        RECT 119.435 129.605 120.395 129.835 ;
        RECT 120.725 129.605 121.685 129.835 ;
        RECT 117.645 129.400 119.365 129.420 ;
        RECT 113.350 128.830 115.085 129.360 ;
        RECT 115.245 128.990 116.205 129.220 ;
        RECT 116.535 128.990 117.495 129.220 ;
        RECT 113.350 127.830 115.195 128.830 ;
        RECT 113.350 126.560 115.085 127.830 ;
        RECT 115.465 127.670 115.985 128.990 ;
        RECT 116.255 127.830 116.485 128.830 ;
        RECT 116.735 127.670 117.255 128.990 ;
        RECT 117.645 128.830 119.385 129.400 ;
        RECT 117.545 127.830 119.385 128.830 ;
        RECT 115.245 127.440 116.205 127.670 ;
        RECT 116.535 127.440 117.495 127.670 ;
        RECT 116.595 127.160 117.435 127.440 ;
        RECT 117.645 127.400 119.385 127.830 ;
        RECT 117.645 127.380 119.365 127.400 ;
        RECT 119.665 127.195 120.185 129.605 ;
        RECT 120.445 127.400 120.675 129.400 ;
        RECT 120.995 127.195 121.515 129.605 ;
        RECT 121.875 129.400 123.765 130.895 ;
        RECT 121.735 128.895 123.765 129.400 ;
        RECT 121.735 128.065 123.625 128.895 ;
        RECT 123.985 128.690 124.505 131.100 ;
        RECT 124.825 128.895 125.055 130.895 ;
        RECT 125.315 128.690 125.835 131.100 ;
        RECT 126.135 130.895 127.855 130.915 ;
        RECT 126.115 130.465 127.855 130.895 ;
        RECT 128.065 130.855 128.905 131.135 ;
        RECT 128.005 130.625 128.965 130.855 ;
        RECT 129.295 130.625 130.255 130.855 ;
        RECT 126.115 129.465 127.955 130.465 ;
        RECT 126.115 128.895 127.855 129.465 ;
        RECT 128.245 129.305 128.765 130.625 ;
        RECT 129.015 129.465 129.245 130.465 ;
        RECT 129.515 129.305 130.035 130.625 ;
        RECT 130.415 130.465 130.955 132.075 ;
        RECT 130.305 129.465 130.955 130.465 ;
        RECT 128.005 129.075 128.965 129.305 ;
        RECT 129.295 129.075 130.255 129.305 ;
        RECT 130.415 128.935 130.955 129.465 ;
        RECT 126.135 128.875 127.855 128.895 ;
        RECT 123.815 128.460 124.775 128.690 ;
        RECT 125.105 128.460 126.065 128.690 ;
        RECT 126.825 128.465 127.515 128.875 ;
        RECT 130.405 128.815 130.955 128.935 ;
        RECT 121.735 127.885 123.620 128.065 ;
        RECT 121.735 127.675 123.625 127.885 ;
        RECT 126.815 127.845 127.515 128.465 ;
        RECT 121.735 127.400 123.620 127.675 ;
        RECT 119.435 127.160 120.395 127.195 ;
        RECT 116.595 126.990 120.395 127.160 ;
        RECT 113.350 125.420 115.105 126.560 ;
        RECT 117.985 126.390 118.675 126.990 ;
        RECT 119.435 126.965 120.395 126.990 ;
        RECT 120.725 126.965 121.685 127.195 ;
        RECT 117.985 125.770 118.685 126.390 ;
        RECT 113.350 125.300 115.095 125.420 ;
        RECT 117.985 125.360 118.675 125.770 ;
        RECT 119.435 125.545 120.395 125.775 ;
        RECT 120.725 125.545 121.685 125.775 ;
        RECT 117.645 125.340 119.365 125.360 ;
        RECT 113.350 124.770 115.085 125.300 ;
        RECT 115.245 124.930 116.205 125.160 ;
        RECT 116.535 124.930 117.495 125.160 ;
        RECT 113.350 123.770 115.195 124.770 ;
        RECT 113.350 123.230 115.085 123.770 ;
        RECT 115.465 123.610 115.985 124.930 ;
        RECT 116.255 123.770 116.485 124.770 ;
        RECT 116.735 123.610 117.255 124.930 ;
        RECT 117.645 124.770 119.385 125.340 ;
        RECT 117.545 123.770 119.385 124.770 ;
        RECT 115.245 123.380 116.205 123.610 ;
        RECT 116.535 123.380 117.495 123.610 ;
        RECT 106.670 122.780 107.520 123.110 ;
        RECT 107.850 123.060 109.000 123.090 ;
        RECT 107.700 122.830 112.700 123.060 ;
        RECT 106.670 122.320 107.540 122.780 ;
        RECT 107.850 122.740 109.000 122.830 ;
        RECT 112.870 122.780 113.180 123.110 ;
        RECT 112.860 122.320 113.180 122.780 ;
        RECT 106.670 121.990 107.520 122.320 ;
        RECT 111.230 122.270 112.500 122.300 ;
        RECT 107.700 122.040 112.700 122.270 ;
        RECT 106.670 121.530 107.540 121.990 ;
        RECT 111.230 121.910 112.500 122.040 ;
        RECT 112.870 121.990 113.180 122.320 ;
        RECT 107.810 121.530 108.990 121.580 ;
        RECT 112.860 121.530 113.180 121.990 ;
        RECT 106.670 121.200 107.520 121.530 ;
        RECT 107.810 121.480 109.000 121.530 ;
        RECT 107.700 121.250 112.700 121.480 ;
        RECT 106.670 120.740 107.540 121.200 ;
        RECT 107.810 121.190 109.000 121.250 ;
        RECT 112.870 121.200 113.180 121.530 ;
        RECT 107.810 121.160 108.990 121.190 ;
        RECT 112.860 120.740 113.180 121.200 ;
        RECT 106.670 120.410 107.520 120.740 ;
        RECT 111.220 120.690 112.500 120.720 ;
        RECT 107.700 120.460 112.700 120.690 ;
        RECT 106.670 119.950 107.540 120.410 ;
        RECT 111.220 120.360 112.500 120.460 ;
        RECT 112.870 120.410 113.180 120.740 ;
        RECT 112.860 119.950 113.180 120.410 ;
        RECT 106.670 119.850 107.520 119.950 ;
        RECT 107.810 119.900 109.010 119.930 ;
        RECT 98.150 117.830 99.020 119.310 ;
        RECT 71.770 99.750 72.600 112.980 ;
        RECT 98.590 102.520 99.010 117.830 ;
        RECT 106.670 117.460 107.420 119.850 ;
        RECT 107.700 119.670 112.700 119.900 ;
        RECT 112.870 119.840 113.180 119.950 ;
        RECT 113.340 122.500 115.085 123.230 ;
        RECT 116.595 123.100 117.435 123.380 ;
        RECT 117.645 123.340 119.385 123.770 ;
        RECT 117.645 123.320 119.365 123.340 ;
        RECT 119.665 123.135 120.185 125.545 ;
        RECT 120.445 123.340 120.675 125.340 ;
        RECT 120.995 123.135 121.515 125.545 ;
        RECT 121.875 125.340 123.620 127.400 ;
        RECT 121.735 124.205 123.620 125.340 ;
        RECT 121.735 123.340 123.625 124.205 ;
        RECT 126.820 123.985 127.510 127.845 ;
        RECT 130.395 127.675 130.955 128.815 ;
        RECT 130.410 124.075 130.955 127.675 ;
        RECT 126.820 123.765 127.515 123.985 ;
        RECT 119.435 123.100 120.395 123.135 ;
        RECT 116.595 122.930 120.395 123.100 ;
        RECT 113.340 121.360 115.105 122.500 ;
        RECT 117.985 122.330 118.675 122.930 ;
        RECT 119.435 122.905 120.395 122.930 ;
        RECT 120.725 122.905 121.685 123.135 ;
        RECT 121.875 122.795 123.625 123.340 ;
        RECT 123.815 123.000 124.775 123.230 ;
        RECT 125.105 123.205 126.065 123.230 ;
        RECT 126.825 123.205 127.515 123.765 ;
        RECT 125.105 123.035 128.905 123.205 ;
        RECT 125.105 123.000 126.065 123.035 ;
        RECT 117.985 121.710 118.685 122.330 ;
        RECT 113.340 121.240 115.095 121.360 ;
        RECT 117.985 121.300 118.675 121.710 ;
        RECT 119.435 121.485 120.395 121.715 ;
        RECT 120.725 121.485 121.685 121.715 ;
        RECT 117.645 121.280 119.365 121.300 ;
        RECT 113.340 120.710 115.085 121.240 ;
        RECT 115.245 120.870 116.205 121.100 ;
        RECT 116.535 120.870 117.495 121.100 ;
        RECT 113.340 119.710 115.195 120.710 ;
        RECT 107.810 119.570 109.010 119.670 ;
        RECT 113.340 118.440 115.085 119.710 ;
        RECT 115.465 119.550 115.985 120.870 ;
        RECT 116.255 119.710 116.485 120.710 ;
        RECT 116.735 119.550 117.255 120.870 ;
        RECT 117.645 120.710 119.385 121.280 ;
        RECT 117.545 119.710 119.385 120.710 ;
        RECT 115.245 119.320 116.205 119.550 ;
        RECT 116.535 119.320 117.495 119.550 ;
        RECT 116.595 119.040 117.435 119.320 ;
        RECT 117.645 119.280 119.385 119.710 ;
        RECT 117.645 119.260 119.365 119.280 ;
        RECT 119.665 119.075 120.185 121.485 ;
        RECT 120.445 119.280 120.675 121.280 ;
        RECT 120.995 119.075 121.515 121.485 ;
        RECT 121.875 121.280 123.765 122.795 ;
        RECT 121.735 120.795 123.765 121.280 ;
        RECT 121.735 119.965 123.625 120.795 ;
        RECT 123.985 120.590 124.505 123.000 ;
        RECT 124.825 120.795 125.055 122.795 ;
        RECT 125.315 120.590 125.835 123.000 ;
        RECT 126.135 122.795 127.855 122.815 ;
        RECT 126.115 122.365 127.855 122.795 ;
        RECT 128.065 122.755 128.905 123.035 ;
        RECT 128.005 122.525 128.965 122.755 ;
        RECT 129.295 122.525 130.255 122.755 ;
        RECT 126.115 121.365 127.955 122.365 ;
        RECT 126.115 120.795 127.855 121.365 ;
        RECT 128.245 121.205 128.765 122.525 ;
        RECT 129.015 121.365 129.245 122.365 ;
        RECT 129.515 121.205 130.035 122.525 ;
        RECT 130.415 122.365 130.955 124.075 ;
        RECT 130.305 121.365 130.955 122.365 ;
        RECT 128.005 120.975 128.965 121.205 ;
        RECT 129.295 120.975 130.255 121.205 ;
        RECT 130.415 120.835 130.955 121.365 ;
        RECT 126.135 120.775 127.855 120.795 ;
        RECT 123.815 120.360 124.775 120.590 ;
        RECT 125.105 120.360 126.065 120.590 ;
        RECT 126.825 120.365 127.515 120.775 ;
        RECT 130.405 120.715 130.955 120.835 ;
        RECT 121.735 119.785 123.620 119.965 ;
        RECT 126.815 119.955 127.515 120.365 ;
        RECT 121.735 119.575 123.625 119.785 ;
        RECT 126.815 119.745 127.520 119.955 ;
        RECT 121.735 119.280 123.620 119.575 ;
        RECT 119.435 119.040 120.395 119.075 ;
        RECT 116.595 118.870 120.395 119.040 ;
        RECT 107.810 117.640 109.010 117.740 ;
        RECT 106.670 117.360 107.520 117.460 ;
        RECT 107.700 117.410 112.700 117.640 ;
        RECT 107.810 117.380 109.010 117.410 ;
        RECT 112.870 117.360 113.180 117.470 ;
        RECT 106.670 116.900 107.540 117.360 ;
        RECT 106.670 116.570 107.520 116.900 ;
        RECT 111.220 116.850 112.500 116.950 ;
        RECT 112.860 116.900 113.180 117.360 ;
        RECT 113.340 117.300 115.105 118.440 ;
        RECT 117.985 118.270 118.675 118.870 ;
        RECT 119.435 118.845 120.395 118.870 ;
        RECT 120.725 118.845 121.685 119.075 ;
        RECT 117.985 117.650 118.685 118.270 ;
        RECT 113.340 117.270 115.095 117.300 ;
        RECT 107.700 116.620 112.700 116.850 ;
        RECT 111.220 116.590 112.500 116.620 ;
        RECT 112.870 116.570 113.180 116.900 ;
        RECT 106.670 116.110 107.540 116.570 ;
        RECT 107.810 116.120 108.990 116.150 ;
        RECT 106.670 115.780 107.520 116.110 ;
        RECT 107.810 116.060 109.000 116.120 ;
        RECT 112.860 116.110 113.180 116.570 ;
        RECT 107.700 115.830 112.700 116.060 ;
        RECT 107.810 115.780 109.000 115.830 ;
        RECT 112.870 115.780 113.180 116.110 ;
        RECT 106.670 115.320 107.540 115.780 ;
        RECT 107.810 115.730 108.990 115.780 ;
        RECT 106.670 114.990 107.520 115.320 ;
        RECT 111.230 115.270 112.500 115.400 ;
        RECT 112.860 115.320 113.180 115.780 ;
        RECT 107.700 115.040 112.700 115.270 ;
        RECT 111.230 115.010 112.500 115.040 ;
        RECT 112.870 114.990 113.180 115.320 ;
        RECT 106.670 114.530 107.540 114.990 ;
        RECT 106.670 114.200 107.520 114.530 ;
        RECT 107.850 114.480 109.000 114.570 ;
        RECT 112.860 114.530 113.180 114.990 ;
        RECT 107.700 114.250 112.700 114.480 ;
        RECT 107.850 114.220 109.000 114.250 ;
        RECT 112.870 114.200 113.180 114.530 ;
        RECT 103.220 113.870 104.480 113.960 ;
        RECT 99.150 102.790 99.450 113.740 ;
        RECT 99.640 113.640 104.640 113.870 ;
        RECT 103.220 113.610 104.480 113.640 ;
        RECT 99.800 113.080 100.880 113.190 ;
        RECT 99.640 112.850 104.640 113.080 ;
        RECT 99.800 112.760 100.880 112.850 ;
        RECT 103.220 112.290 104.480 112.370 ;
        RECT 99.640 112.060 104.640 112.290 ;
        RECT 103.220 112.030 104.480 112.060 ;
        RECT 99.780 111.500 100.880 111.610 ;
        RECT 99.640 111.270 104.640 111.500 ;
        RECT 99.780 111.190 100.880 111.270 ;
        RECT 103.220 110.710 104.480 110.740 ;
        RECT 99.640 110.480 104.640 110.710 ;
        RECT 103.220 110.400 104.480 110.480 ;
        RECT 99.730 109.920 100.880 110.050 ;
        RECT 99.640 109.690 104.640 109.920 ;
        RECT 99.730 109.590 100.880 109.690 ;
        RECT 103.220 109.130 104.480 109.210 ;
        RECT 99.640 108.900 104.640 109.130 ;
        RECT 103.220 108.870 104.480 108.900 ;
        RECT 99.720 108.340 100.880 108.460 ;
        RECT 99.640 108.110 104.640 108.340 ;
        RECT 99.720 108.040 100.880 108.110 ;
        RECT 103.220 107.550 104.480 107.630 ;
        RECT 99.640 107.320 104.640 107.550 ;
        RECT 103.220 107.270 104.480 107.320 ;
        RECT 99.790 106.760 100.880 106.860 ;
        RECT 99.640 106.530 104.640 106.760 ;
        RECT 99.790 106.500 100.880 106.530 ;
        RECT 103.220 105.970 104.480 106.030 ;
        RECT 99.640 105.740 104.640 105.970 ;
        RECT 103.220 105.670 104.480 105.740 ;
        RECT 99.760 105.180 100.880 105.260 ;
        RECT 99.640 104.950 104.640 105.180 ;
        RECT 99.760 104.920 100.880 104.950 ;
        RECT 103.230 104.390 104.490 104.440 ;
        RECT 99.640 104.160 104.640 104.390 ;
        RECT 103.230 104.080 104.490 104.160 ;
        RECT 104.800 103.750 105.100 113.760 ;
        RECT 106.670 113.740 107.540 114.200 ;
        RECT 106.670 113.410 107.520 113.740 ;
        RECT 111.230 113.690 112.510 113.780 ;
        RECT 112.860 113.740 113.180 114.200 ;
        RECT 107.700 113.460 112.700 113.690 ;
        RECT 111.230 113.420 112.510 113.460 ;
        RECT 112.870 113.410 113.180 113.740 ;
        RECT 106.670 112.950 107.540 113.410 ;
        RECT 106.670 112.620 107.520 112.950 ;
        RECT 107.810 112.900 109.000 112.990 ;
        RECT 112.860 112.950 113.180 113.410 ;
        RECT 107.700 112.670 112.700 112.900 ;
        RECT 107.810 112.630 109.000 112.670 ;
        RECT 112.870 112.620 113.180 112.950 ;
        RECT 106.670 112.160 107.540 112.620 ;
        RECT 106.670 111.830 107.520 112.160 ;
        RECT 111.230 112.110 112.500 112.180 ;
        RECT 112.860 112.160 113.180 112.620 ;
        RECT 107.700 111.880 112.700 112.110 ;
        RECT 106.670 111.370 107.540 111.830 ;
        RECT 111.230 111.820 112.500 111.880 ;
        RECT 112.870 111.830 113.180 112.160 ;
        RECT 106.670 111.040 107.520 111.370 ;
        RECT 107.850 111.320 109.000 111.410 ;
        RECT 112.860 111.370 113.180 111.830 ;
        RECT 107.700 111.090 112.700 111.320 ;
        RECT 107.850 111.060 109.000 111.090 ;
        RECT 112.870 111.040 113.180 111.370 ;
        RECT 106.670 110.580 107.540 111.040 ;
        RECT 106.670 110.250 107.520 110.580 ;
        RECT 111.230 110.530 112.490 110.610 ;
        RECT 112.860 110.580 113.180 111.040 ;
        RECT 107.700 110.300 112.700 110.530 ;
        RECT 111.230 110.260 112.490 110.300 ;
        RECT 112.870 110.250 113.180 110.580 ;
        RECT 106.670 109.790 107.540 110.250 ;
        RECT 106.670 109.460 107.520 109.790 ;
        RECT 107.880 109.740 109.000 109.810 ;
        RECT 112.860 109.790 113.180 110.250 ;
        RECT 107.700 109.510 112.700 109.740 ;
        RECT 107.880 109.470 109.000 109.510 ;
        RECT 112.870 109.460 113.180 109.790 ;
        RECT 106.670 109.000 107.540 109.460 ;
        RECT 106.670 108.670 107.520 109.000 ;
        RECT 111.240 108.950 112.500 109.060 ;
        RECT 112.860 109.000 113.180 109.460 ;
        RECT 107.700 108.720 112.700 108.950 ;
        RECT 106.670 108.210 107.540 108.670 ;
        RECT 111.240 108.610 112.500 108.720 ;
        RECT 112.870 108.670 113.180 109.000 ;
        RECT 106.670 107.880 107.520 108.210 ;
        RECT 107.860 108.160 109.010 108.270 ;
        RECT 112.860 108.210 113.180 108.670 ;
        RECT 107.700 107.930 112.700 108.160 ;
        RECT 107.860 107.910 109.010 107.930 ;
        RECT 112.870 107.880 113.180 108.210 ;
        RECT 106.670 107.420 107.540 107.880 ;
        RECT 106.670 107.090 107.520 107.420 ;
        RECT 111.220 107.370 112.550 107.480 ;
        RECT 112.860 107.420 113.180 107.880 ;
        RECT 107.700 107.140 112.700 107.370 ;
        RECT 106.670 106.630 107.540 107.090 ;
        RECT 111.220 107.080 112.550 107.140 ;
        RECT 112.870 107.090 113.180 107.420 ;
        RECT 106.670 106.300 107.520 106.630 ;
        RECT 107.760 106.580 109.000 106.650 ;
        RECT 112.860 106.630 113.180 107.090 ;
        RECT 107.700 106.350 112.700 106.580 ;
        RECT 107.760 106.300 109.000 106.350 ;
        RECT 112.870 106.300 113.180 106.630 ;
        RECT 106.670 105.840 107.540 106.300 ;
        RECT 106.670 105.510 107.520 105.840 ;
        RECT 111.230 105.790 112.510 105.890 ;
        RECT 112.860 105.840 113.180 106.300 ;
        RECT 107.700 105.560 112.700 105.790 ;
        RECT 106.670 105.050 107.540 105.510 ;
        RECT 111.230 105.490 112.510 105.560 ;
        RECT 112.870 105.510 113.180 105.840 ;
        RECT 106.670 104.720 107.520 105.050 ;
        RECT 107.780 105.000 109.000 105.090 ;
        RECT 112.860 105.050 113.180 105.510 ;
        RECT 107.700 104.770 112.700 105.000 ;
        RECT 107.780 104.730 109.000 104.770 ;
        RECT 112.870 104.720 113.180 105.050 ;
        RECT 106.670 104.260 107.540 104.720 ;
        RECT 106.670 103.930 107.520 104.260 ;
        RECT 111.230 104.210 112.510 104.290 ;
        RECT 112.860 104.260 113.180 104.720 ;
        RECT 107.700 103.980 112.700 104.210 ;
        RECT 104.800 103.740 105.760 103.750 ;
        RECT 99.770 103.600 100.890 103.700 ;
        RECT 99.640 103.370 104.640 103.600 ;
        RECT 99.770 103.350 100.890 103.370 ;
        RECT 103.220 102.810 104.480 102.870 ;
        RECT 99.640 102.580 104.640 102.810 ;
        RECT 103.220 102.520 104.480 102.580 ;
        RECT 94.510 101.690 99.010 102.520 ;
        RECT 104.800 102.240 105.980 103.740 ;
        RECT 71.770 95.450 72.340 99.750 ;
        RECT 94.510 96.850 95.410 101.690 ;
        RECT 96.150 100.550 97.060 100.750 ;
        RECT 96.130 100.505 103.100 100.550 ;
        RECT 96.090 100.275 103.100 100.505 ;
        RECT 95.610 97.810 95.900 100.240 ;
        RECT 96.130 100.210 103.100 100.275 ;
        RECT 96.150 100.190 97.060 100.210 ;
        RECT 96.090 99.700 103.090 99.715 ;
        RECT 96.080 98.340 103.120 99.700 ;
        RECT 103.290 98.850 103.580 100.240 ;
        RECT 106.670 99.060 107.540 103.930 ;
        RECT 111.230 103.890 112.510 103.980 ;
        RECT 112.870 103.930 113.180 104.260 ;
        RECT 107.780 103.470 108.990 103.500 ;
        RECT 112.860 103.470 113.180 103.930 ;
        RECT 107.780 103.420 109.000 103.470 ;
        RECT 107.700 103.190 112.700 103.420 ;
        RECT 107.780 103.110 109.000 103.190 ;
        RECT 112.870 103.140 113.180 103.470 ;
        RECT 107.780 103.100 108.990 103.110 ;
        RECT 112.860 102.680 113.180 103.140 ;
        RECT 107.840 102.630 112.680 102.680 ;
        RECT 112.870 102.630 113.180 102.680 ;
        RECT 113.350 117.180 115.095 117.270 ;
        RECT 117.985 117.240 118.675 117.650 ;
        RECT 119.435 117.425 120.395 117.655 ;
        RECT 120.725 117.425 121.685 117.655 ;
        RECT 117.645 117.220 119.365 117.240 ;
        RECT 113.350 116.650 115.085 117.180 ;
        RECT 115.245 116.810 116.205 117.040 ;
        RECT 116.535 116.810 117.495 117.040 ;
        RECT 113.350 115.650 115.195 116.650 ;
        RECT 113.350 114.380 115.085 115.650 ;
        RECT 115.465 115.490 115.985 116.810 ;
        RECT 116.255 115.650 116.485 116.650 ;
        RECT 116.735 115.490 117.255 116.810 ;
        RECT 117.645 116.650 119.385 117.220 ;
        RECT 117.545 115.650 119.385 116.650 ;
        RECT 115.245 115.260 116.205 115.490 ;
        RECT 116.535 115.260 117.495 115.490 ;
        RECT 116.595 114.980 117.435 115.260 ;
        RECT 117.645 115.220 119.385 115.650 ;
        RECT 117.645 115.200 119.365 115.220 ;
        RECT 119.665 115.015 120.185 117.425 ;
        RECT 120.445 115.220 120.675 117.220 ;
        RECT 120.995 115.015 121.515 117.425 ;
        RECT 121.875 117.220 123.620 119.280 ;
        RECT 121.735 116.105 123.620 117.220 ;
        RECT 121.735 115.220 123.625 116.105 ;
        RECT 126.820 115.605 127.520 119.745 ;
        RECT 130.395 119.575 130.955 120.715 ;
        RECT 130.410 115.895 130.955 119.575 ;
        RECT 119.435 114.980 120.395 115.015 ;
        RECT 116.595 114.810 120.395 114.980 ;
        RECT 113.350 113.240 115.105 114.380 ;
        RECT 117.985 114.210 118.675 114.810 ;
        RECT 119.435 114.785 120.395 114.810 ;
        RECT 120.725 114.785 121.685 115.015 ;
        RECT 121.875 114.695 123.625 115.220 ;
        RECT 123.815 114.900 124.775 115.130 ;
        RECT 125.105 115.105 126.065 115.130 ;
        RECT 126.825 115.105 127.515 115.605 ;
        RECT 125.105 114.935 128.905 115.105 ;
        RECT 125.105 114.900 126.065 114.935 ;
        RECT 117.985 113.590 118.685 114.210 ;
        RECT 113.350 113.120 115.095 113.240 ;
        RECT 117.985 113.180 118.675 113.590 ;
        RECT 119.435 113.365 120.395 113.595 ;
        RECT 120.725 113.365 121.685 113.595 ;
        RECT 117.645 113.160 119.365 113.180 ;
        RECT 113.350 112.590 115.085 113.120 ;
        RECT 115.245 112.750 116.205 112.980 ;
        RECT 116.535 112.750 117.495 112.980 ;
        RECT 113.350 111.590 115.195 112.590 ;
        RECT 113.350 110.320 115.085 111.590 ;
        RECT 115.465 111.430 115.985 112.750 ;
        RECT 116.255 111.590 116.485 112.590 ;
        RECT 116.735 111.430 117.255 112.750 ;
        RECT 117.645 112.590 119.385 113.160 ;
        RECT 117.545 111.590 119.385 112.590 ;
        RECT 115.245 111.200 116.205 111.430 ;
        RECT 116.535 111.200 117.495 111.430 ;
        RECT 116.595 110.920 117.435 111.200 ;
        RECT 117.645 111.160 119.385 111.590 ;
        RECT 117.645 111.140 119.365 111.160 ;
        RECT 119.665 110.955 120.185 113.365 ;
        RECT 120.445 111.160 120.675 113.160 ;
        RECT 120.995 110.955 121.515 113.365 ;
        RECT 121.875 113.160 123.765 114.695 ;
        RECT 121.735 112.695 123.765 113.160 ;
        RECT 121.735 111.915 123.625 112.695 ;
        RECT 123.985 112.490 124.505 114.900 ;
        RECT 124.825 112.695 125.055 114.695 ;
        RECT 125.315 112.490 125.835 114.900 ;
        RECT 126.135 114.695 127.855 114.715 ;
        RECT 126.115 114.265 127.855 114.695 ;
        RECT 128.065 114.655 128.905 114.935 ;
        RECT 128.005 114.425 128.965 114.655 ;
        RECT 129.295 114.425 130.255 114.655 ;
        RECT 126.115 113.265 127.955 114.265 ;
        RECT 126.115 112.695 127.855 113.265 ;
        RECT 128.245 113.105 128.765 114.425 ;
        RECT 129.015 113.265 129.245 114.265 ;
        RECT 129.515 113.105 130.035 114.425 ;
        RECT 130.415 114.265 130.955 115.895 ;
        RECT 130.305 113.265 130.955 114.265 ;
        RECT 128.005 112.875 128.965 113.105 ;
        RECT 129.295 112.875 130.255 113.105 ;
        RECT 130.415 112.735 130.955 113.265 ;
        RECT 126.135 112.675 127.855 112.695 ;
        RECT 123.815 112.260 124.775 112.490 ;
        RECT 125.105 112.260 126.065 112.490 ;
        RECT 126.825 112.265 127.515 112.675 ;
        RECT 130.405 112.615 130.955 112.735 ;
        RECT 126.815 111.965 127.515 112.265 ;
        RECT 121.735 111.160 123.630 111.915 ;
        RECT 126.815 111.645 127.520 111.965 ;
        RECT 119.435 110.920 120.395 110.955 ;
        RECT 116.595 110.750 120.395 110.920 ;
        RECT 113.350 109.180 115.105 110.320 ;
        RECT 117.985 110.150 118.675 110.750 ;
        RECT 119.435 110.725 120.395 110.750 ;
        RECT 120.725 110.725 121.685 110.955 ;
        RECT 117.985 109.530 118.685 110.150 ;
        RECT 113.350 109.060 115.095 109.180 ;
        RECT 117.985 109.120 118.675 109.530 ;
        RECT 119.435 109.305 120.395 109.535 ;
        RECT 120.725 109.305 121.685 109.535 ;
        RECT 117.645 109.100 119.365 109.120 ;
        RECT 113.350 108.530 115.085 109.060 ;
        RECT 115.245 108.690 116.205 108.920 ;
        RECT 116.535 108.690 117.495 108.920 ;
        RECT 113.350 107.530 115.195 108.530 ;
        RECT 113.350 106.260 115.085 107.530 ;
        RECT 115.465 107.370 115.985 108.690 ;
        RECT 116.255 107.530 116.485 108.530 ;
        RECT 116.735 107.370 117.255 108.690 ;
        RECT 117.645 108.530 119.385 109.100 ;
        RECT 117.545 107.530 119.385 108.530 ;
        RECT 115.245 107.140 116.205 107.370 ;
        RECT 116.535 107.140 117.495 107.370 ;
        RECT 116.595 106.860 117.435 107.140 ;
        RECT 117.645 107.100 119.385 107.530 ;
        RECT 117.645 107.080 119.365 107.100 ;
        RECT 119.665 106.895 120.185 109.305 ;
        RECT 120.445 107.100 120.675 109.100 ;
        RECT 120.995 106.895 121.515 109.305 ;
        RECT 121.875 109.100 123.630 111.160 ;
        RECT 121.735 107.445 123.630 109.100 ;
        RECT 121.735 107.100 123.625 107.445 ;
        RECT 126.820 107.275 127.520 111.645 ;
        RECT 130.395 111.475 130.955 112.615 ;
        RECT 130.410 107.955 130.955 111.475 ;
        RECT 119.435 106.860 120.395 106.895 ;
        RECT 116.595 106.690 120.395 106.860 ;
        RECT 113.350 105.120 115.105 106.260 ;
        RECT 117.985 106.090 118.675 106.690 ;
        RECT 119.435 106.665 120.395 106.690 ;
        RECT 120.725 106.665 121.685 106.895 ;
        RECT 121.875 106.595 123.625 107.100 ;
        RECT 123.815 106.800 124.775 107.030 ;
        RECT 125.105 107.005 126.065 107.030 ;
        RECT 126.825 107.005 127.515 107.275 ;
        RECT 125.105 106.835 128.905 107.005 ;
        RECT 125.105 106.800 126.065 106.835 ;
        RECT 117.985 105.470 118.685 106.090 ;
        RECT 113.350 105.000 115.095 105.120 ;
        RECT 117.985 105.060 118.675 105.470 ;
        RECT 119.435 105.245 120.395 105.475 ;
        RECT 120.725 105.245 121.685 105.475 ;
        RECT 117.645 105.040 119.365 105.060 ;
        RECT 113.350 104.470 115.085 105.000 ;
        RECT 115.245 104.630 116.205 104.860 ;
        RECT 116.535 104.630 117.495 104.860 ;
        RECT 113.350 103.470 115.195 104.470 ;
        RECT 107.700 102.400 112.700 102.630 ;
        RECT 107.840 102.340 112.680 102.400 ;
        RECT 113.350 102.200 115.085 103.470 ;
        RECT 115.465 103.310 115.985 104.630 ;
        RECT 116.255 103.470 116.485 104.470 ;
        RECT 116.735 103.310 117.255 104.630 ;
        RECT 117.645 104.470 119.385 105.040 ;
        RECT 117.545 103.470 119.385 104.470 ;
        RECT 115.245 103.080 116.205 103.310 ;
        RECT 116.535 103.080 117.495 103.310 ;
        RECT 116.595 102.800 117.435 103.080 ;
        RECT 117.645 103.040 119.385 103.470 ;
        RECT 117.645 103.020 119.365 103.040 ;
        RECT 119.665 102.835 120.185 105.245 ;
        RECT 120.445 103.040 120.675 105.040 ;
        RECT 120.995 102.835 121.515 105.245 ;
        RECT 121.875 105.040 123.765 106.595 ;
        RECT 121.735 104.595 123.765 105.040 ;
        RECT 121.735 103.040 123.625 104.595 ;
        RECT 123.985 104.390 124.505 106.800 ;
        RECT 124.825 104.595 125.055 106.595 ;
        RECT 125.315 104.390 125.835 106.800 ;
        RECT 126.135 106.595 127.855 106.615 ;
        RECT 126.115 106.165 127.855 106.595 ;
        RECT 128.065 106.555 128.905 106.835 ;
        RECT 128.005 106.325 128.965 106.555 ;
        RECT 129.295 106.325 130.255 106.555 ;
        RECT 126.115 105.165 127.955 106.165 ;
        RECT 126.115 104.595 127.855 105.165 ;
        RECT 128.245 105.005 128.765 106.325 ;
        RECT 129.015 105.165 129.245 106.165 ;
        RECT 129.515 105.005 130.035 106.325 ;
        RECT 130.415 106.165 130.955 107.955 ;
        RECT 130.305 105.165 130.955 106.165 ;
        RECT 128.005 104.775 128.965 105.005 ;
        RECT 129.295 104.775 130.255 105.005 ;
        RECT 130.415 104.635 130.955 105.165 ;
        RECT 126.135 104.575 127.855 104.595 ;
        RECT 123.815 104.160 124.775 104.390 ;
        RECT 125.105 104.160 126.065 104.390 ;
        RECT 126.825 104.165 127.515 104.575 ;
        RECT 130.405 104.515 130.955 104.635 ;
        RECT 126.815 103.545 127.515 104.165 ;
        RECT 119.435 102.800 120.395 102.835 ;
        RECT 116.595 102.630 120.395 102.800 ;
        RECT 113.350 101.690 115.105 102.200 ;
        RECT 113.470 101.060 115.105 101.690 ;
        RECT 117.985 102.030 118.675 102.630 ;
        RECT 119.435 102.605 120.395 102.630 ;
        RECT 120.725 102.605 121.685 102.835 ;
        RECT 121.875 102.545 123.625 103.040 ;
        RECT 123.815 102.750 124.775 102.980 ;
        RECT 125.105 102.955 126.065 102.980 ;
        RECT 126.825 102.955 127.515 103.545 ;
        RECT 130.395 103.375 130.955 104.515 ;
        RECT 125.105 102.785 128.905 102.955 ;
        RECT 125.105 102.750 126.065 102.785 ;
        RECT 117.985 101.410 118.685 102.030 ;
        RECT 113.470 100.940 115.095 101.060 ;
        RECT 117.985 101.000 118.675 101.410 ;
        RECT 119.435 101.185 120.395 101.415 ;
        RECT 120.725 101.185 121.685 101.415 ;
        RECT 117.645 100.980 119.365 101.000 ;
        RECT 113.470 100.410 115.085 100.940 ;
        RECT 115.245 100.570 116.205 100.800 ;
        RECT 116.535 100.570 117.495 100.800 ;
        RECT 113.470 99.410 115.195 100.410 ;
        RECT 103.290 97.930 103.590 98.850 ;
        RECT 113.470 97.990 115.085 99.410 ;
        RECT 115.465 99.250 115.985 100.570 ;
        RECT 116.255 99.410 116.485 100.410 ;
        RECT 116.735 99.250 117.255 100.570 ;
        RECT 117.645 100.410 119.385 100.980 ;
        RECT 117.545 99.410 119.385 100.410 ;
        RECT 115.245 99.020 116.205 99.250 ;
        RECT 116.535 99.020 117.495 99.250 ;
        RECT 116.595 98.740 117.435 99.020 ;
        RECT 117.645 98.980 119.385 99.410 ;
        RECT 117.645 98.960 119.365 98.980 ;
        RECT 119.665 98.775 120.185 101.185 ;
        RECT 120.445 98.980 120.675 100.980 ;
        RECT 120.995 98.775 121.515 101.185 ;
        RECT 121.875 100.980 123.765 102.545 ;
        RECT 121.735 100.545 123.765 100.980 ;
        RECT 121.735 98.980 123.625 100.545 ;
        RECT 123.985 100.340 124.505 102.750 ;
        RECT 124.825 100.545 125.055 102.545 ;
        RECT 125.315 100.340 125.835 102.750 ;
        RECT 126.135 102.545 127.855 102.565 ;
        RECT 126.115 102.115 127.855 102.545 ;
        RECT 128.065 102.505 128.905 102.785 ;
        RECT 128.005 102.275 128.965 102.505 ;
        RECT 129.295 102.275 130.255 102.505 ;
        RECT 126.115 101.115 127.955 102.115 ;
        RECT 126.115 100.545 127.855 101.115 ;
        RECT 128.245 100.955 128.765 102.275 ;
        RECT 129.015 101.115 129.245 102.115 ;
        RECT 129.515 100.955 130.035 102.275 ;
        RECT 130.415 102.115 130.955 103.375 ;
        RECT 130.305 101.115 130.955 102.115 ;
        RECT 128.005 100.725 128.965 100.955 ;
        RECT 129.295 100.725 130.255 100.955 ;
        RECT 130.415 100.585 130.955 101.115 ;
        RECT 126.135 100.525 127.855 100.545 ;
        RECT 123.815 100.110 124.775 100.340 ;
        RECT 125.105 100.110 126.065 100.340 ;
        RECT 126.825 100.115 127.515 100.525 ;
        RECT 130.405 100.465 130.955 100.585 ;
        RECT 126.815 99.495 127.515 100.115 ;
        RECT 119.435 98.740 120.395 98.775 ;
        RECT 116.595 98.570 120.395 98.740 ;
        RECT 117.985 98.210 118.675 98.570 ;
        RECT 119.435 98.545 120.395 98.570 ;
        RECT 120.725 98.545 121.685 98.775 ;
        RECT 96.130 97.785 103.100 97.880 ;
        RECT 96.090 97.555 103.100 97.785 ;
        RECT 103.290 97.630 104.010 97.930 ;
        RECT 96.130 97.540 103.100 97.555 ;
        RECT 96.150 97.220 97.060 97.540 ;
        RECT 97.420 96.850 103.040 97.250 ;
        RECT 94.510 96.500 103.040 96.850 ;
        RECT 103.840 96.980 104.010 97.630 ;
        RECT 103.840 96.970 106.240 96.980 ;
        RECT 107.410 96.970 108.110 97.030 ;
        RECT 103.840 96.840 112.930 96.970 ;
        RECT 103.840 96.730 107.630 96.840 ;
        RECT 94.510 96.290 95.410 96.500 ;
        RECT 94.510 95.450 95.000 96.290 ;
        RECT 95.595 96.010 103.535 96.200 ;
        RECT 95.190 95.970 103.535 96.010 ;
        RECT 103.840 95.970 106.240 96.730 ;
        RECT 107.895 96.700 112.930 96.840 ;
        RECT 107.900 96.490 112.930 96.700 ;
        RECT 107.900 96.475 112.900 96.490 ;
        RECT 95.190 95.920 96.170 95.970 ;
        RECT 95.160 95.670 96.170 95.920 ;
        RECT 95.160 95.460 95.390 95.670 ;
        RECT 103.300 95.460 103.535 95.970 ;
        RECT 104.165 95.460 104.555 95.970 ;
        RECT 71.770 95.120 95.000 95.450 ;
        RECT 95.595 95.380 103.095 95.410 ;
        RECT 95.570 95.180 103.095 95.380 ;
        RECT 103.305 95.290 103.535 95.460 ;
        RECT 105.950 95.440 106.240 95.970 ;
        RECT 107.510 96.060 107.740 96.425 ;
        RECT 113.060 96.060 113.290 96.425 ;
        RECT 107.510 95.720 113.290 96.060 ;
        RECT 107.510 95.465 107.740 95.720 ;
        RECT 113.060 95.465 113.290 95.720 ;
        RECT 103.710 95.290 104.090 95.320 ;
        RECT 103.305 95.270 104.090 95.290 ;
        RECT 104.755 95.270 105.755 95.410 ;
        RECT 107.900 95.390 112.900 95.415 ;
        RECT 113.470 95.390 115.090 97.990 ;
        RECT 103.305 95.180 105.755 95.270 ;
        RECT 107.880 95.240 112.900 95.390 ;
        RECT 113.450 95.240 115.090 95.390 ;
        RECT 95.570 95.120 96.350 95.180 ;
        RECT 71.770 94.460 96.350 95.120 ;
        RECT 103.305 95.060 105.730 95.180 ;
        RECT 107.880 94.550 115.090 95.240 ;
        RECT 71.770 67.250 72.340 94.460 ;
        RECT 80.240 93.660 81.470 94.460 ;
        RECT 113.340 94.080 115.090 94.550 ;
        RECT 117.980 97.790 118.675 98.210 ;
        RECT 121.875 98.495 123.625 98.980 ;
        RECT 123.815 98.700 124.775 98.930 ;
        RECT 125.105 98.905 126.065 98.930 ;
        RECT 126.825 98.905 127.515 99.495 ;
        RECT 130.395 99.325 130.955 100.465 ;
        RECT 125.105 98.735 128.905 98.905 ;
        RECT 125.105 98.700 126.065 98.735 ;
        RECT 121.875 98.060 123.765 98.495 ;
        RECT 77.260 91.810 78.510 91.830 ;
        RECT 73.050 91.790 78.510 91.810 ;
        RECT 72.560 91.580 78.510 91.790 ;
        RECT 72.560 91.510 73.280 91.580 ;
        RECT 72.530 91.420 73.280 91.510 ;
        RECT 77.260 91.560 78.510 91.580 ;
        RECT 77.260 91.480 78.560 91.560 ;
        RECT 72.530 82.860 72.860 91.420 ;
        RECT 77.090 91.020 78.090 91.100 ;
        RECT 73.050 90.790 78.090 91.020 ;
        RECT 77.090 90.640 78.090 90.790 ;
        RECT 77.090 87.310 78.060 87.700 ;
        RECT 73.050 87.080 78.060 87.310 ;
        RECT 77.090 86.980 78.060 87.080 ;
        RECT 77.090 86.520 78.030 86.570 ;
        RECT 73.050 86.290 78.050 86.520 ;
        RECT 77.090 86.100 78.030 86.290 ;
        RECT 72.530 82.810 73.370 82.860 ;
        RECT 78.230 82.820 78.560 91.480 ;
        RECT 77.270 82.810 78.560 82.820 ;
        RECT 72.530 82.600 78.560 82.810 ;
        RECT 72.530 81.990 72.860 82.600 ;
        RECT 73.050 82.580 78.560 82.600 ;
        RECT 77.270 82.530 78.560 82.580 ;
        RECT 77.070 82.020 78.020 82.150 ;
        RECT 78.230 82.040 78.560 82.530 ;
        RECT 73.050 81.790 78.050 82.020 ;
        RECT 77.070 81.710 78.020 81.790 ;
        RECT 78.750 81.460 79.140 91.920 ;
        RECT 79.680 81.510 80.320 92.000 ;
        RECT 80.800 81.330 81.190 93.660 ;
        RECT 106.220 93.600 107.150 93.640 ;
        RECT 106.220 93.370 111.230 93.600 ;
        RECT 106.220 93.320 107.150 93.370 ;
        RECT 93.080 92.290 94.810 92.630 ;
        RECT 82.020 91.810 82.680 92.030 ;
        RECT 85.030 91.810 86.830 92.250 ;
        RECT 90.770 92.060 95.770 92.290 ;
        RECT 82.020 91.580 87.050 91.810 ;
        RECT 82.020 91.560 82.680 91.580 ;
        RECT 81.510 91.070 81.845 91.530 ;
        RECT 85.030 91.430 86.830 91.580 ;
        RECT 81.510 87.540 81.840 91.070 ;
        RECT 82.080 91.020 82.900 91.120 ;
        RECT 82.050 90.790 87.050 91.020 ;
        RECT 82.080 90.620 82.900 90.790 ;
        RECT 81.510 87.310 82.830 87.540 ;
        RECT 87.210 87.360 87.540 91.540 ;
        RECT 90.380 91.050 90.610 92.010 ;
        RECT 95.930 91.050 97.040 92.450 ;
        RECT 100.260 92.290 101.780 92.480 ;
        RECT 97.770 92.060 102.770 92.290 ;
        RECT 95.960 91.010 97.040 91.050 ;
        RECT 90.770 90.970 95.770 91.000 ;
        RECT 90.740 90.080 95.790 90.970 ;
        RECT 90.770 90.060 95.770 90.080 ;
        RECT 96.700 90.060 97.040 91.010 ;
        RECT 97.270 90.990 97.620 92.030 ;
        RECT 100.260 91.960 101.780 92.060 ;
        RECT 102.930 91.050 103.160 92.010 ;
        RECT 97.770 90.970 102.770 91.000 ;
        RECT 97.770 90.770 102.800 90.970 ;
        RECT 97.980 90.290 102.800 90.770 ;
        RECT 97.770 90.080 102.800 90.290 ;
        RECT 97.770 90.060 102.770 90.080 ;
        RECT 86.880 87.310 87.540 87.360 ;
        RECT 81.510 87.190 87.540 87.310 ;
        RECT 81.510 87.030 81.840 87.190 ;
        RECT 82.050 87.110 87.540 87.190 ;
        RECT 82.050 87.080 87.050 87.110 ;
        RECT 81.510 86.570 81.845 87.030 ;
        RECT 81.510 82.530 81.840 86.570 ;
        RECT 82.140 86.520 82.860 86.740 ;
        RECT 82.050 86.290 87.050 86.520 ;
        RECT 82.140 86.170 82.860 86.290 ;
        RECT 87.210 86.110 87.540 87.110 ;
        RECT 89.720 90.010 90.580 90.040 ;
        RECT 89.720 89.050 90.610 90.010 ;
        RECT 89.720 89.030 90.580 89.050 ;
        RECT 89.720 88.450 90.040 89.030 ;
        RECT 90.760 89.000 92.650 89.270 ;
        RECT 95.930 89.050 96.160 90.010 ;
        RECT 96.700 89.010 97.610 90.060 ;
        RECT 90.760 88.770 95.770 89.000 ;
        RECT 90.760 88.650 92.650 88.770 ;
        RECT 96.700 88.480 97.040 89.010 ;
        RECT 98.190 89.000 99.710 89.160 ;
        RECT 102.930 89.050 103.160 90.010 ;
        RECT 97.770 88.770 102.770 89.000 ;
        RECT 98.190 88.640 99.710 88.770 ;
        RECT 89.720 86.820 90.050 88.450 ;
        RECT 87.210 85.220 87.870 86.110 ;
        RECT 82.010 82.810 82.630 83.020 ;
        RECT 82.010 82.580 87.050 82.810 ;
        RECT 81.510 82.070 81.845 82.530 ;
        RECT 82.010 82.520 82.630 82.580 ;
        RECT 81.510 82.010 81.840 82.070 ;
        RECT 82.190 82.020 82.910 82.160 ;
        RECT 87.210 82.020 87.540 85.220 ;
        RECT 89.720 84.370 90.040 86.820 ;
        RECT 93.080 86.290 94.810 86.620 ;
        RECT 90.770 86.060 95.770 86.290 ;
        RECT 96.710 86.030 97.030 88.480 ;
        RECT 97.220 86.960 97.610 87.990 ;
        RECT 95.970 86.010 97.030 86.030 ;
        RECT 90.380 85.050 90.610 86.010 ;
        RECT 95.930 85.050 97.030 86.010 ;
        RECT 95.970 85.030 97.030 85.050 ;
        RECT 90.770 84.970 95.770 85.000 ;
        RECT 88.930 84.030 90.040 84.370 ;
        RECT 90.750 84.080 95.800 84.970 ;
        RECT 90.770 84.060 95.770 84.080 ;
        RECT 96.710 84.050 97.030 85.030 ;
        RECT 97.330 85.020 97.610 86.960 ;
        RECT 105.790 87.910 106.070 93.320 ;
        RECT 110.230 92.310 111.180 92.400 ;
        RECT 111.380 92.360 112.530 93.330 ;
        RECT 113.340 92.940 115.105 94.080 ;
        RECT 117.980 93.910 118.670 97.790 ;
        RECT 121.870 96.495 123.765 98.060 ;
        RECT 121.870 94.445 123.625 96.495 ;
        RECT 123.985 96.290 124.505 98.700 ;
        RECT 124.825 96.495 125.055 98.495 ;
        RECT 125.315 96.290 125.835 98.700 ;
        RECT 126.135 98.495 127.855 98.515 ;
        RECT 126.115 98.065 127.855 98.495 ;
        RECT 128.065 98.455 128.905 98.735 ;
        RECT 128.005 98.225 128.965 98.455 ;
        RECT 129.295 98.225 130.255 98.455 ;
        RECT 126.115 97.065 127.955 98.065 ;
        RECT 126.115 96.495 127.855 97.065 ;
        RECT 128.245 96.905 128.765 98.225 ;
        RECT 129.015 97.065 129.245 98.065 ;
        RECT 129.515 96.905 130.035 98.225 ;
        RECT 130.415 98.065 130.955 99.325 ;
        RECT 130.305 97.065 130.955 98.065 ;
        RECT 128.005 96.675 128.965 96.905 ;
        RECT 129.295 96.675 130.255 96.905 ;
        RECT 130.415 96.535 130.955 97.065 ;
        RECT 126.135 96.475 127.855 96.495 ;
        RECT 123.815 96.060 124.775 96.290 ;
        RECT 125.105 96.060 126.065 96.290 ;
        RECT 126.825 96.065 127.515 96.475 ;
        RECT 130.405 96.415 130.955 96.535 ;
        RECT 126.815 95.445 127.515 96.065 ;
        RECT 123.815 94.650 124.775 94.880 ;
        RECT 125.105 94.855 126.065 94.880 ;
        RECT 126.825 94.855 127.515 95.445 ;
        RECT 130.395 95.275 130.955 96.415 ;
        RECT 125.105 94.685 128.905 94.855 ;
        RECT 125.105 94.650 126.065 94.685 ;
        RECT 117.980 93.650 118.685 93.910 ;
        RECT 121.870 93.650 123.765 94.445 ;
        RECT 117.985 93.290 118.685 93.650 ;
        RECT 113.340 92.820 115.095 92.940 ;
        RECT 117.985 92.880 118.675 93.290 ;
        RECT 119.435 93.065 120.395 93.295 ;
        RECT 120.725 93.065 121.685 93.295 ;
        RECT 117.645 92.860 119.365 92.880 ;
        RECT 106.230 92.080 111.240 92.310 ;
        RECT 110.230 92.000 111.180 92.080 ;
        RECT 111.420 92.030 111.810 92.360 ;
        RECT 106.230 91.020 107.150 91.080 ;
        RECT 111.390 91.070 111.810 92.030 ;
        RECT 106.230 91.010 111.230 91.020 ;
        RECT 106.230 90.780 111.240 91.010 ;
        RECT 106.230 90.710 107.150 90.780 ;
        RECT 111.420 90.740 111.810 91.070 ;
        RECT 111.390 89.780 111.810 90.740 ;
        RECT 110.230 89.730 111.180 89.780 ;
        RECT 106.230 89.720 111.230 89.730 ;
        RECT 106.230 89.500 111.240 89.720 ;
        RECT 106.280 89.490 111.240 89.500 ;
        RECT 110.230 89.400 111.180 89.490 ;
        RECT 111.420 89.450 111.810 89.780 ;
        RECT 106.230 88.440 107.160 88.530 ;
        RECT 111.390 88.490 111.810 89.450 ;
        RECT 106.230 88.210 111.240 88.440 ;
        RECT 106.230 88.150 107.160 88.210 ;
        RECT 111.420 88.160 111.810 88.490 ;
        RECT 111.390 87.910 111.810 88.160 ;
        RECT 105.790 87.460 106.160 87.910 ;
        RECT 111.340 87.460 111.810 87.910 ;
        RECT 100.290 86.290 101.810 86.490 ;
        RECT 97.770 86.060 102.770 86.290 ;
        RECT 100.290 85.970 101.810 86.060 ;
        RECT 102.930 85.050 103.160 86.010 ;
        RECT 97.770 84.980 102.770 85.000 ;
        RECT 97.750 84.790 102.790 84.980 ;
        RECT 97.740 84.090 102.790 84.790 ;
        RECT 97.770 84.060 102.770 84.090 ;
        RECT 96.710 84.030 97.580 84.050 ;
        RECT 88.930 84.010 90.590 84.030 ;
        RECT 96.710 84.010 97.600 84.030 ;
        RECT 88.930 83.050 90.610 84.010 ;
        RECT 95.930 83.050 96.160 84.010 ;
        RECT 96.710 83.050 97.610 84.010 ;
        RECT 88.930 83.020 90.520 83.050 ;
        RECT 90.800 83.000 92.520 83.050 ;
        RECT 96.720 83.040 97.580 83.050 ;
        RECT 98.200 83.000 99.720 83.190 ;
        RECT 102.930 83.050 103.160 84.010 ;
        RECT 90.770 82.770 95.770 83.000 ;
        RECT 97.770 82.770 102.770 83.000 ;
        RECT 90.800 82.630 92.520 82.770 ;
        RECT 98.200 82.670 99.720 82.770 ;
        RECT 104.040 82.470 104.620 84.120 ;
        RECT 105.790 83.310 106.070 87.460 ;
        RECT 110.230 87.150 111.170 87.230 ;
        RECT 111.390 87.200 111.810 87.460 ;
        RECT 106.230 87.140 111.230 87.150 ;
        RECT 106.230 86.920 111.240 87.140 ;
        RECT 106.280 86.910 111.240 86.920 ;
        RECT 110.230 86.840 111.170 86.910 ;
        RECT 111.420 86.870 111.810 87.200 ;
        RECT 106.230 85.860 107.150 85.980 ;
        RECT 111.390 85.910 111.810 86.870 ;
        RECT 106.230 85.630 111.240 85.860 ;
        RECT 106.230 85.560 107.150 85.630 ;
        RECT 111.420 85.580 111.810 85.910 ;
        RECT 110.150 84.570 111.250 84.810 ;
        RECT 111.390 84.620 111.810 85.580 ;
        RECT 113.340 92.290 115.085 92.820 ;
        RECT 115.245 92.450 116.205 92.680 ;
        RECT 116.535 92.450 117.495 92.680 ;
        RECT 113.340 91.290 115.195 92.290 ;
        RECT 113.340 90.020 115.085 91.290 ;
        RECT 115.465 91.130 115.985 92.450 ;
        RECT 116.255 91.290 116.485 92.290 ;
        RECT 116.735 91.130 117.255 92.450 ;
        RECT 117.645 92.290 119.385 92.860 ;
        RECT 117.545 91.290 119.385 92.290 ;
        RECT 115.245 90.900 116.205 91.130 ;
        RECT 116.535 90.900 117.495 91.130 ;
        RECT 116.595 90.620 117.435 90.900 ;
        RECT 117.645 90.860 119.385 91.290 ;
        RECT 117.645 90.840 119.365 90.860 ;
        RECT 119.665 90.655 120.185 93.065 ;
        RECT 120.445 90.860 120.675 92.860 ;
        RECT 120.995 90.655 121.515 93.065 ;
        RECT 121.875 92.860 123.765 93.650 ;
        RECT 121.735 92.445 123.765 92.860 ;
        RECT 121.735 90.860 123.625 92.445 ;
        RECT 123.985 92.240 124.505 94.650 ;
        RECT 124.825 92.445 125.055 94.445 ;
        RECT 125.315 92.240 125.835 94.650 ;
        RECT 126.135 94.445 127.855 94.465 ;
        RECT 126.115 94.015 127.855 94.445 ;
        RECT 128.065 94.405 128.905 94.685 ;
        RECT 128.005 94.175 128.965 94.405 ;
        RECT 129.295 94.175 130.255 94.405 ;
        RECT 126.115 93.015 127.955 94.015 ;
        RECT 126.115 92.445 127.855 93.015 ;
        RECT 128.245 92.855 128.765 94.175 ;
        RECT 129.015 93.015 129.245 94.015 ;
        RECT 129.515 92.855 130.035 94.175 ;
        RECT 130.415 94.015 130.955 95.275 ;
        RECT 130.305 93.015 130.955 94.015 ;
        RECT 128.005 92.625 128.965 92.855 ;
        RECT 129.295 92.625 130.255 92.855 ;
        RECT 130.415 92.485 130.955 93.015 ;
        RECT 126.135 92.425 127.855 92.445 ;
        RECT 123.815 92.010 124.775 92.240 ;
        RECT 125.105 92.010 126.065 92.240 ;
        RECT 126.825 92.015 127.515 92.425 ;
        RECT 130.405 92.365 130.955 92.485 ;
        RECT 126.815 91.395 127.515 92.015 ;
        RECT 119.435 90.620 120.395 90.655 ;
        RECT 116.595 90.450 120.395 90.620 ;
        RECT 113.340 88.880 115.105 90.020 ;
        RECT 117.985 89.850 118.675 90.450 ;
        RECT 119.435 90.425 120.395 90.450 ;
        RECT 120.725 90.425 121.685 90.655 ;
        RECT 121.875 90.395 123.625 90.860 ;
        RECT 123.815 90.600 124.775 90.830 ;
        RECT 125.105 90.805 126.065 90.830 ;
        RECT 126.825 90.805 127.515 91.395 ;
        RECT 130.395 91.225 130.955 92.365 ;
        RECT 125.105 90.635 128.905 90.805 ;
        RECT 125.105 90.600 126.065 90.635 ;
        RECT 117.985 89.230 118.685 89.850 ;
        RECT 113.340 88.760 115.095 88.880 ;
        RECT 117.985 88.820 118.675 89.230 ;
        RECT 119.435 89.005 120.395 89.235 ;
        RECT 120.725 89.005 121.685 89.235 ;
        RECT 117.645 88.800 119.365 88.820 ;
        RECT 113.340 88.230 115.085 88.760 ;
        RECT 115.245 88.390 116.205 88.620 ;
        RECT 116.535 88.390 117.495 88.620 ;
        RECT 113.340 87.230 115.195 88.230 ;
        RECT 113.340 85.960 115.085 87.230 ;
        RECT 115.465 87.070 115.985 88.390 ;
        RECT 116.255 87.230 116.485 88.230 ;
        RECT 116.735 87.070 117.255 88.390 ;
        RECT 117.645 88.230 119.385 88.800 ;
        RECT 117.545 87.230 119.385 88.230 ;
        RECT 115.245 86.840 116.205 87.070 ;
        RECT 116.535 86.840 117.495 87.070 ;
        RECT 116.595 86.560 117.435 86.840 ;
        RECT 117.645 86.800 119.385 87.230 ;
        RECT 117.645 86.780 119.365 86.800 ;
        RECT 119.665 86.595 120.185 89.005 ;
        RECT 120.445 86.800 120.675 88.800 ;
        RECT 120.995 86.595 121.515 89.005 ;
        RECT 121.875 88.800 123.765 90.395 ;
        RECT 121.735 88.395 123.765 88.800 ;
        RECT 121.735 86.800 123.625 88.395 ;
        RECT 123.985 88.190 124.505 90.600 ;
        RECT 124.825 88.395 125.055 90.395 ;
        RECT 125.315 88.190 125.835 90.600 ;
        RECT 126.135 90.395 127.855 90.415 ;
        RECT 126.115 89.965 127.855 90.395 ;
        RECT 128.065 90.355 128.905 90.635 ;
        RECT 128.005 90.125 128.965 90.355 ;
        RECT 129.295 90.125 130.255 90.355 ;
        RECT 126.115 88.965 127.955 89.965 ;
        RECT 126.115 88.395 127.855 88.965 ;
        RECT 128.245 88.805 128.765 90.125 ;
        RECT 129.015 88.965 129.245 89.965 ;
        RECT 129.515 88.805 130.035 90.125 ;
        RECT 130.415 89.965 130.955 91.225 ;
        RECT 130.305 88.965 130.955 89.965 ;
        RECT 128.005 88.575 128.965 88.805 ;
        RECT 129.295 88.575 130.255 88.805 ;
        RECT 130.415 88.435 130.955 88.965 ;
        RECT 126.135 88.375 127.855 88.395 ;
        RECT 123.815 87.960 124.775 88.190 ;
        RECT 125.105 87.960 126.065 88.190 ;
        RECT 126.825 87.965 127.515 88.375 ;
        RECT 130.405 88.315 130.955 88.435 ;
        RECT 126.815 87.345 127.515 87.965 ;
        RECT 119.435 86.560 120.395 86.595 ;
        RECT 116.595 86.390 120.395 86.560 ;
        RECT 113.340 84.820 115.105 85.960 ;
        RECT 117.985 85.790 118.675 86.390 ;
        RECT 119.435 86.365 120.395 86.390 ;
        RECT 120.725 86.365 121.685 86.595 ;
        RECT 121.875 86.345 123.625 86.800 ;
        RECT 123.815 86.550 124.775 86.780 ;
        RECT 125.105 86.755 126.065 86.780 ;
        RECT 126.825 86.755 127.515 87.345 ;
        RECT 130.395 87.175 130.955 88.315 ;
        RECT 125.105 86.585 128.905 86.755 ;
        RECT 125.105 86.550 126.065 86.585 ;
        RECT 117.985 85.170 118.685 85.790 ;
        RECT 113.340 84.800 115.095 84.820 ;
        RECT 106.230 84.340 111.250 84.570 ;
        RECT 110.150 84.140 111.250 84.340 ;
        RECT 111.420 84.290 111.810 84.620 ;
        RECT 106.230 83.280 107.150 83.400 ;
        RECT 111.390 83.330 111.810 84.290 ;
        RECT 113.170 84.700 115.095 84.800 ;
        RECT 117.985 84.760 118.675 85.170 ;
        RECT 119.435 84.945 120.395 85.175 ;
        RECT 120.725 84.945 121.685 85.175 ;
        RECT 117.645 84.740 119.365 84.760 ;
        RECT 113.170 84.170 115.085 84.700 ;
        RECT 115.245 84.330 116.205 84.560 ;
        RECT 116.535 84.330 117.495 84.560 ;
        RECT 113.170 84.140 115.195 84.170 ;
        RECT 111.420 83.310 111.810 83.330 ;
        RECT 106.230 83.050 111.250 83.280 ;
        RECT 113.340 83.170 115.195 84.140 ;
        RECT 106.230 82.980 107.150 83.050 ;
        RECT 113.340 82.470 115.085 83.170 ;
        RECT 115.465 83.010 115.985 84.330 ;
        RECT 116.255 83.170 116.485 84.170 ;
        RECT 116.735 83.010 117.255 84.330 ;
        RECT 117.645 84.170 119.385 84.740 ;
        RECT 117.545 83.170 119.385 84.170 ;
        RECT 115.245 82.780 116.205 83.010 ;
        RECT 116.535 82.780 117.495 83.010 ;
        RECT 82.050 81.790 87.050 82.020 ;
        RECT 104.040 81.900 115.085 82.470 ;
        RECT 116.595 82.500 117.435 82.780 ;
        RECT 117.645 82.740 119.385 83.170 ;
        RECT 117.645 82.720 119.365 82.740 ;
        RECT 119.665 82.535 120.185 84.945 ;
        RECT 120.445 82.740 120.675 84.740 ;
        RECT 120.995 82.535 121.515 84.945 ;
        RECT 121.875 84.740 123.765 86.345 ;
        RECT 121.735 84.345 123.765 84.740 ;
        RECT 121.735 82.740 123.625 84.345 ;
        RECT 123.985 84.140 124.505 86.550 ;
        RECT 124.825 84.345 125.055 86.345 ;
        RECT 125.315 84.140 125.835 86.550 ;
        RECT 126.135 86.345 127.855 86.365 ;
        RECT 126.115 85.915 127.855 86.345 ;
        RECT 128.065 86.305 128.905 86.585 ;
        RECT 128.005 86.075 128.965 86.305 ;
        RECT 129.295 86.075 130.255 86.305 ;
        RECT 126.115 84.915 127.955 85.915 ;
        RECT 126.115 84.345 127.855 84.915 ;
        RECT 128.245 84.755 128.765 86.075 ;
        RECT 129.015 84.915 129.245 85.915 ;
        RECT 129.515 84.755 130.035 86.075 ;
        RECT 130.415 85.915 130.955 87.175 ;
        RECT 130.305 84.915 130.955 85.915 ;
        RECT 128.005 84.525 128.965 84.755 ;
        RECT 129.295 84.525 130.255 84.755 ;
        RECT 130.415 84.385 130.955 84.915 ;
        RECT 126.135 84.325 127.855 84.345 ;
        RECT 123.815 83.910 124.775 84.140 ;
        RECT 125.105 83.910 126.065 84.140 ;
        RECT 126.825 83.915 127.515 84.325 ;
        RECT 130.405 84.265 130.955 84.385 ;
        RECT 126.815 83.295 127.515 83.915 ;
        RECT 119.435 82.500 120.395 82.535 ;
        RECT 116.595 82.330 120.395 82.500 ;
        RECT 82.190 81.590 82.910 81.790 ;
        RECT 104.040 81.610 115.105 81.900 ;
        RECT 80.630 80.380 81.310 81.330 ;
        RECT 113.340 80.760 115.105 81.610 ;
        RECT 117.985 81.730 118.675 82.330 ;
        RECT 119.435 82.305 120.395 82.330 ;
        RECT 120.725 82.305 121.685 82.535 ;
        RECT 121.875 82.295 123.625 82.740 ;
        RECT 123.815 82.500 124.775 82.730 ;
        RECT 125.105 82.705 126.065 82.730 ;
        RECT 126.825 82.705 127.515 83.295 ;
        RECT 130.395 83.125 130.955 84.265 ;
        RECT 125.105 82.535 128.905 82.705 ;
        RECT 125.105 82.500 126.065 82.535 ;
        RECT 117.985 81.110 118.685 81.730 ;
        RECT 113.340 80.640 115.095 80.760 ;
        RECT 117.985 80.700 118.675 81.110 ;
        RECT 119.435 80.885 120.395 81.115 ;
        RECT 120.725 80.885 121.685 81.115 ;
        RECT 117.645 80.680 119.365 80.700 ;
        RECT 77.070 79.920 78.020 80.000 ;
        RECT 72.530 79.110 72.860 79.720 ;
        RECT 73.050 79.690 78.050 79.920 ;
        RECT 77.070 79.560 78.020 79.690 ;
        RECT 78.230 79.180 78.560 79.670 ;
        RECT 77.270 79.130 78.560 79.180 ;
        RECT 73.050 79.110 78.560 79.130 ;
        RECT 72.530 78.900 78.560 79.110 ;
        RECT 72.530 78.850 73.370 78.900 ;
        RECT 77.270 78.890 78.560 78.900 ;
        RECT 72.530 70.290 72.860 78.850 ;
        RECT 77.090 75.420 78.030 75.610 ;
        RECT 73.050 75.190 78.050 75.420 ;
        RECT 77.090 75.140 78.030 75.190 ;
        RECT 77.090 74.630 78.060 74.730 ;
        RECT 73.050 74.400 78.060 74.630 ;
        RECT 77.090 74.010 78.060 74.400 ;
        RECT 77.090 70.920 78.090 71.070 ;
        RECT 73.050 70.690 78.090 70.920 ;
        RECT 77.090 70.610 78.090 70.690 ;
        RECT 72.530 70.200 73.280 70.290 ;
        RECT 78.230 70.230 78.560 78.890 ;
        RECT 72.560 70.130 73.280 70.200 ;
        RECT 77.260 70.150 78.560 70.230 ;
        RECT 77.260 70.130 78.510 70.150 ;
        RECT 72.560 69.920 78.510 70.130 ;
        RECT 73.050 69.900 78.510 69.920 ;
        RECT 77.260 69.880 78.510 69.900 ;
        RECT 78.750 69.790 79.140 80.250 ;
        RECT 79.680 69.710 80.320 80.200 ;
        RECT 80.800 68.050 81.190 80.380 ;
        RECT 82.190 79.920 82.910 80.120 ;
        RECT 113.340 80.110 115.085 80.640 ;
        RECT 115.245 80.270 116.205 80.500 ;
        RECT 116.535 80.270 117.495 80.500 ;
        RECT 113.340 80.100 115.195 80.110 ;
        RECT 81.510 79.640 81.840 79.700 ;
        RECT 82.050 79.690 87.050 79.920 ;
        RECT 81.510 79.180 81.845 79.640 ;
        RECT 82.190 79.550 82.910 79.690 ;
        RECT 81.510 75.140 81.840 79.180 ;
        RECT 82.010 79.130 82.630 79.190 ;
        RECT 82.010 78.900 87.050 79.130 ;
        RECT 82.010 78.690 82.630 78.900 ;
        RECT 87.210 76.490 87.540 79.690 ;
        RECT 104.040 79.240 115.195 80.100 ;
        RECT 90.800 78.940 92.520 79.080 ;
        RECT 98.200 78.940 99.720 79.040 ;
        RECT 90.770 78.710 95.770 78.940 ;
        RECT 97.770 78.710 102.770 78.940 ;
        RECT 88.930 78.660 90.520 78.690 ;
        RECT 90.800 78.660 92.520 78.710 ;
        RECT 96.720 78.660 97.580 78.670 ;
        RECT 88.930 77.700 90.610 78.660 ;
        RECT 95.930 77.700 96.160 78.660 ;
        RECT 96.710 77.700 97.610 78.660 ;
        RECT 98.200 78.520 99.720 78.710 ;
        RECT 102.930 77.700 103.160 78.660 ;
        RECT 88.930 77.680 90.590 77.700 ;
        RECT 96.710 77.680 97.600 77.700 ;
        RECT 88.930 77.340 90.040 77.680 ;
        RECT 96.710 77.660 97.580 77.680 ;
        RECT 90.770 77.630 95.770 77.650 ;
        RECT 87.210 75.600 87.870 76.490 ;
        RECT 82.140 75.420 82.860 75.540 ;
        RECT 82.050 75.190 87.050 75.420 ;
        RECT 81.510 74.680 81.845 75.140 ;
        RECT 82.140 74.970 82.860 75.190 ;
        RECT 81.510 74.520 81.840 74.680 ;
        RECT 82.050 74.600 87.050 74.630 ;
        RECT 87.210 74.600 87.540 75.600 ;
        RECT 82.050 74.520 87.540 74.600 ;
        RECT 81.510 74.400 87.540 74.520 ;
        RECT 81.510 74.170 82.830 74.400 ;
        RECT 86.880 74.350 87.540 74.400 ;
        RECT 81.510 70.640 81.840 74.170 ;
        RECT 82.080 70.920 82.900 71.090 ;
        RECT 82.050 70.690 87.050 70.920 ;
        RECT 81.510 70.180 81.845 70.640 ;
        RECT 82.080 70.590 82.900 70.690 ;
        RECT 82.020 70.130 82.680 70.150 ;
        RECT 85.030 70.130 86.830 70.280 ;
        RECT 87.210 70.170 87.540 74.350 ;
        RECT 89.720 74.890 90.040 77.340 ;
        RECT 90.750 76.740 95.800 77.630 ;
        RECT 90.770 76.710 95.770 76.740 ;
        RECT 96.710 76.680 97.030 77.660 ;
        RECT 97.770 77.620 102.770 77.650 ;
        RECT 97.740 76.920 102.790 77.620 ;
        RECT 104.040 77.590 104.620 79.240 ;
        RECT 113.340 79.110 115.195 79.240 ;
        RECT 106.230 78.660 107.150 78.730 ;
        RECT 106.230 78.430 111.250 78.660 ;
        RECT 97.750 76.730 102.790 76.920 ;
        RECT 97.770 76.710 102.770 76.730 ;
        RECT 95.970 76.660 97.030 76.680 ;
        RECT 90.380 75.700 90.610 76.660 ;
        RECT 95.930 75.700 97.030 76.660 ;
        RECT 95.970 75.680 97.030 75.700 ;
        RECT 90.770 75.420 95.770 75.650 ;
        RECT 93.080 75.090 94.810 75.420 ;
        RECT 89.720 73.260 90.050 74.890 ;
        RECT 89.720 72.680 90.040 73.260 ;
        RECT 96.710 73.230 97.030 75.680 ;
        RECT 97.330 74.750 97.610 76.690 ;
        RECT 100.290 75.650 101.810 75.740 ;
        RECT 102.930 75.700 103.160 76.660 ;
        RECT 97.770 75.420 102.770 75.650 ;
        RECT 100.290 75.220 101.810 75.420 ;
        RECT 97.220 73.720 97.610 74.750 ;
        RECT 105.790 74.250 106.070 78.400 ;
        RECT 106.230 78.310 107.150 78.430 ;
        RECT 111.420 78.380 111.810 78.400 ;
        RECT 110.150 77.370 111.250 77.570 ;
        RECT 111.390 77.420 111.810 78.380 ;
        RECT 113.340 77.840 115.085 79.110 ;
        RECT 115.465 78.950 115.985 80.270 ;
        RECT 116.255 79.110 116.485 80.110 ;
        RECT 116.735 78.950 117.255 80.270 ;
        RECT 117.645 80.110 119.385 80.680 ;
        RECT 117.545 79.110 119.385 80.110 ;
        RECT 115.245 78.720 116.205 78.950 ;
        RECT 116.535 78.720 117.495 78.950 ;
        RECT 116.595 78.440 117.435 78.720 ;
        RECT 117.645 78.680 119.385 79.110 ;
        RECT 117.645 78.660 119.365 78.680 ;
        RECT 119.665 78.475 120.185 80.885 ;
        RECT 120.445 78.680 120.675 80.680 ;
        RECT 120.995 78.475 121.515 80.885 ;
        RECT 121.875 80.680 123.765 82.295 ;
        RECT 121.735 80.295 123.765 80.680 ;
        RECT 121.735 78.680 123.625 80.295 ;
        RECT 123.985 80.090 124.505 82.500 ;
        RECT 124.825 80.295 125.055 82.295 ;
        RECT 125.315 80.090 125.835 82.500 ;
        RECT 126.135 82.295 127.855 82.315 ;
        RECT 126.115 81.865 127.855 82.295 ;
        RECT 128.065 82.255 128.905 82.535 ;
        RECT 128.005 82.025 128.965 82.255 ;
        RECT 129.295 82.025 130.255 82.255 ;
        RECT 126.115 80.865 127.955 81.865 ;
        RECT 126.115 80.295 127.855 80.865 ;
        RECT 128.245 80.705 128.765 82.025 ;
        RECT 129.015 80.865 129.245 81.865 ;
        RECT 129.515 80.705 130.035 82.025 ;
        RECT 130.415 81.865 130.955 83.125 ;
        RECT 130.305 80.865 130.955 81.865 ;
        RECT 128.005 80.475 128.965 80.705 ;
        RECT 129.295 80.475 130.255 80.705 ;
        RECT 130.415 80.335 130.955 80.865 ;
        RECT 126.135 80.275 127.855 80.295 ;
        RECT 123.815 79.860 124.775 80.090 ;
        RECT 125.105 79.860 126.065 80.090 ;
        RECT 126.825 79.865 127.515 80.275 ;
        RECT 130.405 80.215 130.955 80.335 ;
        RECT 126.815 79.245 127.515 79.865 ;
        RECT 119.435 78.440 120.395 78.475 ;
        RECT 116.595 78.270 120.395 78.440 ;
        RECT 113.340 77.570 115.105 77.840 ;
        RECT 106.230 77.140 111.250 77.370 ;
        RECT 110.150 76.900 111.250 77.140 ;
        RECT 111.420 77.090 111.810 77.420 ;
        RECT 106.230 76.080 107.150 76.150 ;
        RECT 111.390 76.130 111.810 77.090 ;
        RECT 113.170 76.910 115.105 77.570 ;
        RECT 106.230 75.850 111.240 76.080 ;
        RECT 106.230 75.730 107.150 75.850 ;
        RECT 111.420 75.800 111.810 76.130 ;
        RECT 110.230 74.800 111.170 74.870 ;
        RECT 111.390 74.840 111.810 75.800 ;
        RECT 106.280 74.790 111.240 74.800 ;
        RECT 106.230 74.570 111.240 74.790 ;
        RECT 106.230 74.560 111.230 74.570 ;
        RECT 110.230 74.480 111.170 74.560 ;
        RECT 111.420 74.510 111.810 74.840 ;
        RECT 111.390 74.250 111.810 74.510 ;
        RECT 105.790 73.800 106.160 74.250 ;
        RECT 111.340 73.800 111.810 74.250 ;
        RECT 90.760 72.940 92.650 73.060 ;
        RECT 90.760 72.710 95.770 72.940 ;
        RECT 89.720 72.660 90.580 72.680 ;
        RECT 89.720 71.700 90.610 72.660 ;
        RECT 90.760 72.440 92.650 72.710 ;
        RECT 96.700 72.700 97.040 73.230 ;
        RECT 98.190 72.940 99.710 73.070 ;
        RECT 97.770 72.710 102.770 72.940 ;
        RECT 95.930 71.700 96.160 72.660 ;
        RECT 89.720 71.670 90.580 71.700 ;
        RECT 96.700 71.650 97.610 72.700 ;
        RECT 98.190 72.550 99.710 72.710 ;
        RECT 102.930 71.700 103.160 72.660 ;
        RECT 90.770 71.630 95.770 71.650 ;
        RECT 90.740 70.740 95.790 71.630 ;
        RECT 90.770 70.710 95.770 70.740 ;
        RECT 96.700 70.700 97.040 71.650 ;
        RECT 97.770 71.630 102.770 71.650 ;
        RECT 97.770 71.420 102.800 71.630 ;
        RECT 97.980 70.940 102.800 71.420 ;
        RECT 97.770 70.740 102.800 70.940 ;
        RECT 95.960 70.660 97.040 70.700 ;
        RECT 82.020 69.900 87.050 70.130 ;
        RECT 82.020 69.680 82.680 69.900 ;
        RECT 85.030 69.460 86.830 69.900 ;
        RECT 90.380 69.700 90.610 70.660 ;
        RECT 90.770 69.420 95.770 69.650 ;
        RECT 93.080 69.080 94.810 69.420 ;
        RECT 95.930 69.260 97.040 70.660 ;
        RECT 97.270 69.680 97.620 70.720 ;
        RECT 97.770 70.710 102.770 70.740 ;
        RECT 100.260 69.650 101.780 69.750 ;
        RECT 102.930 69.700 103.160 70.660 ;
        RECT 97.770 69.420 102.770 69.650 ;
        RECT 100.260 69.230 101.780 69.420 ;
        RECT 105.790 68.390 106.070 73.800 ;
        RECT 106.230 73.500 107.160 73.560 ;
        RECT 111.390 73.550 111.810 73.800 ;
        RECT 106.230 73.270 111.240 73.500 ;
        RECT 106.230 73.180 107.160 73.270 ;
        RECT 111.420 73.220 111.810 73.550 ;
        RECT 110.230 72.220 111.180 72.310 ;
        RECT 111.390 72.260 111.810 73.220 ;
        RECT 106.280 72.210 111.240 72.220 ;
        RECT 106.230 71.990 111.240 72.210 ;
        RECT 106.230 71.980 111.230 71.990 ;
        RECT 110.230 71.930 111.180 71.980 ;
        RECT 111.420 71.930 111.810 72.260 ;
        RECT 106.230 70.930 107.150 71.000 ;
        RECT 111.390 70.970 111.810 71.930 ;
        RECT 106.230 70.700 111.240 70.930 ;
        RECT 106.230 70.690 111.230 70.700 ;
        RECT 106.230 70.630 107.150 70.690 ;
        RECT 111.420 70.640 111.810 70.970 ;
        RECT 110.230 69.630 111.180 69.710 ;
        RECT 111.390 69.680 111.810 70.640 ;
        RECT 106.230 69.400 111.240 69.630 ;
        RECT 110.230 69.310 111.180 69.400 ;
        RECT 111.420 69.350 111.810 69.680 ;
        RECT 113.340 76.700 115.105 76.910 ;
        RECT 117.985 77.670 118.675 78.270 ;
        RECT 119.435 78.245 120.395 78.270 ;
        RECT 120.725 78.245 121.685 78.475 ;
        RECT 121.875 78.245 123.625 78.680 ;
        RECT 123.815 78.450 124.775 78.680 ;
        RECT 125.105 78.655 126.065 78.680 ;
        RECT 126.825 78.655 127.515 79.245 ;
        RECT 130.395 79.075 130.955 80.215 ;
        RECT 125.105 78.485 128.905 78.655 ;
        RECT 125.105 78.450 126.065 78.485 ;
        RECT 117.985 77.050 118.685 77.670 ;
        RECT 113.340 76.580 115.095 76.700 ;
        RECT 117.985 76.640 118.675 77.050 ;
        RECT 119.435 76.825 120.395 77.055 ;
        RECT 120.725 76.825 121.685 77.055 ;
        RECT 117.645 76.620 119.365 76.640 ;
        RECT 113.340 76.050 115.085 76.580 ;
        RECT 115.245 76.210 116.205 76.440 ;
        RECT 116.535 76.210 117.495 76.440 ;
        RECT 113.340 75.050 115.195 76.050 ;
        RECT 113.340 73.210 115.085 75.050 ;
        RECT 115.465 74.890 115.985 76.210 ;
        RECT 116.255 75.050 116.485 76.050 ;
        RECT 116.735 74.890 117.255 76.210 ;
        RECT 117.645 76.050 119.385 76.620 ;
        RECT 117.545 75.050 119.385 76.050 ;
        RECT 115.245 74.660 116.205 74.890 ;
        RECT 116.535 74.660 117.495 74.890 ;
        RECT 116.595 74.380 117.435 74.660 ;
        RECT 117.645 74.620 119.385 75.050 ;
        RECT 117.645 74.600 119.365 74.620 ;
        RECT 119.665 74.415 120.185 76.825 ;
        RECT 120.445 74.620 120.675 76.620 ;
        RECT 120.995 74.415 121.515 76.825 ;
        RECT 121.875 76.620 123.765 78.245 ;
        RECT 121.735 76.245 123.765 76.620 ;
        RECT 121.735 74.620 123.625 76.245 ;
        RECT 123.985 76.040 124.505 78.450 ;
        RECT 124.825 76.245 125.055 78.245 ;
        RECT 125.315 76.040 125.835 78.450 ;
        RECT 126.135 78.245 127.855 78.265 ;
        RECT 126.115 77.815 127.855 78.245 ;
        RECT 128.065 78.205 128.905 78.485 ;
        RECT 128.005 77.975 128.965 78.205 ;
        RECT 129.295 77.975 130.255 78.205 ;
        RECT 126.115 76.815 127.955 77.815 ;
        RECT 126.115 76.245 127.855 76.815 ;
        RECT 128.245 76.655 128.765 77.975 ;
        RECT 129.015 76.815 129.245 77.815 ;
        RECT 129.515 76.655 130.035 77.975 ;
        RECT 130.415 77.815 130.955 79.075 ;
        RECT 130.305 76.815 130.955 77.815 ;
        RECT 128.005 76.425 128.965 76.655 ;
        RECT 129.295 76.425 130.255 76.655 ;
        RECT 130.415 76.285 130.955 76.815 ;
        RECT 126.135 76.225 127.855 76.245 ;
        RECT 123.815 75.810 124.775 76.040 ;
        RECT 125.105 75.810 126.065 76.040 ;
        RECT 126.825 75.815 127.515 76.225 ;
        RECT 130.405 76.165 130.955 76.285 ;
        RECT 126.815 75.195 127.515 75.815 ;
        RECT 119.435 74.380 120.395 74.415 ;
        RECT 116.595 74.210 120.395 74.380 ;
        RECT 117.985 73.430 118.675 74.210 ;
        RECT 119.435 74.185 120.395 74.210 ;
        RECT 120.725 74.185 121.685 74.415 ;
        RECT 121.875 74.195 123.625 74.620 ;
        RECT 123.815 74.400 124.775 74.630 ;
        RECT 125.105 74.605 126.065 74.630 ;
        RECT 126.825 74.605 127.515 75.195 ;
        RECT 130.395 75.025 130.955 76.165 ;
        RECT 125.105 74.435 128.905 74.605 ;
        RECT 125.105 74.400 126.065 74.435 ;
        RECT 121.875 73.210 123.765 74.195 ;
        RECT 113.340 73.180 114.710 73.210 ;
        RECT 106.220 68.340 107.150 68.390 ;
        RECT 111.380 68.380 112.530 69.350 ;
        RECT 106.220 68.110 111.230 68.340 ;
        RECT 106.220 68.070 107.150 68.110 ;
        RECT 80.240 67.250 81.470 68.050 ;
        RECT 71.770 66.590 96.350 67.250 ;
        RECT 113.340 67.160 113.960 73.180 ;
        RECT 71.770 66.260 95.000 66.590 ;
        RECT 95.570 66.530 96.350 66.590 ;
        RECT 103.305 66.530 105.730 66.650 ;
        RECT 95.570 66.330 103.095 66.530 ;
        RECT 95.595 66.300 103.095 66.330 ;
        RECT 103.305 66.440 105.755 66.530 ;
        RECT 103.305 66.420 104.090 66.440 ;
        RECT 71.770 65.970 72.340 66.260 ;
        RECT 71.770 65.020 72.510 65.970 ;
        RECT 94.510 65.420 95.000 66.260 ;
        RECT 103.305 66.250 103.535 66.420 ;
        RECT 103.710 66.390 104.090 66.420 ;
        RECT 104.755 66.300 105.755 66.440 ;
        RECT 107.880 66.470 113.960 67.160 ;
        RECT 107.880 66.320 112.900 66.470 ;
        RECT 113.450 66.320 113.960 66.470 ;
        RECT 107.900 66.295 112.900 66.320 ;
        RECT 95.160 66.040 95.390 66.250 ;
        RECT 95.160 65.790 96.170 66.040 ;
        RECT 95.190 65.740 96.170 65.790 ;
        RECT 103.300 65.740 103.535 66.250 ;
        RECT 104.165 65.740 104.555 66.250 ;
        RECT 105.950 65.740 106.240 66.270 ;
        RECT 95.190 65.700 103.535 65.740 ;
        RECT 95.595 65.510 103.535 65.700 ;
        RECT 94.510 65.210 95.410 65.420 ;
        RECT 71.770 64.740 72.710 65.020 ;
        RECT 94.510 64.860 103.040 65.210 ;
        RECT 71.770 44.150 72.510 64.740 ;
        RECT 94.510 60.020 95.410 64.860 ;
        RECT 96.150 64.170 97.060 64.490 ;
        RECT 97.420 64.460 103.040 64.860 ;
        RECT 103.840 64.980 106.240 65.740 ;
        RECT 107.510 65.990 107.740 66.245 ;
        RECT 113.060 65.990 113.290 66.245 ;
        RECT 107.510 65.650 113.290 65.990 ;
        RECT 107.510 65.285 107.740 65.650 ;
        RECT 113.060 65.285 113.290 65.650 ;
        RECT 107.900 65.220 112.900 65.235 ;
        RECT 107.900 65.010 112.930 65.220 ;
        RECT 103.840 64.870 107.630 64.980 ;
        RECT 107.895 64.870 112.930 65.010 ;
        RECT 103.840 64.740 112.930 64.870 ;
        RECT 103.840 64.730 106.240 64.740 ;
        RECT 96.130 64.155 103.100 64.170 ;
        RECT 96.090 63.925 103.100 64.155 ;
        RECT 103.840 64.080 104.010 64.730 ;
        RECT 107.410 64.680 108.110 64.740 ;
        RECT 95.610 61.470 95.900 63.900 ;
        RECT 96.130 63.830 103.100 63.925 ;
        RECT 103.290 63.780 104.010 64.080 ;
        RECT 96.080 62.010 103.120 63.370 ;
        RECT 103.290 62.860 103.590 63.780 ;
        RECT 96.090 61.995 103.090 62.010 ;
        RECT 96.150 61.500 97.060 61.520 ;
        RECT 96.130 61.435 103.100 61.500 ;
        RECT 103.290 61.470 103.580 62.860 ;
        RECT 96.090 61.205 103.100 61.435 ;
        RECT 96.130 61.160 103.100 61.205 ;
        RECT 96.150 60.960 97.060 61.160 ;
        RECT 94.510 59.190 99.010 60.020 ;
        RECT 94.860 58.600 99.010 59.190 ;
        RECT 103.220 59.130 104.480 59.190 ;
        RECT 98.590 46.380 99.010 58.600 ;
        RECT 99.150 47.970 99.450 58.920 ;
        RECT 99.640 58.900 104.640 59.130 ;
        RECT 103.220 58.840 104.480 58.900 ;
        RECT 99.770 58.340 100.890 58.360 ;
        RECT 99.640 58.110 104.640 58.340 ;
        RECT 99.770 58.010 100.890 58.110 ;
        RECT 104.800 57.970 105.980 59.470 ;
        RECT 106.670 59.150 107.540 62.650 ;
        RECT 113.470 60.020 113.960 66.320 ;
        RECT 122.725 72.195 123.765 73.210 ;
        RECT 122.725 70.110 123.625 72.195 ;
        RECT 123.985 71.990 124.505 74.400 ;
        RECT 124.825 72.195 125.055 74.195 ;
        RECT 125.315 71.990 125.835 74.400 ;
        RECT 126.135 74.195 127.855 74.215 ;
        RECT 126.115 73.765 127.855 74.195 ;
        RECT 128.065 74.155 128.905 74.435 ;
        RECT 128.005 73.925 128.965 74.155 ;
        RECT 129.295 73.925 130.255 74.155 ;
        RECT 126.115 72.765 127.955 73.765 ;
        RECT 126.115 72.195 127.855 72.765 ;
        RECT 128.245 72.605 128.765 73.925 ;
        RECT 129.015 72.765 129.245 73.765 ;
        RECT 129.515 72.605 130.035 73.925 ;
        RECT 130.415 73.765 130.955 75.025 ;
        RECT 130.305 72.765 130.955 73.765 ;
        RECT 128.005 72.375 128.965 72.605 ;
        RECT 129.295 72.375 130.255 72.605 ;
        RECT 130.415 72.235 130.955 72.765 ;
        RECT 126.135 72.175 127.855 72.195 ;
        RECT 123.815 71.760 124.775 71.990 ;
        RECT 125.105 71.760 126.065 71.990 ;
        RECT 126.825 71.765 127.515 72.175 ;
        RECT 130.405 72.115 130.955 72.235 ;
        RECT 126.815 71.145 127.515 71.765 ;
        RECT 123.815 70.315 124.775 70.545 ;
        RECT 125.105 70.520 126.065 70.545 ;
        RECT 126.825 70.520 127.515 71.145 ;
        RECT 130.395 70.975 130.955 72.115 ;
        RECT 125.105 70.350 128.905 70.520 ;
        RECT 125.105 70.315 126.065 70.350 ;
        RECT 122.725 68.110 123.765 70.110 ;
        RECT 122.725 65.985 123.625 68.110 ;
        RECT 123.985 67.905 124.505 70.315 ;
        RECT 124.825 68.110 125.055 70.110 ;
        RECT 125.315 67.905 125.835 70.315 ;
        RECT 126.135 70.110 127.855 70.130 ;
        RECT 126.115 69.680 127.855 70.110 ;
        RECT 128.065 70.070 128.905 70.350 ;
        RECT 128.005 69.840 128.965 70.070 ;
        RECT 129.295 69.840 130.255 70.070 ;
        RECT 126.115 68.680 127.955 69.680 ;
        RECT 126.115 68.110 127.855 68.680 ;
        RECT 128.245 68.520 128.765 69.840 ;
        RECT 129.015 68.680 129.245 69.680 ;
        RECT 129.515 68.520 130.035 69.840 ;
        RECT 130.415 69.680 130.955 70.975 ;
        RECT 130.305 68.680 130.955 69.680 ;
        RECT 128.005 68.290 128.965 68.520 ;
        RECT 129.295 68.290 130.255 68.520 ;
        RECT 130.415 68.150 130.955 68.680 ;
        RECT 126.135 68.090 127.855 68.110 ;
        RECT 123.815 67.675 124.775 67.905 ;
        RECT 125.105 67.675 126.065 67.905 ;
        RECT 126.825 67.680 127.515 68.090 ;
        RECT 130.405 68.030 130.955 68.150 ;
        RECT 126.815 67.060 127.515 67.680 ;
        RECT 123.815 66.190 124.775 66.420 ;
        RECT 125.105 66.395 126.065 66.420 ;
        RECT 126.825 66.395 127.515 67.060 ;
        RECT 130.395 66.890 130.955 68.030 ;
        RECT 125.105 66.225 128.905 66.395 ;
        RECT 125.105 66.190 126.065 66.225 ;
        RECT 122.725 63.985 123.765 65.985 ;
        RECT 122.725 62.390 123.625 63.985 ;
        RECT 123.985 63.780 124.505 66.190 ;
        RECT 124.825 63.985 125.055 65.985 ;
        RECT 125.315 63.780 125.835 66.190 ;
        RECT 126.135 65.985 127.855 66.005 ;
        RECT 126.115 65.555 127.855 65.985 ;
        RECT 128.065 65.945 128.905 66.225 ;
        RECT 128.005 65.715 128.965 65.945 ;
        RECT 129.295 65.715 130.255 65.945 ;
        RECT 126.115 64.555 127.955 65.555 ;
        RECT 126.115 63.985 127.855 64.555 ;
        RECT 128.245 64.395 128.765 65.715 ;
        RECT 129.015 64.555 129.245 65.555 ;
        RECT 129.515 64.395 130.035 65.715 ;
        RECT 130.415 65.555 130.955 66.890 ;
        RECT 130.305 64.555 130.955 65.555 ;
        RECT 128.005 64.165 128.965 64.395 ;
        RECT 129.295 64.165 130.255 64.395 ;
        RECT 130.415 64.025 130.955 64.555 ;
        RECT 126.135 63.965 127.855 63.985 ;
        RECT 123.815 63.550 124.775 63.780 ;
        RECT 125.105 63.550 126.065 63.780 ;
        RECT 126.825 63.555 127.515 63.965 ;
        RECT 130.405 63.905 130.955 64.025 ;
        RECT 126.815 62.935 127.515 63.555 ;
        RECT 107.840 59.310 112.680 59.370 ;
        RECT 104.800 57.960 105.760 57.970 ;
        RECT 103.230 57.550 104.490 57.630 ;
        RECT 99.640 57.320 104.640 57.550 ;
        RECT 103.230 57.270 104.490 57.320 ;
        RECT 99.760 56.760 100.880 56.790 ;
        RECT 99.640 56.530 104.640 56.760 ;
        RECT 99.760 56.450 100.880 56.530 ;
        RECT 103.220 55.970 104.480 56.040 ;
        RECT 99.640 55.740 104.640 55.970 ;
        RECT 103.220 55.680 104.480 55.740 ;
        RECT 99.790 55.180 100.880 55.210 ;
        RECT 99.640 54.950 104.640 55.180 ;
        RECT 99.790 54.850 100.880 54.950 ;
        RECT 103.220 54.390 104.480 54.440 ;
        RECT 99.640 54.160 104.640 54.390 ;
        RECT 103.220 54.080 104.480 54.160 ;
        RECT 99.720 53.600 100.880 53.670 ;
        RECT 99.640 53.370 104.640 53.600 ;
        RECT 99.720 53.250 100.880 53.370 ;
        RECT 103.220 52.810 104.480 52.840 ;
        RECT 99.640 52.580 104.640 52.810 ;
        RECT 103.220 52.500 104.480 52.580 ;
        RECT 99.730 52.020 100.880 52.120 ;
        RECT 99.640 51.790 104.640 52.020 ;
        RECT 99.730 51.660 100.880 51.790 ;
        RECT 103.220 51.230 104.480 51.310 ;
        RECT 99.640 51.000 104.640 51.230 ;
        RECT 103.220 50.970 104.480 51.000 ;
        RECT 99.780 50.440 100.880 50.520 ;
        RECT 99.640 50.210 104.640 50.440 ;
        RECT 99.780 50.100 100.880 50.210 ;
        RECT 103.220 49.650 104.480 49.680 ;
        RECT 99.640 49.420 104.640 49.650 ;
        RECT 103.220 49.340 104.480 49.420 ;
        RECT 99.800 48.860 100.880 48.950 ;
        RECT 99.640 48.630 104.640 48.860 ;
        RECT 99.800 48.520 100.880 48.630 ;
        RECT 103.220 48.070 104.480 48.100 ;
        RECT 99.640 47.840 104.640 48.070 ;
        RECT 104.800 47.950 105.100 57.960 ;
        RECT 106.650 57.780 107.540 59.150 ;
        RECT 107.700 59.080 112.700 59.310 ;
        RECT 107.840 59.030 112.680 59.080 ;
        RECT 112.870 59.030 113.180 59.080 ;
        RECT 107.780 58.600 108.990 58.610 ;
        RECT 107.780 58.520 109.000 58.600 ;
        RECT 112.860 58.570 113.180 59.030 ;
        RECT 107.700 58.290 112.700 58.520 ;
        RECT 107.780 58.240 109.000 58.290 ;
        RECT 112.870 58.240 113.180 58.570 ;
        RECT 107.780 58.210 108.990 58.240 ;
        RECT 106.650 57.450 107.520 57.780 ;
        RECT 111.230 57.730 112.510 57.820 ;
        RECT 112.860 57.780 113.180 58.240 ;
        RECT 107.700 57.500 112.700 57.730 ;
        RECT 106.650 56.990 107.540 57.450 ;
        RECT 111.230 57.420 112.510 57.500 ;
        RECT 112.870 57.450 113.180 57.780 ;
        RECT 112.860 56.990 113.180 57.450 ;
        RECT 106.650 56.660 107.520 56.990 ;
        RECT 107.780 56.940 109.000 56.980 ;
        RECT 107.700 56.710 112.700 56.940 ;
        RECT 106.650 56.200 107.540 56.660 ;
        RECT 107.780 56.620 109.000 56.710 ;
        RECT 112.870 56.660 113.180 56.990 ;
        RECT 106.650 55.870 107.520 56.200 ;
        RECT 111.230 56.150 112.510 56.220 ;
        RECT 112.860 56.200 113.180 56.660 ;
        RECT 107.700 55.920 112.700 56.150 ;
        RECT 106.650 55.410 107.540 55.870 ;
        RECT 111.230 55.820 112.510 55.920 ;
        RECT 112.870 55.870 113.180 56.200 ;
        RECT 112.860 55.410 113.180 55.870 ;
        RECT 106.650 55.080 107.520 55.410 ;
        RECT 107.760 55.360 109.000 55.410 ;
        RECT 107.700 55.130 112.700 55.360 ;
        RECT 106.650 54.620 107.540 55.080 ;
        RECT 107.760 55.060 109.000 55.130 ;
        RECT 112.870 55.080 113.180 55.410 ;
        RECT 106.650 54.290 107.520 54.620 ;
        RECT 111.220 54.570 112.550 54.630 ;
        RECT 112.860 54.620 113.180 55.080 ;
        RECT 107.700 54.340 112.700 54.570 ;
        RECT 106.650 53.830 107.540 54.290 ;
        RECT 111.220 54.230 112.550 54.340 ;
        RECT 112.870 54.290 113.180 54.620 ;
        RECT 112.860 53.830 113.180 54.290 ;
        RECT 106.650 53.500 107.520 53.830 ;
        RECT 107.860 53.780 109.010 53.800 ;
        RECT 107.700 53.550 112.700 53.780 ;
        RECT 106.650 53.040 107.540 53.500 ;
        RECT 107.860 53.440 109.010 53.550 ;
        RECT 112.870 53.500 113.180 53.830 ;
        RECT 106.650 52.710 107.520 53.040 ;
        RECT 111.240 52.990 112.500 53.100 ;
        RECT 112.860 53.040 113.180 53.500 ;
        RECT 107.700 52.760 112.700 52.990 ;
        RECT 106.650 52.250 107.540 52.710 ;
        RECT 111.240 52.650 112.500 52.760 ;
        RECT 112.870 52.710 113.180 53.040 ;
        RECT 112.860 52.250 113.180 52.710 ;
        RECT 106.650 51.920 107.520 52.250 ;
        RECT 107.880 52.200 109.000 52.240 ;
        RECT 107.700 51.970 112.700 52.200 ;
        RECT 106.650 51.460 107.540 51.920 ;
        RECT 107.880 51.900 109.000 51.970 ;
        RECT 112.870 51.920 113.180 52.250 ;
        RECT 112.860 51.460 113.180 51.920 ;
        RECT 106.650 51.130 107.520 51.460 ;
        RECT 111.230 51.410 112.490 51.450 ;
        RECT 107.700 51.180 112.700 51.410 ;
        RECT 106.650 50.670 107.540 51.130 ;
        RECT 111.230 51.100 112.490 51.180 ;
        RECT 112.870 51.130 113.180 51.460 ;
        RECT 112.860 50.670 113.180 51.130 ;
        RECT 106.650 50.340 107.520 50.670 ;
        RECT 107.850 50.620 109.000 50.650 ;
        RECT 107.700 50.390 112.700 50.620 ;
        RECT 106.650 49.880 107.540 50.340 ;
        RECT 107.850 50.300 109.000 50.390 ;
        RECT 112.870 50.340 113.180 50.670 ;
        RECT 106.650 49.550 107.520 49.880 ;
        RECT 111.230 49.830 112.500 49.890 ;
        RECT 112.860 49.880 113.180 50.340 ;
        RECT 107.700 49.600 112.700 49.830 ;
        RECT 106.650 49.090 107.540 49.550 ;
        RECT 111.230 49.530 112.500 49.600 ;
        RECT 112.870 49.550 113.180 49.880 ;
        RECT 112.860 49.090 113.180 49.550 ;
        RECT 106.650 48.760 107.520 49.090 ;
        RECT 107.810 49.040 109.000 49.080 ;
        RECT 107.700 48.810 112.700 49.040 ;
        RECT 106.650 48.300 107.540 48.760 ;
        RECT 107.810 48.720 109.000 48.810 ;
        RECT 112.870 48.760 113.180 49.090 ;
        RECT 112.860 48.300 113.180 48.760 ;
        RECT 106.650 47.970 107.520 48.300 ;
        RECT 111.230 48.250 112.510 48.290 ;
        RECT 107.700 48.020 112.700 48.250 ;
        RECT 103.220 47.750 104.480 47.840 ;
        RECT 106.650 47.510 107.540 47.970 ;
        RECT 111.230 47.930 112.510 48.020 ;
        RECT 112.870 47.970 113.180 48.300 ;
        RECT 112.860 47.510 113.180 47.970 ;
        RECT 106.650 47.180 107.520 47.510 ;
        RECT 107.850 47.460 109.000 47.490 ;
        RECT 107.700 47.230 112.700 47.460 ;
        RECT 106.650 46.720 107.540 47.180 ;
        RECT 107.850 47.140 109.000 47.230 ;
        RECT 112.870 47.180 113.180 47.510 ;
        RECT 112.860 46.720 113.180 47.180 ;
        RECT 106.650 46.390 107.520 46.720 ;
        RECT 111.230 46.670 112.500 46.700 ;
        RECT 107.700 46.440 112.700 46.670 ;
        RECT 106.650 45.930 107.540 46.390 ;
        RECT 111.230 46.310 112.500 46.440 ;
        RECT 112.870 46.390 113.180 46.720 ;
        RECT 107.810 45.930 108.990 45.980 ;
        RECT 112.860 45.930 113.180 46.390 ;
        RECT 106.650 45.600 107.520 45.930 ;
        RECT 107.810 45.880 109.000 45.930 ;
        RECT 107.700 45.650 112.700 45.880 ;
        RECT 106.650 45.140 107.540 45.600 ;
        RECT 107.810 45.590 109.000 45.650 ;
        RECT 112.870 45.600 113.180 45.930 ;
        RECT 107.810 45.560 108.990 45.590 ;
        RECT 112.860 45.140 113.180 45.600 ;
        RECT 106.650 44.810 107.520 45.140 ;
        RECT 111.220 45.090 112.500 45.120 ;
        RECT 107.700 44.860 112.700 45.090 ;
        RECT 106.650 44.350 107.540 44.810 ;
        RECT 111.220 44.760 112.500 44.860 ;
        RECT 112.870 44.810 113.180 45.140 ;
        RECT 112.860 44.350 113.180 44.810 ;
        RECT 106.650 44.250 107.520 44.350 ;
        RECT 107.810 44.300 109.010 44.330 ;
        RECT 70.530 43.210 70.950 43.680 ;
        RECT 106.650 42.480 107.500 44.250 ;
        RECT 107.700 44.070 112.700 44.300 ;
        RECT 112.870 44.240 113.180 44.350 ;
        RECT 107.810 43.970 109.010 44.070 ;
        RECT 113.350 43.530 113.960 60.020 ;
        RECT 121.090 61.430 123.625 62.390 ;
        RECT 126.820 62.620 127.510 62.935 ;
        RECT 130.395 62.765 130.955 63.905 ;
        RECT 126.820 62.130 127.515 62.620 ;
        RECT 123.815 61.635 124.775 61.865 ;
        RECT 125.105 61.840 126.065 61.865 ;
        RECT 126.825 61.840 127.515 62.130 ;
        RECT 125.105 61.670 128.905 61.840 ;
        RECT 125.105 61.635 126.065 61.670 ;
        RECT 121.090 59.430 123.765 61.430 ;
        RECT 121.090 58.600 123.625 59.430 ;
        RECT 123.985 59.225 124.505 61.635 ;
        RECT 124.825 59.430 125.055 61.430 ;
        RECT 125.315 59.225 125.835 61.635 ;
        RECT 126.135 61.430 127.855 61.450 ;
        RECT 126.115 61.000 127.855 61.430 ;
        RECT 128.065 61.390 128.905 61.670 ;
        RECT 128.005 61.160 128.965 61.390 ;
        RECT 129.295 61.160 130.255 61.390 ;
        RECT 126.115 60.000 127.955 61.000 ;
        RECT 126.115 59.430 127.855 60.000 ;
        RECT 128.245 59.840 128.765 61.160 ;
        RECT 129.015 60.000 129.245 61.000 ;
        RECT 129.515 59.840 130.035 61.160 ;
        RECT 130.415 61.000 130.955 62.765 ;
        RECT 130.305 60.000 130.955 61.000 ;
        RECT 128.005 59.610 128.965 59.840 ;
        RECT 129.295 59.610 130.255 59.840 ;
        RECT 130.415 59.470 130.955 60.000 ;
        RECT 126.135 59.410 127.855 59.430 ;
        RECT 123.815 58.995 124.775 59.225 ;
        RECT 125.105 58.995 126.065 59.225 ;
        RECT 121.090 58.420 123.620 58.600 ;
        RECT 121.090 58.210 123.625 58.420 ;
        RECT 106.100 41.050 107.610 42.480 ;
        RECT 122.450 39.110 123.420 58.210 ;
        RECT 126.660 55.180 127.660 59.410 ;
        RECT 130.405 59.350 130.955 59.470 ;
        RECT 130.395 58.210 130.955 59.350 ;
        RECT 126.020 53.440 128.170 55.180 ;
        RECT 27.920 36.910 30.100 38.880 ;
        RECT 121.860 36.000 123.930 39.110 ;
        RECT 122.450 35.860 123.420 36.000 ;
      LAYER via ;
        RECT 26.690 197.680 28.310 198.820 ;
        RECT 71.850 196.940 73.110 199.640 ;
        RECT 130.250 196.900 131.060 199.620 ;
        RECT 106.460 195.730 107.380 196.330 ;
        RECT 30.850 191.880 32.260 192.700 ;
        RECT 62.430 191.630 69.580 193.040 ;
        RECT 107.890 194.330 108.960 194.610 ;
        RECT 111.280 193.530 112.460 193.820 ;
        RECT 107.890 192.720 108.950 193.000 ;
        RECT 63.610 185.960 65.950 189.220 ;
        RECT 28.850 182.230 29.250 183.000 ;
        RECT 27.470 173.340 27.940 174.480 ;
        RECT 18.460 152.970 19.050 154.890 ;
        RECT 34.110 182.510 35.010 182.810 ;
        RECT 35.790 182.550 36.080 182.830 ;
        RECT 29.550 180.900 29.820 181.380 ;
        RECT 35.240 180.870 35.510 181.350 ;
        RECT 34.150 178.090 34.940 178.440 ;
        RECT 34.250 177.020 34.990 177.480 ;
        RECT 34.180 173.590 34.970 173.900 ;
        RECT 35.800 178.100 36.090 178.380 ;
        RECT 36.740 181.760 37.210 182.130 ;
        RECT 36.750 177.070 37.210 177.630 ;
        RECT 36.760 172.680 37.250 173.140 ;
        RECT 37.850 182.540 38.140 182.820 ;
        RECT 37.850 178.010 38.140 178.290 ;
        RECT 37.840 173.520 38.130 173.800 ;
        RECT 39.240 182.510 39.810 182.870 ;
        RECT 39.060 181.630 39.560 181.990 ;
        RECT 38.540 180.870 38.810 181.350 ;
        RECT 47.790 181.580 49.510 181.860 ;
        RECT 44.220 180.890 44.490 181.370 ;
        RECT 55.280 181.540 56.610 181.850 ;
        RECT 46.070 180.470 46.850 181.380 ;
        RECT 44.250 178.530 44.740 179.300 ;
        RECT 39.220 177.910 39.790 178.370 ;
        RECT 39.130 173.540 39.820 173.930 ;
        RECT 48.060 179.820 49.210 180.380 ;
        RECT 63.280 181.290 64.050 181.550 ;
        RECT 58.440 179.770 59.590 180.330 ;
        RECT 50.160 178.050 51.680 178.390 ;
        RECT 46.740 176.630 47.010 177.540 ;
        RECT 57.380 178.210 58.710 178.520 ;
        RECT 54.300 176.660 54.570 177.500 ;
        RECT 67.260 179.900 68.150 180.380 ;
        RECT 70.250 179.880 70.640 180.360 ;
        RECT 63.280 178.680 64.100 178.980 ;
        RECT 67.280 177.420 68.080 177.690 ;
        RECT 62.820 176.720 63.080 177.080 ;
        RECT 68.350 176.730 68.610 177.090 ;
        RECT 47.780 175.560 49.610 175.890 ;
        RECT 55.280 175.490 56.610 175.800 ;
        RECT 48.060 173.810 49.210 174.370 ;
        RECT 58.390 173.760 59.540 174.320 ;
        RECT 39.040 172.610 39.620 172.970 ;
        RECT 42.170 172.450 43.590 173.030 ;
        RECT 50.190 172.010 51.690 172.460 ;
        RECT 53.070 172.340 53.920 173.310 ;
        RECT 54.320 172.640 54.580 173.480 ;
        RECT 57.390 172.200 58.720 172.510 ;
        RECT 63.260 176.090 64.100 176.390 ;
        RECT 67.270 174.860 68.110 175.130 ;
        RECT 63.270 173.570 64.070 173.830 ;
        RECT 67.270 172.250 68.120 172.530 ;
        RECT 68.790 171.320 69.420 172.130 ;
        RECT 63.280 170.970 64.090 171.230 ;
        RECT 71.850 185.810 72.650 189.410 ;
        RECT 111.280 191.980 112.440 192.260 ;
        RECT 107.930 191.180 108.950 191.440 ;
        RECT 98.650 183.090 98.940 184.490 ;
        RECT 96.880 178.840 98.800 179.790 ;
        RECT 103.270 190.560 104.430 190.830 ;
        RECT 99.860 189.720 100.820 190.040 ;
        RECT 103.260 188.980 104.420 189.250 ;
        RECT 99.840 188.150 100.800 188.460 ;
        RECT 103.260 187.350 104.430 187.620 ;
        RECT 99.800 186.550 100.830 186.890 ;
        RECT 103.260 185.800 104.430 186.090 ;
        RECT 99.780 184.980 100.830 185.320 ;
        RECT 103.270 184.230 104.410 184.500 ;
        RECT 99.830 183.440 100.830 183.730 ;
        RECT 103.270 182.620 104.410 182.890 ;
        RECT 99.820 181.890 100.800 182.150 ;
        RECT 103.270 181.030 104.410 181.300 ;
        RECT 111.270 190.390 112.440 190.650 ;
        RECT 107.930 189.580 108.950 189.840 ;
        RECT 111.290 188.770 112.430 189.040 ;
        RECT 107.930 188.020 108.950 188.280 ;
        RECT 111.280 187.220 112.440 187.480 ;
        RECT 107.940 186.430 108.950 186.690 ;
        RECT 111.300 185.620 112.450 185.880 ;
        RECT 107.910 184.860 108.950 185.130 ;
        RECT 111.320 184.040 112.450 184.320 ;
        RECT 107.820 183.240 108.950 183.520 ;
        RECT 111.300 182.470 112.410 182.750 ;
        RECT 107.870 181.700 108.940 181.960 ;
        RECT 111.310 180.870 112.350 181.150 ;
        RECT 99.840 180.310 100.810 180.600 ;
        RECT 103.270 179.510 104.400 179.780 ;
        RECT 104.980 179.260 105.900 180.490 ;
        RECT 107.840 180.070 108.950 180.350 ;
        RECT 96.190 177.170 97.000 177.590 ;
        RECT 101.380 175.460 102.900 176.370 ;
        RECT 111.370 179.280 112.410 179.560 ;
        RECT 113.390 185.450 113.700 186.180 ;
        RECT 126.880 187.960 127.430 188.725 ;
        RECT 123.435 186.175 123.705 186.625 ;
        RECT 123.985 186.965 124.505 187.465 ;
        RECT 129.515 186.165 130.035 186.645 ;
        RECT 130.455 186.995 130.905 187.465 ;
        RECT 106.790 176.150 107.400 176.970 ;
        RECT 96.200 174.190 97.010 174.610 ;
        RECT 111.920 172.660 113.210 172.920 ;
        RECT 121.750 177.790 122.950 179.420 ;
        RECT 123.435 178.075 123.705 178.525 ;
        RECT 123.985 178.865 124.505 179.365 ;
        RECT 129.515 178.065 130.035 178.545 ;
        RECT 130.455 178.895 130.905 179.365 ;
        RECT 68.910 168.580 70.200 168.840 ;
        RECT 53.190 166.890 54.000 167.310 ;
        RECT 58.370 165.130 59.890 166.040 ;
        RECT 63.780 164.530 64.390 165.350 ;
        RECT 53.180 163.910 53.990 164.330 ;
        RECT 55.640 157.010 55.930 158.410 ;
        RECT 60.260 161.720 61.390 161.990 ;
        RECT 56.830 160.900 57.800 161.190 ;
        RECT 61.970 161.010 62.890 162.240 ;
        RECT 68.360 161.940 69.400 162.220 ;
        RECT 64.830 161.150 65.940 161.430 ;
        RECT 60.260 160.200 61.400 160.470 ;
        RECT 56.810 159.350 57.790 159.610 ;
        RECT 60.260 158.610 61.400 158.880 ;
        RECT 56.820 157.770 57.820 158.060 ;
        RECT 60.260 157.000 61.400 157.270 ;
        RECT 56.770 156.180 57.820 156.520 ;
        RECT 60.250 155.410 61.420 155.700 ;
        RECT 56.790 154.610 57.820 154.950 ;
        RECT 60.250 153.880 61.420 154.150 ;
        RECT 56.830 153.040 57.790 153.350 ;
        RECT 60.250 152.250 61.410 152.520 ;
        RECT 56.850 151.460 57.810 151.780 ;
        RECT 60.260 150.670 61.420 150.940 ;
        RECT 68.300 160.350 69.340 160.630 ;
        RECT 64.860 159.540 65.930 159.800 ;
        RECT 68.290 158.750 69.400 159.030 ;
        RECT 64.810 157.980 65.940 158.260 ;
        RECT 68.310 157.180 69.440 157.460 ;
        RECT 64.900 156.370 65.940 156.640 ;
        RECT 68.290 155.620 69.440 155.880 ;
        RECT 64.930 154.810 65.940 155.070 ;
        RECT 68.270 154.020 69.430 154.280 ;
        RECT 64.920 153.220 65.940 153.480 ;
        RECT 68.280 152.460 69.420 152.730 ;
        RECT 64.920 151.660 65.940 151.920 ;
        RECT 68.260 150.850 69.430 151.110 ;
        RECT 64.920 150.060 65.940 150.320 ;
        RECT 60.370 147.940 61.350 149.180 ;
        RECT 68.270 149.240 69.430 149.520 ;
        RECT 64.880 148.500 65.940 148.780 ;
        RECT 68.270 147.680 69.450 147.970 ;
        RECT 70.380 155.320 70.690 156.050 ;
        RECT 64.880 146.890 65.950 147.170 ;
        RECT 63.790 146.080 64.440 146.690 ;
        RECT 20.760 141.810 21.380 142.430 ;
        RECT 19.140 131.410 19.660 131.800 ;
        RECT 19.340 130.380 19.710 130.730 ;
        RECT 59.840 129.920 60.950 130.250 ;
        RECT 18.820 120.450 19.630 121.490 ;
        RECT 71.860 158.500 72.260 159.270 ;
        RECT 77.190 167.600 77.980 167.910 ;
        RECT 77.260 164.020 78.000 164.480 ;
        RECT 77.160 163.060 77.950 163.410 ;
        RECT 72.560 160.120 72.830 160.600 ;
        RECT 78.250 160.150 78.520 160.630 ;
        RECT 77.120 158.690 78.020 158.990 ;
        RECT 78.810 163.120 79.100 163.400 ;
        RECT 78.800 158.670 79.090 158.950 ;
        RECT 79.770 168.360 80.260 168.820 ;
        RECT 79.760 163.870 80.220 164.430 ;
        RECT 79.750 159.370 80.220 159.740 ;
        RECT 106.290 170.270 107.100 170.530 ;
        RECT 82.050 168.530 82.630 168.890 ;
        RECT 85.180 168.470 86.600 169.050 ;
        RECT 93.200 169.040 94.700 169.490 ;
        RECT 80.850 167.700 81.140 167.980 ;
        RECT 80.860 163.210 81.150 163.490 ;
        RECT 80.860 158.680 81.150 158.960 ;
        RECT 82.140 167.570 82.830 167.960 ;
        RECT 96.080 168.190 96.930 169.160 ;
        RECT 100.400 168.990 101.730 169.300 ;
        RECT 91.070 167.130 92.220 167.690 ;
        RECT 97.330 168.020 97.590 168.860 ;
        RECT 101.400 167.180 102.550 167.740 ;
        RECT 82.230 163.130 82.800 163.590 ;
        RECT 81.550 160.150 81.820 160.630 ;
        RECT 90.790 165.610 92.620 165.940 ;
        RECT 98.290 165.700 99.620 166.010 ;
        RECT 89.750 163.960 90.020 164.870 ;
        RECT 87.260 162.200 87.750 162.970 ;
        RECT 93.170 163.110 94.690 163.450 ;
        RECT 97.310 164.000 97.580 164.840 ;
        RECT 87.230 160.130 87.500 160.610 ;
        RECT 82.070 159.510 82.570 159.870 ;
        RECT 82.250 158.630 82.820 158.990 ;
        RECT 89.080 160.120 89.860 161.030 ;
        RECT 91.070 161.120 92.220 161.680 ;
        RECT 111.800 169.370 112.430 170.180 ;
        RECT 110.280 168.970 111.130 169.250 ;
        RECT 106.280 167.670 107.080 167.930 ;
        RECT 110.280 166.370 111.120 166.640 ;
        RECT 106.270 165.110 107.110 165.410 ;
        RECT 105.830 164.420 106.090 164.780 ;
        RECT 111.360 164.410 111.620 164.770 ;
        RECT 100.390 162.980 101.720 163.290 ;
        RECT 101.450 161.170 102.600 161.730 ;
        RECT 90.800 159.640 92.520 159.920 ;
        RECT 98.290 159.650 99.620 159.960 ;
        RECT 110.290 163.810 111.090 164.080 ;
        RECT 106.290 162.520 107.110 162.820 ;
        RECT 110.270 161.120 111.160 161.600 ;
        RECT 123.435 169.975 123.705 170.425 ;
        RECT 123.985 170.765 124.505 171.265 ;
        RECT 129.515 169.965 130.035 170.445 ;
        RECT 130.455 170.795 130.905 171.265 ;
        RECT 117.090 165.150 119.290 166.910 ;
        RECT 113.260 161.140 113.650 161.620 ;
        RECT 114.595 160.490 115.045 160.960 ;
        RECT 115.465 161.310 115.985 161.790 ;
        RECT 106.290 159.950 107.060 160.210 ;
        RECT 120.995 160.490 121.515 160.990 ;
        RECT 123.435 161.875 123.705 162.325 ;
        RECT 121.795 161.330 122.065 161.780 ;
        RECT 123.985 162.665 124.505 163.165 ;
        RECT 129.515 161.865 130.035 162.345 ;
        RECT 130.455 162.695 130.905 163.165 ;
        RECT 118.050 158.050 118.620 158.820 ;
        RECT 71.860 154.950 72.260 155.720 ;
        RECT 77.120 155.230 78.020 155.530 ;
        RECT 78.800 155.270 79.090 155.550 ;
        RECT 72.560 153.620 72.830 154.100 ;
        RECT 78.250 153.590 78.520 154.070 ;
        RECT 77.160 150.810 77.950 151.160 ;
        RECT 77.260 149.740 78.000 150.200 ;
        RECT 77.190 146.310 77.980 146.620 ;
        RECT 78.810 150.820 79.100 151.100 ;
        RECT 79.750 154.480 80.220 154.850 ;
        RECT 79.760 149.790 80.220 150.350 ;
        RECT 79.770 145.400 80.260 145.860 ;
        RECT 114.595 155.950 115.045 156.420 ;
        RECT 115.465 156.770 115.985 157.250 ;
        RECT 80.860 155.260 81.150 155.540 ;
        RECT 80.860 150.730 81.150 151.010 ;
        RECT 80.850 146.240 81.140 146.520 ;
        RECT 82.250 155.230 82.820 155.590 ;
        RECT 82.070 154.350 82.570 154.710 ;
        RECT 81.550 153.590 81.820 154.070 ;
        RECT 120.995 155.950 121.515 156.450 ;
        RECT 121.795 156.790 122.065 157.240 ;
        RECT 90.800 154.300 92.520 154.580 ;
        RECT 87.230 153.610 87.500 154.090 ;
        RECT 98.290 154.260 99.620 154.570 ;
        RECT 89.080 153.190 89.860 154.100 ;
        RECT 87.260 151.250 87.750 152.020 ;
        RECT 82.230 150.630 82.800 151.090 ;
        RECT 82.140 146.260 82.830 146.650 ;
        RECT 91.070 152.540 92.220 153.100 ;
        RECT 106.290 154.010 107.060 154.270 ;
        RECT 101.450 152.490 102.600 153.050 ;
        RECT 93.170 150.770 94.690 151.110 ;
        RECT 89.750 149.350 90.020 150.260 ;
        RECT 100.390 150.930 101.720 151.240 ;
        RECT 97.310 149.380 97.580 150.220 ;
        RECT 110.270 152.620 111.160 153.100 ;
        RECT 113.260 152.600 113.650 153.080 ;
        RECT 106.290 151.400 107.110 151.700 ;
        RECT 110.290 150.140 111.090 150.410 ;
        RECT 105.830 149.440 106.090 149.800 ;
        RECT 111.360 149.450 111.620 149.810 ;
        RECT 90.790 148.280 92.620 148.610 ;
        RECT 98.290 148.210 99.620 148.520 ;
        RECT 91.070 146.530 92.220 147.090 ;
        RECT 101.400 146.480 102.550 147.040 ;
        RECT 82.050 145.330 82.630 145.690 ;
        RECT 85.180 145.170 86.600 145.750 ;
        RECT 93.200 144.730 94.700 145.180 ;
        RECT 96.080 145.060 96.930 146.030 ;
        RECT 97.330 145.360 97.590 146.200 ;
        RECT 100.400 144.920 101.730 145.230 ;
        RECT 106.270 148.810 107.110 149.110 ;
        RECT 110.280 147.580 111.120 147.850 ;
        RECT 106.280 146.290 107.080 146.550 ;
        RECT 110.280 144.970 111.130 145.250 ;
        RECT 114.595 151.890 115.045 152.360 ;
        RECT 115.465 152.710 115.985 153.190 ;
        RECT 123.435 153.775 123.705 154.225 ;
        RECT 120.995 151.890 121.515 152.390 ;
        RECT 123.985 154.565 124.505 155.065 ;
        RECT 121.795 152.730 122.065 153.180 ;
        RECT 129.515 153.765 130.035 154.245 ;
        RECT 130.455 154.595 130.905 155.065 ;
        RECT 114.595 147.830 115.045 148.300 ;
        RECT 115.465 148.650 115.985 149.130 ;
        RECT 120.995 147.830 121.515 148.330 ;
        RECT 121.795 148.670 122.065 149.120 ;
        RECT 111.800 144.040 112.430 144.850 ;
        RECT 106.290 143.690 107.100 143.950 ;
        RECT 114.595 143.770 115.045 144.240 ;
        RECT 115.465 144.590 115.985 145.070 ;
        RECT 123.435 145.675 123.705 146.125 ;
        RECT 120.995 143.770 121.515 144.270 ;
        RECT 123.985 146.465 124.505 146.965 ;
        RECT 121.795 144.610 122.065 145.060 ;
        RECT 129.515 145.665 130.035 146.145 ;
        RECT 130.455 146.495 130.905 146.965 ;
        RECT 111.920 141.300 113.210 141.560 ;
        RECT 96.200 139.610 97.010 140.030 ;
        RECT 114.595 139.710 115.045 140.180 ;
        RECT 115.465 140.530 115.985 141.010 ;
        RECT 101.380 137.850 102.900 138.760 ;
        RECT 106.790 137.250 107.400 138.070 ;
        RECT 96.190 136.630 97.000 137.050 ;
        RECT 98.650 129.730 98.940 131.130 ;
        RECT 18.810 105.630 19.770 106.460 ;
        RECT 59.850 96.980 60.960 97.310 ;
        RECT 19.350 96.500 19.720 96.850 ;
        RECT 19.150 95.430 19.670 95.820 ;
        RECT 20.770 84.800 21.390 85.420 ;
        RECT 63.970 80.070 64.440 81.020 ;
        RECT 64.890 80.060 65.960 80.340 ;
        RECT 60.380 78.050 61.360 79.290 ;
        RECT 18.470 72.340 19.060 74.260 ;
        RECT 68.280 79.260 69.460 79.550 ;
        RECT 64.890 78.450 65.950 78.730 ;
        RECT 68.280 77.710 69.440 77.990 ;
        RECT 64.930 76.910 65.950 77.170 ;
        RECT 55.650 68.820 55.940 70.220 ;
        RECT 60.270 76.290 61.430 76.560 ;
        RECT 56.860 75.450 57.820 75.770 ;
        RECT 60.260 74.710 61.420 74.980 ;
        RECT 56.840 73.880 57.800 74.190 ;
        RECT 60.260 73.080 61.430 73.350 ;
        RECT 56.800 72.280 57.830 72.620 ;
        RECT 60.260 71.530 61.430 71.820 ;
        RECT 56.780 70.710 57.830 71.050 ;
        RECT 60.270 69.960 61.410 70.230 ;
        RECT 56.830 69.170 57.830 69.460 ;
        RECT 60.270 68.350 61.410 68.620 ;
        RECT 56.820 67.620 57.800 67.880 ;
        RECT 60.270 66.760 61.410 67.030 ;
        RECT 68.270 76.120 69.440 76.380 ;
        RECT 64.930 75.310 65.950 75.570 ;
        RECT 68.290 74.500 69.430 74.770 ;
        RECT 64.930 73.750 65.950 74.010 ;
        RECT 68.280 72.950 69.440 73.210 ;
        RECT 64.940 72.160 65.950 72.420 ;
        RECT 68.300 71.350 69.450 71.610 ;
        RECT 64.910 70.590 65.950 70.860 ;
        RECT 68.320 69.770 69.450 70.050 ;
        RECT 64.820 68.970 65.950 69.250 ;
        RECT 68.300 68.200 69.410 68.480 ;
        RECT 64.870 67.430 65.940 67.690 ;
        RECT 68.310 66.600 69.350 66.880 ;
        RECT 56.840 66.040 57.810 66.330 ;
        RECT 60.270 65.240 61.400 65.510 ;
        RECT 61.980 64.990 62.900 66.220 ;
        RECT 53.190 62.900 54.000 63.320 ;
        RECT 58.380 61.190 59.900 62.100 ;
        RECT 64.840 65.800 65.950 66.080 ;
        RECT 68.370 65.010 69.410 65.290 ;
        RECT 70.390 71.180 70.700 71.910 ;
        RECT 63.790 61.880 64.400 62.700 ;
        RECT 53.200 59.920 54.010 60.340 ;
        RECT 68.920 58.390 70.210 58.650 ;
        RECT 27.480 52.750 27.950 53.890 ;
        RECT 27.090 41.380 27.980 43.850 ;
        RECT 28.860 44.230 29.260 45.000 ;
        RECT 34.190 53.330 34.980 53.640 ;
        RECT 34.260 49.750 35.000 50.210 ;
        RECT 34.160 48.790 34.950 49.140 ;
        RECT 29.560 45.850 29.830 46.330 ;
        RECT 35.250 45.880 35.520 46.360 ;
        RECT 34.120 44.420 35.020 44.720 ;
        RECT 35.810 48.850 36.100 49.130 ;
        RECT 35.800 44.400 36.090 44.680 ;
        RECT 36.770 54.090 37.260 54.550 ;
        RECT 36.760 49.600 37.220 50.160 ;
        RECT 36.750 45.100 37.220 45.470 ;
        RECT 63.290 56.000 64.100 56.260 ;
        RECT 39.050 54.260 39.630 54.620 ;
        RECT 42.180 54.200 43.600 54.780 ;
        RECT 50.200 54.770 51.700 55.220 ;
        RECT 37.850 53.430 38.140 53.710 ;
        RECT 37.860 48.940 38.150 49.220 ;
        RECT 37.860 44.410 38.150 44.690 ;
        RECT 39.140 53.300 39.830 53.690 ;
        RECT 53.080 53.920 53.930 54.890 ;
        RECT 57.400 54.720 58.730 55.030 ;
        RECT 48.070 52.860 49.220 53.420 ;
        RECT 54.330 53.750 54.590 54.590 ;
        RECT 58.400 52.910 59.550 53.470 ;
        RECT 39.230 48.860 39.800 49.320 ;
        RECT 38.550 45.880 38.820 46.360 ;
        RECT 47.790 51.340 49.620 51.670 ;
        RECT 55.290 51.430 56.620 51.740 ;
        RECT 46.750 49.690 47.020 50.600 ;
        RECT 44.260 47.930 44.750 48.700 ;
        RECT 50.170 48.840 51.690 49.180 ;
        RECT 54.310 49.730 54.580 50.570 ;
        RECT 44.230 45.860 44.500 46.340 ;
        RECT 39.070 45.240 39.570 45.600 ;
        RECT 39.250 44.360 39.820 44.720 ;
        RECT 46.080 45.850 46.860 46.760 ;
        RECT 48.070 46.850 49.220 47.410 ;
        RECT 68.800 55.100 69.430 55.910 ;
        RECT 67.280 54.700 68.130 54.980 ;
        RECT 63.280 53.400 64.080 53.660 ;
        RECT 67.280 52.100 68.120 52.370 ;
        RECT 63.270 50.840 64.110 51.140 ;
        RECT 62.830 50.150 63.090 50.510 ;
        RECT 68.360 50.140 68.620 50.500 ;
        RECT 57.390 48.710 58.720 49.020 ;
        RECT 58.450 46.900 59.600 47.460 ;
        RECT 47.800 45.370 49.520 45.650 ;
        RECT 55.290 45.380 56.620 45.690 ;
        RECT 67.290 49.540 68.090 49.810 ;
        RECT 63.290 48.250 64.110 48.550 ;
        RECT 67.270 46.850 68.160 47.330 ;
        RECT 70.260 46.870 70.650 47.350 ;
        RECT 63.290 45.680 64.060 45.940 ;
        RECT 103.270 134.440 104.400 134.710 ;
        RECT 99.840 133.620 100.810 133.910 ;
        RECT 104.980 133.730 105.900 134.960 ;
        RECT 103.270 132.920 104.410 133.190 ;
        RECT 99.820 132.070 100.800 132.330 ;
        RECT 103.270 131.330 104.410 131.600 ;
        RECT 99.830 130.490 100.830 130.780 ;
        RECT 103.270 129.720 104.410 129.990 ;
        RECT 99.780 128.900 100.830 129.240 ;
        RECT 103.260 128.130 104.430 128.420 ;
        RECT 99.800 127.330 100.830 127.670 ;
        RECT 103.260 126.600 104.430 126.870 ;
        RECT 99.840 125.760 100.800 126.070 ;
        RECT 103.260 124.970 104.420 125.240 ;
        RECT 99.860 124.180 100.820 124.500 ;
        RECT 103.270 123.390 104.430 123.660 ;
        RECT 120.995 139.710 121.515 140.210 ;
        RECT 121.795 140.550 122.065 141.000 ;
        RECT 111.370 134.660 112.410 134.940 ;
        RECT 107.840 133.870 108.950 134.150 ;
        RECT 111.310 133.070 112.350 133.350 ;
        RECT 107.870 132.260 108.940 132.520 ;
        RECT 111.300 131.470 112.410 131.750 ;
        RECT 107.820 130.700 108.950 130.980 ;
        RECT 111.320 129.900 112.450 130.180 ;
        RECT 107.910 129.090 108.950 129.360 ;
        RECT 111.300 128.340 112.450 128.600 ;
        RECT 107.940 127.530 108.950 127.790 ;
        RECT 111.280 126.740 112.440 127.000 ;
        RECT 107.930 125.940 108.950 126.200 ;
        RECT 111.290 125.180 112.430 125.450 ;
        RECT 107.930 124.380 108.950 124.640 ;
        RECT 111.270 123.570 112.440 123.830 ;
        RECT 114.570 134.390 115.310 136.010 ;
        RECT 123.435 137.575 123.705 138.025 ;
        RECT 123.985 138.365 124.505 138.865 ;
        RECT 129.515 137.565 130.035 138.045 ;
        RECT 130.455 138.395 130.905 138.865 ;
        RECT 114.595 131.590 115.045 132.060 ;
        RECT 115.465 132.410 115.985 132.890 ;
        RECT 120.995 131.590 121.515 132.090 ;
        RECT 121.795 132.430 122.065 132.880 ;
        RECT 129.930 134.400 130.800 135.980 ;
        RECT 113.390 128.040 113.700 128.770 ;
        RECT 114.595 127.530 115.045 128.000 ;
        RECT 115.465 128.350 115.985 128.830 ;
        RECT 123.435 129.475 123.705 129.925 ;
        RECT 120.995 127.530 121.515 128.030 ;
        RECT 123.985 130.265 124.505 130.765 ;
        RECT 121.795 128.370 122.065 128.820 ;
        RECT 129.515 129.465 130.035 129.945 ;
        RECT 130.455 130.295 130.905 130.765 ;
        RECT 114.595 123.470 115.045 123.940 ;
        RECT 115.465 124.290 115.985 124.770 ;
        RECT 107.930 122.780 108.950 123.040 ;
        RECT 111.280 121.960 112.440 122.240 ;
        RECT 107.890 121.220 108.950 121.500 ;
        RECT 111.280 120.400 112.460 120.690 ;
        RECT 98.250 117.980 98.890 119.160 ;
        RECT 107.890 119.610 108.960 119.890 ;
        RECT 120.995 123.470 121.515 123.970 ;
        RECT 121.795 124.310 122.065 124.760 ;
        RECT 114.595 119.410 115.045 119.880 ;
        RECT 115.465 120.230 115.985 120.710 ;
        RECT 123.435 121.375 123.705 121.825 ;
        RECT 120.995 119.410 121.515 119.910 ;
        RECT 123.985 122.165 124.505 122.665 ;
        RECT 121.795 120.250 122.065 120.700 ;
        RECT 129.515 121.365 130.035 121.845 ;
        RECT 130.455 122.195 130.905 122.665 ;
        RECT 107.890 117.420 108.960 117.700 ;
        RECT 111.280 116.620 112.460 116.910 ;
        RECT 122.130 117.900 123.300 119.230 ;
        RECT 107.890 115.810 108.950 116.090 ;
        RECT 111.280 115.070 112.440 115.350 ;
        RECT 107.930 114.270 108.950 114.530 ;
        RECT 98.650 106.180 98.940 107.580 ;
        RECT 103.270 113.650 104.430 113.920 ;
        RECT 99.860 112.810 100.820 113.130 ;
        RECT 103.260 112.070 104.420 112.340 ;
        RECT 99.840 111.240 100.800 111.550 ;
        RECT 103.260 110.440 104.430 110.710 ;
        RECT 99.800 109.640 100.830 109.980 ;
        RECT 103.260 108.890 104.430 109.180 ;
        RECT 99.780 108.070 100.830 108.410 ;
        RECT 103.270 107.320 104.410 107.590 ;
        RECT 99.830 106.530 100.830 106.820 ;
        RECT 103.270 105.710 104.410 105.980 ;
        RECT 99.820 104.980 100.800 105.240 ;
        RECT 103.270 104.120 104.410 104.390 ;
        RECT 111.270 113.480 112.440 113.740 ;
        RECT 107.930 112.670 108.950 112.930 ;
        RECT 111.290 111.860 112.430 112.130 ;
        RECT 107.930 111.110 108.950 111.370 ;
        RECT 111.280 110.310 112.440 110.570 ;
        RECT 107.940 109.520 108.950 109.780 ;
        RECT 111.300 108.710 112.450 108.970 ;
        RECT 107.910 107.950 108.950 108.220 ;
        RECT 111.320 107.130 112.450 107.410 ;
        RECT 107.820 106.330 108.950 106.610 ;
        RECT 111.300 105.560 112.410 105.840 ;
        RECT 107.870 104.790 108.940 105.050 ;
        RECT 111.310 103.960 112.350 104.240 ;
        RECT 99.840 103.400 100.810 103.690 ;
        RECT 103.270 102.600 104.400 102.870 ;
        RECT 104.980 102.350 105.900 103.580 ;
        RECT 96.190 100.260 97.000 100.680 ;
        RECT 101.380 98.550 102.900 99.460 ;
        RECT 107.840 103.160 108.950 103.440 ;
        RECT 111.370 102.370 112.410 102.650 ;
        RECT 114.595 115.350 115.045 115.820 ;
        RECT 115.465 116.170 115.985 116.650 ;
        RECT 120.995 115.350 121.515 115.850 ;
        RECT 121.795 116.190 122.065 116.640 ;
        RECT 114.595 111.290 115.045 111.760 ;
        RECT 115.465 112.110 115.985 112.590 ;
        RECT 123.435 113.275 123.705 113.725 ;
        RECT 120.995 111.290 121.515 111.790 ;
        RECT 123.985 114.065 124.505 114.565 ;
        RECT 121.795 112.130 122.065 112.580 ;
        RECT 129.515 113.265 130.035 113.745 ;
        RECT 130.455 114.095 130.905 114.565 ;
        RECT 113.390 108.540 113.700 109.270 ;
        RECT 114.595 107.230 115.045 107.700 ;
        RECT 115.465 108.050 115.985 108.530 ;
        RECT 120.995 107.230 121.515 107.730 ;
        RECT 121.795 108.070 122.065 108.520 ;
        RECT 114.595 103.170 115.045 103.640 ;
        RECT 115.465 103.990 115.985 104.470 ;
        RECT 123.435 105.175 123.705 105.625 ;
        RECT 120.995 103.170 121.515 103.670 ;
        RECT 123.985 105.965 124.505 106.465 ;
        RECT 121.795 104.010 122.065 104.460 ;
        RECT 129.515 105.165 130.035 105.645 ;
        RECT 130.455 105.995 130.905 106.465 ;
        RECT 106.790 99.240 107.400 100.060 ;
        RECT 114.595 99.110 115.045 99.580 ;
        RECT 115.465 99.930 115.985 100.410 ;
        RECT 123.435 101.125 123.705 101.575 ;
        RECT 120.995 99.110 121.515 99.610 ;
        RECT 123.985 101.915 124.505 102.415 ;
        RECT 121.795 99.950 122.065 100.400 ;
        RECT 129.515 101.115 130.035 101.595 ;
        RECT 130.455 101.945 130.905 102.415 ;
        RECT 96.200 97.280 97.010 97.700 ;
        RECT 111.920 95.750 113.210 96.010 ;
        RECT 71.860 81.590 72.260 82.360 ;
        RECT 77.190 90.690 77.980 91.000 ;
        RECT 77.260 87.110 78.000 87.570 ;
        RECT 77.160 86.150 77.950 86.500 ;
        RECT 72.560 83.210 72.830 83.690 ;
        RECT 78.250 83.240 78.520 83.720 ;
        RECT 77.120 81.780 78.020 82.080 ;
        RECT 78.810 86.210 79.100 86.490 ;
        RECT 78.800 81.760 79.090 82.040 ;
        RECT 79.770 91.450 80.260 91.910 ;
        RECT 79.760 86.960 80.220 87.520 ;
        RECT 79.750 82.460 80.220 82.830 ;
        RECT 106.290 93.360 107.100 93.620 ;
        RECT 82.050 91.620 82.630 91.980 ;
        RECT 85.180 91.560 86.600 92.140 ;
        RECT 93.200 92.130 94.700 92.580 ;
        RECT 80.850 90.790 81.140 91.070 ;
        RECT 80.860 86.300 81.150 86.580 ;
        RECT 80.860 81.770 81.150 82.050 ;
        RECT 82.140 90.660 82.830 91.050 ;
        RECT 96.080 91.280 96.930 92.250 ;
        RECT 100.400 92.080 101.730 92.390 ;
        RECT 91.070 90.220 92.220 90.780 ;
        RECT 97.330 91.110 97.590 91.950 ;
        RECT 101.400 90.270 102.550 90.830 ;
        RECT 82.230 86.220 82.800 86.680 ;
        RECT 81.550 83.240 81.820 83.720 ;
        RECT 90.790 88.700 92.620 89.030 ;
        RECT 98.290 88.790 99.620 89.100 ;
        RECT 89.750 87.050 90.020 87.960 ;
        RECT 87.260 85.290 87.750 86.060 ;
        RECT 93.170 86.200 94.690 86.540 ;
        RECT 97.310 87.090 97.580 87.930 ;
        RECT 87.230 83.220 87.500 83.700 ;
        RECT 82.070 82.600 82.570 82.960 ;
        RECT 82.250 81.720 82.820 82.080 ;
        RECT 89.080 83.210 89.860 84.120 ;
        RECT 91.070 84.210 92.220 84.770 ;
        RECT 111.800 92.460 112.430 93.270 ;
        RECT 123.435 97.075 123.705 97.525 ;
        RECT 123.985 97.865 124.505 98.365 ;
        RECT 129.515 97.065 130.035 97.545 ;
        RECT 130.455 97.895 130.905 98.365 ;
        RECT 110.280 92.060 111.130 92.340 ;
        RECT 106.280 90.760 107.080 91.020 ;
        RECT 110.280 89.460 111.120 89.730 ;
        RECT 106.270 88.200 107.110 88.500 ;
        RECT 105.830 87.510 106.090 87.870 ;
        RECT 111.360 87.500 111.620 87.860 ;
        RECT 100.390 86.070 101.720 86.380 ;
        RECT 101.450 84.260 102.600 84.820 ;
        RECT 90.800 82.730 92.520 83.010 ;
        RECT 98.290 82.740 99.620 83.050 ;
        RECT 110.290 86.900 111.090 87.170 ;
        RECT 106.290 85.610 107.110 85.910 ;
        RECT 110.270 84.210 111.160 84.690 ;
        RECT 114.595 90.990 115.045 91.460 ;
        RECT 115.465 91.810 115.985 92.290 ;
        RECT 123.435 93.025 123.705 93.475 ;
        RECT 120.995 90.990 121.515 91.490 ;
        RECT 123.985 93.815 124.505 94.315 ;
        RECT 121.795 91.830 122.065 92.280 ;
        RECT 129.515 93.015 130.035 93.495 ;
        RECT 130.455 93.845 130.905 94.315 ;
        RECT 114.595 86.930 115.045 87.400 ;
        RECT 115.465 87.750 115.985 88.230 ;
        RECT 123.435 88.975 123.705 89.425 ;
        RECT 120.995 86.930 121.515 87.430 ;
        RECT 123.985 89.765 124.505 90.265 ;
        RECT 121.795 87.770 122.065 88.220 ;
        RECT 129.515 88.965 130.035 89.445 ;
        RECT 130.455 89.795 130.905 90.265 ;
        RECT 113.260 84.230 113.650 84.710 ;
        RECT 106.290 83.040 107.060 83.300 ;
        RECT 114.595 82.870 115.045 83.340 ;
        RECT 115.465 83.690 115.985 84.170 ;
        RECT 123.435 84.925 123.705 85.375 ;
        RECT 120.995 82.870 121.515 83.370 ;
        RECT 123.985 85.715 124.505 86.215 ;
        RECT 121.795 83.710 122.065 84.160 ;
        RECT 129.515 84.915 130.035 85.395 ;
        RECT 130.455 85.745 130.905 86.215 ;
        RECT 71.860 79.350 72.260 80.120 ;
        RECT 77.120 79.630 78.020 79.930 ;
        RECT 78.800 79.670 79.090 79.950 ;
        RECT 72.560 78.020 72.830 78.500 ;
        RECT 78.250 77.990 78.520 78.470 ;
        RECT 77.160 75.210 77.950 75.560 ;
        RECT 77.260 74.140 78.000 74.600 ;
        RECT 77.190 70.710 77.980 71.020 ;
        RECT 78.810 75.220 79.100 75.500 ;
        RECT 79.750 78.880 80.220 79.250 ;
        RECT 79.760 74.190 80.220 74.750 ;
        RECT 79.770 69.800 80.260 70.260 ;
        RECT 80.860 79.660 81.150 79.940 ;
        RECT 80.860 75.130 81.150 75.410 ;
        RECT 80.850 70.640 81.140 70.920 ;
        RECT 82.250 79.630 82.820 79.990 ;
        RECT 82.070 78.750 82.570 79.110 ;
        RECT 81.550 77.990 81.820 78.470 ;
        RECT 90.800 78.700 92.520 78.980 ;
        RECT 87.230 78.010 87.500 78.490 ;
        RECT 98.290 78.660 99.620 78.970 ;
        RECT 89.080 77.590 89.860 78.500 ;
        RECT 87.260 75.650 87.750 76.420 ;
        RECT 82.230 75.030 82.800 75.490 ;
        RECT 82.140 70.660 82.830 71.050 ;
        RECT 91.070 76.940 92.220 77.500 ;
        RECT 114.595 78.810 115.045 79.280 ;
        RECT 115.465 79.630 115.985 80.110 ;
        RECT 106.290 78.410 107.060 78.670 ;
        RECT 101.450 76.890 102.600 77.450 ;
        RECT 93.170 75.170 94.690 75.510 ;
        RECT 89.750 73.750 90.020 74.660 ;
        RECT 100.390 75.330 101.720 75.640 ;
        RECT 97.310 73.780 97.580 74.620 ;
        RECT 110.270 77.020 111.160 77.500 ;
        RECT 123.435 80.875 123.705 81.325 ;
        RECT 120.995 78.810 121.515 79.310 ;
        RECT 123.985 81.665 124.505 82.165 ;
        RECT 121.795 79.650 122.065 80.100 ;
        RECT 129.515 80.865 130.035 81.345 ;
        RECT 130.455 81.695 130.905 82.165 ;
        RECT 113.260 77.000 113.650 77.480 ;
        RECT 106.290 75.800 107.110 76.100 ;
        RECT 110.290 74.540 111.090 74.810 ;
        RECT 105.830 73.840 106.090 74.200 ;
        RECT 111.360 73.850 111.620 74.210 ;
        RECT 90.790 72.680 92.620 73.010 ;
        RECT 98.290 72.610 99.620 72.920 ;
        RECT 91.070 70.930 92.220 71.490 ;
        RECT 101.400 70.880 102.550 71.440 ;
        RECT 82.050 69.730 82.630 70.090 ;
        RECT 85.180 69.570 86.600 70.150 ;
        RECT 93.200 69.130 94.700 69.580 ;
        RECT 96.080 69.460 96.930 70.430 ;
        RECT 97.330 69.760 97.590 70.600 ;
        RECT 100.400 69.320 101.730 69.630 ;
        RECT 106.270 73.210 107.110 73.510 ;
        RECT 110.280 71.980 111.120 72.250 ;
        RECT 106.280 70.690 107.080 70.950 ;
        RECT 110.280 69.370 111.130 69.650 ;
        RECT 123.435 76.825 123.705 77.275 ;
        RECT 114.595 74.750 115.045 75.220 ;
        RECT 115.465 75.570 115.985 76.050 ;
        RECT 120.995 74.750 121.515 75.250 ;
        RECT 123.985 77.615 124.505 78.115 ;
        RECT 129.515 76.815 130.035 77.295 ;
        RECT 130.455 77.645 130.905 78.115 ;
        RECT 121.795 75.590 122.065 76.040 ;
        RECT 118.050 73.520 118.610 74.110 ;
        RECT 111.800 68.440 112.430 69.250 ;
        RECT 106.290 68.090 107.100 68.350 ;
        RECT 111.920 65.700 113.210 65.960 ;
        RECT 96.200 64.010 97.010 64.430 ;
        RECT 101.380 62.250 102.900 63.160 ;
        RECT 106.790 61.650 107.400 62.470 ;
        RECT 96.190 61.030 97.000 61.450 ;
        RECT 95.110 58.730 98.650 59.820 ;
        RECT 98.650 54.130 98.940 55.530 ;
        RECT 103.270 58.840 104.400 59.110 ;
        RECT 99.840 58.020 100.810 58.310 ;
        RECT 104.980 58.130 105.900 59.360 ;
        RECT 123.435 72.775 123.705 73.225 ;
        RECT 123.985 73.565 124.505 74.065 ;
        RECT 129.515 72.765 130.035 73.245 ;
        RECT 130.455 73.595 130.905 74.065 ;
        RECT 123.435 68.690 123.705 69.140 ;
        RECT 123.985 69.480 124.505 69.980 ;
        RECT 129.515 68.680 130.035 69.160 ;
        RECT 130.455 69.510 130.905 69.980 ;
        RECT 123.435 64.565 123.705 65.015 ;
        RECT 123.985 65.355 124.505 65.855 ;
        RECT 129.515 64.555 130.035 65.035 ;
        RECT 130.455 65.385 130.905 65.855 ;
        RECT 126.870 63.055 127.455 63.825 ;
        RECT 103.270 57.320 104.410 57.590 ;
        RECT 99.820 56.470 100.800 56.730 ;
        RECT 103.270 55.730 104.410 56.000 ;
        RECT 99.830 54.890 100.830 55.180 ;
        RECT 103.270 54.120 104.410 54.390 ;
        RECT 99.780 53.300 100.830 53.640 ;
        RECT 103.260 52.530 104.430 52.820 ;
        RECT 99.800 51.730 100.830 52.070 ;
        RECT 103.260 51.000 104.430 51.270 ;
        RECT 99.840 50.160 100.800 50.470 ;
        RECT 103.260 49.370 104.420 49.640 ;
        RECT 99.860 48.580 100.820 48.900 ;
        RECT 103.270 47.790 104.430 48.060 ;
        RECT 111.370 59.060 112.410 59.340 ;
        RECT 107.840 58.270 108.950 58.550 ;
        RECT 111.310 57.470 112.350 57.750 ;
        RECT 107.870 56.660 108.940 56.920 ;
        RECT 111.300 55.870 112.410 56.150 ;
        RECT 107.820 55.100 108.950 55.380 ;
        RECT 111.320 54.300 112.450 54.580 ;
        RECT 107.910 53.490 108.950 53.760 ;
        RECT 111.300 52.740 112.450 53.000 ;
        RECT 107.940 51.930 108.950 52.190 ;
        RECT 111.280 51.140 112.440 51.400 ;
        RECT 107.930 50.340 108.950 50.600 ;
        RECT 111.290 49.580 112.430 49.850 ;
        RECT 107.930 48.780 108.950 49.040 ;
        RECT 111.270 47.970 112.440 48.230 ;
        RECT 107.930 47.180 108.950 47.440 ;
        RECT 111.280 46.360 112.440 46.640 ;
        RECT 107.890 45.620 108.950 45.900 ;
        RECT 111.280 44.800 112.460 45.090 ;
        RECT 107.890 44.010 108.960 44.290 ;
        RECT 121.400 58.600 122.600 62.050 ;
        RECT 123.435 60.010 123.705 60.460 ;
        RECT 123.985 60.800 124.505 61.300 ;
        RECT 129.515 60.000 130.035 60.480 ;
        RECT 130.455 60.830 130.905 61.300 ;
        RECT 113.390 52.440 113.700 53.170 ;
        RECT 106.260 41.260 107.440 42.310 ;
        RECT 126.230 53.680 127.970 55.000 ;
        RECT 28.130 37.230 29.930 38.610 ;
        RECT 122.080 36.240 123.730 38.900 ;
      LAYER met2 ;
        RECT 26.470 198.720 28.630 199.050 ;
        RECT 26.470 197.650 70.980 198.720 ;
        RECT 26.470 197.400 28.630 197.650 ;
        RECT 70.460 196.355 70.970 197.650 ;
        RECT 71.670 196.690 73.270 199.800 ;
        RECT 101.780 197.730 104.760 198.080 ;
        RECT 74.400 197.715 104.760 197.730 ;
        RECT 73.705 197.350 104.760 197.715 ;
        RECT 73.705 197.205 74.885 197.350 ;
        RECT 73.705 196.410 74.215 197.205 ;
        RECT 101.780 196.790 104.760 197.350 ;
        RECT 130.110 196.690 131.170 199.800 ;
        RECT 73.705 196.355 74.000 196.410 ;
        RECT 31.050 195.715 70.050 196.140 ;
        RECT 70.460 195.845 74.000 196.355 ;
        RECT 106.270 196.140 107.580 196.490 ;
        RECT 31.050 192.890 31.475 195.715 ;
        RECT 65.795 195.710 70.050 195.715 ;
        RECT 74.500 195.710 108.250 196.140 ;
        RECT 69.620 194.995 70.050 195.710 ;
        RECT 74.285 195.220 75.370 195.710 ;
        RECT 106.270 195.580 107.580 195.710 ;
        RECT 74.285 194.995 74.715 195.220 ;
        RECT 69.620 194.565 74.715 194.995 ;
        RECT 107.810 194.640 109.010 194.650 ;
        RECT 107.810 194.300 112.700 194.640 ;
        RECT 107.810 194.290 109.010 194.300 ;
        RECT 111.220 193.850 112.500 193.860 ;
        RECT 107.850 193.510 112.690 193.850 ;
        RECT 111.220 193.500 112.500 193.510 ;
        RECT 30.720 191.780 32.420 192.890 ;
        RECT 62.050 191.280 69.880 193.340 ;
        RECT 107.810 193.030 108.990 193.060 ;
        RECT 107.810 192.690 112.690 193.030 ;
        RECT 107.810 192.640 108.990 192.690 ;
        RECT 111.230 192.270 112.500 192.310 ;
        RECT 107.860 191.930 112.700 192.270 ;
        RECT 111.230 191.920 112.500 191.930 ;
        RECT 107.850 191.470 109.000 191.480 ;
        RECT 107.850 191.130 112.690 191.470 ;
        RECT 99.790 190.530 104.630 190.870 ;
        RECT 103.220 190.520 104.480 190.530 ;
        RECT 107.830 190.340 112.670 190.680 ;
        RECT 99.800 190.050 100.880 190.100 ;
        RECT 99.800 189.710 104.650 190.050 ;
        RECT 107.810 189.890 109.000 189.900 ;
        RECT 63.180 185.310 72.930 189.680 ;
        RECT 99.800 189.670 100.880 189.710 ;
        RECT 107.810 189.550 112.650 189.890 ;
        RECT 107.810 189.540 109.000 189.550 ;
        RECT 99.810 188.940 104.650 189.280 ;
        RECT 107.800 188.740 112.640 189.080 ;
        RECT 99.780 188.480 100.880 188.520 ;
        RECT 99.780 188.140 104.660 188.480 ;
        RECT 99.780 188.100 100.880 188.140 ;
        RECT 107.850 187.980 112.690 188.320 ;
        RECT 107.850 187.970 109.000 187.980 ;
        RECT 126.810 187.860 127.510 188.780 ;
        RECT 99.750 187.310 104.590 187.650 ;
        RECT 107.850 187.170 112.690 187.510 ;
        RECT 99.730 186.880 100.880 186.960 ;
        RECT 123.945 186.935 130.935 187.505 ;
        RECT 99.730 186.540 104.570 186.880 ;
        RECT 99.730 186.500 100.880 186.540 ;
        RECT 107.880 186.380 112.720 186.720 ;
        RECT 99.690 185.780 104.530 186.120 ;
        RECT 113.350 185.970 113.770 186.230 ;
        RECT 123.395 186.125 130.095 186.695 ;
        RECT 111.230 185.920 113.770 185.970 ;
        RECT 107.860 185.580 113.770 185.920 ;
        RECT 111.230 185.510 113.770 185.580 ;
        RECT 113.350 185.370 113.770 185.510 ;
        RECT 99.720 185.320 100.880 185.370 ;
        RECT 99.710 184.980 104.550 185.320 ;
        RECT 106.210 185.190 106.540 185.210 ;
        RECT 106.210 185.180 108.940 185.190 ;
        RECT 106.210 185.170 109.010 185.180 ;
        RECT 99.720 184.950 100.880 184.980 ;
        RECT 106.210 184.830 112.700 185.170 ;
        RECT 106.210 184.820 109.010 184.830 ;
        RECT 98.580 183.830 99.010 184.570 ;
        RECT 106.210 184.540 106.540 184.820 ;
        RECT 103.220 184.530 106.540 184.540 ;
        RECT 99.700 184.190 106.540 184.530 ;
        RECT 103.220 184.180 106.540 184.190 ;
        RECT 103.690 184.170 106.540 184.180 ;
        RECT 106.210 184.150 106.540 184.170 ;
        RECT 107.810 184.020 112.650 184.360 ;
        RECT 98.580 183.760 100.890 183.830 ;
        RECT 98.580 183.420 104.640 183.760 ;
        RECT 98.580 183.350 100.890 183.420 ;
        RECT 28.770 182.910 29.320 183.080 ;
        RECT 28.760 182.880 35.100 182.910 ;
        RECT 35.720 182.880 38.240 182.890 ;
        RECT 39.180 182.880 39.900 183.000 ;
        RECT 98.580 182.980 99.010 183.350 ;
        RECT 107.760 183.220 112.600 183.560 ;
        RECT 107.760 183.210 109.000 183.220 ;
        RECT 103.220 182.930 104.480 182.940 ;
        RECT 28.760 182.510 39.900 182.880 ;
        RECT 99.760 182.590 104.600 182.930 ;
        RECT 111.230 182.760 112.510 182.800 ;
        RECT 103.220 182.580 104.480 182.590 ;
        RECT 28.760 182.460 35.100 182.510 ;
        RECT 35.720 182.490 38.240 182.510 ;
        RECT 28.760 182.390 35.060 182.460 ;
        RECT 39.180 182.430 39.900 182.510 ;
        RECT 107.730 182.420 112.570 182.760 ;
        RECT 111.230 182.400 112.510 182.420 ;
        RECT 28.770 182.120 29.320 182.390 ;
        RECT 36.630 182.040 37.570 182.340 ;
        RECT 99.740 182.170 100.890 182.220 ;
        RECT 38.990 182.040 39.620 182.070 ;
        RECT 36.630 181.640 39.620 182.040 ;
        RECT 36.630 181.580 37.570 181.640 ;
        RECT 38.990 181.600 39.620 181.640 ;
        RECT 29.520 180.800 44.520 181.440 ;
        RECT 45.920 181.270 47.030 181.570 ;
        RECT 47.720 181.530 49.640 181.960 ;
        RECT 55.230 181.430 56.690 181.910 ;
        RECT 99.740 181.830 104.600 182.170 ;
        RECT 107.780 181.650 112.620 181.990 ;
        RECT 45.920 180.900 61.250 181.270 ;
        RECT 63.220 181.190 64.140 181.610 ;
        RECT 103.230 181.340 104.490 181.350 ;
        RECT 99.800 181.000 104.640 181.340 ;
        RECT 103.230 180.990 104.490 181.000 ;
        RECT 45.920 180.220 47.030 180.900 ;
        RECT 52.180 180.510 56.160 180.520 ;
        RECT 47.740 179.620 59.780 180.510 ;
        RECT 60.750 180.500 61.250 180.900 ;
        RECT 107.750 180.820 112.590 181.160 ;
        RECT 67.140 179.790 70.760 180.450 ;
        RECT 99.770 180.270 104.610 180.610 ;
        RECT 99.770 180.260 100.890 180.270 ;
        RECT 67.140 179.780 68.240 179.790 ;
        RECT 34.080 178.420 35.020 178.490 ;
        RECT 44.200 178.480 49.590 179.370 ;
        RECT 50.070 178.610 53.620 178.620 ;
        RECT 63.220 178.610 64.140 179.030 ;
        RECT 96.550 178.820 98.980 180.040 ;
        RECT 99.750 179.440 104.590 179.780 ;
        RECT 104.800 179.150 105.980 180.650 ;
        RECT 107.780 180.370 108.990 180.410 ;
        RECT 107.780 180.030 112.640 180.370 ;
        RECT 107.780 180.010 108.990 180.030 ;
        RECT 107.840 179.250 112.680 179.590 ;
        RECT 121.570 178.820 123.140 179.560 ;
        RECT 123.945 178.835 130.935 179.405 ;
        RECT 34.080 178.380 36.160 178.420 ;
        RECT 34.080 178.350 38.150 178.380 ;
        RECT 39.130 178.350 39.850 178.420 ;
        RECT 34.080 178.070 39.860 178.350 ;
        RECT 34.080 178.050 36.160 178.070 ;
        RECT 34.080 178.020 35.020 178.050 ;
        RECT 37.800 177.980 39.860 178.070 ;
        RECT 39.130 177.850 39.850 177.980 ;
        RECT 50.070 177.970 56.640 178.610 ;
        RECT 57.320 178.120 58.780 178.600 ;
        RECT 96.550 178.590 123.140 178.820 ;
        RECT 50.070 177.950 53.620 177.970 ;
        RECT 36.650 177.620 37.310 177.740 ;
        RECT 34.330 177.610 37.310 177.620 ;
        RECT 34.080 177.220 37.310 177.610 ;
        RECT 34.080 176.890 35.050 177.220 ;
        RECT 36.650 176.940 37.310 177.220 ;
        RECT 46.710 177.570 53.410 177.580 ;
        RECT 46.710 176.610 54.780 177.570 ;
        RECT 67.190 177.330 68.200 177.790 ;
        RECT 93.920 177.660 97.030 178.000 ;
        RECT 98.410 177.740 123.140 178.590 ;
        RECT 123.395 178.025 130.095 178.595 ;
        RECT 62.780 176.680 68.660 177.130 ;
        RECT 46.710 176.600 47.340 176.610 ;
        RECT 52.910 176.600 54.780 176.610 ;
        RECT 57.360 176.430 58.710 176.550 ;
        RECT 47.860 176.360 58.710 176.430 ;
        RECT 47.740 176.060 58.710 176.360 ;
        RECT 47.740 175.360 49.670 176.060 ;
        RECT 57.360 175.970 58.710 176.060 ;
        RECT 63.210 176.020 64.150 176.450 ;
        RECT 55.200 175.420 56.660 175.900 ;
        RECT 47.750 175.320 49.640 175.360 ;
        RECT 59.210 174.790 64.140 175.660 ;
        RECT 93.920 175.440 97.060 177.660 ;
        RECT 121.570 177.580 123.140 177.740 ;
        RECT 67.200 174.770 68.200 175.230 ;
        RECT 27.350 174.360 40.800 174.600 ;
        RECT 51.440 174.500 59.790 174.530 ;
        RECT 27.350 173.210 28.040 174.360 ;
        RECT 40.530 174.190 40.800 174.360 ;
        RECT 34.080 173.850 35.080 173.950 ;
        RECT 39.070 173.880 39.890 173.970 ;
        RECT 40.530 173.910 47.570 174.190 ;
        RECT 41.610 173.900 47.570 173.910 ;
        RECT 34.080 173.840 36.140 173.850 ;
        RECT 37.800 173.840 39.890 173.880 ;
        RECT 34.080 173.530 39.890 173.840 ;
        RECT 34.080 173.480 36.140 173.530 ;
        RECT 37.800 173.510 39.890 173.530 ;
        RECT 39.070 173.470 39.890 173.510 ;
        RECT 36.680 173.040 37.330 173.200 ;
        RECT 42.010 173.040 46.980 173.620 ;
        RECT 36.680 172.640 46.980 173.040 ;
        RECT 47.230 173.290 47.570 173.900 ;
        RECT 47.790 173.870 59.790 174.500 ;
        RECT 96.150 174.130 97.060 175.440 ;
        RECT 98.030 176.580 102.950 176.710 ;
        RECT 98.030 175.340 103.040 176.580 ;
        RECT 106.670 175.960 112.900 177.200 ;
        RECT 101.200 175.260 103.040 175.340 ;
        RECT 47.790 173.600 52.770 173.870 ;
        RECT 54.810 173.630 59.790 173.870 ;
        RECT 52.920 173.290 54.030 173.470 ;
        RECT 47.230 172.790 54.030 173.290 ;
        RECT 36.680 172.590 37.330 172.640 ;
        RECT 38.940 172.310 46.980 172.640 ;
        RECT 46.330 171.490 46.970 172.310 ;
        RECT 50.070 171.950 51.800 172.500 ;
        RECT 52.920 172.140 54.030 172.790 ;
        RECT 54.250 172.560 54.680 173.570 ;
        RECT 63.220 173.510 64.140 173.880 ;
        RECT 92.230 173.270 93.910 173.850 ;
        RECT 87.770 172.860 104.570 173.270 ;
        RECT 57.300 172.110 58.760 172.590 ;
        RECT 67.220 172.180 68.170 172.610 ;
        RECT 87.760 172.560 104.570 172.860 ;
        RECT 46.330 171.480 56.620 171.490 ;
        RECT 46.330 170.920 62.840 171.480 ;
        RECT 63.210 170.940 64.150 171.310 ;
        RECT 55.160 170.580 62.840 170.920 ;
        RECT 68.400 170.770 69.870 172.240 ;
        RECT 87.760 170.930 92.310 172.560 ;
        RECT 111.760 172.340 113.340 173.380 ;
        RECT 98.170 170.580 105.850 170.920 ;
        RECT 123.945 170.735 130.935 171.305 ;
        RECT 44.750 168.940 49.300 170.570 ;
        RECT 89.340 170.020 105.850 170.580 ;
        RECT 106.220 170.190 107.160 170.560 ;
        RECT 89.340 170.010 99.630 170.020 ;
        RECT 89.340 169.190 89.980 170.010 ;
        RECT 44.750 168.640 61.560 168.940 ;
        RECT 44.760 168.230 61.560 168.640 ;
        RECT 49.220 167.650 50.900 168.230 ;
        RECT 68.750 168.120 70.330 169.160 ;
        RECT 79.690 168.860 80.340 168.910 ;
        RECT 81.950 168.860 89.990 169.190 ;
        RECT 93.080 169.000 94.810 169.550 ;
        RECT 79.690 168.460 89.990 168.860 ;
        RECT 79.690 168.300 80.340 168.460 ;
        RECT 77.090 167.970 79.150 168.020 ;
        RECT 82.080 167.990 82.900 168.030 ;
        RECT 80.810 167.970 82.900 167.990 ;
        RECT 77.090 167.660 82.900 167.970 ;
        RECT 85.020 167.880 89.990 168.460 ;
        RECT 95.930 168.030 97.040 169.360 ;
        RECT 97.260 167.930 97.690 168.940 ;
        RECT 100.310 168.910 101.770 169.390 ;
        RECT 110.230 168.890 111.180 169.320 ;
        RECT 111.410 169.260 112.880 170.730 ;
        RECT 123.395 169.925 130.095 170.495 ;
        RECT 77.090 167.650 79.150 167.660 ;
        RECT 77.090 167.550 78.090 167.650 ;
        RECT 80.810 167.620 82.900 167.660 ;
        RECT 82.080 167.530 82.900 167.620 ;
        RECT 90.800 167.630 95.780 167.900 ;
        RECT 97.820 167.630 102.800 167.870 ;
        RECT 53.140 166.060 54.050 167.370 ;
        RECT 90.800 167.000 102.800 167.630 ;
        RECT 106.230 167.620 107.150 167.990 ;
        RECT 94.450 166.970 102.800 167.000 ;
        RECT 58.190 166.160 60.030 166.240 ;
        RECT 50.910 163.840 54.050 166.060 ;
        RECT 55.020 164.920 60.030 166.160 ;
        RECT 90.760 166.140 92.650 166.180 ;
        RECT 55.020 164.790 59.940 164.920 ;
        RECT 63.660 164.300 69.890 165.540 ;
        RECT 90.750 165.440 92.680 166.140 ;
        RECT 98.210 165.600 99.670 166.080 ;
        RECT 102.220 165.840 107.150 166.710 ;
        RECT 110.210 166.270 111.210 166.730 ;
        RECT 100.370 165.440 101.720 165.530 ;
        RECT 90.750 165.140 101.720 165.440 ;
        RECT 90.870 165.070 101.720 165.140 ;
        RECT 100.370 164.950 101.720 165.070 ;
        RECT 106.220 165.050 107.160 165.480 ;
        RECT 89.720 164.890 90.350 164.900 ;
        RECT 95.920 164.890 97.790 164.900 ;
        RECT 77.090 164.280 78.060 164.610 ;
        RECT 79.660 164.280 80.320 164.560 ;
        RECT 77.090 163.890 80.320 164.280 ;
        RECT 89.720 163.930 97.790 164.890 ;
        RECT 116.950 164.850 119.550 167.100 ;
        RECT 105.790 164.370 111.670 164.820 ;
        RECT 89.720 163.920 96.420 163.930 ;
        RECT 77.340 163.880 80.320 163.890 ;
        RECT 50.910 163.500 54.020 163.840 ;
        RECT 79.660 163.760 80.320 163.880 ;
        RECT 110.200 163.710 111.210 164.170 ;
        RECT 82.140 163.520 82.860 163.650 ;
        RECT 93.080 163.530 96.630 163.550 ;
        RECT 77.090 163.450 78.030 163.480 ;
        RECT 77.090 163.430 79.170 163.450 ;
        RECT 80.810 163.430 82.870 163.520 ;
        RECT 77.090 163.150 82.870 163.430 ;
        RECT 77.090 163.120 81.160 163.150 ;
        RECT 77.090 163.080 79.170 163.120 ;
        RECT 82.140 163.080 82.860 163.150 ;
        RECT 77.090 163.010 78.030 163.080 ;
        RECT 56.740 161.720 61.580 162.060 ;
        RECT 56.760 161.230 57.880 161.240 ;
        RECT 56.760 160.890 61.600 161.230 ;
        RECT 61.790 160.850 62.970 162.350 ;
        RECT 64.830 161.910 69.670 162.250 ;
        RECT 87.210 162.130 92.600 163.020 ;
        RECT 93.080 162.890 99.650 163.530 ;
        RECT 100.330 162.900 101.790 163.380 ;
        RECT 93.080 162.880 96.630 162.890 ;
        RECT 106.230 162.470 107.150 162.890 ;
        RECT 123.945 162.635 130.935 163.205 ;
        RECT 64.770 161.470 65.980 161.490 ;
        RECT 64.770 161.130 69.630 161.470 ;
        RECT 64.770 161.090 65.980 161.130 ;
        RECT 60.220 160.500 61.480 160.510 ;
        RECT 56.790 160.160 61.630 160.500 ;
        RECT 64.740 160.340 69.580 160.680 ;
        RECT 60.220 160.150 61.480 160.160 ;
        RECT 72.530 160.060 87.530 160.700 ;
        RECT 88.930 159.930 90.040 161.280 ;
        RECT 90.750 160.990 102.790 161.880 ;
        RECT 110.150 161.710 111.250 161.720 ;
        RECT 110.150 161.050 113.770 161.710 ;
        RECT 115.405 161.260 122.105 161.830 ;
        RECT 123.395 161.825 130.095 162.395 ;
        RECT 95.190 160.980 99.170 160.990 ;
        RECT 114.565 160.450 121.555 161.020 ;
        RECT 79.640 159.860 80.580 159.920 ;
        RECT 82.000 159.860 82.630 159.900 ;
        RECT 56.730 159.330 61.590 159.670 ;
        RECT 64.770 159.510 69.610 159.850 ;
        RECT 79.640 159.460 82.630 159.860 ;
        RECT 90.730 159.540 92.650 159.970 ;
        RECT 98.240 159.590 99.700 160.070 ;
        RECT 106.230 159.890 107.150 160.310 ;
        RECT 56.730 159.280 57.880 159.330 ;
        RECT 71.780 159.110 72.330 159.380 ;
        RECT 79.640 159.160 80.580 159.460 ;
        RECT 82.000 159.430 82.630 159.460 ;
        RECT 68.220 159.080 69.500 159.100 ;
        RECT 60.210 158.910 61.470 158.920 ;
        RECT 56.750 158.570 61.590 158.910 ;
        RECT 64.720 158.740 69.560 159.080 ;
        RECT 71.770 159.040 78.070 159.110 ;
        RECT 71.770 158.990 78.110 159.040 ;
        RECT 78.730 158.990 81.250 159.010 ;
        RECT 82.190 158.990 82.910 159.070 ;
        RECT 68.220 158.700 69.500 158.740 ;
        RECT 71.770 158.620 82.910 158.990 ;
        RECT 71.770 158.590 78.110 158.620 ;
        RECT 78.730 158.610 81.250 158.620 ;
        RECT 60.210 158.560 61.470 158.570 ;
        RECT 55.570 158.150 56.000 158.520 ;
        RECT 71.780 158.420 72.330 158.590 ;
        RECT 82.190 158.500 82.910 158.620 ;
        RECT 64.750 158.280 65.990 158.290 ;
        RECT 55.570 158.080 57.880 158.150 ;
        RECT 55.570 157.740 61.630 158.080 ;
        RECT 64.750 157.940 69.590 158.280 ;
        RECT 117.990 158.000 118.690 158.870 ;
        RECT 55.570 157.670 57.880 157.740 ;
        RECT 55.570 156.930 56.000 157.670 ;
        RECT 63.200 157.330 63.530 157.350 ;
        RECT 60.680 157.320 63.530 157.330 ;
        RECT 60.210 157.310 63.530 157.320 ;
        RECT 56.690 156.970 63.530 157.310 ;
        RECT 64.800 157.140 69.640 157.480 ;
        RECT 60.210 156.960 63.530 156.970 ;
        RECT 63.200 156.680 63.530 156.960 ;
        RECT 115.405 156.720 122.105 157.290 ;
        RECT 63.200 156.670 66.000 156.680 ;
        RECT 56.710 156.520 57.870 156.550 ;
        RECT 56.700 156.180 61.540 156.520 ;
        RECT 63.200 156.330 69.690 156.670 ;
        RECT 63.200 156.320 66.000 156.330 ;
        RECT 63.200 156.310 65.930 156.320 ;
        RECT 63.200 156.290 63.530 156.310 ;
        RECT 56.710 156.130 57.870 156.180 ;
        RECT 70.340 155.990 70.760 156.130 ;
        RECT 68.220 155.920 70.760 155.990 ;
        RECT 56.680 155.380 61.520 155.720 ;
        RECT 64.850 155.580 70.760 155.920 ;
        RECT 114.565 155.910 121.555 156.480 ;
        RECT 71.780 155.630 72.330 155.800 ;
        RECT 68.220 155.530 70.760 155.580 ;
        RECT 70.340 155.270 70.760 155.530 ;
        RECT 71.770 155.600 78.110 155.630 ;
        RECT 78.730 155.600 81.250 155.610 ;
        RECT 82.190 155.600 82.910 155.720 ;
        RECT 71.770 155.230 82.910 155.600 ;
        RECT 71.770 155.180 78.110 155.230 ;
        RECT 78.730 155.210 81.250 155.230 ;
        RECT 18.360 152.870 19.120 155.020 ;
        RECT 56.720 154.960 57.870 155.000 ;
        RECT 56.720 154.620 61.560 154.960 ;
        RECT 64.870 154.780 69.710 155.120 ;
        RECT 71.770 155.110 78.070 155.180 ;
        RECT 82.190 155.150 82.910 155.230 ;
        RECT 71.780 154.840 72.330 155.110 ;
        RECT 79.640 154.760 80.580 155.060 ;
        RECT 82.000 154.760 82.630 154.790 ;
        RECT 56.720 154.540 57.870 154.620 ;
        RECT 79.640 154.360 82.630 154.760 ;
        RECT 56.740 153.850 61.580 154.190 ;
        RECT 64.840 153.990 69.680 154.330 ;
        RECT 79.640 154.300 80.580 154.360 ;
        RECT 82.000 154.320 82.630 154.360 ;
        RECT 64.840 153.520 65.990 153.530 ;
        RECT 72.530 153.520 87.530 154.160 ;
        RECT 56.770 153.360 57.870 153.400 ;
        RECT 56.770 153.020 61.650 153.360 ;
        RECT 64.840 153.180 69.680 153.520 ;
        RECT 56.770 152.980 57.870 153.020 ;
        RECT 88.930 152.940 90.040 154.290 ;
        RECT 90.730 154.250 92.650 154.680 ;
        RECT 98.240 154.150 99.700 154.630 ;
        RECT 123.945 154.535 130.935 155.105 ;
        RECT 106.230 153.910 107.150 154.330 ;
        RECT 123.395 153.725 130.095 154.295 ;
        RECT 95.190 153.230 99.170 153.240 ;
        RECT 56.800 152.220 61.640 152.560 ;
        RECT 64.790 152.420 69.630 152.760 ;
        RECT 90.750 152.340 102.790 153.230 ;
        RECT 110.150 152.510 113.770 153.170 ;
        RECT 115.405 152.660 122.105 153.230 ;
        RECT 110.150 152.500 111.250 152.510 ;
        RECT 64.800 151.950 65.990 151.960 ;
        RECT 56.790 151.790 57.870 151.830 ;
        RECT 56.790 151.450 61.640 151.790 ;
        RECT 64.800 151.610 69.640 151.950 ;
        RECT 64.800 151.600 65.990 151.610 ;
        RECT 56.790 151.400 57.870 151.450 ;
        RECT 60.210 150.970 61.470 150.980 ;
        RECT 56.780 150.630 61.620 150.970 ;
        RECT 64.820 150.820 69.660 151.160 ;
        RECT 77.090 151.140 78.030 151.210 ;
        RECT 87.210 151.200 92.600 152.090 ;
        RECT 114.565 151.850 121.555 152.420 ;
        RECT 93.080 151.330 96.630 151.340 ;
        RECT 106.230 151.330 107.150 151.750 ;
        RECT 77.090 151.100 79.170 151.140 ;
        RECT 77.090 151.070 81.160 151.100 ;
        RECT 82.140 151.070 82.860 151.140 ;
        RECT 77.090 150.790 82.870 151.070 ;
        RECT 77.090 150.770 79.170 150.790 ;
        RECT 77.090 150.740 78.030 150.770 ;
        RECT 80.810 150.700 82.870 150.790 ;
        RECT 82.140 150.570 82.860 150.700 ;
        RECT 93.080 150.690 99.650 151.330 ;
        RECT 100.330 150.840 101.790 151.320 ;
        RECT 93.080 150.670 96.630 150.690 ;
        RECT 64.840 150.030 69.680 150.370 ;
        RECT 79.660 150.340 80.320 150.460 ;
        RECT 77.340 150.330 80.320 150.340 ;
        RECT 64.840 150.020 65.990 150.030 ;
        RECT 77.090 149.940 80.320 150.330 ;
        RECT 77.090 149.610 78.060 149.940 ;
        RECT 79.660 149.660 80.320 149.940 ;
        RECT 89.720 150.290 96.420 150.300 ;
        RECT 68.220 149.570 69.490 149.580 ;
        RECT 60.200 147.820 61.460 149.320 ;
        RECT 64.850 149.230 69.690 149.570 ;
        RECT 89.720 149.330 97.790 150.290 ;
        RECT 110.200 150.050 111.210 150.510 ;
        RECT 105.790 149.400 111.670 149.850 ;
        RECT 89.720 149.320 90.350 149.330 ;
        RECT 95.920 149.320 97.790 149.330 ;
        RECT 68.220 149.190 69.490 149.230 ;
        RECT 100.370 149.150 101.720 149.270 ;
        RECT 90.870 149.080 101.720 149.150 ;
        RECT 64.800 148.810 65.980 148.860 ;
        RECT 64.800 148.470 69.680 148.810 ;
        RECT 90.750 148.780 101.720 149.080 ;
        RECT 64.800 148.440 65.980 148.470 ;
        RECT 90.750 148.080 92.680 148.780 ;
        RECT 100.370 148.690 101.720 148.780 ;
        RECT 106.220 148.740 107.160 149.170 ;
        RECT 98.210 148.140 99.670 148.620 ;
        RECT 115.405 148.600 122.105 149.170 ;
        RECT 90.760 148.040 92.650 148.080 ;
        RECT 68.210 147.990 69.490 148.000 ;
        RECT 64.840 147.650 69.680 147.990 ;
        RECT 68.210 147.640 69.490 147.650 ;
        RECT 102.220 147.510 107.150 148.380 ;
        RECT 110.210 147.490 111.210 147.950 ;
        RECT 114.565 147.790 121.555 148.360 ;
        RECT 94.450 147.220 102.800 147.250 ;
        RECT 64.800 147.200 66.000 147.210 ;
        RECT 64.800 146.860 69.690 147.200 ;
        RECT 64.800 146.850 66.000 146.860 ;
        RECT 63.700 146.460 64.540 146.820 ;
        RECT 77.090 146.570 78.090 146.670 ;
        RECT 82.080 146.600 82.900 146.690 ;
        RECT 77.090 146.560 79.150 146.570 ;
        RECT 80.810 146.560 82.900 146.600 ;
        RECT 69.500 146.460 70.170 146.530 ;
        RECT 63.700 145.960 70.170 146.460 ;
        RECT 77.090 146.250 82.900 146.560 ;
        RECT 90.800 146.590 102.800 147.220 ;
        RECT 77.090 146.200 79.150 146.250 ;
        RECT 80.810 146.230 82.900 146.250 ;
        RECT 82.080 146.190 82.900 146.230 ;
        RECT 69.500 145.810 70.170 145.960 ;
        RECT 79.690 145.760 80.340 145.920 ;
        RECT 85.020 145.760 89.990 146.340 ;
        RECT 90.800 146.320 95.780 146.590 ;
        RECT 97.820 146.350 102.800 146.590 ;
        RECT 79.690 145.360 89.990 145.760 ;
        RECT 79.690 145.310 80.340 145.360 ;
        RECT 81.950 145.030 89.990 145.360 ;
        RECT 89.340 144.210 89.980 145.030 ;
        RECT 93.080 144.670 94.810 145.220 ;
        RECT 95.930 144.860 97.040 146.190 ;
        RECT 97.260 145.280 97.690 146.290 ;
        RECT 106.230 146.230 107.150 146.600 ;
        RECT 123.945 146.435 130.935 147.005 ;
        RECT 123.395 145.625 130.095 146.195 ;
        RECT 100.310 144.830 101.770 145.310 ;
        RECT 110.230 144.900 111.180 145.330 ;
        RECT 89.340 144.200 99.630 144.210 ;
        RECT 89.340 143.640 105.850 144.200 ;
        RECT 106.220 143.660 107.160 144.030 ;
        RECT 98.170 143.300 105.850 143.640 ;
        RECT 111.410 143.490 112.880 144.960 ;
        RECT 115.405 144.540 122.105 145.110 ;
        RECT 114.565 143.730 121.555 144.300 ;
        RECT 20.730 141.810 21.410 142.430 ;
        RECT 19.090 131.340 19.700 131.830 ;
        RECT 20.760 131.070 21.380 141.810 ;
        RECT 87.760 141.660 92.310 143.290 ;
        RECT 87.760 141.360 104.570 141.660 ;
        RECT 87.770 140.950 104.570 141.360 ;
        RECT 92.230 140.370 93.910 140.950 ;
        RECT 111.760 140.840 113.340 141.880 ;
        RECT 115.405 140.480 122.105 141.050 ;
        RECT 96.150 138.780 97.060 140.090 ;
        RECT 114.565 139.670 121.555 140.240 ;
        RECT 101.200 138.880 103.040 138.960 ;
        RECT 93.920 136.560 97.060 138.780 ;
        RECT 98.030 137.640 103.040 138.880 ;
        RECT 123.945 138.335 130.935 138.905 ;
        RECT 98.030 137.510 102.950 137.640 ;
        RECT 106.670 137.020 112.900 138.260 ;
        RECT 123.395 137.525 130.095 138.095 ;
        RECT 93.920 136.220 97.030 136.560 ;
        RECT 99.750 134.440 104.590 134.780 ;
        RECT 99.770 133.950 100.890 133.960 ;
        RECT 99.770 133.610 104.610 133.950 ;
        RECT 104.800 133.570 105.980 135.070 ;
        RECT 107.840 134.630 112.680 134.970 ;
        RECT 114.510 134.210 130.960 136.120 ;
        RECT 107.780 134.190 108.990 134.210 ;
        RECT 129.770 134.200 130.960 134.210 ;
        RECT 107.780 133.850 112.640 134.190 ;
        RECT 107.780 133.810 108.990 133.850 ;
        RECT 103.230 133.220 104.490 133.230 ;
        RECT 99.800 132.880 104.640 133.220 ;
        RECT 107.750 133.060 112.590 133.400 ;
        RECT 103.230 132.870 104.490 132.880 ;
        RECT 99.740 132.050 104.600 132.390 ;
        RECT 107.780 132.230 112.620 132.570 ;
        RECT 115.405 132.360 122.105 132.930 ;
        RECT 99.740 132.000 100.890 132.050 ;
        RECT 111.230 131.800 112.510 131.820 ;
        RECT 103.220 131.630 104.480 131.640 ;
        RECT 99.760 131.290 104.600 131.630 ;
        RECT 107.730 131.460 112.570 131.800 ;
        RECT 114.565 131.550 121.555 132.120 ;
        RECT 111.230 131.420 112.510 131.460 ;
        RECT 103.220 131.280 104.480 131.290 ;
        RECT 19.810 130.820 21.380 131.070 ;
        RECT 19.260 130.670 21.380 130.820 ;
        RECT 98.580 130.870 99.010 131.240 ;
        RECT 107.760 131.000 109.000 131.010 ;
        RECT 98.580 130.800 100.890 130.870 ;
        RECT 19.260 130.280 19.810 130.670 ;
        RECT 98.580 130.460 104.640 130.800 ;
        RECT 107.760 130.660 112.600 131.000 ;
        RECT 98.580 130.390 100.890 130.460 ;
        RECT 59.800 129.880 60.990 130.320 ;
        RECT 98.580 129.650 99.010 130.390 ;
        RECT 123.945 130.235 130.935 130.805 ;
        RECT 106.210 130.050 106.540 130.070 ;
        RECT 103.690 130.040 106.540 130.050 ;
        RECT 103.220 130.030 106.540 130.040 ;
        RECT 99.700 129.690 106.540 130.030 ;
        RECT 107.810 129.860 112.650 130.200 ;
        RECT 103.220 129.680 106.540 129.690 ;
        RECT 106.210 129.400 106.540 129.680 ;
        RECT 123.395 129.425 130.095 129.995 ;
        RECT 106.210 129.390 109.010 129.400 ;
        RECT 99.720 129.240 100.880 129.270 ;
        RECT 99.710 128.900 104.550 129.240 ;
        RECT 106.210 129.050 112.700 129.390 ;
        RECT 106.210 129.040 109.010 129.050 ;
        RECT 106.210 129.030 108.940 129.040 ;
        RECT 106.210 129.010 106.540 129.030 ;
        RECT 99.720 128.850 100.880 128.900 ;
        RECT 113.350 128.710 113.770 128.850 ;
        RECT 111.230 128.640 113.770 128.710 ;
        RECT 99.690 128.100 104.530 128.440 ;
        RECT 107.860 128.300 113.770 128.640 ;
        RECT 115.405 128.300 122.105 128.870 ;
        RECT 111.230 128.250 113.770 128.300 ;
        RECT 113.350 127.990 113.770 128.250 ;
        RECT 99.730 127.680 100.880 127.720 ;
        RECT 99.730 127.340 104.570 127.680 ;
        RECT 107.880 127.500 112.720 127.840 ;
        RECT 114.565 127.490 121.555 128.060 ;
        RECT 99.730 127.260 100.880 127.340 ;
        RECT 99.750 126.570 104.590 126.910 ;
        RECT 107.850 126.710 112.690 127.050 ;
        RECT 107.850 126.240 109.000 126.250 ;
        RECT 99.780 126.080 100.880 126.120 ;
        RECT 99.780 125.740 104.660 126.080 ;
        RECT 107.850 125.900 112.690 126.240 ;
        RECT 99.780 125.700 100.880 125.740 ;
        RECT 99.810 124.940 104.650 125.280 ;
        RECT 107.800 125.140 112.640 125.480 ;
        RECT 107.810 124.670 109.000 124.680 ;
        RECT 99.800 124.510 100.880 124.550 ;
        RECT 99.800 124.170 104.650 124.510 ;
        RECT 107.810 124.330 112.650 124.670 ;
        RECT 107.810 124.320 109.000 124.330 ;
        RECT 115.405 124.240 122.105 124.810 ;
        RECT 99.800 124.120 100.880 124.170 ;
        RECT 103.220 123.690 104.480 123.700 ;
        RECT 99.790 123.350 104.630 123.690 ;
        RECT 107.830 123.540 112.670 123.880 ;
        RECT 114.565 123.430 121.555 124.000 ;
        RECT 107.850 122.750 112.690 123.090 ;
        RECT 107.850 122.740 109.000 122.750 ;
        RECT 111.230 122.290 112.500 122.300 ;
        RECT 107.860 121.950 112.700 122.290 ;
        RECT 123.945 122.135 130.935 122.705 ;
        RECT 111.230 121.910 112.500 121.950 ;
        RECT 18.560 120.230 19.840 121.600 ;
        RECT 107.810 121.530 108.990 121.580 ;
        RECT 107.810 121.190 112.690 121.530 ;
        RECT 123.395 121.325 130.095 121.895 ;
        RECT 107.810 121.160 108.990 121.190 ;
        RECT 111.220 120.710 112.500 120.720 ;
        RECT 107.850 120.370 112.690 120.710 ;
        RECT 111.220 120.360 112.500 120.370 ;
        RECT 115.405 120.180 122.105 120.750 ;
        RECT 107.810 119.920 109.010 119.930 ;
        RECT 107.810 119.580 112.700 119.920 ;
        RECT 107.810 119.570 109.010 119.580 ;
        RECT 114.565 119.370 121.555 119.940 ;
        RECT 98.150 119.140 99.020 119.310 ;
        RECT 121.970 119.140 123.460 119.360 ;
        RECT 98.150 117.990 123.460 119.140 ;
        RECT 98.150 117.830 99.020 117.990 ;
        RECT 121.970 117.790 123.460 117.990 ;
        RECT 107.810 117.730 109.010 117.740 ;
        RECT 107.810 117.390 112.700 117.730 ;
        RECT 107.810 117.380 109.010 117.390 ;
        RECT 111.220 116.940 112.500 116.950 ;
        RECT 107.850 116.600 112.690 116.940 ;
        RECT 111.220 116.590 112.500 116.600 ;
        RECT 107.810 116.120 108.990 116.150 ;
        RECT 115.405 116.120 122.105 116.690 ;
        RECT 107.810 115.780 112.690 116.120 ;
        RECT 107.810 115.730 108.990 115.780 ;
        RECT 111.230 115.360 112.500 115.400 ;
        RECT 107.860 115.020 112.700 115.360 ;
        RECT 114.565 115.310 121.555 115.880 ;
        RECT 111.230 115.010 112.500 115.020 ;
        RECT 107.850 114.560 109.000 114.570 ;
        RECT 107.850 114.220 112.690 114.560 ;
        RECT 123.945 114.035 130.935 114.605 ;
        RECT 99.790 113.620 104.630 113.960 ;
        RECT 103.220 113.610 104.480 113.620 ;
        RECT 107.830 113.430 112.670 113.770 ;
        RECT 123.395 113.225 130.095 113.795 ;
        RECT 99.800 113.140 100.880 113.190 ;
        RECT 99.800 112.800 104.650 113.140 ;
        RECT 107.810 112.980 109.000 112.990 ;
        RECT 99.800 112.760 100.880 112.800 ;
        RECT 107.810 112.640 112.650 112.980 ;
        RECT 107.810 112.630 109.000 112.640 ;
        RECT 99.810 112.030 104.650 112.370 ;
        RECT 107.800 111.830 112.640 112.170 ;
        RECT 115.405 112.060 122.105 112.630 ;
        RECT 99.780 111.570 100.880 111.610 ;
        RECT 99.780 111.230 104.660 111.570 ;
        RECT 99.780 111.190 100.880 111.230 ;
        RECT 107.850 111.070 112.690 111.410 ;
        RECT 114.565 111.250 121.555 111.820 ;
        RECT 107.850 111.060 109.000 111.070 ;
        RECT 99.750 110.400 104.590 110.740 ;
        RECT 107.850 110.260 112.690 110.600 ;
        RECT 99.730 109.970 100.880 110.050 ;
        RECT 99.730 109.630 104.570 109.970 ;
        RECT 99.730 109.590 100.880 109.630 ;
        RECT 107.880 109.470 112.720 109.810 ;
        RECT 99.690 108.870 104.530 109.210 ;
        RECT 113.350 109.060 113.770 109.320 ;
        RECT 111.230 109.010 113.770 109.060 ;
        RECT 107.860 108.670 113.770 109.010 ;
        RECT 111.230 108.600 113.770 108.670 ;
        RECT 113.350 108.460 113.770 108.600 ;
        RECT 99.720 108.410 100.880 108.460 ;
        RECT 99.710 108.070 104.550 108.410 ;
        RECT 106.210 108.280 106.540 108.300 ;
        RECT 106.210 108.270 108.940 108.280 ;
        RECT 106.210 108.260 109.010 108.270 ;
        RECT 99.720 108.040 100.880 108.070 ;
        RECT 106.210 107.920 112.700 108.260 ;
        RECT 115.405 108.000 122.105 108.570 ;
        RECT 106.210 107.910 109.010 107.920 ;
        RECT 98.580 106.920 99.010 107.660 ;
        RECT 106.210 107.630 106.540 107.910 ;
        RECT 103.220 107.620 106.540 107.630 ;
        RECT 99.700 107.280 106.540 107.620 ;
        RECT 103.220 107.270 106.540 107.280 ;
        RECT 103.690 107.260 106.540 107.270 ;
        RECT 106.210 107.240 106.540 107.260 ;
        RECT 107.810 107.110 112.650 107.450 ;
        RECT 114.565 107.190 121.555 107.760 ;
        RECT 98.580 106.850 100.890 106.920 ;
        RECT 18.560 105.450 19.960 106.670 ;
        RECT 98.580 106.510 104.640 106.850 ;
        RECT 98.580 106.440 100.890 106.510 ;
        RECT 98.580 106.070 99.010 106.440 ;
        RECT 107.760 106.310 112.600 106.650 ;
        RECT 107.760 106.300 109.000 106.310 ;
        RECT 103.220 106.020 104.480 106.030 ;
        RECT 99.760 105.680 104.600 106.020 ;
        RECT 123.945 105.935 130.935 106.505 ;
        RECT 111.230 105.850 112.510 105.890 ;
        RECT 103.220 105.670 104.480 105.680 ;
        RECT 107.730 105.510 112.570 105.850 ;
        RECT 111.230 105.490 112.510 105.510 ;
        RECT 99.740 105.260 100.890 105.310 ;
        RECT 99.740 104.920 104.600 105.260 ;
        RECT 123.395 105.125 130.095 105.695 ;
        RECT 107.780 104.740 112.620 105.080 ;
        RECT 103.230 104.430 104.490 104.440 ;
        RECT 99.800 104.090 104.640 104.430 ;
        RECT 103.230 104.080 104.490 104.090 ;
        RECT 107.750 103.910 112.590 104.250 ;
        RECT 115.405 103.940 122.105 104.510 ;
        RECT 99.770 103.360 104.610 103.700 ;
        RECT 99.770 103.350 100.890 103.360 ;
        RECT 99.750 102.530 104.590 102.870 ;
        RECT 104.800 102.240 105.980 103.740 ;
        RECT 107.780 103.460 108.990 103.500 ;
        RECT 107.780 103.120 112.640 103.460 ;
        RECT 114.565 103.130 121.555 103.700 ;
        RECT 107.780 103.100 108.990 103.120 ;
        RECT 107.840 102.340 112.680 102.680 ;
        RECT 123.945 101.885 130.935 102.455 ;
        RECT 93.920 100.750 97.030 101.090 ;
        RECT 123.395 101.075 130.095 101.645 ;
        RECT 93.920 98.530 97.060 100.750 ;
        RECT 19.270 96.560 19.820 96.950 ;
        RECT 59.810 96.910 61.000 97.350 ;
        RECT 96.150 97.220 97.060 98.530 ;
        RECT 98.030 99.670 102.950 99.800 ;
        RECT 98.030 98.430 103.040 99.670 ;
        RECT 106.670 99.050 112.900 100.290 ;
        RECT 115.405 99.880 122.105 100.450 ;
        RECT 114.565 99.070 121.555 99.640 ;
        RECT 101.200 98.350 103.040 98.430 ;
        RECT 123.945 97.835 130.935 98.405 ;
        RECT 123.395 97.025 130.095 97.595 ;
        RECT 19.270 96.410 21.390 96.560 ;
        RECT 19.820 96.160 21.390 96.410 ;
        RECT 92.230 96.360 93.910 96.940 ;
        RECT 19.100 95.400 19.710 95.890 ;
        RECT 20.770 85.420 21.390 96.160 ;
        RECT 87.770 95.950 104.570 96.360 ;
        RECT 87.760 95.650 104.570 95.950 ;
        RECT 87.760 94.020 92.310 95.650 ;
        RECT 111.760 95.430 113.340 96.470 ;
        RECT 98.170 93.670 105.850 94.010 ;
        RECT 89.340 93.110 105.850 93.670 ;
        RECT 106.220 93.280 107.160 93.650 ;
        RECT 89.340 93.100 99.630 93.110 ;
        RECT 89.340 92.280 89.980 93.100 ;
        RECT 79.690 91.950 80.340 92.000 ;
        RECT 81.950 91.950 89.990 92.280 ;
        RECT 93.080 92.090 94.810 92.640 ;
        RECT 79.690 91.550 89.990 91.950 ;
        RECT 79.690 91.390 80.340 91.550 ;
        RECT 77.090 91.060 79.150 91.110 ;
        RECT 82.080 91.080 82.900 91.120 ;
        RECT 80.810 91.060 82.900 91.080 ;
        RECT 77.090 90.750 82.900 91.060 ;
        RECT 85.020 90.970 89.990 91.550 ;
        RECT 95.930 91.120 97.040 92.450 ;
        RECT 97.260 91.020 97.690 92.030 ;
        RECT 100.310 92.000 101.770 92.480 ;
        RECT 110.230 91.980 111.180 92.410 ;
        RECT 111.410 92.350 112.880 93.820 ;
        RECT 123.945 93.785 130.935 94.355 ;
        RECT 123.395 92.975 130.095 93.545 ;
        RECT 115.405 91.760 122.105 92.330 ;
        RECT 77.090 90.740 79.150 90.750 ;
        RECT 77.090 90.640 78.090 90.740 ;
        RECT 80.810 90.710 82.900 90.750 ;
        RECT 82.080 90.620 82.900 90.710 ;
        RECT 90.800 90.720 95.780 90.990 ;
        RECT 97.820 90.720 102.800 90.960 ;
        RECT 90.800 90.090 102.800 90.720 ;
        RECT 106.230 90.710 107.150 91.080 ;
        RECT 114.565 90.950 121.555 91.520 ;
        RECT 94.450 90.060 102.800 90.090 ;
        RECT 90.760 89.230 92.650 89.270 ;
        RECT 90.750 88.530 92.680 89.230 ;
        RECT 98.210 88.690 99.670 89.170 ;
        RECT 102.220 88.930 107.150 89.800 ;
        RECT 110.210 89.360 111.210 89.820 ;
        RECT 123.945 89.735 130.935 90.305 ;
        RECT 123.395 88.925 130.095 89.495 ;
        RECT 100.370 88.530 101.720 88.620 ;
        RECT 90.750 88.230 101.720 88.530 ;
        RECT 90.870 88.160 101.720 88.230 ;
        RECT 100.370 88.040 101.720 88.160 ;
        RECT 106.220 88.140 107.160 88.570 ;
        RECT 89.720 87.980 90.350 87.990 ;
        RECT 95.920 87.980 97.790 87.990 ;
        RECT 77.090 87.370 78.060 87.700 ;
        RECT 79.660 87.370 80.320 87.650 ;
        RECT 77.090 86.980 80.320 87.370 ;
        RECT 89.720 87.020 97.790 87.980 ;
        RECT 105.790 87.460 111.670 87.910 ;
        RECT 115.405 87.700 122.105 88.270 ;
        RECT 89.720 87.010 96.420 87.020 ;
        RECT 77.340 86.970 80.320 86.980 ;
        RECT 79.660 86.850 80.320 86.970 ;
        RECT 110.200 86.800 111.210 87.260 ;
        RECT 114.565 86.890 121.555 87.460 ;
        RECT 82.140 86.610 82.860 86.740 ;
        RECT 93.080 86.620 96.630 86.640 ;
        RECT 77.090 86.540 78.030 86.570 ;
        RECT 77.090 86.520 79.170 86.540 ;
        RECT 80.810 86.520 82.870 86.610 ;
        RECT 77.090 86.240 82.870 86.520 ;
        RECT 77.090 86.210 81.160 86.240 ;
        RECT 77.090 86.170 79.170 86.210 ;
        RECT 82.140 86.170 82.860 86.240 ;
        RECT 77.090 86.100 78.030 86.170 ;
        RECT 20.740 84.800 21.420 85.420 ;
        RECT 87.210 85.220 92.600 86.110 ;
        RECT 93.080 85.980 99.650 86.620 ;
        RECT 100.330 85.990 101.790 86.470 ;
        RECT 93.080 85.970 96.630 85.980 ;
        RECT 106.230 85.560 107.150 85.980 ;
        RECT 123.945 85.685 130.935 86.255 ;
        RECT 72.530 83.150 87.530 83.790 ;
        RECT 88.930 83.020 90.040 84.370 ;
        RECT 90.750 84.080 102.790 84.970 ;
        RECT 123.395 84.875 130.095 85.445 ;
        RECT 110.150 84.800 111.250 84.810 ;
        RECT 110.150 84.140 113.770 84.800 ;
        RECT 95.190 84.070 99.170 84.080 ;
        RECT 115.405 83.640 122.105 84.210 ;
        RECT 79.640 82.950 80.580 83.010 ;
        RECT 82.000 82.950 82.630 82.990 ;
        RECT 79.640 82.550 82.630 82.950 ;
        RECT 90.730 82.630 92.650 83.060 ;
        RECT 98.240 82.680 99.700 83.160 ;
        RECT 106.230 82.980 107.150 83.400 ;
        RECT 114.565 82.830 121.555 83.400 ;
        RECT 71.780 82.200 72.330 82.470 ;
        RECT 79.640 82.250 80.580 82.550 ;
        RECT 82.000 82.520 82.630 82.550 ;
        RECT 71.770 82.130 78.070 82.200 ;
        RECT 71.770 82.080 78.110 82.130 ;
        RECT 78.730 82.080 81.250 82.100 ;
        RECT 82.190 82.080 82.910 82.160 ;
        RECT 69.500 81.150 70.070 82.010 ;
        RECT 71.770 81.710 82.910 82.080 ;
        RECT 71.770 81.680 78.110 81.710 ;
        RECT 78.730 81.700 81.250 81.710 ;
        RECT 71.780 81.510 72.330 81.680 ;
        RECT 82.190 81.590 82.910 81.710 ;
        RECT 123.945 81.635 130.935 82.205 ;
        RECT 63.890 80.650 70.070 81.150 ;
        RECT 123.395 80.825 130.095 81.395 ;
        RECT 63.890 80.610 70.060 80.650 ;
        RECT 63.890 79.930 64.520 80.610 ;
        RECT 64.810 80.370 66.010 80.380 ;
        RECT 64.810 80.030 69.700 80.370 ;
        RECT 71.780 80.030 72.330 80.200 ;
        RECT 64.810 80.020 66.010 80.030 ;
        RECT 71.770 80.000 78.110 80.030 ;
        RECT 78.730 80.000 81.250 80.010 ;
        RECT 82.190 80.000 82.910 80.120 ;
        RECT 71.770 79.630 82.910 80.000 ;
        RECT 68.220 79.580 69.500 79.590 ;
        RECT 71.770 79.580 78.110 79.630 ;
        RECT 78.730 79.610 81.250 79.630 ;
        RECT 60.210 77.910 61.470 79.410 ;
        RECT 64.850 79.240 69.690 79.580 ;
        RECT 71.770 79.510 78.070 79.580 ;
        RECT 82.190 79.550 82.910 79.630 ;
        RECT 115.405 79.580 122.105 80.150 ;
        RECT 71.780 79.240 72.330 79.510 ;
        RECT 68.220 79.230 69.500 79.240 ;
        RECT 79.640 79.160 80.580 79.460 ;
        RECT 82.000 79.160 82.630 79.190 ;
        RECT 64.810 78.760 65.990 78.790 ;
        RECT 79.640 78.760 82.630 79.160 ;
        RECT 64.810 78.420 69.690 78.760 ;
        RECT 79.640 78.700 80.580 78.760 ;
        RECT 82.000 78.720 82.630 78.760 ;
        RECT 64.810 78.370 65.990 78.420 ;
        RECT 68.230 78.000 69.500 78.040 ;
        RECT 64.860 77.660 69.700 78.000 ;
        RECT 72.530 77.920 87.530 78.560 ;
        RECT 68.230 77.650 69.500 77.660 ;
        RECT 88.930 77.340 90.040 78.690 ;
        RECT 90.730 78.650 92.650 79.080 ;
        RECT 98.240 78.550 99.700 79.030 ;
        RECT 114.565 78.770 121.555 79.340 ;
        RECT 106.230 78.310 107.150 78.730 ;
        RECT 95.190 77.630 99.170 77.640 ;
        RECT 64.850 77.200 66.000 77.210 ;
        RECT 64.850 76.860 69.690 77.200 ;
        RECT 90.750 76.740 102.790 77.630 ;
        RECT 123.945 77.585 130.935 78.155 ;
        RECT 110.150 76.910 113.770 77.570 ;
        RECT 110.150 76.900 111.250 76.910 ;
        RECT 123.395 76.775 130.095 77.345 ;
        RECT 56.790 76.260 61.630 76.600 ;
        RECT 60.220 76.250 61.480 76.260 ;
        RECT 64.830 76.070 69.670 76.410 ;
        RECT 56.800 75.780 57.880 75.830 ;
        RECT 56.800 75.440 61.650 75.780 ;
        RECT 64.810 75.620 66.000 75.630 ;
        RECT 56.800 75.400 57.880 75.440 ;
        RECT 64.810 75.280 69.650 75.620 ;
        RECT 77.090 75.540 78.030 75.610 ;
        RECT 87.210 75.600 92.600 76.490 ;
        RECT 93.080 75.730 96.630 75.740 ;
        RECT 106.230 75.730 107.150 76.150 ;
        RECT 77.090 75.500 79.170 75.540 ;
        RECT 77.090 75.470 81.160 75.500 ;
        RECT 82.140 75.470 82.860 75.540 ;
        RECT 64.810 75.270 66.000 75.280 ;
        RECT 77.090 75.190 82.870 75.470 ;
        RECT 77.090 75.170 79.170 75.190 ;
        RECT 77.090 75.140 78.030 75.170 ;
        RECT 80.810 75.100 82.870 75.190 ;
        RECT 56.810 74.670 61.650 75.010 ;
        RECT 82.140 74.970 82.860 75.100 ;
        RECT 93.080 75.090 99.650 75.730 ;
        RECT 100.330 75.240 101.790 75.720 ;
        RECT 115.405 75.520 122.105 76.090 ;
        RECT 93.080 75.070 96.630 75.090 ;
        RECT 64.800 74.470 69.640 74.810 ;
        RECT 79.660 74.740 80.320 74.860 ;
        RECT 77.340 74.730 80.320 74.740 ;
        RECT 18.370 72.210 19.130 74.360 ;
        RECT 77.090 74.340 80.320 74.730 ;
        RECT 56.780 74.210 57.880 74.250 ;
        RECT 56.780 73.870 61.660 74.210 ;
        RECT 56.780 73.830 57.880 73.870 ;
        RECT 64.850 73.710 69.690 74.050 ;
        RECT 77.090 74.010 78.060 74.340 ;
        RECT 79.660 74.060 80.320 74.340 ;
        RECT 89.720 74.690 96.420 74.700 ;
        RECT 89.720 73.730 97.790 74.690 ;
        RECT 110.200 74.450 111.210 74.910 ;
        RECT 114.565 74.710 121.555 75.280 ;
        RECT 105.790 73.800 111.670 74.250 ;
        RECT 89.720 73.720 90.350 73.730 ;
        RECT 95.920 73.720 97.790 73.730 ;
        RECT 64.850 73.700 66.000 73.710 ;
        RECT 100.370 73.550 101.720 73.670 ;
        RECT 90.870 73.480 101.720 73.550 ;
        RECT 56.750 73.040 61.590 73.380 ;
        RECT 64.850 72.900 69.690 73.240 ;
        RECT 90.750 73.180 101.720 73.480 ;
        RECT 56.730 72.610 57.880 72.690 ;
        RECT 56.730 72.270 61.570 72.610 ;
        RECT 90.750 72.480 92.680 73.180 ;
        RECT 100.370 73.090 101.720 73.180 ;
        RECT 106.220 73.140 107.160 73.570 ;
        RECT 117.990 73.430 118.690 74.200 ;
        RECT 123.945 73.535 130.935 74.105 ;
        RECT 98.210 72.540 99.670 73.020 ;
        RECT 56.730 72.230 57.880 72.270 ;
        RECT 64.880 72.110 69.720 72.450 ;
        RECT 90.760 72.440 92.650 72.480 ;
        RECT 56.690 71.510 61.530 71.850 ;
        RECT 70.350 71.700 70.770 71.960 ;
        RECT 102.220 71.910 107.150 72.780 ;
        RECT 123.395 72.725 130.095 73.295 ;
        RECT 110.210 71.890 111.210 72.350 ;
        RECT 68.230 71.650 70.770 71.700 ;
        RECT 64.860 71.310 70.770 71.650 ;
        RECT 94.450 71.620 102.800 71.650 ;
        RECT 68.230 71.240 70.770 71.310 ;
        RECT 70.350 71.100 70.770 71.240 ;
        RECT 56.720 71.050 57.880 71.100 ;
        RECT 56.710 70.710 61.550 71.050 ;
        RECT 77.090 70.970 78.090 71.070 ;
        RECT 82.080 71.000 82.900 71.090 ;
        RECT 77.090 70.960 79.150 70.970 ;
        RECT 80.810 70.960 82.900 71.000 ;
        RECT 63.210 70.920 63.540 70.940 ;
        RECT 63.210 70.910 65.940 70.920 ;
        RECT 63.210 70.900 66.010 70.910 ;
        RECT 56.720 70.680 57.880 70.710 ;
        RECT 63.210 70.560 69.700 70.900 ;
        RECT 77.090 70.650 82.900 70.960 ;
        RECT 90.800 70.990 102.800 71.620 ;
        RECT 77.090 70.600 79.150 70.650 ;
        RECT 80.810 70.630 82.900 70.650 ;
        RECT 82.080 70.590 82.900 70.630 ;
        RECT 63.210 70.550 66.010 70.560 ;
        RECT 55.580 69.560 56.010 70.300 ;
        RECT 63.210 70.270 63.540 70.550 ;
        RECT 60.220 70.260 63.540 70.270 ;
        RECT 56.700 69.920 63.540 70.260 ;
        RECT 79.690 70.160 80.340 70.320 ;
        RECT 85.020 70.160 89.990 70.740 ;
        RECT 90.800 70.720 95.780 70.990 ;
        RECT 97.820 70.750 102.800 70.990 ;
        RECT 60.220 69.910 63.540 69.920 ;
        RECT 60.690 69.900 63.540 69.910 ;
        RECT 63.210 69.880 63.540 69.900 ;
        RECT 64.810 69.750 69.650 70.090 ;
        RECT 79.690 69.760 89.990 70.160 ;
        RECT 79.690 69.710 80.340 69.760 ;
        RECT 55.580 69.490 57.890 69.560 ;
        RECT 55.580 69.150 61.640 69.490 ;
        RECT 81.950 69.430 89.990 69.760 ;
        RECT 55.580 69.080 57.890 69.150 ;
        RECT 55.580 68.710 56.010 69.080 ;
        RECT 64.760 68.950 69.600 69.290 ;
        RECT 64.760 68.940 66.000 68.950 ;
        RECT 60.220 68.660 61.480 68.670 ;
        RECT 56.760 68.320 61.600 68.660 ;
        RECT 89.340 68.610 89.980 69.430 ;
        RECT 93.080 69.070 94.810 69.620 ;
        RECT 95.930 69.260 97.050 70.590 ;
        RECT 97.260 69.680 97.690 70.690 ;
        RECT 106.230 70.630 107.150 71.000 ;
        RECT 100.310 69.230 101.770 69.710 ;
        RECT 110.230 69.300 111.180 69.730 ;
        RECT 123.945 69.450 130.935 70.020 ;
        RECT 89.340 68.600 99.630 68.610 ;
        RECT 68.230 68.490 69.510 68.530 ;
        RECT 60.220 68.310 61.480 68.320 ;
        RECT 64.730 68.150 69.570 68.490 ;
        RECT 68.230 68.130 69.510 68.150 ;
        RECT 89.340 68.040 105.850 68.600 ;
        RECT 106.220 68.060 107.160 68.430 ;
        RECT 56.740 67.900 57.890 67.950 ;
        RECT 56.740 67.560 61.600 67.900 ;
        RECT 64.780 67.380 69.620 67.720 ;
        RECT 98.170 67.700 105.850 68.040 ;
        RECT 111.410 67.890 112.880 69.360 ;
        RECT 123.395 68.640 130.095 69.210 ;
        RECT 60.230 67.070 61.490 67.080 ;
        RECT 56.800 66.730 61.640 67.070 ;
        RECT 60.230 66.720 61.490 66.730 ;
        RECT 64.750 66.550 69.590 66.890 ;
        RECT 56.770 66.000 61.610 66.340 ;
        RECT 56.770 65.990 57.890 66.000 ;
        RECT 56.750 65.170 61.590 65.510 ;
        RECT 61.800 64.880 62.980 66.380 ;
        RECT 64.780 66.100 65.990 66.140 ;
        RECT 64.780 65.760 69.640 66.100 ;
        RECT 87.760 66.060 92.310 67.690 ;
        RECT 87.760 65.760 104.570 66.060 ;
        RECT 64.780 65.740 65.990 65.760 ;
        RECT 87.770 65.350 104.570 65.760 ;
        RECT 64.840 64.980 69.680 65.320 ;
        RECT 92.230 64.770 93.910 65.350 ;
        RECT 111.760 65.240 113.340 66.280 ;
        RECT 123.945 65.325 130.935 65.895 ;
        RECT 123.395 64.515 130.095 65.085 ;
        RECT 50.920 63.390 54.030 63.730 ;
        RECT 50.920 61.170 54.060 63.390 ;
        RECT 96.150 63.180 97.060 64.490 ;
        RECT 101.200 63.280 103.040 63.360 ;
        RECT 53.150 59.860 54.060 61.170 ;
        RECT 55.030 62.310 59.950 62.440 ;
        RECT 55.030 61.070 60.040 62.310 ;
        RECT 63.670 61.690 69.900 62.930 ;
        RECT 58.200 60.990 60.040 61.070 ;
        RECT 93.920 60.960 97.060 63.180 ;
        RECT 98.030 62.040 103.040 63.280 ;
        RECT 126.810 62.975 127.510 63.935 ;
        RECT 98.030 61.910 102.950 62.040 ;
        RECT 106.670 61.420 112.900 62.660 ;
        RECT 93.920 60.620 97.030 60.960 ;
        RECT 97.870 60.520 98.830 60.530 ;
        RECT 121.090 60.520 122.870 62.390 ;
        RECT 123.945 60.770 130.935 61.340 ;
        RECT 97.870 60.020 122.870 60.520 ;
        RECT 94.860 59.630 122.870 60.020 ;
        RECT 123.395 59.960 130.095 60.530 ;
        RECT 49.230 59.000 50.910 59.580 ;
        RECT 44.770 58.590 61.570 59.000 ;
        RECT 44.760 58.290 61.570 58.590 ;
        RECT 44.760 56.660 49.310 58.290 ;
        RECT 68.760 58.070 70.340 59.110 ;
        RECT 94.860 58.600 99.230 59.630 ;
        RECT 99.750 58.840 104.590 59.180 ;
        RECT 99.770 58.350 100.890 58.360 ;
        RECT 99.770 58.010 104.610 58.350 ;
        RECT 104.800 57.970 105.980 59.470 ;
        RECT 107.840 59.030 112.680 59.370 ;
        RECT 107.780 58.590 108.990 58.610 ;
        RECT 107.780 58.250 112.640 58.590 ;
        RECT 107.780 58.210 108.990 58.250 ;
        RECT 121.090 58.210 122.870 59.630 ;
        RECT 103.230 57.620 104.490 57.630 ;
        RECT 99.800 57.280 104.640 57.620 ;
        RECT 107.750 57.460 112.590 57.800 ;
        RECT 103.230 57.270 104.490 57.280 ;
        RECT 55.170 56.310 62.850 56.650 ;
        RECT 46.340 55.750 62.850 56.310 ;
        RECT 63.220 55.920 64.160 56.290 ;
        RECT 46.340 55.740 56.630 55.750 ;
        RECT 46.340 54.920 46.980 55.740 ;
        RECT 36.690 54.590 37.340 54.640 ;
        RECT 38.950 54.590 46.990 54.920 ;
        RECT 50.080 54.730 51.810 55.280 ;
        RECT 36.690 54.190 46.990 54.590 ;
        RECT 52.930 54.440 54.040 55.090 ;
        RECT 36.690 54.030 37.340 54.190 ;
        RECT 27.360 52.870 28.050 54.020 ;
        RECT 34.090 53.700 36.150 53.750 ;
        RECT 39.080 53.720 39.900 53.760 ;
        RECT 37.810 53.700 39.900 53.720 ;
        RECT 34.090 53.390 39.900 53.700 ;
        RECT 42.020 53.610 46.990 54.190 ;
        RECT 47.240 53.940 54.040 54.440 ;
        RECT 34.090 53.380 36.150 53.390 ;
        RECT 34.090 53.280 35.090 53.380 ;
        RECT 37.810 53.350 39.900 53.390 ;
        RECT 39.080 53.260 39.900 53.350 ;
        RECT 47.240 53.330 47.580 53.940 ;
        RECT 52.930 53.760 54.040 53.940 ;
        RECT 54.260 53.660 54.690 54.670 ;
        RECT 57.310 54.640 58.770 55.120 ;
        RECT 67.230 54.620 68.180 55.050 ;
        RECT 68.410 54.990 69.880 56.460 ;
        RECT 99.740 56.450 104.600 56.790 ;
        RECT 107.780 56.630 112.620 56.970 ;
        RECT 99.740 56.400 100.890 56.450 ;
        RECT 111.230 56.200 112.510 56.220 ;
        RECT 103.220 56.030 104.480 56.040 ;
        RECT 99.760 55.690 104.600 56.030 ;
        RECT 107.730 55.860 112.570 56.200 ;
        RECT 111.230 55.820 112.510 55.860 ;
        RECT 103.220 55.680 104.480 55.690 ;
        RECT 98.580 55.270 99.010 55.640 ;
        RECT 107.760 55.400 109.000 55.410 ;
        RECT 98.580 55.200 100.890 55.270 ;
        RECT 98.580 54.860 104.640 55.200 ;
        RECT 107.760 55.060 112.600 55.400 ;
        RECT 98.580 54.790 100.890 54.860 ;
        RECT 98.580 54.050 99.010 54.790 ;
        RECT 106.210 54.450 106.540 54.470 ;
        RECT 103.690 54.440 106.540 54.450 ;
        RECT 103.220 54.430 106.540 54.440 ;
        RECT 99.700 54.090 106.540 54.430 ;
        RECT 107.810 54.260 112.650 54.600 ;
        RECT 103.220 54.080 106.540 54.090 ;
        RECT 106.210 53.800 106.540 54.080 ;
        RECT 106.210 53.790 109.010 53.800 ;
        RECT 41.620 53.320 47.580 53.330 ;
        RECT 40.540 53.040 47.580 53.320 ;
        RECT 47.800 53.360 52.780 53.630 ;
        RECT 54.820 53.360 59.800 53.600 ;
        RECT 40.540 52.870 40.810 53.040 ;
        RECT 27.360 52.630 40.810 52.870 ;
        RECT 47.800 52.730 59.800 53.360 ;
        RECT 63.230 53.350 64.150 53.720 ;
        RECT 99.720 53.640 100.880 53.670 ;
        RECT 99.710 53.300 104.550 53.640 ;
        RECT 106.210 53.450 112.700 53.790 ;
        RECT 106.210 53.440 109.010 53.450 ;
        RECT 126.020 53.440 128.170 55.180 ;
        RECT 106.210 53.430 108.940 53.440 ;
        RECT 106.210 53.410 106.540 53.430 ;
        RECT 99.720 53.250 100.880 53.300 ;
        RECT 113.350 53.110 113.770 53.250 ;
        RECT 111.230 53.040 113.770 53.110 ;
        RECT 51.450 52.700 59.800 52.730 ;
        RECT 99.690 52.500 104.530 52.840 ;
        RECT 107.860 52.700 113.770 53.040 ;
        RECT 111.230 52.650 113.770 52.700 ;
        RECT 47.760 51.870 49.650 51.910 ;
        RECT 47.750 51.170 49.680 51.870 ;
        RECT 55.210 51.330 56.670 51.810 ;
        RECT 59.220 51.570 64.150 52.440 ;
        RECT 67.210 52.000 68.210 52.460 ;
        RECT 113.350 52.390 113.770 52.650 ;
        RECT 99.730 52.080 100.880 52.120 ;
        RECT 99.730 51.740 104.570 52.080 ;
        RECT 107.880 51.900 112.720 52.240 ;
        RECT 99.730 51.660 100.880 51.740 ;
        RECT 57.370 51.170 58.720 51.260 ;
        RECT 47.750 50.870 58.720 51.170 ;
        RECT 47.870 50.800 58.720 50.870 ;
        RECT 57.370 50.680 58.720 50.800 ;
        RECT 63.220 50.780 64.160 51.210 ;
        RECT 99.750 50.970 104.590 51.310 ;
        RECT 107.850 51.110 112.690 51.450 ;
        RECT 107.850 50.640 109.000 50.650 ;
        RECT 46.720 50.620 47.350 50.630 ;
        RECT 52.920 50.620 54.790 50.630 ;
        RECT 34.090 50.010 35.060 50.340 ;
        RECT 36.660 50.010 37.320 50.290 ;
        RECT 34.090 49.620 37.320 50.010 ;
        RECT 46.720 49.660 54.790 50.620 ;
        RECT 62.790 50.100 68.670 50.550 ;
        RECT 99.780 50.480 100.880 50.520 ;
        RECT 99.780 50.140 104.660 50.480 ;
        RECT 107.850 50.300 112.690 50.640 ;
        RECT 99.780 50.100 100.880 50.140 ;
        RECT 46.720 49.650 53.420 49.660 ;
        RECT 34.340 49.610 37.320 49.620 ;
        RECT 36.660 49.490 37.320 49.610 ;
        RECT 67.200 49.440 68.210 49.900 ;
        RECT 39.140 49.250 39.860 49.380 ;
        RECT 99.810 49.340 104.650 49.680 ;
        RECT 107.800 49.540 112.640 49.880 ;
        RECT 50.080 49.260 53.630 49.280 ;
        RECT 34.090 49.180 35.030 49.210 ;
        RECT 34.090 49.160 36.170 49.180 ;
        RECT 37.810 49.160 39.870 49.250 ;
        RECT 34.090 48.880 39.870 49.160 ;
        RECT 34.090 48.850 38.160 48.880 ;
        RECT 34.090 48.810 36.170 48.850 ;
        RECT 39.140 48.810 39.860 48.880 ;
        RECT 34.090 48.740 35.030 48.810 ;
        RECT 44.210 47.860 49.600 48.750 ;
        RECT 50.080 48.620 56.650 49.260 ;
        RECT 57.330 48.630 58.790 49.110 ;
        RECT 107.810 49.070 109.000 49.080 ;
        RECT 99.800 48.910 100.880 48.950 ;
        RECT 50.080 48.610 53.630 48.620 ;
        RECT 63.230 48.200 64.150 48.620 ;
        RECT 99.800 48.570 104.650 48.910 ;
        RECT 107.810 48.730 112.650 49.070 ;
        RECT 107.810 48.720 109.000 48.730 ;
        RECT 99.800 48.520 100.880 48.570 ;
        RECT 103.220 48.090 104.480 48.100 ;
        RECT 99.790 47.750 104.630 48.090 ;
        RECT 107.830 47.940 112.670 48.280 ;
        RECT 29.530 45.790 44.530 46.430 ;
        RECT 45.930 46.330 47.040 47.010 ;
        RECT 47.750 46.720 59.790 47.610 ;
        RECT 67.150 47.440 68.250 47.450 ;
        RECT 67.150 46.780 70.770 47.440 ;
        RECT 107.850 47.150 112.690 47.490 ;
        RECT 107.850 47.140 109.000 47.150 ;
        RECT 52.190 46.710 56.170 46.720 ;
        RECT 60.760 46.330 61.260 46.730 ;
        RECT 111.230 46.690 112.500 46.700 ;
        RECT 107.860 46.350 112.700 46.690 ;
        RECT 45.930 45.960 61.260 46.330 ;
        RECT 111.230 46.310 112.500 46.350 ;
        RECT 45.930 45.660 47.040 45.960 ;
        RECT 36.640 45.590 37.580 45.650 ;
        RECT 39.000 45.590 39.630 45.630 ;
        RECT 36.640 45.190 39.630 45.590 ;
        RECT 47.730 45.270 49.650 45.700 ;
        RECT 55.240 45.320 56.700 45.800 ;
        RECT 63.230 45.620 64.150 46.040 ;
        RECT 107.810 45.930 108.990 45.980 ;
        RECT 107.810 45.590 112.690 45.930 ;
        RECT 107.810 45.560 108.990 45.590 ;
        RECT 28.780 44.840 29.330 45.110 ;
        RECT 36.640 44.890 37.580 45.190 ;
        RECT 39.000 45.160 39.630 45.190 ;
        RECT 111.220 45.110 112.500 45.120 ;
        RECT 28.770 44.770 35.070 44.840 ;
        RECT 28.770 44.720 35.110 44.770 ;
        RECT 35.730 44.720 38.250 44.740 ;
        RECT 39.190 44.720 39.910 44.800 ;
        RECT 107.850 44.770 112.690 45.110 ;
        RECT 111.220 44.760 112.500 44.770 ;
        RECT 28.770 44.350 39.910 44.720 ;
        RECT 28.770 44.320 35.110 44.350 ;
        RECT 35.730 44.340 38.250 44.350 ;
        RECT 28.780 44.150 29.330 44.320 ;
        RECT 39.190 44.230 39.910 44.350 ;
        RECT 107.810 44.320 109.010 44.330 ;
        RECT 26.950 40.390 28.210 44.140 ;
        RECT 107.810 43.980 112.700 44.320 ;
        RECT 107.810 43.970 109.010 43.980 ;
        RECT 106.100 42.470 107.610 42.480 ;
        RECT 68.610 41.050 107.610 42.470 ;
        RECT 103.210 40.390 104.510 40.760 ;
        RECT 26.950 39.720 104.510 40.390 ;
        RECT 26.950 39.710 104.020 39.720 ;
        RECT 26.950 39.700 28.210 39.710 ;
        RECT 27.920 36.910 30.100 38.880 ;
        RECT 121.860 36.000 123.930 39.110 ;
      LAYER via2 ;
        RECT 71.850 196.940 73.110 199.640 ;
        RECT 102.090 196.920 104.560 197.860 ;
        RECT 130.250 196.900 131.060 199.620 ;
        RECT 107.890 194.330 108.960 194.610 ;
        RECT 111.280 193.530 112.460 193.820 ;
        RECT 62.430 191.630 69.580 193.040 ;
        RECT 107.890 192.720 108.950 193.000 ;
        RECT 111.280 191.980 112.440 192.260 ;
        RECT 107.930 191.180 108.950 191.460 ;
        RECT 103.270 190.560 104.430 190.840 ;
        RECT 111.270 190.390 112.440 190.670 ;
        RECT 99.860 189.720 100.820 190.040 ;
        RECT 107.930 189.580 108.950 189.860 ;
        RECT 103.260 188.980 104.420 189.260 ;
        RECT 111.280 188.770 112.430 189.060 ;
        RECT 99.840 188.150 100.800 188.460 ;
        RECT 107.930 188.020 108.950 188.300 ;
        RECT 126.880 187.960 127.430 188.725 ;
        RECT 103.260 187.350 104.430 187.640 ;
        RECT 111.280 187.220 112.440 187.500 ;
        RECT 99.800 186.550 100.830 186.890 ;
        RECT 107.940 186.430 108.950 186.720 ;
        RECT 103.260 185.800 104.430 186.090 ;
        RECT 111.290 185.620 112.450 185.920 ;
        RECT 99.780 184.980 100.830 185.320 ;
        RECT 107.910 184.860 108.950 185.150 ;
        RECT 103.270 184.230 104.410 184.510 ;
        RECT 111.320 184.040 112.450 184.320 ;
        RECT 99.830 183.440 100.830 183.730 ;
        RECT 107.820 183.240 108.950 183.520 ;
        RECT 103.270 182.620 104.410 182.900 ;
        RECT 111.300 182.470 112.410 182.750 ;
        RECT 47.820 181.560 49.580 181.910 ;
        RECT 55.340 181.460 56.580 181.850 ;
        RECT 99.820 181.890 100.800 182.180 ;
        RECT 107.870 181.700 108.940 181.980 ;
        RECT 46.070 180.470 46.850 181.380 ;
        RECT 60.790 180.590 61.200 181.220 ;
        RECT 63.260 181.240 64.090 181.550 ;
        RECT 103.270 181.030 104.410 181.310 ;
        RECT 111.310 180.870 112.350 181.150 ;
        RECT 52.290 179.680 52.740 180.470 ;
        RECT 59.270 179.700 59.740 180.420 ;
        RECT 67.290 179.950 68.140 180.320 ;
        RECT 99.840 180.310 100.810 180.600 ;
        RECT 47.910 178.620 49.440 179.260 ;
        RECT 63.280 178.670 64.110 178.980 ;
        RECT 103.290 179.490 104.420 179.770 ;
        RECT 104.980 179.260 105.900 180.490 ;
        RECT 107.840 180.070 108.950 180.350 ;
        RECT 111.370 179.280 112.410 179.560 ;
        RECT 50.150 178.060 51.730 178.410 ;
        RECT 55.340 178.040 56.600 178.520 ;
        RECT 57.360 178.200 58.750 178.550 ;
        RECT 54.280 176.660 54.570 177.510 ;
        RECT 67.260 177.390 68.120 177.730 ;
        RECT 57.480 176.010 58.610 176.510 ;
        RECT 63.280 176.080 64.110 176.390 ;
        RECT 47.830 175.570 49.600 175.870 ;
        RECT 55.300 175.450 56.540 175.840 ;
        RECT 94.030 175.740 94.490 177.560 ;
        RECT 59.270 174.850 59.720 175.550 ;
        RECT 63.280 174.920 64.090 175.580 ;
        RECT 67.260 174.850 68.110 175.150 ;
        RECT 52.260 173.650 52.760 174.430 ;
        RECT 59.250 173.680 59.720 174.400 ;
        RECT 98.140 175.520 99.170 176.560 ;
        RECT 111.810 176.110 112.770 177.030 ;
        RECT 63.270 173.550 64.060 173.840 ;
        RECT 50.180 172.060 51.760 172.410 ;
        RECT 53.050 172.270 53.700 172.970 ;
        RECT 54.290 172.610 54.610 173.510 ;
        RECT 57.380 172.210 58.710 172.510 ;
        RECT 67.270 172.230 68.120 172.590 ;
        RECT 50.600 171.050 51.740 171.400 ;
        RECT 55.370 170.820 56.440 171.330 ;
        RECT 62.160 170.680 62.770 171.380 ;
        RECT 63.290 170.950 64.100 171.260 ;
        RECT 68.810 170.930 69.810 172.130 ;
        RECT 87.970 171.160 92.020 172.830 ;
        RECT 103.370 172.700 104.360 173.150 ;
        RECT 111.820 172.410 112.790 173.290 ;
        RECT 44.960 168.670 49.010 170.340 ;
        RECT 93.610 170.100 94.750 170.450 ;
        RECT 98.380 170.170 99.450 170.680 ;
        RECT 105.170 170.120 105.780 170.820 ;
        RECT 106.300 170.240 107.110 170.550 ;
        RECT 60.360 168.350 61.350 168.800 ;
        RECT 68.810 168.210 69.780 169.090 ;
        RECT 93.190 169.090 94.770 169.440 ;
        RECT 96.060 168.530 96.710 169.230 ;
        RECT 111.820 169.370 112.820 170.570 ;
        RECT 100.390 168.990 101.720 169.290 ;
        RECT 110.280 168.910 111.130 169.270 ;
        RECT 97.300 167.990 97.620 168.890 ;
        RECT 95.270 167.070 95.770 167.850 ;
        RECT 102.260 167.100 102.730 167.820 ;
        RECT 106.280 167.660 107.070 167.950 ;
        RECT 51.020 163.940 51.480 165.760 ;
        RECT 55.130 164.940 56.160 165.980 ;
        RECT 90.840 165.630 92.610 165.930 ;
        RECT 68.800 164.470 69.760 165.390 ;
        RECT 98.310 165.660 99.550 166.050 ;
        RECT 102.280 165.950 102.730 166.650 ;
        RECT 106.290 165.920 107.100 166.580 ;
        RECT 110.270 166.350 111.120 166.650 ;
        RECT 100.490 164.990 101.620 165.490 ;
        RECT 106.290 165.110 107.120 165.420 ;
        RECT 117.090 165.150 119.290 166.910 ;
        RECT 97.290 163.990 97.580 164.840 ;
        RECT 110.270 163.770 111.130 164.110 ;
        RECT 93.160 163.090 94.740 163.440 ;
        RECT 98.350 162.980 99.610 163.460 ;
        RECT 100.370 162.950 101.760 163.300 ;
        RECT 60.280 161.730 61.410 162.010 ;
        RECT 56.830 160.900 57.800 161.190 ;
        RECT 61.970 161.010 62.890 162.240 ;
        RECT 68.360 161.940 69.400 162.220 ;
        RECT 90.920 162.240 92.450 162.880 ;
        RECT 106.290 162.520 107.120 162.830 ;
        RECT 64.830 161.150 65.940 161.430 ;
        RECT 60.260 160.190 61.400 160.470 ;
        RECT 68.300 160.350 69.340 160.630 ;
        RECT 89.080 160.120 89.860 161.030 ;
        RECT 95.300 161.030 95.750 161.820 ;
        RECT 102.280 161.080 102.750 161.800 ;
        RECT 110.300 161.180 111.150 161.550 ;
        RECT 56.810 159.320 57.790 159.610 ;
        RECT 64.860 159.520 65.930 159.800 ;
        RECT 90.830 159.590 92.590 159.940 ;
        RECT 98.350 159.650 99.590 160.040 ;
        RECT 106.270 159.950 107.100 160.260 ;
        RECT 60.260 158.600 61.400 158.880 ;
        RECT 68.290 158.750 69.400 159.030 ;
        RECT 56.820 157.770 57.820 158.060 ;
        RECT 64.810 157.980 65.940 158.260 ;
        RECT 118.050 158.050 118.620 158.820 ;
        RECT 60.260 156.990 61.400 157.270 ;
        RECT 68.310 157.180 69.440 157.460 ;
        RECT 56.770 156.180 57.820 156.520 ;
        RECT 64.900 156.350 65.940 156.640 ;
        RECT 60.250 155.410 61.420 155.700 ;
        RECT 68.280 155.580 69.440 155.880 ;
        RECT 18.460 152.970 19.050 154.890 ;
        RECT 56.790 154.610 57.820 154.950 ;
        RECT 64.930 154.780 65.940 155.070 ;
        RECT 60.250 153.860 61.420 154.150 ;
        RECT 68.270 154.000 69.430 154.280 ;
        RECT 90.830 154.280 92.590 154.630 ;
        RECT 98.350 154.180 99.590 154.570 ;
        RECT 56.830 153.040 57.790 153.350 ;
        RECT 64.920 153.200 65.940 153.480 ;
        RECT 89.080 153.190 89.860 154.100 ;
        RECT 106.270 153.960 107.100 154.270 ;
        RECT 60.250 152.240 61.410 152.520 ;
        RECT 68.270 152.440 69.420 152.730 ;
        RECT 95.300 152.400 95.750 153.190 ;
        RECT 102.280 152.420 102.750 153.140 ;
        RECT 110.300 152.670 111.150 153.040 ;
        RECT 56.850 151.460 57.810 151.780 ;
        RECT 64.920 151.640 65.940 151.920 ;
        RECT 90.920 151.340 92.450 151.980 ;
        RECT 106.290 151.390 107.120 151.700 ;
        RECT 60.260 150.660 61.420 150.940 ;
        RECT 68.260 150.830 69.430 151.110 ;
        RECT 93.160 150.780 94.740 151.130 ;
        RECT 98.350 150.760 99.610 151.240 ;
        RECT 100.370 150.920 101.760 151.270 ;
        RECT 64.920 150.040 65.940 150.320 ;
        RECT 68.270 149.240 69.430 149.520 ;
        RECT 97.290 149.380 97.580 150.230 ;
        RECT 110.270 150.110 111.130 150.450 ;
        RECT 60.370 147.940 61.350 149.180 ;
        RECT 64.880 148.500 65.940 148.780 ;
        RECT 100.490 148.730 101.620 149.230 ;
        RECT 106.290 148.800 107.120 149.110 ;
        RECT 90.840 148.290 92.610 148.590 ;
        RECT 98.310 148.170 99.550 148.560 ;
        RECT 68.270 147.680 69.450 147.970 ;
        RECT 102.280 147.570 102.730 148.270 ;
        RECT 106.290 147.640 107.100 148.300 ;
        RECT 110.270 147.570 111.120 147.870 ;
        RECT 64.880 146.890 65.950 147.170 ;
        RECT 69.590 145.930 70.110 146.460 ;
        RECT 95.270 146.370 95.770 147.150 ;
        RECT 102.260 146.400 102.730 147.120 ;
        RECT 106.280 146.270 107.070 146.560 ;
        RECT 93.190 144.780 94.770 145.130 ;
        RECT 96.060 144.990 96.710 145.690 ;
        RECT 97.300 145.330 97.620 146.230 ;
        RECT 100.390 144.930 101.720 145.230 ;
        RECT 110.280 144.950 111.130 145.310 ;
        RECT 93.610 143.770 94.750 144.120 ;
        RECT 98.380 143.540 99.450 144.050 ;
        RECT 105.170 143.400 105.780 144.100 ;
        RECT 106.300 143.670 107.110 143.980 ;
        RECT 111.820 143.650 112.820 144.850 ;
        RECT 19.170 131.450 19.630 131.780 ;
        RECT 87.970 141.390 92.020 143.060 ;
        RECT 103.370 141.070 104.360 141.520 ;
        RECT 111.820 140.930 112.790 141.810 ;
        RECT 94.030 136.660 94.490 138.480 ;
        RECT 98.140 137.660 99.170 138.700 ;
        RECT 111.810 137.190 112.770 138.110 ;
        RECT 103.290 134.450 104.420 134.730 ;
        RECT 99.840 133.620 100.810 133.910 ;
        RECT 104.980 133.730 105.900 134.960 ;
        RECT 111.370 134.660 112.410 134.940 ;
        RECT 107.840 133.870 108.950 134.150 ;
        RECT 103.270 132.910 104.410 133.190 ;
        RECT 111.310 133.070 112.350 133.350 ;
        RECT 99.820 132.040 100.800 132.330 ;
        RECT 107.870 132.240 108.940 132.520 ;
        RECT 103.270 131.320 104.410 131.600 ;
        RECT 111.300 131.470 112.410 131.750 ;
        RECT 19.340 130.380 19.710 130.730 ;
        RECT 99.830 130.490 100.830 130.780 ;
        RECT 107.820 130.700 108.950 130.980 ;
        RECT 59.930 129.920 60.880 130.250 ;
        RECT 103.270 129.710 104.410 129.990 ;
        RECT 111.320 129.900 112.450 130.180 ;
        RECT 99.780 128.900 100.830 129.240 ;
        RECT 107.910 129.070 108.950 129.360 ;
        RECT 103.260 128.130 104.430 128.420 ;
        RECT 111.290 128.300 112.450 128.600 ;
        RECT 99.800 127.330 100.830 127.670 ;
        RECT 107.940 127.500 108.950 127.790 ;
        RECT 103.260 126.580 104.430 126.870 ;
        RECT 111.280 126.720 112.440 127.000 ;
        RECT 99.840 125.760 100.800 126.070 ;
        RECT 107.930 125.920 108.950 126.200 ;
        RECT 103.260 124.960 104.420 125.240 ;
        RECT 111.280 125.160 112.430 125.450 ;
        RECT 99.860 124.180 100.820 124.500 ;
        RECT 107.930 124.360 108.950 124.640 ;
        RECT 103.270 123.380 104.430 123.660 ;
        RECT 111.270 123.550 112.440 123.830 ;
        RECT 107.930 122.760 108.950 123.040 ;
        RECT 111.280 121.960 112.440 122.240 ;
        RECT 18.820 120.450 19.630 121.490 ;
        RECT 107.890 121.220 108.950 121.500 ;
        RECT 111.280 120.400 112.460 120.690 ;
        RECT 107.890 119.610 108.960 119.890 ;
        RECT 107.890 117.420 108.960 117.700 ;
        RECT 111.280 116.620 112.460 116.910 ;
        RECT 107.890 115.810 108.950 116.090 ;
        RECT 111.280 115.070 112.440 115.350 ;
        RECT 107.930 114.270 108.950 114.550 ;
        RECT 103.270 113.650 104.430 113.930 ;
        RECT 111.270 113.480 112.440 113.760 ;
        RECT 99.860 112.810 100.820 113.130 ;
        RECT 107.930 112.670 108.950 112.950 ;
        RECT 103.260 112.070 104.420 112.350 ;
        RECT 111.280 111.860 112.430 112.150 ;
        RECT 99.840 111.240 100.800 111.550 ;
        RECT 107.930 111.110 108.950 111.390 ;
        RECT 103.260 110.440 104.430 110.730 ;
        RECT 111.280 110.310 112.440 110.590 ;
        RECT 99.800 109.640 100.830 109.980 ;
        RECT 107.940 109.520 108.950 109.810 ;
        RECT 103.260 108.890 104.430 109.180 ;
        RECT 111.290 108.710 112.450 109.010 ;
        RECT 99.780 108.070 100.830 108.410 ;
        RECT 107.910 107.950 108.950 108.240 ;
        RECT 103.270 107.320 104.410 107.600 ;
        RECT 111.320 107.130 112.450 107.410 ;
        RECT 18.810 105.630 19.770 106.460 ;
        RECT 99.830 106.530 100.830 106.820 ;
        RECT 107.820 106.330 108.950 106.610 ;
        RECT 103.270 105.710 104.410 105.990 ;
        RECT 111.300 105.560 112.410 105.840 ;
        RECT 99.820 104.980 100.800 105.270 ;
        RECT 107.870 104.790 108.940 105.070 ;
        RECT 103.270 104.120 104.410 104.400 ;
        RECT 111.310 103.960 112.350 104.240 ;
        RECT 99.840 103.400 100.810 103.690 ;
        RECT 103.290 102.580 104.420 102.860 ;
        RECT 104.980 102.350 105.900 103.580 ;
        RECT 107.840 103.160 108.950 103.440 ;
        RECT 111.370 102.370 112.410 102.650 ;
        RECT 94.030 98.830 94.490 100.650 ;
        RECT 59.940 96.980 60.890 97.310 ;
        RECT 98.140 98.610 99.170 99.650 ;
        RECT 111.810 99.200 112.770 100.120 ;
        RECT 19.350 96.500 19.720 96.850 ;
        RECT 19.180 95.450 19.640 95.780 ;
        RECT 87.970 94.250 92.020 95.920 ;
        RECT 103.370 95.790 104.360 96.240 ;
        RECT 111.820 95.500 112.790 96.380 ;
        RECT 93.610 93.190 94.750 93.540 ;
        RECT 98.380 93.260 99.450 93.770 ;
        RECT 105.170 93.210 105.780 93.910 ;
        RECT 106.300 93.330 107.110 93.640 ;
        RECT 93.190 92.180 94.770 92.530 ;
        RECT 96.060 91.620 96.710 92.320 ;
        RECT 111.820 92.460 112.820 93.660 ;
        RECT 100.390 92.080 101.720 92.380 ;
        RECT 110.280 92.000 111.130 92.360 ;
        RECT 97.300 91.080 97.620 91.980 ;
        RECT 95.270 90.160 95.770 90.940 ;
        RECT 102.260 90.190 102.730 90.910 ;
        RECT 106.280 90.750 107.070 91.040 ;
        RECT 90.840 88.720 92.610 89.020 ;
        RECT 98.310 88.750 99.550 89.140 ;
        RECT 102.280 89.040 102.730 89.740 ;
        RECT 106.290 89.010 107.100 89.670 ;
        RECT 110.270 89.440 111.120 89.740 ;
        RECT 100.490 88.080 101.620 88.580 ;
        RECT 106.290 88.200 107.120 88.510 ;
        RECT 97.290 87.080 97.580 87.930 ;
        RECT 110.270 86.860 111.130 87.200 ;
        RECT 93.160 86.180 94.740 86.530 ;
        RECT 98.350 86.070 99.610 86.550 ;
        RECT 100.370 86.040 101.760 86.390 ;
        RECT 90.920 85.330 92.450 85.970 ;
        RECT 106.290 85.610 107.120 85.920 ;
        RECT 89.080 83.210 89.860 84.120 ;
        RECT 95.300 84.120 95.750 84.910 ;
        RECT 102.280 84.170 102.750 84.890 ;
        RECT 110.300 84.270 111.150 84.640 ;
        RECT 90.830 82.680 92.590 83.030 ;
        RECT 98.350 82.740 99.590 83.130 ;
        RECT 106.270 83.040 107.100 83.350 ;
        RECT 69.580 80.710 70.000 81.910 ;
        RECT 64.890 80.060 65.960 80.340 ;
        RECT 60.380 78.050 61.360 79.290 ;
        RECT 68.280 79.260 69.460 79.550 ;
        RECT 64.890 78.450 65.950 78.730 ;
        RECT 68.280 77.710 69.440 77.990 ;
        RECT 90.830 78.680 92.590 79.030 ;
        RECT 98.350 78.580 99.590 78.970 ;
        RECT 89.080 77.590 89.860 78.500 ;
        RECT 106.270 78.360 107.100 78.670 ;
        RECT 64.930 76.910 65.950 77.190 ;
        RECT 95.300 76.800 95.750 77.590 ;
        RECT 102.280 76.820 102.750 77.540 ;
        RECT 110.300 77.070 111.150 77.440 ;
        RECT 60.270 76.290 61.430 76.570 ;
        RECT 68.270 76.120 69.440 76.400 ;
        RECT 56.860 75.450 57.820 75.770 ;
        RECT 90.920 75.740 92.450 76.380 ;
        RECT 106.290 75.790 107.120 76.100 ;
        RECT 64.930 75.310 65.950 75.590 ;
        RECT 93.160 75.180 94.740 75.530 ;
        RECT 98.350 75.160 99.610 75.640 ;
        RECT 100.370 75.320 101.760 75.670 ;
        RECT 60.260 74.710 61.420 74.990 ;
        RECT 68.280 74.500 69.430 74.790 ;
        RECT 18.470 72.340 19.060 74.260 ;
        RECT 56.840 73.880 57.800 74.190 ;
        RECT 64.930 73.750 65.950 74.030 ;
        RECT 97.290 73.780 97.580 74.630 ;
        RECT 110.270 74.510 111.130 74.850 ;
        RECT 60.260 73.080 61.430 73.370 ;
        RECT 68.280 72.950 69.440 73.230 ;
        RECT 100.490 73.130 101.620 73.630 ;
        RECT 106.290 73.200 107.120 73.510 ;
        RECT 118.050 73.520 118.610 74.110 ;
        RECT 90.840 72.690 92.610 72.990 ;
        RECT 56.800 72.280 57.830 72.620 ;
        RECT 98.310 72.570 99.550 72.960 ;
        RECT 64.940 72.160 65.950 72.450 ;
        RECT 102.280 71.970 102.730 72.670 ;
        RECT 106.290 72.040 107.100 72.700 ;
        RECT 60.260 71.530 61.430 71.820 ;
        RECT 110.270 71.970 111.120 72.270 ;
        RECT 68.290 71.350 69.450 71.650 ;
        RECT 56.780 70.710 57.830 71.050 ;
        RECT 64.910 70.590 65.950 70.880 ;
        RECT 95.270 70.770 95.770 71.550 ;
        RECT 60.270 69.960 61.410 70.240 ;
        RECT 102.260 70.800 102.730 71.520 ;
        RECT 106.280 70.670 107.070 70.960 ;
        RECT 68.320 69.770 69.450 70.050 ;
        RECT 56.830 69.170 57.830 69.460 ;
        RECT 64.820 68.970 65.950 69.250 ;
        RECT 60.270 68.350 61.410 68.630 ;
        RECT 93.190 69.180 94.770 69.530 ;
        RECT 96.060 69.390 96.710 70.090 ;
        RECT 97.300 69.730 97.620 70.630 ;
        RECT 100.390 69.330 101.720 69.630 ;
        RECT 110.280 69.350 111.130 69.710 ;
        RECT 68.300 68.200 69.410 68.480 ;
        RECT 93.610 68.170 94.750 68.520 ;
        RECT 56.820 67.620 57.800 67.910 ;
        RECT 98.380 67.940 99.450 68.450 ;
        RECT 105.170 67.800 105.780 68.500 ;
        RECT 106.300 68.070 107.110 68.380 ;
        RECT 111.820 68.050 112.820 69.250 ;
        RECT 64.870 67.430 65.940 67.710 ;
        RECT 60.270 66.760 61.410 67.040 ;
        RECT 68.310 66.600 69.350 66.880 ;
        RECT 56.840 66.040 57.810 66.330 ;
        RECT 60.290 65.220 61.420 65.500 ;
        RECT 61.980 64.990 62.900 66.220 ;
        RECT 64.840 65.800 65.950 66.080 ;
        RECT 87.970 65.790 92.020 67.460 ;
        RECT 103.370 65.470 104.360 65.920 ;
        RECT 68.370 65.010 69.410 65.290 ;
        RECT 111.820 65.330 112.790 66.210 ;
        RECT 51.030 61.470 51.490 63.290 ;
        RECT 55.140 61.250 56.170 62.290 ;
        RECT 68.810 61.840 69.770 62.760 ;
        RECT 94.030 61.060 94.490 62.880 ;
        RECT 98.140 62.060 99.170 63.100 ;
        RECT 126.870 63.055 127.455 63.825 ;
        RECT 111.810 61.590 112.770 62.510 ;
        RECT 44.970 56.890 49.020 58.560 ;
        RECT 60.370 58.430 61.360 58.880 ;
        RECT 68.820 58.140 69.790 59.020 ;
        RECT 103.290 58.850 104.420 59.130 ;
        RECT 99.840 58.020 100.810 58.310 ;
        RECT 104.980 58.130 105.900 59.360 ;
        RECT 111.370 59.060 112.410 59.340 ;
        RECT 107.840 58.270 108.950 58.550 ;
        RECT 103.270 57.310 104.410 57.590 ;
        RECT 111.310 57.470 112.350 57.750 ;
        RECT 50.610 55.830 51.750 56.180 ;
        RECT 55.380 55.900 56.450 56.410 ;
        RECT 62.170 55.850 62.780 56.550 ;
        RECT 99.820 56.440 100.800 56.730 ;
        RECT 107.870 56.640 108.940 56.920 ;
        RECT 63.300 55.970 64.110 56.280 ;
        RECT 50.190 54.820 51.770 55.170 ;
        RECT 53.060 54.260 53.710 54.960 ;
        RECT 68.820 55.100 69.820 56.300 ;
        RECT 103.270 55.720 104.410 56.000 ;
        RECT 111.300 55.870 112.410 56.150 ;
        RECT 57.390 54.720 58.720 55.020 ;
        RECT 67.280 54.640 68.130 55.000 ;
        RECT 99.830 54.890 100.830 55.180 ;
        RECT 107.820 55.100 108.950 55.380 ;
        RECT 54.300 53.720 54.620 54.620 ;
        RECT 103.270 54.110 104.410 54.390 ;
        RECT 111.320 54.300 112.450 54.580 ;
        RECT 52.270 52.800 52.770 53.580 ;
        RECT 59.260 52.830 59.730 53.550 ;
        RECT 63.280 53.390 64.070 53.680 ;
        RECT 99.780 53.300 100.830 53.640 ;
        RECT 107.910 53.470 108.950 53.760 ;
        RECT 126.230 53.680 127.970 55.000 ;
        RECT 103.260 52.530 104.430 52.820 ;
        RECT 111.290 52.700 112.450 53.000 ;
        RECT 47.840 51.360 49.610 51.660 ;
        RECT 55.310 51.390 56.550 51.780 ;
        RECT 59.280 51.680 59.730 52.380 ;
        RECT 63.290 51.650 64.100 52.310 ;
        RECT 67.270 52.080 68.120 52.380 ;
        RECT 99.800 51.730 100.830 52.070 ;
        RECT 107.940 51.900 108.950 52.190 ;
        RECT 57.490 50.720 58.620 51.220 ;
        RECT 63.290 50.840 64.120 51.150 ;
        RECT 103.260 50.980 104.430 51.270 ;
        RECT 111.280 51.120 112.440 51.400 ;
        RECT 54.290 49.720 54.580 50.570 ;
        RECT 99.840 50.160 100.800 50.470 ;
        RECT 107.930 50.320 108.950 50.600 ;
        RECT 67.270 49.500 68.130 49.840 ;
        RECT 103.260 49.360 104.420 49.640 ;
        RECT 111.280 49.560 112.430 49.850 ;
        RECT 50.160 48.820 51.740 49.170 ;
        RECT 55.350 48.710 56.610 49.190 ;
        RECT 57.370 48.680 58.760 49.030 ;
        RECT 47.920 47.970 49.450 48.610 ;
        RECT 63.290 48.250 64.120 48.560 ;
        RECT 99.860 48.580 100.820 48.900 ;
        RECT 107.930 48.760 108.950 49.040 ;
        RECT 103.270 47.780 104.430 48.060 ;
        RECT 111.270 47.950 112.440 48.230 ;
        RECT 46.080 45.850 46.860 46.760 ;
        RECT 52.300 46.760 52.750 47.550 ;
        RECT 59.280 46.810 59.750 47.530 ;
        RECT 67.300 46.910 68.150 47.280 ;
        RECT 107.930 47.160 108.950 47.440 ;
        RECT 60.800 46.010 61.210 46.640 ;
        RECT 111.280 46.360 112.440 46.640 ;
        RECT 47.830 45.320 49.590 45.670 ;
        RECT 55.350 45.380 56.590 45.770 ;
        RECT 63.270 45.680 64.100 45.990 ;
        RECT 107.890 45.620 108.950 45.900 ;
        RECT 111.280 44.800 112.460 45.090 ;
        RECT 107.890 44.010 108.960 44.290 ;
        RECT 69.020 41.130 69.860 42.210 ;
        RECT 103.430 39.860 104.410 40.590 ;
        RECT 28.130 37.230 29.930 38.610 ;
        RECT 122.080 36.240 123.730 38.900 ;
      LAYER met3 ;
        RECT 71.670 196.690 73.270 199.800 ;
        RECT 101.780 196.790 104.760 198.080 ;
        RECT 62.050 191.280 69.880 193.340 ;
        RECT 45.920 180.220 47.030 181.570 ;
        RECT 47.730 180.990 49.650 182.070 ;
        RECT 47.730 175.530 49.640 180.990 ;
        RECT 55.250 180.840 56.640 181.930 ;
        RECT 50.060 171.940 51.810 178.500 ;
        RECT 52.230 173.620 52.800 180.510 ;
        RECT 52.710 171.810 53.820 173.140 ;
        RECT 54.250 172.560 54.780 177.570 ;
        RECT 44.710 168.620 49.300 170.570 ;
        RECT 50.530 169.320 51.800 171.640 ;
        RECT 55.260 170.690 56.630 180.840 ;
        RECT 57.250 178.070 58.860 178.690 ;
        RECT 57.350 177.380 58.750 178.070 ;
        RECT 57.370 172.910 58.740 177.380 ;
        RECT 59.210 173.630 59.780 180.520 ;
        RECT 57.370 172.690 58.750 172.910 ;
        RECT 57.260 172.070 58.850 172.690 ;
        RECT 57.370 171.810 58.750 172.070 ;
        RECT 50.880 169.090 51.800 169.320 ;
        RECT 18.360 152.870 19.120 155.020 ;
        RECT 18.610 132.620 19.110 152.870 ;
        RECT 36.200 146.760 49.600 168.620 ;
        RECT 50.890 167.520 51.800 169.090 ;
        RECT 60.750 168.990 61.250 181.380 ;
        RECT 63.220 172.900 64.140 181.580 ;
        RECT 67.240 180.380 68.160 181.540 ;
        RECT 67.190 179.850 68.250 180.380 ;
        RECT 67.240 177.780 68.160 179.850 ;
        RECT 67.180 177.320 68.200 177.780 ;
        RECT 67.240 175.240 68.160 177.320 ;
        RECT 67.170 174.740 68.210 175.240 ;
        RECT 50.910 163.500 51.800 167.520 ;
        RECT 54.700 160.510 56.240 166.150 ;
        RECT 56.610 150.290 57.870 162.160 ;
        RECT 60.190 160.980 61.550 168.990 ;
        RECT 62.050 162.400 62.840 171.480 ;
        RECT 63.210 170.680 64.140 172.900 ;
        RECT 67.240 172.670 68.160 174.740 ;
        RECT 67.230 170.450 68.160 172.670 ;
        RECT 68.780 172.240 69.880 191.280 ;
        RECT 79.210 172.880 92.610 194.740 ;
        RECT 103.210 192.690 104.500 196.790 ;
        RECT 130.110 196.690 131.170 199.800 ;
        RECT 107.810 194.620 109.010 194.650 ;
        RECT 107.730 194.290 109.010 194.620 ;
        RECT 93.920 173.980 94.810 178.000 ;
        RECT 97.710 175.350 99.250 180.990 ;
        RECT 99.620 179.340 100.880 191.210 ;
        RECT 103.220 180.520 104.480 192.690 ;
        RECT 68.720 164.310 69.880 172.240 ;
        RECT 87.720 170.930 92.310 172.880 ;
        RECT 93.900 172.410 94.810 173.980 ;
        RECT 103.200 172.510 104.560 180.520 ;
        RECT 104.900 179.100 106.080 180.600 ;
        RECT 107.730 179.210 109.000 194.290 ;
        RECT 111.230 193.860 112.500 194.600 ;
        RECT 111.220 193.500 112.500 193.860 ;
        RECT 111.230 179.190 112.500 193.500 ;
        RECT 93.890 172.180 94.810 172.410 ;
        RECT 60.210 147.830 61.470 160.980 ;
        RECT 61.890 160.900 63.070 162.400 ;
        RECT 60.750 147.820 61.250 147.830 ;
        RECT 64.720 147.210 65.990 162.290 ;
        RECT 68.220 148.000 69.490 162.310 ;
        RECT 88.930 159.930 90.040 170.930 ;
        RECT 93.540 169.860 94.810 172.180 ;
        RECT 95.340 169.690 96.820 170.660 ;
        RECT 90.740 160.510 92.650 165.970 ;
        RECT 93.070 163.000 94.820 169.560 ;
        RECT 95.340 168.350 96.830 169.690 ;
        RECT 95.240 160.990 95.810 167.880 ;
        RECT 90.740 159.430 92.660 160.510 ;
        RECT 96.380 158.260 96.830 168.350 ;
        RECT 97.260 163.930 97.790 168.940 ;
        RECT 98.270 160.660 99.640 170.810 ;
        RECT 105.060 170.020 105.850 179.100 ;
        RECT 100.380 169.430 101.760 169.690 ;
        RECT 100.270 168.810 101.860 169.430 ;
        RECT 100.380 168.590 101.760 168.810 ;
        RECT 106.220 168.600 107.150 170.820 ;
        RECT 110.240 168.830 111.170 171.050 ;
        RECT 111.730 169.240 112.890 177.190 ;
        RECT 100.380 164.120 101.750 168.590 ;
        RECT 100.360 163.430 101.760 164.120 ;
        RECT 100.260 162.810 101.870 163.430 ;
        RECT 102.220 160.980 102.790 167.870 ;
        RECT 98.260 159.570 99.650 160.660 ;
        RECT 106.230 159.920 107.150 168.600 ;
        RECT 110.250 166.760 111.170 168.830 ;
        RECT 110.180 166.260 111.220 166.760 ;
        RECT 110.250 164.180 111.170 166.260 ;
        RECT 110.190 163.720 111.210 164.180 ;
        RECT 110.250 161.650 111.170 163.720 ;
        RECT 110.200 161.120 111.260 161.650 ;
        RECT 110.250 159.960 111.170 161.120 ;
        RECT 68.210 147.640 69.490 148.000 ;
        RECT 64.720 146.880 66.000 147.210 ;
        RECT 68.220 146.900 69.490 147.640 ;
        RECT 64.800 146.850 66.000 146.880 ;
        RECT 69.500 145.810 70.170 146.530 ;
        RECT 20.320 145.220 69.120 145.520 ;
        RECT 20.320 132.820 20.620 145.220 ;
        RECT 30.420 145.210 69.120 145.220 ;
        RECT 30.420 145.200 60.800 145.210 ;
        RECT 30.420 145.020 30.890 145.200 ;
        RECT 43.170 145.020 43.630 145.200 ;
        RECT 45.630 145.170 60.800 145.200 ;
        RECT 61.700 145.170 69.120 145.210 ;
        RECT 45.630 145.110 53.690 145.170 ;
        RECT 53.230 145.040 53.690 145.110 ;
        RECT 20.920 144.720 30.010 144.900 ;
        RECT 45.240 144.720 45.540 144.740 ;
        RECT 20.920 144.710 49.220 144.720 ;
        RECT 52.840 144.710 53.140 144.750 ;
        RECT 60.840 144.710 61.380 144.840 ;
        RECT 20.920 144.690 52.380 144.710 ;
        RECT 52.840 144.690 68.350 144.710 ;
        RECT 20.920 144.600 68.350 144.690 ;
        RECT 20.920 144.590 21.490 144.600 ;
        RECT 20.920 133.340 21.220 144.590 ;
        RECT 22.810 144.360 23.360 144.600 ;
        RECT 29.640 144.420 68.350 144.600 ;
        RECT 48.920 144.410 68.350 144.420 ;
        RECT 52.080 144.390 52.950 144.410 ;
        RECT 20.920 133.080 21.260 133.340 ;
        RECT 20.320 132.380 20.660 132.820 ;
        RECT 19.090 131.340 19.700 131.830 ;
        RECT 19.260 130.280 19.810 130.820 ;
        RECT 18.560 120.230 19.840 121.600 ;
        RECT 20.320 115.270 20.620 132.380 ;
        RECT 20.960 131.940 21.260 133.080 ;
        RECT 20.920 131.830 21.260 131.940 ;
        RECT 20.920 131.330 21.420 131.830 ;
        RECT 22.420 131.350 28.820 143.210 ;
        RECT 30.030 131.350 36.430 143.210 ;
        RECT 37.630 131.360 44.030 143.220 ;
        RECT 45.240 131.350 51.640 143.210 ;
        RECT 52.840 131.350 59.240 143.210 ;
        RECT 60.450 131.350 66.850 143.210 ;
        RECT 20.920 116.080 21.220 131.330 ;
        RECT 35.960 130.820 36.370 130.830 ;
        RECT 22.820 130.810 36.990 130.820 ;
        RECT 22.820 130.440 53.370 130.810 ;
        RECT 22.820 130.430 36.990 130.440 ;
        RECT 59.800 130.030 60.990 130.320 ;
        RECT 22.820 129.660 60.990 130.030 ;
        RECT 22.820 129.640 29.040 129.660 ;
        RECT 22.420 117.350 28.820 129.210 ;
        RECT 30.020 117.350 36.420 129.210 ;
        RECT 37.620 117.350 44.020 129.210 ;
        RECT 45.230 117.360 51.630 129.220 ;
        RECT 52.840 117.370 59.240 129.230 ;
        RECT 60.450 117.380 66.850 129.240 ;
        RECT 30.420 116.150 30.880 116.160 ;
        RECT 29.870 116.140 30.890 116.150 ;
        RECT 20.920 116.070 21.380 116.080 ;
        RECT 20.920 116.060 21.670 116.070 ;
        RECT 29.870 116.060 31.190 116.140 ;
        RECT 36.310 116.120 43.630 116.140 ;
        RECT 36.310 116.080 46.100 116.120 ;
        RECT 60.860 116.080 61.350 116.090 ;
        RECT 68.050 116.080 68.350 144.410 ;
        RECT 36.310 116.060 53.090 116.080 ;
        RECT 20.920 116.000 22.800 116.060 ;
        RECT 29.870 116.050 53.720 116.060 ;
        RECT 60.790 116.050 68.350 116.080 ;
        RECT 29.870 116.040 68.350 116.050 ;
        RECT 29.410 116.000 68.350 116.040 ;
        RECT 20.920 115.710 68.350 116.000 ;
        RECT 20.920 115.700 30.880 115.710 ;
        RECT 31.200 115.700 68.350 115.710 ;
        RECT 20.920 115.630 29.910 115.700 ;
        RECT 31.200 115.640 37.080 115.700 ;
        RECT 22.790 115.590 29.910 115.630 ;
        RECT 30.260 115.270 30.880 115.400 ;
        RECT 20.320 115.180 30.880 115.270 ;
        RECT 43.150 115.200 53.690 115.400 ;
        RECT 68.820 115.200 69.120 145.170 ;
        RECT 43.150 115.190 69.120 115.200 ;
        RECT 37.410 115.180 69.120 115.190 ;
        RECT 20.320 114.880 69.120 115.180 ;
        RECT 20.330 112.050 69.130 112.350 ;
        RECT 20.330 111.960 30.890 112.050 ;
        RECT 37.420 112.040 69.130 112.050 ;
        RECT 18.560 105.450 19.960 106.670 ;
        RECT 19.270 96.410 19.820 96.950 ;
        RECT 19.100 95.400 19.710 95.890 ;
        RECT 20.330 94.850 20.630 111.960 ;
        RECT 30.270 111.830 30.890 111.960 ;
        RECT 43.160 112.030 69.130 112.040 ;
        RECT 43.160 111.830 53.700 112.030 ;
        RECT 22.800 111.600 29.920 111.640 ;
        RECT 20.930 111.530 29.920 111.600 ;
        RECT 31.210 111.530 37.090 111.590 ;
        RECT 20.930 111.520 30.890 111.530 ;
        RECT 31.210 111.520 68.360 111.530 ;
        RECT 20.930 111.230 68.360 111.520 ;
        RECT 20.930 111.170 22.810 111.230 ;
        RECT 29.420 111.190 68.360 111.230 ;
        RECT 29.880 111.180 68.360 111.190 ;
        RECT 29.880 111.170 53.730 111.180 ;
        RECT 20.930 111.160 21.680 111.170 ;
        RECT 20.930 111.150 21.390 111.160 ;
        RECT 20.930 95.900 21.230 111.150 ;
        RECT 29.880 111.090 31.200 111.170 ;
        RECT 36.320 111.150 53.100 111.170 ;
        RECT 60.800 111.150 68.360 111.180 ;
        RECT 36.320 111.110 46.110 111.150 ;
        RECT 60.870 111.140 61.360 111.150 ;
        RECT 36.320 111.090 43.640 111.110 ;
        RECT 29.880 111.080 30.900 111.090 ;
        RECT 30.430 111.070 30.890 111.080 ;
        RECT 22.430 98.020 28.830 109.880 ;
        RECT 30.030 98.020 36.430 109.880 ;
        RECT 37.630 98.020 44.030 109.880 ;
        RECT 45.240 98.010 51.640 109.870 ;
        RECT 52.850 98.000 59.250 109.860 ;
        RECT 60.460 97.990 66.860 109.850 ;
        RECT 22.830 97.570 29.050 97.590 ;
        RECT 22.830 97.200 61.000 97.570 ;
        RECT 59.810 96.910 61.000 97.200 ;
        RECT 22.830 96.790 37.000 96.800 ;
        RECT 22.830 96.420 53.380 96.790 ;
        RECT 22.830 96.410 37.000 96.420 ;
        RECT 35.970 96.400 36.380 96.410 ;
        RECT 20.930 95.400 21.430 95.900 ;
        RECT 20.930 95.290 21.270 95.400 ;
        RECT 18.620 74.360 19.120 94.610 ;
        RECT 20.330 94.410 20.670 94.850 ;
        RECT 20.330 82.010 20.630 94.410 ;
        RECT 20.970 94.150 21.270 95.290 ;
        RECT 20.930 93.890 21.270 94.150 ;
        RECT 20.930 82.640 21.230 93.890 ;
        RECT 22.430 84.020 28.830 95.880 ;
        RECT 30.040 84.020 36.440 95.880 ;
        RECT 37.640 84.010 44.040 95.870 ;
        RECT 45.250 84.020 51.650 95.880 ;
        RECT 52.850 84.020 59.250 95.880 ;
        RECT 60.460 84.020 66.860 95.880 ;
        RECT 20.930 82.630 21.500 82.640 ;
        RECT 22.820 82.630 23.370 82.870 ;
        RECT 52.090 82.820 52.960 82.840 ;
        RECT 68.060 82.820 68.360 111.150 ;
        RECT 48.930 82.810 68.360 82.820 ;
        RECT 29.650 82.630 68.360 82.810 ;
        RECT 20.930 82.540 68.360 82.630 ;
        RECT 20.930 82.520 52.390 82.540 ;
        RECT 52.850 82.520 68.360 82.540 ;
        RECT 20.930 82.510 49.230 82.520 ;
        RECT 20.930 82.330 30.020 82.510 ;
        RECT 45.250 82.490 45.550 82.510 ;
        RECT 52.850 82.480 53.150 82.520 ;
        RECT 60.850 82.390 61.390 82.520 ;
        RECT 30.430 82.030 30.900 82.210 ;
        RECT 43.180 82.030 43.640 82.210 ;
        RECT 53.240 82.120 53.700 82.190 ;
        RECT 45.640 82.060 53.700 82.120 ;
        RECT 68.830 82.060 69.130 112.030 ;
        RECT 45.640 82.030 60.810 82.060 ;
        RECT 30.430 82.020 60.810 82.030 ;
        RECT 61.710 82.020 69.130 82.060 ;
        RECT 30.430 82.010 69.130 82.020 ;
        RECT 69.700 82.010 70.050 145.810 ;
        RECT 88.930 143.290 90.040 154.290 ;
        RECT 90.740 153.710 92.660 154.790 ;
        RECT 90.740 148.250 92.650 153.710 ;
        RECT 93.070 144.660 94.820 151.220 ;
        RECT 95.240 146.340 95.810 153.230 ;
        RECT 96.380 145.860 96.830 155.960 ;
        RECT 98.260 153.560 99.650 154.650 ;
        RECT 95.720 145.840 96.830 145.860 ;
        RECT 95.310 144.530 96.830 145.840 ;
        RECT 97.260 145.280 97.790 150.290 ;
        RECT 87.720 141.340 92.310 143.290 ;
        RECT 93.540 142.040 94.810 144.360 ;
        RECT 95.310 143.950 96.810 144.530 ;
        RECT 98.270 143.410 99.640 153.560 ;
        RECT 100.260 150.790 101.870 151.410 ;
        RECT 100.360 150.100 101.760 150.790 ;
        RECT 100.380 145.630 101.750 150.100 ;
        RECT 102.220 146.350 102.790 153.240 ;
        RECT 100.380 145.410 101.760 145.630 ;
        RECT 106.230 145.620 107.150 154.300 ;
        RECT 110.250 153.100 111.170 154.260 ;
        RECT 110.200 152.570 111.260 153.100 ;
        RECT 110.250 150.500 111.170 152.570 ;
        RECT 110.190 150.040 111.210 150.500 ;
        RECT 110.250 147.960 111.170 150.040 ;
        RECT 110.180 147.460 111.220 147.960 ;
        RECT 100.270 144.790 101.860 145.410 ;
        RECT 100.380 144.530 101.760 144.790 ;
        RECT 93.890 141.810 94.810 142.040 ;
        RECT 79.210 119.480 92.610 141.340 ;
        RECT 93.900 140.240 94.810 141.810 ;
        RECT 93.920 136.220 94.810 140.240 ;
        RECT 97.710 133.230 99.250 138.870 ;
        RECT 99.620 123.010 100.880 134.880 ;
        RECT 103.200 133.700 104.560 141.710 ;
        RECT 105.060 135.120 105.850 144.200 ;
        RECT 106.220 143.400 107.150 145.620 ;
        RECT 110.250 145.390 111.170 147.460 ;
        RECT 110.240 143.170 111.170 145.390 ;
        RECT 111.720 138.260 112.890 169.240 ;
        RECT 116.950 164.850 119.550 167.100 ;
        RECT 111.730 137.030 112.890 138.260 ;
        RECT 103.220 120.230 104.480 133.700 ;
        RECT 104.900 133.620 106.080 135.120 ;
        RECT 107.730 119.930 109.000 135.010 ;
        RECT 111.230 120.720 112.500 135.030 ;
        RECT 111.220 120.360 112.500 120.720 ;
        RECT 107.730 119.600 109.010 119.930 ;
        RECT 111.230 119.620 112.500 120.360 ;
        RECT 107.810 119.570 109.010 119.600 ;
        RECT 79.210 95.970 92.610 117.830 ;
        RECT 107.810 117.710 109.010 117.740 ;
        RECT 103.010 117.080 104.470 117.410 ;
        RECT 107.730 117.380 109.010 117.710 ;
        RECT 103.010 115.830 104.480 117.080 ;
        RECT 93.920 97.070 94.810 101.090 ;
        RECT 97.710 98.440 99.250 104.080 ;
        RECT 99.620 102.430 100.880 114.300 ;
        RECT 103.220 103.610 104.480 115.830 ;
        RECT 87.720 94.020 92.310 95.970 ;
        RECT 93.900 95.500 94.810 97.070 ;
        RECT 103.200 95.600 104.560 103.610 ;
        RECT 104.900 102.190 106.080 103.690 ;
        RECT 107.730 102.300 109.000 117.380 ;
        RECT 111.230 116.950 112.500 117.690 ;
        RECT 111.220 116.590 112.500 116.950 ;
        RECT 111.230 102.280 112.500 116.590 ;
        RECT 93.890 95.270 94.810 95.500 ;
        RECT 88.930 83.020 90.040 94.020 ;
        RECT 93.540 92.950 94.810 95.270 ;
        RECT 95.400 92.780 96.820 93.820 ;
        RECT 90.740 83.600 92.650 89.060 ;
        RECT 93.070 86.090 94.820 92.650 ;
        RECT 95.400 91.540 96.830 92.780 ;
        RECT 95.720 91.450 96.830 91.540 ;
        RECT 95.240 84.080 95.810 90.970 ;
        RECT 90.740 82.520 92.660 83.600 ;
        RECT 20.330 81.710 69.130 82.010 ;
        RECT 69.500 80.650 70.070 82.010 ;
        RECT 96.380 81.350 96.830 91.450 ;
        RECT 97.260 87.020 97.790 92.030 ;
        RECT 98.270 83.750 99.640 93.900 ;
        RECT 105.060 93.110 105.850 102.190 ;
        RECT 100.380 92.520 101.760 92.780 ;
        RECT 100.270 91.900 101.860 92.520 ;
        RECT 100.380 91.680 101.760 91.900 ;
        RECT 106.220 91.690 107.150 93.910 ;
        RECT 110.240 91.920 111.170 94.140 ;
        RECT 100.380 87.210 101.750 91.680 ;
        RECT 100.360 86.520 101.760 87.210 ;
        RECT 100.260 85.900 101.870 86.520 ;
        RECT 102.220 84.070 102.790 90.960 ;
        RECT 98.260 82.660 99.650 83.750 ;
        RECT 106.230 83.010 107.150 91.690 ;
        RECT 110.250 89.850 111.170 91.920 ;
        RECT 111.730 90.350 112.890 100.280 ;
        RECT 110.180 89.350 111.220 89.850 ;
        RECT 110.250 87.270 111.170 89.350 ;
        RECT 110.190 86.810 111.210 87.270 ;
        RECT 110.250 84.740 111.170 86.810 ;
        RECT 110.200 84.210 111.260 84.740 ;
        RECT 110.250 83.050 111.170 84.210 ;
        RECT 69.690 80.610 70.060 80.650 ;
        RECT 18.370 72.210 19.130 74.360 ;
        RECT 36.210 58.610 49.610 80.470 ;
        RECT 64.810 80.350 66.010 80.380 ;
        RECT 64.730 80.020 66.010 80.350 ;
        RECT 60.760 79.400 61.260 79.410 ;
        RECT 50.920 59.710 51.810 63.730 ;
        RECT 54.710 61.080 56.250 66.720 ;
        RECT 56.620 65.070 57.880 76.940 ;
        RECT 60.220 66.250 61.480 79.400 ;
        RECT 44.720 56.660 49.310 58.610 ;
        RECT 50.900 58.140 51.810 59.710 ;
        RECT 60.200 58.240 61.560 66.250 ;
        RECT 61.900 64.830 63.080 66.330 ;
        RECT 64.730 64.940 66.000 80.020 ;
        RECT 68.230 79.590 69.500 80.330 ;
        RECT 68.220 79.230 69.500 79.590 ;
        RECT 68.230 64.920 69.500 79.230 ;
        RECT 88.930 67.690 90.040 78.690 ;
        RECT 90.740 78.110 92.660 79.190 ;
        RECT 90.740 72.650 92.650 78.110 ;
        RECT 93.070 69.060 94.820 75.620 ;
        RECT 95.240 70.740 95.810 77.630 ;
        RECT 96.380 70.270 96.830 80.360 ;
        RECT 98.260 77.960 99.650 79.050 ;
        RECT 87.720 65.740 92.310 67.690 ;
        RECT 93.540 66.440 94.810 68.760 ;
        RECT 95.480 66.900 96.910 70.270 ;
        RECT 97.260 69.680 97.790 74.690 ;
        RECT 98.270 67.810 99.640 77.960 ;
        RECT 100.260 75.190 101.870 75.810 ;
        RECT 100.360 74.500 101.760 75.190 ;
        RECT 100.380 70.030 101.750 74.500 ;
        RECT 102.220 70.750 102.790 77.640 ;
        RECT 100.380 69.810 101.760 70.030 ;
        RECT 106.230 70.020 107.150 78.700 ;
        RECT 110.250 77.500 111.170 78.660 ;
        RECT 110.200 76.970 111.260 77.500 ;
        RECT 110.250 74.900 111.170 76.970 ;
        RECT 110.190 74.440 111.210 74.900 ;
        RECT 110.250 72.360 111.170 74.440 ;
        RECT 110.180 71.860 111.220 72.360 ;
        RECT 100.270 69.190 101.860 69.810 ;
        RECT 100.380 68.930 101.760 69.190 ;
        RECT 93.890 66.210 94.810 66.440 ;
        RECT 50.890 57.910 51.810 58.140 ;
        RECT 50.540 55.590 51.810 57.910 ;
        RECT 45.930 45.660 47.040 47.010 ;
        RECT 47.740 46.240 49.650 51.700 ;
        RECT 50.070 48.730 51.820 55.290 ;
        RECT 52.720 54.090 53.830 55.420 ;
        RECT 52.240 46.720 52.810 53.610 ;
        RECT 54.260 49.660 54.790 54.670 ;
        RECT 55.270 46.390 56.640 56.540 ;
        RECT 57.380 55.160 58.760 55.420 ;
        RECT 57.270 54.540 58.860 55.160 ;
        RECT 57.380 54.320 58.760 54.540 ;
        RECT 57.380 49.850 58.750 54.320 ;
        RECT 57.360 49.160 58.760 49.850 ;
        RECT 57.260 48.540 58.870 49.160 ;
        RECT 59.220 46.710 59.790 53.600 ;
        RECT 47.740 45.160 49.660 46.240 ;
        RECT 55.260 45.300 56.650 46.390 ;
        RECT 60.760 45.850 61.260 58.240 ;
        RECT 62.060 55.750 62.850 64.830 ;
        RECT 68.730 60.470 69.890 62.920 ;
        RECT 63.220 54.330 64.150 56.550 ;
        RECT 67.240 54.560 68.170 56.780 ;
        RECT 68.730 54.990 69.990 60.470 ;
        RECT 63.230 45.650 64.150 54.330 ;
        RECT 67.250 52.490 68.170 54.560 ;
        RECT 67.180 51.990 68.220 52.490 ;
        RECT 67.250 49.910 68.170 51.990 ;
        RECT 67.190 49.450 68.210 49.910 ;
        RECT 67.250 47.380 68.170 49.450 ;
        RECT 67.200 46.850 68.260 47.380 ;
        RECT 67.250 45.690 68.170 46.850 ;
        RECT 68.820 41.030 69.990 54.990 ;
        RECT 79.210 43.880 92.610 65.740 ;
        RECT 93.900 64.640 94.810 66.210 ;
        RECT 93.920 60.620 94.810 64.640 ;
        RECT 97.710 57.630 99.250 63.270 ;
        RECT 99.620 47.410 100.880 59.280 ;
        RECT 103.200 58.100 104.560 66.110 ;
        RECT 105.060 59.520 105.850 68.600 ;
        RECT 106.220 67.800 107.150 70.020 ;
        RECT 110.250 69.790 111.170 71.860 ;
        RECT 110.240 67.570 111.170 69.790 ;
        RECT 111.730 71.360 112.880 90.350 ;
        RECT 117.990 73.430 118.690 158.870 ;
        RECT 111.730 61.430 112.890 71.360 ;
        RECT 126.815 62.940 127.510 188.780 ;
        RECT 138.490 115.740 157.280 117.410 ;
        RECT 103.220 49.300 104.480 58.100 ;
        RECT 104.900 58.020 106.080 59.520 ;
        RECT 103.220 40.760 104.510 49.300 ;
        RECT 107.730 44.330 109.000 59.410 ;
        RECT 111.230 45.120 112.500 59.430 ;
        RECT 126.020 53.440 128.170 55.180 ;
        RECT 111.220 44.760 112.500 45.120 ;
        RECT 107.730 44.000 109.010 44.330 ;
        RECT 111.230 44.020 112.500 44.760 ;
        RECT 107.810 43.970 109.010 44.000 ;
        RECT 103.210 39.720 104.510 40.760 ;
        RECT 27.920 36.910 30.100 38.880 ;
        RECT 121.860 36.000 123.930 39.110 ;
      LAYER via3 ;
        RECT 71.850 196.940 73.110 199.640 ;
        RECT 130.250 196.900 131.060 199.620 ;
        RECT 44.940 168.650 49.050 170.430 ;
        RECT 36.340 168.200 49.460 168.520 ;
        RECT 54.860 160.710 56.010 161.590 ;
        RECT 97.870 179.910 99.020 180.790 ;
        RECT 79.350 172.980 92.470 173.300 ;
        RECT 87.950 171.070 92.060 172.850 ;
        RECT 95.570 168.710 96.610 170.420 ;
        RECT 18.670 132.680 19.040 133.070 ;
        RECT 30.460 145.060 30.850 145.460 ;
        RECT 43.210 145.060 43.600 145.460 ;
        RECT 45.670 145.110 46.060 145.460 ;
        RECT 53.270 145.070 53.660 145.470 ;
        RECT 22.850 144.420 23.310 144.870 ;
        RECT 60.920 144.490 61.330 144.810 ;
        RECT 20.330 132.410 20.650 132.790 ;
        RECT 19.170 131.450 19.630 131.780 ;
        RECT 19.340 130.380 19.710 130.730 ;
        RECT 18.820 120.450 19.630 121.490 ;
        RECT 20.960 131.380 21.380 131.790 ;
        RECT 22.560 131.450 28.680 131.770 ;
        RECT 30.170 131.450 36.290 131.770 ;
        RECT 37.770 131.460 43.890 131.780 ;
        RECT 45.380 131.450 51.500 131.770 ;
        RECT 52.980 131.450 59.100 131.770 ;
        RECT 60.590 131.450 66.710 131.770 ;
        RECT 22.860 130.470 23.970 130.790 ;
        RECT 35.990 130.460 36.360 130.800 ;
        RECT 43.580 130.460 43.950 130.800 ;
        RECT 45.310 130.460 45.680 130.800 ;
        RECT 52.920 130.460 53.310 130.780 ;
        RECT 22.860 129.680 23.970 130.000 ;
        RECT 28.310 129.690 28.710 130.010 ;
        RECT 60.550 129.690 60.950 130.010 ;
        RECT 22.560 128.790 28.680 129.110 ;
        RECT 30.160 128.790 36.280 129.110 ;
        RECT 37.760 128.790 43.880 129.110 ;
        RECT 45.370 128.800 51.490 129.120 ;
        RECT 52.980 128.810 59.100 129.130 ;
        RECT 60.590 128.820 66.710 129.140 ;
        RECT 22.830 115.600 23.240 115.990 ;
        RECT 60.890 115.750 61.350 116.070 ;
        RECT 30.460 114.900 30.840 115.330 ;
        RECT 43.200 114.930 43.580 115.360 ;
        RECT 45.660 114.910 46.040 115.340 ;
        RECT 53.270 114.920 53.650 115.350 ;
        RECT 18.810 105.630 19.770 106.460 ;
        RECT 19.350 96.500 19.720 96.850 ;
        RECT 19.180 95.450 19.640 95.780 ;
        RECT 30.470 111.900 30.850 112.330 ;
        RECT 43.210 111.870 43.590 112.300 ;
        RECT 45.670 111.890 46.050 112.320 ;
        RECT 53.280 111.880 53.660 112.310 ;
        RECT 22.840 111.240 23.250 111.630 ;
        RECT 60.900 111.160 61.360 111.480 ;
        RECT 22.570 98.120 28.690 98.440 ;
        RECT 30.170 98.120 36.290 98.440 ;
        RECT 37.770 98.120 43.890 98.440 ;
        RECT 45.380 98.110 51.500 98.430 ;
        RECT 52.990 98.100 59.110 98.420 ;
        RECT 60.600 98.090 66.720 98.410 ;
        RECT 22.870 97.230 23.980 97.550 ;
        RECT 28.320 97.220 28.720 97.540 ;
        RECT 60.560 97.220 60.960 97.540 ;
        RECT 22.870 96.440 23.980 96.760 ;
        RECT 36.000 96.430 36.370 96.770 ;
        RECT 43.590 96.430 43.960 96.770 ;
        RECT 45.320 96.430 45.690 96.770 ;
        RECT 52.930 96.450 53.320 96.770 ;
        RECT 20.970 95.440 21.390 95.850 ;
        RECT 22.570 95.460 28.690 95.780 ;
        RECT 18.680 94.160 19.050 94.550 ;
        RECT 20.340 94.440 20.660 94.820 ;
        RECT 30.180 95.460 36.300 95.780 ;
        RECT 37.780 95.450 43.900 95.770 ;
        RECT 45.390 95.460 51.510 95.780 ;
        RECT 52.990 95.460 59.110 95.780 ;
        RECT 60.600 95.460 66.720 95.780 ;
        RECT 22.860 82.360 23.320 82.810 ;
        RECT 60.930 82.420 61.340 82.740 ;
        RECT 30.470 81.770 30.860 82.170 ;
        RECT 43.220 81.770 43.610 82.170 ;
        RECT 45.680 81.770 46.070 82.120 ;
        RECT 53.280 81.760 53.670 82.160 ;
        RECT 87.950 141.370 92.060 143.150 ;
        RECT 95.520 144.090 96.690 145.540 ;
        RECT 79.350 140.920 92.470 141.240 ;
        RECT 97.870 133.430 99.020 134.310 ;
        RECT 117.090 165.150 119.290 166.910 ;
        RECT 103.340 121.850 104.350 123.080 ;
        RECT 103.200 116.060 104.280 117.180 ;
        RECT 97.870 103.000 99.020 103.880 ;
        RECT 79.350 96.070 92.470 96.390 ;
        RECT 87.950 94.160 92.060 95.940 ;
        RECT 95.590 91.920 96.550 93.530 ;
        RECT 54.870 65.640 56.020 66.520 ;
        RECT 36.350 58.710 49.470 59.030 ;
        RECT 44.950 56.800 49.060 58.580 ;
        RECT 87.950 65.770 92.060 67.550 ;
        RECT 95.690 67.190 96.740 69.950 ;
        RECT 79.350 65.320 92.470 65.640 ;
        RECT 97.870 57.830 99.020 58.710 ;
        RECT 138.630 116.010 139.460 117.210 ;
        RECT 156.630 115.830 157.020 117.270 ;
        RECT 126.230 53.680 127.970 55.000 ;
        RECT 28.130 37.230 29.930 38.610 ;
        RECT 122.080 36.240 123.730 38.900 ;
      LAYER met4 ;
        RECT 3.990 223.220 4.290 224.760 ;
        RECT 7.670 223.220 7.970 224.760 ;
        RECT 11.350 223.220 11.650 224.760 ;
        RECT 15.030 223.220 15.330 224.760 ;
        RECT 18.710 223.220 19.010 224.760 ;
        RECT 22.390 223.220 22.690 224.760 ;
        RECT 26.070 223.220 26.370 224.760 ;
        RECT 29.750 223.220 30.050 224.760 ;
        RECT 33.430 223.220 33.730 224.760 ;
        RECT 37.110 223.220 37.410 224.760 ;
        RECT 40.790 223.220 41.090 224.760 ;
        RECT 44.470 223.220 44.770 224.760 ;
        RECT 48.150 223.220 48.450 224.760 ;
        RECT 51.830 223.220 52.130 224.760 ;
        RECT 55.510 223.220 55.810 224.760 ;
        RECT 59.190 223.220 59.490 224.760 ;
        RECT 62.870 223.220 63.170 224.760 ;
        RECT 66.550 223.220 66.850 224.760 ;
        RECT 70.230 223.220 70.530 224.760 ;
        RECT 73.910 223.220 74.210 224.760 ;
        RECT 77.590 223.220 77.890 224.760 ;
        RECT 81.270 223.220 81.570 224.760 ;
        RECT 84.950 223.220 85.250 224.760 ;
        RECT 88.630 223.220 88.930 224.760 ;
        RECT 2.970 223.170 89.590 223.220 ;
        RECT 2.970 223.160 147.870 223.170 ;
        RECT 2.970 221.620 147.890 223.160 ;
        RECT 48.080 221.610 51.530 221.620 ;
        RECT 88.700 221.610 147.890 221.620 ;
        RECT 146.390 220.700 147.890 221.610 ;
        RECT 112.380 199.800 146.390 199.810 ;
        RECT 13.980 196.720 146.390 199.800 ;
        RECT 13.980 196.690 131.180 196.720 ;
        RECT 129.330 196.680 131.180 196.690 ;
        RECT 79.600 182.500 92.220 194.350 ;
        RECT 79.600 180.950 95.140 182.500 ;
        RECT 79.600 179.730 99.200 180.950 ;
        RECT 79.600 179.710 95.140 179.730 ;
        RECT 79.600 174.730 92.220 179.710 ;
        RECT 79.240 173.410 91.450 173.550 ;
        RECT 79.240 173.380 92.310 173.410 ;
        RECT 79.240 172.900 92.550 173.380 ;
        RECT 79.240 172.890 92.310 172.900 ;
        RECT 87.760 170.880 92.310 172.890 ;
        RECT 44.750 168.610 49.300 170.620 ;
        RECT 36.230 168.600 49.300 168.610 ;
        RECT 36.230 168.120 49.540 168.600 ;
        RECT 95.340 168.350 96.820 170.660 ;
        RECT 36.230 168.090 49.300 168.120 ;
        RECT 36.230 167.950 48.440 168.090 ;
        RECT 36.590 161.790 49.210 166.770 ;
        RECT 95.800 166.430 96.820 168.350 ;
        RECT 116.950 166.430 119.550 167.100 ;
        RECT 95.800 165.470 119.550 166.430 ;
        RECT 116.950 164.850 119.550 165.470 ;
        RECT 36.590 161.770 52.130 161.790 ;
        RECT 36.590 160.550 56.190 161.770 ;
        RECT 36.590 159.000 52.130 160.550 ;
        RECT 36.590 147.150 49.210 159.000 ;
        RECT 22.810 144.360 23.350 144.900 ;
        RECT 22.810 143.210 23.110 144.360 ;
        RECT 22.810 142.820 23.350 143.210 ;
        RECT 30.430 142.820 30.890 145.520 ;
        RECT 43.170 142.830 43.630 145.530 ;
        RECT 45.630 144.420 46.090 145.520 ;
        RECT 45.630 143.210 45.930 144.420 ;
        RECT 22.810 133.200 28.430 142.820 ;
        RECT 30.420 133.200 36.040 142.820 ;
        RECT 38.020 133.210 43.640 142.830 ;
        RECT 45.630 142.820 46.090 143.210 ;
        RECT 53.230 142.820 53.690 145.520 ;
        RECT 95.310 144.880 96.810 145.840 ;
        RECT 60.840 142.820 61.380 144.840 ;
        RECT 74.480 144.500 96.810 144.880 ;
        RECT 45.630 133.200 51.250 142.820 ;
        RECT 53.230 133.200 58.850 142.820 ;
        RECT 60.840 133.200 66.460 142.820 ;
        RECT 18.610 132.880 19.070 133.120 ;
        RECT 18.610 132.380 20.880 132.880 ;
        RECT 35.970 131.850 36.370 131.860 ;
        RECT 19.090 131.340 21.480 131.830 ;
        RECT 22.480 131.370 28.760 131.850 ;
        RECT 30.090 131.370 36.370 131.850 ;
        RECT 37.690 131.380 43.970 131.860 ;
        RECT 60.510 131.850 60.990 131.880 ;
        RECT 20.360 131.330 21.480 131.340 ;
        RECT 19.260 130.430 24.000 130.820 ;
        RECT 19.260 130.280 19.810 130.430 ;
        RECT 20.370 129.640 24.000 130.030 ;
        RECT 28.280 129.190 28.760 131.370 ;
        RECT 35.970 129.190 36.370 131.370 ;
        RECT 43.560 129.190 43.960 131.380 ;
        RECT 22.480 128.710 28.760 129.190 ;
        RECT 30.080 128.710 36.370 129.190 ;
        RECT 37.680 128.710 43.960 129.190 ;
        RECT 45.290 131.370 51.580 131.850 ;
        RECT 52.900 131.370 59.180 131.850 ;
        RECT 60.510 131.370 66.790 131.850 ;
        RECT 45.290 129.200 45.690 131.370 ;
        RECT 52.910 130.810 53.310 131.370 ;
        RECT 52.910 130.440 53.320 130.810 ;
        RECT 52.910 129.210 53.310 130.440 ;
        RECT 60.510 129.220 60.990 131.370 ;
        RECT 45.290 128.720 51.570 129.200 ;
        RECT 52.900 128.730 59.180 129.210 ;
        RECT 60.510 128.740 66.790 129.220 ;
        RECT 52.910 128.720 53.310 128.730 ;
        RECT 18.560 120.760 19.840 121.600 ;
        RECT 18.560 120.230 19.850 120.760 ;
        RECT 19.470 114.830 19.850 120.230 ;
        RECT 22.810 117.740 28.430 127.360 ;
        RECT 30.410 117.740 36.030 127.360 ;
        RECT 38.010 117.740 43.630 127.360 ;
        RECT 45.620 117.750 51.240 127.370 ;
        RECT 53.230 117.760 58.850 127.380 ;
        RECT 60.820 117.760 66.450 127.390 ;
        RECT 22.810 116.640 23.350 117.740 ;
        RECT 22.800 115.570 23.350 116.640 ;
        RECT 30.420 114.870 30.880 117.740 ;
        RECT 43.160 114.880 43.620 117.740 ;
        RECT 45.620 114.880 46.080 117.750 ;
        RECT 53.230 114.880 53.690 117.760 ;
        RECT 60.840 116.360 61.380 117.760 ;
        RECT 60.840 115.700 61.390 116.360 ;
        RECT 19.470 114.450 29.360 114.830 ;
        RECT 19.470 114.390 19.850 114.450 ;
        RECT 28.980 114.250 29.360 114.450 ;
        RECT 74.480 114.250 74.860 144.500 ;
        RECT 95.310 143.950 96.810 144.500 ;
        RECT 87.760 141.330 92.310 143.340 ;
        RECT 79.240 141.320 92.310 141.330 ;
        RECT 79.240 140.840 92.550 141.320 ;
        RECT 79.240 140.810 92.310 140.840 ;
        RECT 79.240 140.670 91.450 140.810 ;
        RECT 79.600 134.510 92.220 139.490 ;
        RECT 79.600 134.490 95.140 134.510 ;
        RECT 79.600 133.270 99.200 134.490 ;
        RECT 79.600 131.720 95.140 133.270 ;
        RECT 79.600 119.870 92.220 131.720 ;
        RECT 98.930 126.030 101.170 126.130 ;
        RECT 98.730 124.130 133.670 126.030 ;
        RECT 98.930 120.620 101.170 124.130 ;
        RECT 103.240 123.260 133.650 123.270 ;
        RECT 103.240 121.700 142.910 123.260 ;
        RECT 131.790 121.690 142.910 121.700 ;
        RECT 98.930 119.050 133.600 120.620 ;
        RECT 28.980 113.870 74.860 114.250 ;
        RECT 29.330 112.950 68.080 113.120 ;
        RECT 29.330 112.660 74.990 112.950 ;
        RECT 29.330 112.540 30.150 112.660 ;
        RECT 31.190 112.650 74.990 112.660 ;
        RECT 31.190 112.540 42.870 112.650 ;
        RECT 43.930 112.540 45.330 112.650 ;
        RECT 46.390 112.540 52.940 112.650 ;
        RECT 54.000 112.550 74.990 112.650 ;
        RECT 54.000 112.540 67.470 112.550 ;
        RECT 22.210 111.960 24.090 112.390 ;
        RECT 22.210 111.900 22.510 111.960 ;
        RECT 19.510 111.870 19.990 111.880 ;
        RECT 22.180 111.870 22.510 111.900 ;
        RECT 19.510 111.440 22.510 111.870 ;
        RECT 23.660 111.900 24.090 111.960 ;
        RECT 23.660 111.865 24.100 111.900 ;
        RECT 29.330 111.865 29.750 112.540 ;
        RECT 19.510 106.670 19.990 111.440 ;
        RECT 22.810 110.590 23.360 111.660 ;
        RECT 23.660 111.445 29.750 111.865 ;
        RECT 18.560 105.610 19.990 106.670 ;
        RECT 22.820 109.490 23.360 110.590 ;
        RECT 30.430 109.490 30.890 112.360 ;
        RECT 43.170 109.490 43.630 112.350 ;
        RECT 18.560 105.450 19.960 105.610 ;
        RECT 22.820 99.870 28.440 109.490 ;
        RECT 30.420 99.870 36.040 109.490 ;
        RECT 38.020 99.870 43.640 109.490 ;
        RECT 45.630 109.480 46.090 112.350 ;
        RECT 45.630 99.860 51.250 109.480 ;
        RECT 53.240 109.470 53.700 112.350 ;
        RECT 73.640 112.060 74.990 112.550 ;
        RECT 60.850 110.870 61.400 111.530 ;
        RECT 60.850 109.470 61.390 110.870 ;
        RECT 53.240 99.850 58.860 109.470 ;
        RECT 60.830 99.840 66.460 109.470 ;
        RECT 22.490 98.040 28.770 98.520 ;
        RECT 30.090 98.040 36.380 98.520 ;
        RECT 37.690 98.040 43.970 98.520 ;
        RECT 20.380 97.200 24.010 97.590 ;
        RECT 19.270 96.800 19.820 96.950 ;
        RECT 19.270 96.410 24.010 96.800 ;
        RECT 20.370 95.890 21.490 95.900 ;
        RECT 19.100 95.400 21.490 95.890 ;
        RECT 28.290 95.860 28.770 98.040 ;
        RECT 35.980 95.860 36.380 98.040 ;
        RECT 22.490 95.380 28.770 95.860 ;
        RECT 30.100 95.380 36.380 95.860 ;
        RECT 43.570 95.850 43.970 98.040 ;
        RECT 45.300 98.030 51.580 98.510 ;
        RECT 52.920 98.500 53.320 98.510 ;
        RECT 45.300 95.860 45.700 98.030 ;
        RECT 52.910 98.020 59.190 98.500 ;
        RECT 52.920 96.790 53.320 98.020 ;
        RECT 60.520 98.010 66.800 98.490 ;
        RECT 52.920 96.420 53.330 96.790 ;
        RECT 52.920 95.860 53.320 96.420 ;
        RECT 60.520 95.860 61.000 98.010 ;
        RECT 35.980 95.370 36.380 95.380 ;
        RECT 37.700 95.370 43.980 95.850 ;
        RECT 45.300 95.380 51.590 95.860 ;
        RECT 52.910 95.380 59.190 95.860 ;
        RECT 60.520 95.380 66.800 95.860 ;
        RECT 60.520 95.350 61.000 95.380 ;
        RECT 18.620 94.350 20.890 94.850 ;
        RECT 18.620 94.110 19.080 94.350 ;
        RECT 22.820 84.410 28.440 94.030 ;
        RECT 30.430 84.410 36.050 94.030 ;
        RECT 22.820 84.020 23.360 84.410 ;
        RECT 22.820 82.870 23.120 84.020 ;
        RECT 22.820 82.330 23.360 82.870 ;
        RECT 30.440 81.710 30.900 84.410 ;
        RECT 38.030 84.400 43.650 94.020 ;
        RECT 45.640 84.410 51.260 94.030 ;
        RECT 53.240 84.410 58.860 94.030 ;
        RECT 60.850 84.410 66.470 94.030 ;
        RECT 74.260 92.120 74.990 112.060 ;
        RECT 79.600 105.590 92.220 117.440 ;
        RECT 98.930 114.510 101.170 119.050 ;
        RECT 103.010 117.400 104.470 117.410 ;
        RECT 103.010 115.830 139.650 117.400 ;
        RECT 98.930 112.470 133.530 114.510 ;
        RECT 142.030 112.115 142.905 121.690 ;
        RECT 139.790 111.240 142.905 112.115 ;
        RECT 79.600 104.040 95.140 105.590 ;
        RECT 79.600 102.820 99.200 104.040 ;
        RECT 79.600 102.800 95.140 102.820 ;
        RECT 79.600 97.820 92.220 102.800 ;
        RECT 79.240 96.500 91.450 96.640 ;
        RECT 79.240 96.470 92.310 96.500 ;
        RECT 79.240 95.990 92.550 96.470 ;
        RECT 79.240 95.980 92.310 95.990 ;
        RECT 87.760 93.970 92.310 95.980 ;
        RECT 95.400 92.120 96.820 93.820 ;
        RECT 74.240 91.540 96.820 92.120 ;
        RECT 74.240 91.210 96.800 91.540 ;
        RECT 43.180 81.700 43.640 84.400 ;
        RECT 45.640 84.020 46.100 84.410 ;
        RECT 45.640 82.810 45.940 84.020 ;
        RECT 45.640 81.710 46.100 82.810 ;
        RECT 53.240 81.710 53.700 84.410 ;
        RECT 60.850 82.390 61.390 84.410 ;
        RECT 36.600 68.230 49.220 80.080 ;
        RECT 36.600 66.680 52.140 68.230 ;
        RECT 95.480 67.820 96.910 70.270 ;
        RECT 36.600 65.460 56.200 66.680 ;
        RECT 87.760 65.730 92.310 67.740 ;
        RECT 95.430 66.640 115.430 67.820 ;
        RECT 79.240 65.720 92.310 65.730 ;
        RECT 36.600 65.440 52.140 65.460 ;
        RECT 36.600 60.460 49.220 65.440 ;
        RECT 79.240 65.240 92.550 65.720 ;
        RECT 79.240 65.210 92.310 65.240 ;
        RECT 79.240 65.070 91.450 65.210 ;
        RECT 36.240 59.140 48.450 59.280 ;
        RECT 36.240 59.110 49.310 59.140 ;
        RECT 36.240 58.630 49.550 59.110 ;
        RECT 79.600 58.910 92.220 63.890 ;
        RECT 79.600 58.890 95.140 58.910 ;
        RECT 36.240 58.620 49.310 58.630 ;
        RECT 44.760 56.610 49.310 58.620 ;
        RECT 79.600 57.670 99.200 58.890 ;
        RECT 79.600 56.120 95.140 57.670 ;
        RECT 79.600 44.270 92.220 56.120 ;
        RECT 114.500 55.270 115.430 66.640 ;
        RECT 114.500 55.180 128.020 55.270 ;
        RECT 114.500 54.550 128.170 55.180 ;
        RECT 114.590 54.510 128.170 54.550 ;
        RECT 126.020 53.440 128.170 54.510 ;
        RECT 2.500 36.000 132.290 39.110 ;
        RECT 139.790 5.040 140.665 111.240 ;
        RECT 134.345 4.165 140.665 5.040 ;
        RECT 134.345 2.495 135.220 4.165 ;
        RECT 134.355 1.000 135.205 2.495 ;
        RECT 156.535 1.000 157.130 117.850 ;
  END
END tt_um_devinatkin_dual_oscillator
END LIBRARY

