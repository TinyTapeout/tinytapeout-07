MACRO tt_um_brucemack_sb_mixer
  CLASS BLOCK ;
  FOREIGN tt_um_brucemack_sb_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 20.000000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.435600 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 243.321594 ;
    ANTENNADIFFAREA 112.550797 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 62.015 203.875 62.185 204.065 ;
        RECT 63.395 203.875 63.565 204.065 ;
        RECT 68.915 203.875 69.085 204.065 ;
        RECT 74.430 203.925 74.550 204.035 ;
        RECT 75.355 203.875 75.525 204.065 ;
        RECT 80.875 203.875 81.045 204.065 ;
        RECT 86.395 203.875 86.565 204.065 ;
        RECT 88.235 203.875 88.405 204.065 ;
        RECT 91.915 203.875 92.085 204.065 ;
        RECT 94.205 203.875 94.375 204.065 ;
        RECT 95.595 203.875 95.765 204.065 ;
        RECT 61.875 203.065 63.245 203.875 ;
        RECT 63.255 203.065 68.765 203.875 ;
        RECT 68.775 203.065 74.285 203.875 ;
        RECT 74.765 203.005 75.195 203.790 ;
        RECT 75.215 203.065 80.725 203.875 ;
        RECT 80.735 203.065 86.245 203.875 ;
        RECT 86.255 203.065 87.625 203.875 ;
        RECT 87.645 203.005 88.075 203.790 ;
        RECT 88.095 203.065 91.765 203.875 ;
        RECT 91.775 203.065 93.145 203.875 ;
        RECT 93.155 203.095 94.525 203.875 ;
        RECT 94.535 203.065 95.905 203.875 ;
      LAYER nwell ;
        RECT 61.680 199.845 96.100 202.675 ;
      LAYER pwell ;
        RECT 61.875 198.645 63.245 199.455 ;
        RECT 63.255 198.645 68.765 199.455 ;
        RECT 68.775 198.645 74.285 199.455 ;
        RECT 74.765 198.730 75.195 199.515 ;
        RECT 75.675 199.325 76.605 199.555 ;
        RECT 75.675 198.645 78.425 199.325 ;
        RECT 78.905 198.645 80.255 199.555 ;
        RECT 80.285 198.645 81.635 199.555 ;
        RECT 81.655 198.645 83.485 199.455 ;
        RECT 84.050 199.325 84.970 199.555 ;
        RECT 84.050 198.645 87.515 199.325 ;
        RECT 87.635 198.645 93.145 199.455 ;
        RECT 93.155 198.645 94.525 199.455 ;
        RECT 94.535 198.645 95.905 199.455 ;
        RECT 62.015 198.435 62.185 198.645 ;
        RECT 63.395 198.435 63.565 198.645 ;
        RECT 68.915 198.435 69.085 198.645 ;
        RECT 70.750 198.485 70.870 198.595 ;
        RECT 73.515 198.435 73.685 198.625 ;
        RECT 74.430 198.485 74.550 198.595 ;
        RECT 75.350 198.485 75.470 198.595 ;
        RECT 77.650 198.435 77.820 198.625 ;
        RECT 78.115 198.435 78.285 198.645 ;
        RECT 78.570 198.485 78.690 198.595 ;
        RECT 79.035 198.455 79.205 198.645 ;
        RECT 81.335 198.455 81.505 198.645 ;
        RECT 81.795 198.455 81.965 198.645 ;
        RECT 83.630 198.485 83.750 198.595 ;
        RECT 87.315 198.455 87.485 198.645 ;
        RECT 87.775 198.455 87.945 198.645 ;
        RECT 88.235 198.435 88.405 198.625 ;
        RECT 93.295 198.455 93.465 198.645 ;
        RECT 93.765 198.480 93.925 198.590 ;
        RECT 95.595 198.435 95.765 198.645 ;
        RECT 61.875 197.625 63.245 198.435 ;
        RECT 63.255 197.625 68.765 198.435 ;
        RECT 68.775 197.625 70.605 198.435 ;
        RECT 71.085 197.755 73.825 198.435 ;
        RECT 74.075 197.525 77.965 198.435 ;
        RECT 77.975 197.755 87.585 198.435 ;
        RECT 82.485 197.535 83.415 197.755 ;
        RECT 86.245 197.525 87.585 197.755 ;
        RECT 87.645 197.565 88.075 198.350 ;
        RECT 88.095 197.625 93.605 198.435 ;
        RECT 94.535 197.625 95.905 198.435 ;
      LAYER nwell ;
        RECT 61.680 194.405 96.100 197.235 ;
      LAYER pwell ;
        RECT 61.875 193.205 63.245 194.015 ;
        RECT 63.255 193.205 68.765 194.015 ;
        RECT 68.775 193.205 74.285 194.015 ;
        RECT 74.765 193.290 75.195 194.075 ;
        RECT 75.215 193.205 77.045 194.015 ;
        RECT 77.095 193.885 78.435 194.115 ;
        RECT 81.265 193.885 82.195 194.105 ;
        RECT 77.095 193.205 86.705 193.885 ;
        RECT 86.715 193.205 92.225 194.015 ;
        RECT 92.235 193.205 94.065 194.015 ;
        RECT 94.535 193.205 95.905 194.015 ;
        RECT 62.015 192.995 62.185 193.205 ;
        RECT 63.395 192.995 63.565 193.205 ;
        RECT 68.915 192.995 69.085 193.205 ;
        RECT 74.435 193.155 74.605 193.185 ;
        RECT 74.430 193.045 74.605 193.155 ;
        RECT 74.435 192.995 74.605 193.045 ;
        RECT 75.355 193.015 75.525 193.205 ;
        RECT 79.955 192.995 80.125 193.185 ;
        RECT 85.475 192.995 85.645 193.185 ;
        RECT 86.395 193.015 86.565 193.205 ;
        RECT 86.855 193.015 87.025 193.205 ;
        RECT 87.310 193.045 87.430 193.155 ;
        RECT 88.235 192.995 88.405 193.185 ;
        RECT 92.375 193.015 92.545 193.205 ;
        RECT 93.765 193.040 93.925 193.150 ;
        RECT 94.210 193.045 94.330 193.155 ;
        RECT 95.595 192.995 95.765 193.205 ;
        RECT 61.875 192.185 63.245 192.995 ;
        RECT 63.255 192.185 68.765 192.995 ;
        RECT 68.775 192.185 74.285 192.995 ;
        RECT 74.295 192.185 79.805 192.995 ;
        RECT 79.815 192.185 85.325 192.995 ;
        RECT 85.335 192.185 87.165 192.995 ;
        RECT 87.645 192.125 88.075 192.910 ;
        RECT 88.095 192.185 93.605 192.995 ;
        RECT 94.535 192.185 95.905 192.995 ;
      LAYER nwell ;
        RECT 61.680 188.965 96.100 191.795 ;
      LAYER pwell ;
        RECT 61.875 187.765 63.245 188.575 ;
        RECT 63.255 187.765 68.765 188.575 ;
        RECT 68.775 187.765 74.285 188.575 ;
        RECT 74.765 187.850 75.195 188.635 ;
        RECT 75.215 187.765 80.725 188.575 ;
        RECT 80.735 187.765 86.245 188.575 ;
        RECT 86.255 187.765 91.765 188.575 ;
        RECT 91.775 187.765 94.525 188.575 ;
        RECT 94.535 187.765 95.905 188.575 ;
        RECT 62.015 187.555 62.185 187.765 ;
        RECT 63.395 187.555 63.565 187.765 ;
        RECT 68.915 187.555 69.085 187.765 ;
        RECT 74.435 187.715 74.605 187.745 ;
        RECT 74.430 187.605 74.605 187.715 ;
        RECT 74.435 187.555 74.605 187.605 ;
        RECT 75.355 187.575 75.525 187.765 ;
        RECT 79.955 187.555 80.125 187.745 ;
        RECT 80.875 187.575 81.045 187.765 ;
        RECT 85.475 187.555 85.645 187.745 ;
        RECT 86.395 187.575 86.565 187.765 ;
        RECT 87.310 187.605 87.430 187.715 ;
        RECT 88.235 187.555 88.405 187.745 ;
        RECT 91.915 187.575 92.085 187.765 ;
        RECT 93.765 187.600 93.925 187.710 ;
        RECT 95.595 187.555 95.765 187.765 ;
        RECT 61.875 186.745 63.245 187.555 ;
        RECT 63.255 186.745 68.765 187.555 ;
        RECT 68.775 186.745 74.285 187.555 ;
        RECT 74.295 186.745 79.805 187.555 ;
        RECT 79.815 186.745 85.325 187.555 ;
        RECT 85.335 186.745 87.165 187.555 ;
        RECT 87.645 186.685 88.075 187.470 ;
        RECT 88.095 186.745 93.605 187.555 ;
        RECT 94.535 186.745 95.905 187.555 ;
      LAYER nwell ;
        RECT 61.680 183.525 96.100 186.355 ;
      LAYER pwell ;
        RECT 61.875 182.325 63.245 183.135 ;
        RECT 63.255 182.325 68.765 183.135 ;
        RECT 68.775 182.325 74.285 183.135 ;
        RECT 74.765 182.410 75.195 183.195 ;
        RECT 75.215 182.325 80.725 183.135 ;
        RECT 80.735 182.325 86.245 183.135 ;
        RECT 86.255 182.325 91.765 183.135 ;
        RECT 91.775 182.325 94.525 183.135 ;
        RECT 94.535 182.325 95.905 183.135 ;
        RECT 62.015 182.115 62.185 182.325 ;
        RECT 63.395 182.115 63.565 182.325 ;
        RECT 68.915 182.115 69.085 182.325 ;
        RECT 74.435 182.275 74.605 182.305 ;
        RECT 74.430 182.165 74.605 182.275 ;
        RECT 74.435 182.115 74.605 182.165 ;
        RECT 75.355 182.135 75.525 182.325 ;
        RECT 79.955 182.115 80.125 182.305 ;
        RECT 80.875 182.135 81.045 182.325 ;
        RECT 85.475 182.115 85.645 182.305 ;
        RECT 86.395 182.135 86.565 182.325 ;
        RECT 87.310 182.165 87.430 182.275 ;
        RECT 88.235 182.115 88.405 182.305 ;
        RECT 91.915 182.135 92.085 182.325 ;
        RECT 93.765 182.160 93.925 182.270 ;
        RECT 95.595 182.115 95.765 182.325 ;
        RECT 61.875 181.305 63.245 182.115 ;
        RECT 63.255 181.305 68.765 182.115 ;
        RECT 68.775 181.305 74.285 182.115 ;
        RECT 74.295 181.305 79.805 182.115 ;
        RECT 79.815 181.305 85.325 182.115 ;
        RECT 85.335 181.305 87.165 182.115 ;
        RECT 87.645 181.245 88.075 182.030 ;
        RECT 88.095 181.305 93.605 182.115 ;
        RECT 94.535 181.305 95.905 182.115 ;
      LAYER nwell ;
        RECT 61.680 178.085 96.100 180.915 ;
      LAYER pwell ;
        RECT 61.875 176.885 63.245 177.695 ;
        RECT 63.255 176.885 68.765 177.695 ;
        RECT 68.775 176.885 74.285 177.695 ;
        RECT 74.765 176.970 75.195 177.755 ;
        RECT 75.215 176.885 80.725 177.695 ;
        RECT 80.735 176.885 86.245 177.695 ;
        RECT 86.255 176.885 91.765 177.695 ;
        RECT 91.775 176.885 94.525 177.695 ;
        RECT 94.535 176.885 95.905 177.695 ;
        RECT 62.015 176.675 62.185 176.885 ;
        RECT 63.395 176.675 63.565 176.885 ;
        RECT 68.915 176.675 69.085 176.885 ;
        RECT 74.435 176.835 74.605 176.865 ;
        RECT 74.430 176.725 74.605 176.835 ;
        RECT 74.435 176.675 74.605 176.725 ;
        RECT 75.355 176.695 75.525 176.885 ;
        RECT 79.955 176.675 80.125 176.865 ;
        RECT 80.875 176.695 81.045 176.885 ;
        RECT 85.475 176.675 85.645 176.865 ;
        RECT 86.395 176.695 86.565 176.885 ;
        RECT 87.310 176.725 87.430 176.835 ;
        RECT 88.235 176.675 88.405 176.865 ;
        RECT 91.915 176.695 92.085 176.885 ;
        RECT 93.765 176.720 93.925 176.830 ;
        RECT 95.595 176.675 95.765 176.885 ;
        RECT 61.875 175.865 63.245 176.675 ;
        RECT 63.255 175.865 68.765 176.675 ;
        RECT 68.775 175.865 74.285 176.675 ;
        RECT 74.295 175.865 79.805 176.675 ;
        RECT 79.815 175.865 85.325 176.675 ;
        RECT 85.335 175.865 87.165 176.675 ;
        RECT 87.645 175.805 88.075 176.590 ;
        RECT 88.095 175.865 93.605 176.675 ;
        RECT 94.535 175.865 95.905 176.675 ;
      LAYER nwell ;
        RECT 61.680 172.645 96.100 175.475 ;
      LAYER pwell ;
        RECT 61.875 171.445 63.245 172.255 ;
        RECT 63.255 171.445 68.765 172.255 ;
        RECT 68.775 171.445 74.285 172.255 ;
        RECT 74.765 171.530 75.195 172.315 ;
        RECT 75.215 171.445 80.725 172.255 ;
        RECT 80.735 171.445 86.245 172.255 ;
        RECT 86.255 171.445 87.625 172.255 ;
        RECT 87.645 171.530 88.075 172.315 ;
        RECT 88.095 171.445 93.605 172.255 ;
        RECT 94.535 171.445 95.905 172.255 ;
        RECT 62.015 171.255 62.185 171.445 ;
        RECT 63.395 171.255 63.565 171.445 ;
        RECT 68.915 171.255 69.085 171.445 ;
        RECT 74.430 171.285 74.550 171.395 ;
        RECT 75.355 171.255 75.525 171.445 ;
        RECT 80.875 171.255 81.045 171.445 ;
        RECT 86.395 171.255 86.565 171.445 ;
        RECT 88.235 171.255 88.405 171.445 ;
        RECT 93.765 171.290 93.925 171.400 ;
        RECT 95.595 171.255 95.765 171.445 ;
        RECT 110.740 63.630 126.560 65.640 ;
        RECT 136.490 63.630 152.310 65.640 ;
        RECT 110.750 53.990 122.850 57.950 ;
        RECT 99.620 50.650 106.130 53.000 ;
        RECT 130.170 49.150 134.130 61.250 ;
        RECT 110.830 44.150 122.930 48.110 ;
      LAYER nwell ;
        RECT 128.980 39.930 130.585 42.530 ;
      LAYER pwell ;
        RECT 130.875 41.275 131.785 42.100 ;
        RECT 130.875 41.170 131.975 41.275 ;
        RECT 131.805 41.105 131.975 41.170 ;
        RECT 130.915 40.135 131.700 40.565 ;
      LAYER nwell ;
        RECT 134.980 39.930 136.585 42.530 ;
      LAYER pwell ;
        RECT 136.875 41.275 137.785 42.100 ;
        RECT 136.875 41.170 137.975 41.275 ;
        RECT 137.805 41.105 137.975 41.170 ;
        RECT 136.915 40.135 137.700 40.565 ;
        RECT 110.830 35.190 122.930 39.150 ;
        RECT 129.620 37.060 131.660 39.100 ;
        RECT 143.300 35.600 154.130 47.700 ;
        RECT 149.060 35.120 150.630 35.600 ;
        RECT 151.370 35.130 152.940 35.600 ;
        RECT 99.620 31.470 106.130 33.820 ;
        RECT 110.830 26.230 122.930 30.190 ;
        RECT 130.170 22.050 134.130 34.150 ;
        RECT 132.100 20.940 132.880 22.050 ;
        RECT 142.740 21.230 143.450 22.900 ;
        RECT 142.740 20.880 144.210 21.230 ;
        RECT 144.980 20.880 146.630 21.220 ;
        RECT 147.420 20.880 148.730 21.210 ;
        RECT 149.520 20.880 151.230 21.200 ;
        RECT 111.940 17.670 137.760 18.360 ;
        RECT 141.530 17.670 152.360 20.880 ;
        RECT 111.940 17.050 152.360 17.670 ;
        RECT 111.940 16.350 137.760 17.050 ;
        RECT 141.530 13.780 152.360 17.050 ;
      LAYER li1 ;
        RECT 61.870 203.895 95.910 204.065 ;
        RECT 61.955 203.145 63.165 203.895 ;
        RECT 63.335 203.350 68.680 203.895 ;
        RECT 68.855 203.350 74.200 203.895 ;
        RECT 61.955 202.605 62.475 203.145 ;
        RECT 62.645 202.435 63.165 202.975 ;
        RECT 64.920 202.520 65.260 203.350 ;
        RECT 61.955 201.345 63.165 202.435 ;
        RECT 66.740 201.780 67.090 203.030 ;
        RECT 70.440 202.520 70.780 203.350 ;
        RECT 74.835 203.170 75.125 203.895 ;
        RECT 75.295 203.350 80.640 203.895 ;
        RECT 80.815 203.350 86.160 203.895 ;
        RECT 72.260 201.780 72.610 203.030 ;
        RECT 76.880 202.520 77.220 203.350 ;
        RECT 63.335 201.345 68.680 201.780 ;
        RECT 68.855 201.345 74.200 201.780 ;
        RECT 74.835 201.345 75.125 202.510 ;
        RECT 78.700 201.780 79.050 203.030 ;
        RECT 82.400 202.520 82.740 203.350 ;
        RECT 86.335 203.145 87.545 203.895 ;
        RECT 87.715 203.170 88.005 203.895 ;
        RECT 84.220 201.780 84.570 203.030 ;
        RECT 86.335 202.605 86.855 203.145 ;
        RECT 88.175 203.125 91.685 203.895 ;
        RECT 91.855 203.145 93.065 203.895 ;
        RECT 93.235 203.220 93.495 203.725 ;
        RECT 93.675 203.515 94.005 203.895 ;
        RECT 94.185 203.345 94.355 203.725 ;
        RECT 87.025 202.435 87.545 202.975 ;
        RECT 88.175 202.605 89.825 203.125 ;
        RECT 75.295 201.345 80.640 201.780 ;
        RECT 80.815 201.345 86.160 201.780 ;
        RECT 86.335 201.345 87.545 202.435 ;
        RECT 87.715 201.345 88.005 202.510 ;
        RECT 89.995 202.435 91.685 202.955 ;
        RECT 91.855 202.605 92.375 203.145 ;
        RECT 92.545 202.435 93.065 202.975 ;
        RECT 88.175 201.345 91.685 202.435 ;
        RECT 91.855 201.345 93.065 202.435 ;
        RECT 93.235 202.420 93.415 203.220 ;
        RECT 93.690 203.175 94.355 203.345 ;
        RECT 93.690 202.920 93.860 203.175 ;
        RECT 94.615 203.145 95.825 203.895 ;
        RECT 93.585 202.590 93.860 202.920 ;
        RECT 94.085 202.625 94.425 202.995 ;
        RECT 93.690 202.445 93.860 202.590 ;
        RECT 93.235 201.515 93.505 202.420 ;
        RECT 93.690 202.275 94.365 202.445 ;
        RECT 93.675 201.345 94.005 202.105 ;
        RECT 94.185 201.515 94.365 202.275 ;
        RECT 94.615 202.435 95.135 202.975 ;
        RECT 95.305 202.605 95.825 203.145 ;
        RECT 94.615 201.345 95.825 202.435 ;
        RECT 61.870 201.175 95.910 201.345 ;
        RECT 61.955 200.085 63.165 201.175 ;
        RECT 63.335 200.740 68.680 201.175 ;
        RECT 68.855 200.740 74.200 201.175 ;
        RECT 61.955 199.375 62.475 199.915 ;
        RECT 62.645 199.545 63.165 200.085 ;
        RECT 61.955 198.625 63.165 199.375 ;
        RECT 64.920 199.170 65.260 200.000 ;
        RECT 66.740 199.490 67.090 200.740 ;
        RECT 70.440 199.170 70.780 200.000 ;
        RECT 72.260 199.490 72.610 200.740 ;
        RECT 74.835 200.010 75.125 201.175 ;
        RECT 75.775 200.120 76.080 200.905 ;
        RECT 76.260 200.705 76.945 201.175 ;
        RECT 76.255 200.185 76.950 200.495 ;
        RECT 63.335 198.625 68.680 199.170 ;
        RECT 68.855 198.625 74.200 199.170 ;
        RECT 74.835 198.625 75.125 199.350 ;
        RECT 75.775 199.315 75.950 200.120 ;
        RECT 77.125 200.015 77.410 200.960 ;
        RECT 77.585 200.725 77.915 201.175 ;
        RECT 78.085 200.555 78.255 200.985 ;
        RECT 76.550 199.865 77.410 200.015 ;
        RECT 76.125 199.845 77.410 199.865 ;
        RECT 77.580 200.325 78.255 200.555 ;
        RECT 76.125 199.485 77.110 199.845 ;
        RECT 77.580 199.675 77.815 200.325 ;
        RECT 75.775 198.795 76.015 199.315 ;
        RECT 76.940 199.150 77.110 199.485 ;
        RECT 77.280 199.345 77.815 199.675 ;
        RECT 77.595 199.195 77.815 199.345 ;
        RECT 77.985 199.305 78.285 200.155 ;
        RECT 79.015 200.035 79.245 201.175 ;
        RECT 79.415 200.025 79.745 201.005 ;
        RECT 79.915 200.035 80.125 201.175 ;
        RECT 80.415 200.035 80.625 201.175 ;
        RECT 78.995 199.615 79.325 199.865 ;
        RECT 76.185 198.625 76.580 199.120 ;
        RECT 76.940 198.955 77.315 199.150 ;
        RECT 77.145 198.810 77.315 198.955 ;
        RECT 77.595 198.820 77.835 199.195 ;
        RECT 78.005 198.625 78.340 199.130 ;
        RECT 79.015 198.625 79.245 199.445 ;
        RECT 79.495 199.425 79.745 200.025 ;
        RECT 80.795 200.025 81.125 201.005 ;
        RECT 81.295 200.035 81.525 201.175 ;
        RECT 81.735 200.085 83.405 201.175 ;
        RECT 79.415 198.795 79.745 199.425 ;
        RECT 79.915 198.625 80.125 199.445 ;
        RECT 80.415 198.625 80.625 199.445 ;
        RECT 80.795 199.425 81.045 200.025 ;
        RECT 81.215 199.615 81.545 199.865 ;
        RECT 80.795 198.795 81.125 199.425 ;
        RECT 81.295 198.625 81.525 199.445 ;
        RECT 81.735 199.395 82.485 199.915 ;
        RECT 82.655 199.565 83.405 200.085 ;
        RECT 84.035 200.035 84.420 201.005 ;
        RECT 84.590 200.715 84.915 201.175 ;
        RECT 85.435 200.545 85.715 201.005 ;
        RECT 84.590 200.325 85.715 200.545 ;
        RECT 81.735 198.625 83.405 199.395 ;
        RECT 84.035 199.365 84.315 200.035 ;
        RECT 84.590 199.865 85.040 200.325 ;
        RECT 85.905 200.155 86.305 201.005 ;
        RECT 86.705 200.715 86.975 201.175 ;
        RECT 87.145 200.545 87.430 201.005 ;
        RECT 87.715 200.740 93.060 201.175 ;
        RECT 84.485 199.535 85.040 199.865 ;
        RECT 85.210 199.595 86.305 200.155 ;
        RECT 84.590 199.425 85.040 199.535 ;
        RECT 84.035 198.795 84.420 199.365 ;
        RECT 84.590 199.255 85.715 199.425 ;
        RECT 84.590 198.625 84.915 199.085 ;
        RECT 85.435 198.795 85.715 199.255 ;
        RECT 85.905 198.795 86.305 199.595 ;
        RECT 86.475 200.325 87.430 200.545 ;
        RECT 86.475 199.425 86.685 200.325 ;
        RECT 86.855 199.595 87.545 200.155 ;
        RECT 86.475 199.255 87.430 199.425 ;
        RECT 86.705 198.625 86.975 199.085 ;
        RECT 87.145 198.795 87.430 199.255 ;
        RECT 89.300 199.170 89.640 200.000 ;
        RECT 91.120 199.490 91.470 200.740 ;
        RECT 93.235 200.085 94.445 201.175 ;
        RECT 93.235 199.375 93.755 199.915 ;
        RECT 93.925 199.545 94.445 200.085 ;
        RECT 94.615 200.085 95.825 201.175 ;
        RECT 94.615 199.545 95.135 200.085 ;
        RECT 95.305 199.375 95.825 199.915 ;
        RECT 87.715 198.625 93.060 199.170 ;
        RECT 93.235 198.625 94.445 199.375 ;
        RECT 94.615 198.625 95.825 199.375 ;
        RECT 61.870 198.455 95.910 198.625 ;
        RECT 61.955 197.705 63.165 198.455 ;
        RECT 63.335 197.910 68.680 198.455 ;
        RECT 61.955 197.165 62.475 197.705 ;
        RECT 62.645 196.995 63.165 197.535 ;
        RECT 64.920 197.080 65.260 197.910 ;
        RECT 68.855 197.685 70.525 198.455 ;
        RECT 71.215 197.975 71.495 198.455 ;
        RECT 71.665 197.805 71.925 198.195 ;
        RECT 72.100 197.975 72.355 198.455 ;
        RECT 72.525 197.805 72.820 198.195 ;
        RECT 73.000 197.975 73.275 198.455 ;
        RECT 73.445 197.955 73.745 198.285 ;
        RECT 74.130 197.985 74.415 198.455 ;
        RECT 61.955 195.905 63.165 196.995 ;
        RECT 66.740 196.340 67.090 197.590 ;
        RECT 68.855 197.165 69.605 197.685 ;
        RECT 71.170 197.635 72.820 197.805 ;
        RECT 69.775 196.995 70.525 197.515 ;
        RECT 63.335 195.905 68.680 196.340 ;
        RECT 68.855 195.905 70.525 196.995 ;
        RECT 71.170 197.125 71.575 197.635 ;
        RECT 71.745 197.295 72.885 197.465 ;
        RECT 71.170 196.955 71.925 197.125 ;
        RECT 71.210 195.905 71.495 196.775 ;
        RECT 71.665 196.705 71.925 196.955 ;
        RECT 72.715 197.045 72.885 197.295 ;
        RECT 73.055 197.215 73.405 197.785 ;
        RECT 73.575 197.045 73.745 197.955 ;
        RECT 74.585 197.815 74.915 198.285 ;
        RECT 75.085 197.985 75.255 198.455 ;
        RECT 75.425 197.815 75.755 198.285 ;
        RECT 75.925 197.985 76.095 198.455 ;
        RECT 76.265 197.815 76.595 198.285 ;
        RECT 76.765 197.985 76.935 198.455 ;
        RECT 77.105 197.815 77.435 198.285 ;
        RECT 72.715 196.875 73.745 197.045 ;
        RECT 71.665 196.535 72.785 196.705 ;
        RECT 71.665 196.075 71.925 196.535 ;
        RECT 72.100 195.905 72.355 196.365 ;
        RECT 72.525 196.075 72.785 196.535 ;
        RECT 72.955 195.905 73.265 196.705 ;
        RECT 73.435 196.075 73.745 196.875 ;
        RECT 73.915 197.635 77.435 197.815 ;
        RECT 77.605 197.635 77.880 198.455 ;
        RECT 78.060 197.905 78.315 198.195 ;
        RECT 78.485 198.075 78.815 198.455 ;
        RECT 78.060 197.735 78.810 197.905 ;
        RECT 73.915 197.095 74.315 197.635 ;
        RECT 74.485 197.265 75.850 197.465 ;
        RECT 76.170 197.265 77.830 197.465 ;
        RECT 73.915 196.795 75.675 197.095 ;
        RECT 74.080 196.245 74.495 196.625 ;
        RECT 74.665 196.415 74.835 196.795 ;
        RECT 75.005 196.245 75.335 196.605 ;
        RECT 75.505 196.415 75.675 196.795 ;
        RECT 75.845 196.875 77.880 197.085 ;
        RECT 78.060 196.915 78.410 197.565 ;
        RECT 75.845 196.245 76.175 196.875 ;
        RECT 74.080 196.075 76.175 196.245 ;
        RECT 76.345 195.905 76.595 196.705 ;
        RECT 76.765 196.075 76.935 196.875 ;
        RECT 77.105 195.905 77.435 196.705 ;
        RECT 77.605 196.075 77.880 196.875 ;
        RECT 78.580 196.745 78.810 197.735 ;
        RECT 78.060 196.575 78.810 196.745 ;
        RECT 78.060 196.075 78.315 196.575 ;
        RECT 78.485 195.905 78.815 196.405 ;
        RECT 78.985 196.075 79.155 198.195 ;
        RECT 79.515 198.095 79.845 198.455 ;
        RECT 80.015 198.065 80.510 198.235 ;
        RECT 80.715 198.065 81.570 198.235 ;
        RECT 79.385 196.875 79.845 197.925 ;
        RECT 79.325 196.090 79.650 196.875 ;
        RECT 80.015 196.705 80.185 198.065 ;
        RECT 80.355 197.155 80.705 197.775 ;
        RECT 80.875 197.555 81.230 197.775 ;
        RECT 80.875 196.965 81.045 197.555 ;
        RECT 81.400 197.355 81.570 198.065 ;
        RECT 82.445 197.995 82.775 198.455 ;
        RECT 82.985 198.095 83.335 198.265 ;
        RECT 81.775 197.525 82.565 197.775 ;
        RECT 82.985 197.705 83.245 198.095 ;
        RECT 83.555 198.005 84.505 198.285 ;
        RECT 84.675 198.015 84.865 198.455 ;
        RECT 85.035 198.075 86.105 198.245 ;
        RECT 82.735 197.355 82.905 197.535 ;
        RECT 80.015 196.535 80.410 196.705 ;
        RECT 80.580 196.575 81.045 196.965 ;
        RECT 81.215 197.185 82.905 197.355 ;
        RECT 80.240 196.405 80.410 196.535 ;
        RECT 81.215 196.405 81.385 197.185 ;
        RECT 83.075 197.015 83.245 197.705 ;
        RECT 81.745 196.845 83.245 197.015 ;
        RECT 83.435 197.045 83.645 197.835 ;
        RECT 83.815 197.215 84.165 197.835 ;
        RECT 84.335 197.225 84.505 198.005 ;
        RECT 85.035 197.845 85.205 198.075 ;
        RECT 84.675 197.675 85.205 197.845 ;
        RECT 84.675 197.395 84.895 197.675 ;
        RECT 85.375 197.505 85.615 197.905 ;
        RECT 84.335 197.055 84.740 197.225 ;
        RECT 85.075 197.135 85.615 197.505 ;
        RECT 85.785 197.720 86.105 198.075 ;
        RECT 86.350 197.995 86.655 198.455 ;
        RECT 86.825 197.745 87.075 198.275 ;
        RECT 85.785 197.545 86.110 197.720 ;
        RECT 85.785 197.245 86.700 197.545 ;
        RECT 85.960 197.215 86.700 197.245 ;
        RECT 83.435 196.885 84.110 197.045 ;
        RECT 84.570 196.965 84.740 197.055 ;
        RECT 83.435 196.875 84.400 196.885 ;
        RECT 83.075 196.705 83.245 196.845 ;
        RECT 79.820 195.905 80.070 196.365 ;
        RECT 80.240 196.075 80.490 196.405 ;
        RECT 80.705 196.075 81.385 196.405 ;
        RECT 81.555 196.505 82.630 196.675 ;
        RECT 83.075 196.535 83.635 196.705 ;
        RECT 83.940 196.585 84.400 196.875 ;
        RECT 84.570 196.795 85.790 196.965 ;
        RECT 81.555 196.165 81.725 196.505 ;
        RECT 81.960 195.905 82.290 196.335 ;
        RECT 82.460 196.165 82.630 196.505 ;
        RECT 82.925 195.905 83.295 196.365 ;
        RECT 83.465 196.075 83.635 196.535 ;
        RECT 84.570 196.415 84.740 196.795 ;
        RECT 85.960 196.625 86.130 197.215 ;
        RECT 86.870 197.095 87.075 197.745 ;
        RECT 87.245 197.700 87.495 198.455 ;
        RECT 87.715 197.730 88.005 198.455 ;
        RECT 88.175 197.910 93.520 198.455 ;
        RECT 83.870 196.075 84.740 196.415 ;
        RECT 85.330 196.455 86.130 196.625 ;
        RECT 84.910 195.905 85.160 196.365 ;
        RECT 85.330 196.165 85.500 196.455 ;
        RECT 85.680 195.905 86.010 196.285 ;
        RECT 86.350 195.905 86.655 197.045 ;
        RECT 86.825 196.215 87.075 197.095 ;
        RECT 89.760 197.080 90.100 197.910 ;
        RECT 94.615 197.705 95.825 198.455 ;
        RECT 87.245 195.905 87.495 197.045 ;
        RECT 87.715 195.905 88.005 197.070 ;
        RECT 91.580 196.340 91.930 197.590 ;
        RECT 94.615 196.995 95.135 197.535 ;
        RECT 95.305 197.165 95.825 197.705 ;
        RECT 88.175 195.905 93.520 196.340 ;
        RECT 94.615 195.905 95.825 196.995 ;
        RECT 61.870 195.735 95.910 195.905 ;
        RECT 61.955 194.645 63.165 195.735 ;
        RECT 63.335 195.300 68.680 195.735 ;
        RECT 68.855 195.300 74.200 195.735 ;
        RECT 61.955 193.935 62.475 194.475 ;
        RECT 62.645 194.105 63.165 194.645 ;
        RECT 61.955 193.185 63.165 193.935 ;
        RECT 64.920 193.730 65.260 194.560 ;
        RECT 66.740 194.050 67.090 195.300 ;
        RECT 70.440 193.730 70.780 194.560 ;
        RECT 72.260 194.050 72.610 195.300 ;
        RECT 74.835 194.570 75.125 195.735 ;
        RECT 75.295 194.645 76.965 195.735 ;
        RECT 75.295 193.955 76.045 194.475 ;
        RECT 76.215 194.125 76.965 194.645 ;
        RECT 77.185 194.595 77.435 195.735 ;
        RECT 77.605 194.545 77.855 195.425 ;
        RECT 78.025 194.595 78.330 195.735 ;
        RECT 78.670 195.355 79.000 195.735 ;
        RECT 79.180 195.185 79.350 195.475 ;
        RECT 79.520 195.275 79.770 195.735 ;
        RECT 78.550 195.015 79.350 195.185 ;
        RECT 79.940 195.225 80.810 195.565 ;
        RECT 63.335 193.185 68.680 193.730 ;
        RECT 68.855 193.185 74.200 193.730 ;
        RECT 74.835 193.185 75.125 193.910 ;
        RECT 75.295 193.185 76.965 193.955 ;
        RECT 77.185 193.185 77.435 193.940 ;
        RECT 77.605 193.895 77.810 194.545 ;
        RECT 78.550 194.425 78.720 195.015 ;
        RECT 79.940 194.845 80.110 195.225 ;
        RECT 81.045 195.105 81.215 195.565 ;
        RECT 81.385 195.275 81.755 195.735 ;
        RECT 82.050 195.135 82.220 195.475 ;
        RECT 82.390 195.305 82.720 195.735 ;
        RECT 82.955 195.135 83.125 195.475 ;
        RECT 78.890 194.675 80.110 194.845 ;
        RECT 80.280 194.765 80.740 195.055 ;
        RECT 81.045 194.935 81.605 195.105 ;
        RECT 82.050 194.965 83.125 195.135 ;
        RECT 83.295 195.235 83.975 195.565 ;
        RECT 84.190 195.235 84.440 195.565 ;
        RECT 84.610 195.275 84.860 195.735 ;
        RECT 81.435 194.795 81.605 194.935 ;
        RECT 80.280 194.755 81.245 194.765 ;
        RECT 79.940 194.585 80.110 194.675 ;
        RECT 80.570 194.595 81.245 194.755 ;
        RECT 77.980 194.395 78.720 194.425 ;
        RECT 77.980 194.095 78.895 194.395 ;
        RECT 78.570 193.920 78.895 194.095 ;
        RECT 77.605 193.365 77.855 193.895 ;
        RECT 78.025 193.185 78.330 193.645 ;
        RECT 78.575 193.565 78.895 193.920 ;
        RECT 79.065 194.135 79.605 194.505 ;
        RECT 79.940 194.415 80.345 194.585 ;
        RECT 79.065 193.735 79.305 194.135 ;
        RECT 79.785 193.965 80.005 194.245 ;
        RECT 79.475 193.795 80.005 193.965 ;
        RECT 79.475 193.565 79.645 193.795 ;
        RECT 80.175 193.635 80.345 194.415 ;
        RECT 80.515 193.805 80.865 194.425 ;
        RECT 81.035 193.805 81.245 194.595 ;
        RECT 81.435 194.625 82.935 194.795 ;
        RECT 81.435 193.935 81.605 194.625 ;
        RECT 83.295 194.455 83.465 195.235 ;
        RECT 84.270 195.105 84.440 195.235 ;
        RECT 81.775 194.285 83.465 194.455 ;
        RECT 83.635 194.675 84.100 195.065 ;
        RECT 84.270 194.935 84.665 195.105 ;
        RECT 81.775 194.105 81.945 194.285 ;
        RECT 78.575 193.395 79.645 193.565 ;
        RECT 79.815 193.185 80.005 193.625 ;
        RECT 80.175 193.355 81.125 193.635 ;
        RECT 81.435 193.545 81.695 193.935 ;
        RECT 82.115 193.865 82.905 194.115 ;
        RECT 81.345 193.375 81.695 193.545 ;
        RECT 81.905 193.185 82.235 193.645 ;
        RECT 83.110 193.575 83.280 194.285 ;
        RECT 83.635 194.085 83.805 194.675 ;
        RECT 83.450 193.865 83.805 194.085 ;
        RECT 83.975 193.865 84.325 194.485 ;
        RECT 84.495 193.575 84.665 194.935 ;
        RECT 85.030 194.765 85.355 195.550 ;
        RECT 84.835 193.715 85.295 194.765 ;
        RECT 83.110 193.405 83.965 193.575 ;
        RECT 84.170 193.405 84.665 193.575 ;
        RECT 84.835 193.185 85.165 193.545 ;
        RECT 85.525 193.445 85.695 195.565 ;
        RECT 85.865 195.235 86.195 195.735 ;
        RECT 86.365 195.065 86.620 195.565 ;
        RECT 86.795 195.300 92.140 195.735 ;
        RECT 85.870 194.895 86.620 195.065 ;
        RECT 85.870 193.905 86.100 194.895 ;
        RECT 86.270 194.075 86.620 194.725 ;
        RECT 85.870 193.735 86.620 193.905 ;
        RECT 85.865 193.185 86.195 193.565 ;
        RECT 86.365 193.445 86.620 193.735 ;
        RECT 88.380 193.730 88.720 194.560 ;
        RECT 90.200 194.050 90.550 195.300 ;
        RECT 92.315 194.645 93.985 195.735 ;
        RECT 92.315 193.955 93.065 194.475 ;
        RECT 93.235 194.125 93.985 194.645 ;
        RECT 94.615 194.645 95.825 195.735 ;
        RECT 94.615 194.105 95.135 194.645 ;
        RECT 86.795 193.185 92.140 193.730 ;
        RECT 92.315 193.185 93.985 193.955 ;
        RECT 95.305 193.935 95.825 194.475 ;
        RECT 94.615 193.185 95.825 193.935 ;
        RECT 61.870 193.015 95.910 193.185 ;
        RECT 61.955 192.265 63.165 193.015 ;
        RECT 63.335 192.470 68.680 193.015 ;
        RECT 68.855 192.470 74.200 193.015 ;
        RECT 74.375 192.470 79.720 193.015 ;
        RECT 79.895 192.470 85.240 193.015 ;
        RECT 61.955 191.725 62.475 192.265 ;
        RECT 62.645 191.555 63.165 192.095 ;
        RECT 64.920 191.640 65.260 192.470 ;
        RECT 61.955 190.465 63.165 191.555 ;
        RECT 66.740 190.900 67.090 192.150 ;
        RECT 70.440 191.640 70.780 192.470 ;
        RECT 72.260 190.900 72.610 192.150 ;
        RECT 75.960 191.640 76.300 192.470 ;
        RECT 77.780 190.900 78.130 192.150 ;
        RECT 81.480 191.640 81.820 192.470 ;
        RECT 85.415 192.245 87.085 193.015 ;
        RECT 87.715 192.290 88.005 193.015 ;
        RECT 88.175 192.470 93.520 193.015 ;
        RECT 83.300 190.900 83.650 192.150 ;
        RECT 85.415 191.725 86.165 192.245 ;
        RECT 86.335 191.555 87.085 192.075 ;
        RECT 89.760 191.640 90.100 192.470 ;
        RECT 94.615 192.265 95.825 193.015 ;
        RECT 63.335 190.465 68.680 190.900 ;
        RECT 68.855 190.465 74.200 190.900 ;
        RECT 74.375 190.465 79.720 190.900 ;
        RECT 79.895 190.465 85.240 190.900 ;
        RECT 85.415 190.465 87.085 191.555 ;
        RECT 87.715 190.465 88.005 191.630 ;
        RECT 91.580 190.900 91.930 192.150 ;
        RECT 94.615 191.555 95.135 192.095 ;
        RECT 95.305 191.725 95.825 192.265 ;
        RECT 88.175 190.465 93.520 190.900 ;
        RECT 94.615 190.465 95.825 191.555 ;
        RECT 61.870 190.295 95.910 190.465 ;
        RECT 61.955 189.205 63.165 190.295 ;
        RECT 63.335 189.860 68.680 190.295 ;
        RECT 68.855 189.860 74.200 190.295 ;
        RECT 61.955 188.495 62.475 189.035 ;
        RECT 62.645 188.665 63.165 189.205 ;
        RECT 61.955 187.745 63.165 188.495 ;
        RECT 64.920 188.290 65.260 189.120 ;
        RECT 66.740 188.610 67.090 189.860 ;
        RECT 70.440 188.290 70.780 189.120 ;
        RECT 72.260 188.610 72.610 189.860 ;
        RECT 74.835 189.130 75.125 190.295 ;
        RECT 75.295 189.860 80.640 190.295 ;
        RECT 80.815 189.860 86.160 190.295 ;
        RECT 86.335 189.860 91.680 190.295 ;
        RECT 63.335 187.745 68.680 188.290 ;
        RECT 68.855 187.745 74.200 188.290 ;
        RECT 74.835 187.745 75.125 188.470 ;
        RECT 76.880 188.290 77.220 189.120 ;
        RECT 78.700 188.610 79.050 189.860 ;
        RECT 82.400 188.290 82.740 189.120 ;
        RECT 84.220 188.610 84.570 189.860 ;
        RECT 87.920 188.290 88.260 189.120 ;
        RECT 89.740 188.610 90.090 189.860 ;
        RECT 91.855 189.205 94.445 190.295 ;
        RECT 91.855 188.515 93.065 189.035 ;
        RECT 93.235 188.685 94.445 189.205 ;
        RECT 94.615 189.205 95.825 190.295 ;
        RECT 94.615 188.665 95.135 189.205 ;
        RECT 75.295 187.745 80.640 188.290 ;
        RECT 80.815 187.745 86.160 188.290 ;
        RECT 86.335 187.745 91.680 188.290 ;
        RECT 91.855 187.745 94.445 188.515 ;
        RECT 95.305 188.495 95.825 189.035 ;
        RECT 94.615 187.745 95.825 188.495 ;
        RECT 61.870 187.575 95.910 187.745 ;
        RECT 61.955 186.825 63.165 187.575 ;
        RECT 63.335 187.030 68.680 187.575 ;
        RECT 68.855 187.030 74.200 187.575 ;
        RECT 74.375 187.030 79.720 187.575 ;
        RECT 79.895 187.030 85.240 187.575 ;
        RECT 61.955 186.285 62.475 186.825 ;
        RECT 62.645 186.115 63.165 186.655 ;
        RECT 64.920 186.200 65.260 187.030 ;
        RECT 61.955 185.025 63.165 186.115 ;
        RECT 66.740 185.460 67.090 186.710 ;
        RECT 70.440 186.200 70.780 187.030 ;
        RECT 72.260 185.460 72.610 186.710 ;
        RECT 75.960 186.200 76.300 187.030 ;
        RECT 77.780 185.460 78.130 186.710 ;
        RECT 81.480 186.200 81.820 187.030 ;
        RECT 85.415 186.805 87.085 187.575 ;
        RECT 87.715 186.850 88.005 187.575 ;
        RECT 88.175 187.030 93.520 187.575 ;
        RECT 83.300 185.460 83.650 186.710 ;
        RECT 85.415 186.285 86.165 186.805 ;
        RECT 86.335 186.115 87.085 186.635 ;
        RECT 89.760 186.200 90.100 187.030 ;
        RECT 94.615 186.825 95.825 187.575 ;
        RECT 63.335 185.025 68.680 185.460 ;
        RECT 68.855 185.025 74.200 185.460 ;
        RECT 74.375 185.025 79.720 185.460 ;
        RECT 79.895 185.025 85.240 185.460 ;
        RECT 85.415 185.025 87.085 186.115 ;
        RECT 87.715 185.025 88.005 186.190 ;
        RECT 91.580 185.460 91.930 186.710 ;
        RECT 94.615 186.115 95.135 186.655 ;
        RECT 95.305 186.285 95.825 186.825 ;
        RECT 88.175 185.025 93.520 185.460 ;
        RECT 94.615 185.025 95.825 186.115 ;
        RECT 61.870 184.855 95.910 185.025 ;
        RECT 61.955 183.765 63.165 184.855 ;
        RECT 63.335 184.420 68.680 184.855 ;
        RECT 68.855 184.420 74.200 184.855 ;
        RECT 61.955 183.055 62.475 183.595 ;
        RECT 62.645 183.225 63.165 183.765 ;
        RECT 61.955 182.305 63.165 183.055 ;
        RECT 64.920 182.850 65.260 183.680 ;
        RECT 66.740 183.170 67.090 184.420 ;
        RECT 70.440 182.850 70.780 183.680 ;
        RECT 72.260 183.170 72.610 184.420 ;
        RECT 74.835 183.690 75.125 184.855 ;
        RECT 75.295 184.420 80.640 184.855 ;
        RECT 80.815 184.420 86.160 184.855 ;
        RECT 86.335 184.420 91.680 184.855 ;
        RECT 63.335 182.305 68.680 182.850 ;
        RECT 68.855 182.305 74.200 182.850 ;
        RECT 74.835 182.305 75.125 183.030 ;
        RECT 76.880 182.850 77.220 183.680 ;
        RECT 78.700 183.170 79.050 184.420 ;
        RECT 82.400 182.850 82.740 183.680 ;
        RECT 84.220 183.170 84.570 184.420 ;
        RECT 87.920 182.850 88.260 183.680 ;
        RECT 89.740 183.170 90.090 184.420 ;
        RECT 91.855 183.765 94.445 184.855 ;
        RECT 91.855 183.075 93.065 183.595 ;
        RECT 93.235 183.245 94.445 183.765 ;
        RECT 94.615 183.765 95.825 184.855 ;
        RECT 94.615 183.225 95.135 183.765 ;
        RECT 75.295 182.305 80.640 182.850 ;
        RECT 80.815 182.305 86.160 182.850 ;
        RECT 86.335 182.305 91.680 182.850 ;
        RECT 91.855 182.305 94.445 183.075 ;
        RECT 95.305 183.055 95.825 183.595 ;
        RECT 94.615 182.305 95.825 183.055 ;
        RECT 61.870 182.135 95.910 182.305 ;
        RECT 61.955 181.385 63.165 182.135 ;
        RECT 63.335 181.590 68.680 182.135 ;
        RECT 68.855 181.590 74.200 182.135 ;
        RECT 74.375 181.590 79.720 182.135 ;
        RECT 79.895 181.590 85.240 182.135 ;
        RECT 61.955 180.845 62.475 181.385 ;
        RECT 62.645 180.675 63.165 181.215 ;
        RECT 64.920 180.760 65.260 181.590 ;
        RECT 61.955 179.585 63.165 180.675 ;
        RECT 66.740 180.020 67.090 181.270 ;
        RECT 70.440 180.760 70.780 181.590 ;
        RECT 72.260 180.020 72.610 181.270 ;
        RECT 75.960 180.760 76.300 181.590 ;
        RECT 77.780 180.020 78.130 181.270 ;
        RECT 81.480 180.760 81.820 181.590 ;
        RECT 85.415 181.365 87.085 182.135 ;
        RECT 87.715 181.410 88.005 182.135 ;
        RECT 88.175 181.590 93.520 182.135 ;
        RECT 83.300 180.020 83.650 181.270 ;
        RECT 85.415 180.845 86.165 181.365 ;
        RECT 86.335 180.675 87.085 181.195 ;
        RECT 89.760 180.760 90.100 181.590 ;
        RECT 94.615 181.385 95.825 182.135 ;
        RECT 63.335 179.585 68.680 180.020 ;
        RECT 68.855 179.585 74.200 180.020 ;
        RECT 74.375 179.585 79.720 180.020 ;
        RECT 79.895 179.585 85.240 180.020 ;
        RECT 85.415 179.585 87.085 180.675 ;
        RECT 87.715 179.585 88.005 180.750 ;
        RECT 91.580 180.020 91.930 181.270 ;
        RECT 94.615 180.675 95.135 181.215 ;
        RECT 95.305 180.845 95.825 181.385 ;
        RECT 88.175 179.585 93.520 180.020 ;
        RECT 94.615 179.585 95.825 180.675 ;
        RECT 61.870 179.415 95.910 179.585 ;
        RECT 61.955 178.325 63.165 179.415 ;
        RECT 63.335 178.980 68.680 179.415 ;
        RECT 68.855 178.980 74.200 179.415 ;
        RECT 61.955 177.615 62.475 178.155 ;
        RECT 62.645 177.785 63.165 178.325 ;
        RECT 61.955 176.865 63.165 177.615 ;
        RECT 64.920 177.410 65.260 178.240 ;
        RECT 66.740 177.730 67.090 178.980 ;
        RECT 70.440 177.410 70.780 178.240 ;
        RECT 72.260 177.730 72.610 178.980 ;
        RECT 74.835 178.250 75.125 179.415 ;
        RECT 75.295 178.980 80.640 179.415 ;
        RECT 80.815 178.980 86.160 179.415 ;
        RECT 86.335 178.980 91.680 179.415 ;
        RECT 63.335 176.865 68.680 177.410 ;
        RECT 68.855 176.865 74.200 177.410 ;
        RECT 74.835 176.865 75.125 177.590 ;
        RECT 76.880 177.410 77.220 178.240 ;
        RECT 78.700 177.730 79.050 178.980 ;
        RECT 82.400 177.410 82.740 178.240 ;
        RECT 84.220 177.730 84.570 178.980 ;
        RECT 87.920 177.410 88.260 178.240 ;
        RECT 89.740 177.730 90.090 178.980 ;
        RECT 91.855 178.325 94.445 179.415 ;
        RECT 91.855 177.635 93.065 178.155 ;
        RECT 93.235 177.805 94.445 178.325 ;
        RECT 94.615 178.325 95.825 179.415 ;
        RECT 94.615 177.785 95.135 178.325 ;
        RECT 75.295 176.865 80.640 177.410 ;
        RECT 80.815 176.865 86.160 177.410 ;
        RECT 86.335 176.865 91.680 177.410 ;
        RECT 91.855 176.865 94.445 177.635 ;
        RECT 95.305 177.615 95.825 178.155 ;
        RECT 94.615 176.865 95.825 177.615 ;
        RECT 61.870 176.695 95.910 176.865 ;
        RECT 61.955 175.945 63.165 176.695 ;
        RECT 63.335 176.150 68.680 176.695 ;
        RECT 68.855 176.150 74.200 176.695 ;
        RECT 74.375 176.150 79.720 176.695 ;
        RECT 79.895 176.150 85.240 176.695 ;
        RECT 61.955 175.405 62.475 175.945 ;
        RECT 62.645 175.235 63.165 175.775 ;
        RECT 64.920 175.320 65.260 176.150 ;
        RECT 61.955 174.145 63.165 175.235 ;
        RECT 66.740 174.580 67.090 175.830 ;
        RECT 70.440 175.320 70.780 176.150 ;
        RECT 72.260 174.580 72.610 175.830 ;
        RECT 75.960 175.320 76.300 176.150 ;
        RECT 77.780 174.580 78.130 175.830 ;
        RECT 81.480 175.320 81.820 176.150 ;
        RECT 85.415 175.925 87.085 176.695 ;
        RECT 87.715 175.970 88.005 176.695 ;
        RECT 88.175 176.150 93.520 176.695 ;
        RECT 83.300 174.580 83.650 175.830 ;
        RECT 85.415 175.405 86.165 175.925 ;
        RECT 86.335 175.235 87.085 175.755 ;
        RECT 89.760 175.320 90.100 176.150 ;
        RECT 94.615 175.945 95.825 176.695 ;
        RECT 63.335 174.145 68.680 174.580 ;
        RECT 68.855 174.145 74.200 174.580 ;
        RECT 74.375 174.145 79.720 174.580 ;
        RECT 79.895 174.145 85.240 174.580 ;
        RECT 85.415 174.145 87.085 175.235 ;
        RECT 87.715 174.145 88.005 175.310 ;
        RECT 91.580 174.580 91.930 175.830 ;
        RECT 94.615 175.235 95.135 175.775 ;
        RECT 95.305 175.405 95.825 175.945 ;
        RECT 88.175 174.145 93.520 174.580 ;
        RECT 94.615 174.145 95.825 175.235 ;
        RECT 61.870 173.975 95.910 174.145 ;
        RECT 61.955 172.885 63.165 173.975 ;
        RECT 63.335 173.540 68.680 173.975 ;
        RECT 68.855 173.540 74.200 173.975 ;
        RECT 61.955 172.175 62.475 172.715 ;
        RECT 62.645 172.345 63.165 172.885 ;
        RECT 61.955 171.425 63.165 172.175 ;
        RECT 64.920 171.970 65.260 172.800 ;
        RECT 66.740 172.290 67.090 173.540 ;
        RECT 70.440 171.970 70.780 172.800 ;
        RECT 72.260 172.290 72.610 173.540 ;
        RECT 74.835 172.810 75.125 173.975 ;
        RECT 75.295 173.540 80.640 173.975 ;
        RECT 80.815 173.540 86.160 173.975 ;
        RECT 63.335 171.425 68.680 171.970 ;
        RECT 68.855 171.425 74.200 171.970 ;
        RECT 74.835 171.425 75.125 172.150 ;
        RECT 76.880 171.970 77.220 172.800 ;
        RECT 78.700 172.290 79.050 173.540 ;
        RECT 82.400 171.970 82.740 172.800 ;
        RECT 84.220 172.290 84.570 173.540 ;
        RECT 86.335 172.885 87.545 173.975 ;
        RECT 86.335 172.175 86.855 172.715 ;
        RECT 87.025 172.345 87.545 172.885 ;
        RECT 87.715 172.810 88.005 173.975 ;
        RECT 88.175 173.540 93.520 173.975 ;
        RECT 75.295 171.425 80.640 171.970 ;
        RECT 80.815 171.425 86.160 171.970 ;
        RECT 86.335 171.425 87.545 172.175 ;
        RECT 87.715 171.425 88.005 172.150 ;
        RECT 89.760 171.970 90.100 172.800 ;
        RECT 91.580 172.290 91.930 173.540 ;
        RECT 94.615 172.885 95.825 173.975 ;
        RECT 94.615 172.345 95.135 172.885 ;
        RECT 95.305 172.175 95.825 172.715 ;
        RECT 88.175 171.425 93.520 171.970 ;
        RECT 94.615 171.425 95.825 172.175 ;
        RECT 61.870 171.255 95.910 171.425 ;
        RECT 110.920 65.290 126.380 65.460 ;
        RECT 110.920 63.980 111.090 65.290 ;
        RECT 111.570 64.460 113.730 64.810 ;
        RECT 123.570 64.460 125.730 64.810 ;
        RECT 111.410 63.980 112.110 64.080 ;
        RECT 126.210 63.980 126.380 65.290 ;
        RECT 110.920 63.810 126.380 63.980 ;
        RECT 136.670 65.290 152.130 65.460 ;
        RECT 136.670 63.980 136.840 65.290 ;
        RECT 151.960 65.050 152.130 65.290 ;
        RECT 137.320 64.460 139.480 64.810 ;
        RECT 149.320 64.460 151.480 64.810 ;
        RECT 151.860 64.250 152.260 65.050 ;
        RECT 151.960 63.980 152.130 64.250 ;
        RECT 136.670 63.810 152.130 63.980 ;
        RECT 111.410 63.620 112.110 63.810 ;
        RECT 130.350 60.900 133.950 61.070 ;
        RECT 110.930 57.600 122.670 57.770 ;
        RECT 110.930 57.250 111.100 57.600 ;
        RECT 110.790 54.720 111.190 57.250 ;
        RECT 111.780 57.030 121.820 57.200 ;
        RECT 111.440 54.970 111.610 56.970 ;
        RECT 121.990 54.970 122.160 56.970 ;
        RECT 111.780 54.740 121.820 54.910 ;
        RECT 110.930 54.340 111.100 54.720 ;
        RECT 122.500 54.340 122.670 57.600 ;
        RECT 110.930 54.170 122.670 54.340 ;
        RECT 103.720 52.820 104.820 52.910 ;
        RECT 99.800 52.650 105.950 52.820 ;
        RECT 99.800 51.000 99.970 52.650 ;
        RECT 103.720 52.560 104.820 52.650 ;
        RECT 100.450 51.480 102.610 52.170 ;
        RECT 103.140 51.480 105.300 52.170 ;
        RECT 105.780 51.000 105.950 52.650 ;
        RECT 99.800 50.830 105.950 51.000 ;
        RECT 130.350 49.500 130.520 60.900 ;
        RECT 131.150 60.390 133.150 60.560 ;
        RECT 130.920 50.180 131.090 60.220 ;
        RECT 133.210 50.180 133.380 60.220 ;
        RECT 131.150 49.840 133.150 50.010 ;
        RECT 131.100 49.500 133.100 49.560 ;
        RECT 133.780 49.500 133.950 60.900 ;
        RECT 130.350 49.330 133.950 49.500 ;
        RECT 131.100 49.240 133.100 49.330 ;
        RECT 111.010 47.760 122.750 47.930 ;
        RECT 111.010 47.360 111.180 47.760 ;
        RECT 110.890 44.880 111.280 47.360 ;
        RECT 111.860 47.190 121.900 47.360 ;
        RECT 111.520 45.130 111.690 47.130 ;
        RECT 122.070 45.130 122.240 47.130 ;
        RECT 111.860 44.900 121.900 45.070 ;
        RECT 111.010 44.500 111.180 44.880 ;
        RECT 122.580 44.500 122.750 47.760 ;
        RECT 111.010 44.330 122.750 44.500 ;
        RECT 143.480 47.350 153.950 47.520 ;
        RECT 129.085 41.510 129.255 42.340 ;
        RECT 129.425 41.780 131.635 42.010 ;
        RECT 129.425 41.680 130.405 41.780 ;
        RECT 131.005 41.680 131.635 41.780 ;
        RECT 129.085 41.300 130.395 41.510 ;
        RECT 129.085 40.960 129.255 41.300 ;
        RECT 130.575 41.280 130.815 41.610 ;
        RECT 131.805 41.510 131.975 42.340 ;
        RECT 130.985 41.280 131.975 41.510 ;
        RECT 131.805 40.960 131.975 41.280 ;
        RECT 135.085 41.510 135.255 42.340 ;
        RECT 135.425 41.780 137.635 42.010 ;
        RECT 135.425 41.680 136.405 41.780 ;
        RECT 137.005 41.680 137.635 41.780 ;
        RECT 135.085 41.300 136.395 41.510 ;
        RECT 135.085 40.960 135.255 41.300 ;
        RECT 136.575 41.280 136.815 41.610 ;
        RECT 137.805 41.510 137.975 42.340 ;
        RECT 136.985 41.280 137.975 41.510 ;
        RECT 137.805 40.960 137.975 41.280 ;
        RECT 129.085 40.495 129.255 40.580 ;
        RECT 131.805 40.495 131.975 40.580 ;
        RECT 129.085 40.205 130.420 40.495 ;
        RECT 131.080 40.205 131.975 40.495 ;
        RECT 129.085 40.120 129.255 40.205 ;
        RECT 131.805 40.120 131.975 40.205 ;
        RECT 135.085 40.495 135.255 40.580 ;
        RECT 137.805 40.495 137.975 40.580 ;
        RECT 135.085 40.205 136.420 40.495 ;
        RECT 137.080 40.205 137.975 40.495 ;
        RECT 135.085 40.120 135.255 40.205 ;
        RECT 137.805 40.120 137.975 40.205 ;
        RECT 111.010 38.800 122.750 38.970 ;
        RECT 111.010 38.430 111.180 38.800 ;
        RECT 110.900 35.940 111.250 38.430 ;
        RECT 111.860 38.230 121.900 38.400 ;
        RECT 111.520 36.170 111.690 38.170 ;
        RECT 122.070 36.170 122.240 38.170 ;
        RECT 111.860 35.940 121.900 36.110 ;
        RECT 111.010 35.540 111.180 35.940 ;
        RECT 122.580 35.540 122.750 38.800 ;
        RECT 129.800 38.750 131.480 38.920 ;
        RECT 129.800 37.410 129.970 38.750 ;
        RECT 131.310 38.510 131.480 38.750 ;
        RECT 130.370 37.730 130.910 38.430 ;
        RECT 131.250 37.680 131.560 38.510 ;
        RECT 131.310 37.410 131.480 37.680 ;
        RECT 129.800 37.240 131.480 37.410 ;
        RECT 143.480 35.950 143.650 47.350 ;
        RECT 144.280 46.840 146.280 47.010 ;
        RECT 146.570 46.840 148.570 47.010 ;
        RECT 148.860 46.840 150.860 47.010 ;
        RECT 151.150 46.840 153.150 47.010 ;
        RECT 144.050 36.630 144.220 46.670 ;
        RECT 146.340 36.630 146.510 46.670 ;
        RECT 148.630 36.630 148.800 46.670 ;
        RECT 150.920 36.630 151.090 46.670 ;
        RECT 153.210 36.630 153.380 46.670 ;
        RECT 153.780 41.960 153.950 47.350 ;
        RECT 153.660 40.420 154.040 41.960 ;
        RECT 144.280 36.290 146.280 36.460 ;
        RECT 146.570 36.290 148.570 36.460 ;
        RECT 148.860 36.290 150.860 36.460 ;
        RECT 151.150 36.290 153.150 36.460 ;
        RECT 153.780 35.950 153.950 40.420 ;
        RECT 143.480 35.780 153.950 35.950 ;
        RECT 111.010 35.370 122.750 35.540 ;
        RECT 130.940 33.970 133.120 34.090 ;
        RECT 130.350 33.800 133.950 33.970 ;
        RECT 99.800 33.470 105.950 33.640 ;
        RECT 99.800 31.820 99.970 33.470 ;
        RECT 100.450 32.300 102.610 32.990 ;
        RECT 103.140 32.300 105.300 32.990 ;
        RECT 103.910 31.820 105.210 31.940 ;
        RECT 105.780 31.820 105.950 33.470 ;
        RECT 99.800 31.650 105.950 31.820 ;
        RECT 103.910 31.540 105.210 31.650 ;
        RECT 111.010 29.840 122.750 30.010 ;
        RECT 111.010 29.400 111.180 29.840 ;
        RECT 110.950 27.040 111.280 29.400 ;
        RECT 111.860 29.270 121.900 29.440 ;
        RECT 111.520 27.210 111.690 29.210 ;
        RECT 122.070 27.210 122.240 29.210 ;
        RECT 111.010 26.580 111.180 27.040 ;
        RECT 111.860 26.980 121.900 27.150 ;
        RECT 122.580 26.580 122.750 29.840 ;
        RECT 111.010 26.410 122.750 26.580 ;
        RECT 130.350 22.400 130.520 33.800 ;
        RECT 130.940 33.710 133.120 33.800 ;
        RECT 131.150 33.290 133.150 33.460 ;
        RECT 130.920 23.080 131.090 33.120 ;
        RECT 133.210 23.080 133.380 33.120 ;
        RECT 131.150 22.740 133.150 22.910 ;
        RECT 133.780 22.400 133.950 33.800 ;
        RECT 130.350 22.230 133.950 22.400 ;
        RECT 141.710 20.530 152.180 20.700 ;
        RECT 113.630 18.180 114.840 18.310 ;
        RECT 112.120 18.010 137.580 18.180 ;
        RECT 112.120 16.700 112.290 18.010 ;
        RECT 113.630 17.890 114.840 18.010 ;
        RECT 112.770 17.180 114.930 17.530 ;
        RECT 134.770 17.180 136.930 17.530 ;
        RECT 137.410 16.700 137.580 18.010 ;
        RECT 112.120 16.530 137.580 16.700 ;
        RECT 141.710 14.130 141.880 20.530 ;
        RECT 142.510 20.020 144.510 20.190 ;
        RECT 144.800 20.020 146.800 20.190 ;
        RECT 147.090 20.020 149.090 20.190 ;
        RECT 149.380 20.020 151.380 20.190 ;
        RECT 142.280 14.810 142.450 19.850 ;
        RECT 144.570 14.810 144.740 19.850 ;
        RECT 146.860 14.810 147.030 19.850 ;
        RECT 149.150 14.810 149.320 19.850 ;
        RECT 151.440 14.810 151.610 19.850 ;
        RECT 152.010 18.370 152.180 20.530 ;
        RECT 151.940 14.900 152.340 18.370 ;
        RECT 142.510 14.470 144.510 14.640 ;
        RECT 144.800 14.470 146.800 14.640 ;
        RECT 147.090 14.470 149.090 14.640 ;
        RECT 149.380 14.470 151.380 14.640 ;
        RECT 152.010 14.130 152.180 14.900 ;
        RECT 141.710 13.960 152.180 14.130 ;
      LAYER met1 ;
        RECT 61.870 203.740 96.710 204.220 ;
        RECT 93.220 203.340 93.540 203.600 ;
        RECT 93.310 202.860 93.450 203.340 ;
        RECT 94.155 202.860 94.445 202.905 ;
        RECT 93.310 202.720 94.445 202.860 ;
        RECT 94.155 202.675 94.445 202.720 ;
        RECT 85.860 201.840 86.180 201.900 ;
        RECT 93.235 201.840 93.525 201.885 ;
        RECT 85.860 201.700 93.525 201.840 ;
        RECT 85.860 201.640 86.180 201.700 ;
        RECT 93.235 201.655 93.525 201.700 ;
        RECT 61.870 201.020 95.910 201.500 ;
        RECT 76.200 200.280 76.520 200.540 ;
        RECT 78.975 199.615 79.265 199.845 ;
        RECT 81.275 199.800 81.565 199.845 ;
        RECT 84.035 199.800 84.325 199.845 ;
        RECT 81.275 199.660 84.325 199.800 ;
        RECT 81.275 199.615 81.565 199.660 ;
        RECT 84.035 199.615 84.325 199.660 ;
        RECT 85.400 199.800 85.720 199.860 ;
        RECT 86.795 199.800 87.085 199.845 ;
        RECT 85.400 199.660 87.085 199.800 ;
        RECT 77.580 199.460 77.900 199.520 ;
        RECT 78.055 199.460 78.345 199.505 ;
        RECT 79.050 199.460 79.190 199.615 ;
        RECT 85.400 199.600 85.720 199.660 ;
        RECT 86.795 199.615 87.085 199.660 ;
        RECT 77.580 199.320 79.190 199.460 ;
        RECT 77.580 199.260 77.900 199.320 ;
        RECT 78.055 199.275 78.345 199.320 ;
        RECT 75.740 198.920 76.060 199.180 ;
        RECT 79.435 199.120 79.725 199.165 ;
        RECT 79.880 199.120 80.200 199.180 ;
        RECT 79.435 198.980 80.200 199.120 ;
        RECT 79.435 198.935 79.725 198.980 ;
        RECT 79.880 198.920 80.200 198.980 ;
        RECT 80.800 198.920 81.120 199.180 ;
        RECT 61.870 198.300 96.710 198.780 ;
        RECT 75.740 198.100 76.060 198.160 ;
        RECT 73.070 197.960 76.060 198.100 ;
        RECT 67.000 197.760 67.320 197.820 ;
        RECT 73.070 197.805 73.210 197.960 ;
        RECT 75.740 197.900 76.060 197.960 ;
        RECT 76.200 197.900 76.520 198.160 ;
        RECT 84.020 198.100 84.340 198.160 ;
        RECT 78.130 197.960 84.340 198.100 ;
        RECT 71.155 197.760 71.445 197.805 ;
        RECT 67.000 197.620 71.445 197.760 ;
        RECT 67.000 197.560 67.320 197.620 ;
        RECT 71.155 197.575 71.445 197.620 ;
        RECT 72.995 197.575 73.285 197.805 ;
        RECT 73.900 197.560 74.220 197.820 ;
        RECT 75.295 197.420 75.585 197.465 ;
        RECT 76.290 197.420 76.430 197.900 ;
        RECT 75.295 197.280 76.430 197.420 ;
        RECT 75.295 197.235 75.585 197.280 ;
        RECT 76.290 197.080 76.430 197.280 ;
        RECT 77.580 197.220 77.900 197.480 ;
        RECT 78.130 197.465 78.270 197.960 ;
        RECT 84.020 197.900 84.340 197.960 ;
        RECT 79.435 197.760 79.725 197.805 ;
        RECT 80.800 197.760 81.120 197.820 ;
        RECT 79.435 197.620 81.120 197.760 ;
        RECT 79.435 197.575 79.725 197.620 ;
        RECT 80.800 197.560 81.120 197.620 ;
        RECT 81.715 197.760 82.365 197.805 ;
        RECT 85.315 197.760 85.605 197.805 ;
        RECT 85.860 197.760 86.180 197.820 ;
        RECT 81.715 197.620 86.180 197.760 ;
        RECT 81.715 197.575 82.365 197.620 ;
        RECT 85.015 197.575 85.605 197.620 ;
        RECT 78.055 197.235 78.345 197.465 ;
        RECT 78.520 197.420 78.810 197.465 ;
        RECT 80.355 197.420 80.645 197.465 ;
        RECT 83.935 197.420 84.225 197.465 ;
        RECT 78.520 197.280 84.225 197.420 ;
        RECT 78.520 197.235 78.810 197.280 ;
        RECT 80.355 197.235 80.645 197.280 ;
        RECT 83.935 197.235 84.225 197.280 ;
        RECT 85.015 197.260 85.305 197.575 ;
        RECT 85.860 197.560 86.180 197.620 ;
        RECT 85.400 197.080 85.720 197.140 ;
        RECT 86.320 197.080 86.640 197.140 ;
        RECT 86.795 197.080 87.085 197.125 ;
        RECT 76.290 196.940 87.085 197.080 ;
        RECT 85.400 196.880 85.720 196.940 ;
        RECT 86.320 196.880 86.640 196.940 ;
        RECT 86.795 196.895 87.085 196.940 ;
        RECT 78.925 196.740 79.215 196.785 ;
        RECT 80.815 196.740 81.105 196.785 ;
        RECT 83.935 196.740 84.225 196.785 ;
        RECT 78.925 196.600 84.225 196.740 ;
        RECT 78.925 196.555 79.215 196.600 ;
        RECT 80.815 196.555 81.105 196.600 ;
        RECT 83.935 196.555 84.225 196.600 ;
        RECT 61.870 195.580 95.910 196.060 ;
        RECT 77.580 195.180 77.900 195.440 ;
        RECT 79.880 195.180 80.200 195.440 ;
        RECT 79.970 194.700 80.110 195.180 ;
        RECT 80.455 195.040 80.745 195.085 ;
        RECT 83.575 195.040 83.865 195.085 ;
        RECT 85.465 195.040 85.755 195.085 ;
        RECT 80.455 194.900 85.755 195.040 ;
        RECT 80.455 194.855 80.745 194.900 ;
        RECT 83.575 194.855 83.865 194.900 ;
        RECT 85.465 194.855 85.755 194.900 ;
        RECT 84.955 194.700 85.245 194.745 ;
        RECT 79.970 194.560 85.245 194.700 ;
        RECT 84.955 194.515 85.245 194.560 ;
        RECT 86.320 194.500 86.640 194.760 ;
        RECT 79.375 194.065 79.665 194.380 ;
        RECT 80.455 194.360 80.745 194.405 ;
        RECT 84.035 194.360 84.325 194.405 ;
        RECT 85.870 194.360 86.160 194.405 ;
        RECT 80.455 194.220 86.160 194.360 ;
        RECT 80.455 194.175 80.745 194.220 ;
        RECT 84.035 194.175 84.325 194.220 ;
        RECT 85.870 194.175 86.160 194.220 ;
        RECT 79.075 194.020 79.665 194.065 ;
        RECT 82.315 194.020 82.965 194.065 ;
        RECT 79.075 193.880 86.090 194.020 ;
        RECT 79.075 193.835 79.365 193.880 ;
        RECT 82.315 193.835 82.965 193.880 ;
        RECT 85.950 193.740 86.090 193.880 ;
        RECT 85.860 193.480 86.180 193.740 ;
        RECT 61.870 192.860 96.710 193.340 ;
        RECT 61.870 190.140 95.910 190.620 ;
        RECT 61.870 187.420 96.710 187.900 ;
        RECT 61.870 184.700 95.910 185.180 ;
        RECT 61.870 181.980 96.710 182.460 ;
        RECT 61.870 179.260 95.910 179.740 ;
        RECT 61.870 176.540 96.710 177.020 ;
        RECT 61.870 173.820 95.910 174.300 ;
        RECT 61.870 171.100 96.710 171.580 ;
        RECT 109.270 64.900 110.040 65.510 ;
        RECT 109.270 64.330 113.800 64.900 ;
        RECT 123.660 64.760 139.600 65.050 ;
        RECT 149.680 64.980 151.000 65.030 ;
        RECT 123.595 64.510 139.600 64.760 ;
        RECT 109.270 63.740 110.040 64.330 ;
        RECT 123.660 64.300 139.600 64.510 ;
        RECT 149.290 64.310 151.630 64.980 ;
        RECT 111.370 63.130 112.200 64.140 ;
        RECT 111.510 62.710 111.960 63.130 ;
        RECT 112.190 60.585 113.120 60.610 ;
        RECT 131.320 60.590 132.890 64.300 ;
        RECT 149.680 64.260 151.000 64.310 ;
        RECT 151.770 64.170 152.480 65.160 ;
        RECT 108.705 59.655 113.120 60.585 ;
        RECT 131.170 60.360 133.130 60.590 ;
        RECT 130.890 60.070 131.120 60.200 ;
        RECT 104.190 53.520 104.600 53.800 ;
        RECT 103.660 52.500 104.910 53.520 ;
        RECT 98.140 52.330 99.120 52.370 ;
        RECT 98.130 51.360 102.660 52.330 ;
        RECT 108.705 52.310 109.635 59.655 ;
        RECT 112.190 58.260 113.120 59.655 ;
        RECT 110.570 56.530 111.250 57.310 ;
        RECT 111.990 57.230 121.630 58.260 ;
        RECT 111.800 57.000 121.800 57.230 ;
        RECT 109.900 55.190 111.250 56.530 ;
        RECT 110.570 54.640 111.250 55.190 ;
        RECT 111.410 54.990 111.640 56.950 ;
        RECT 111.990 56.890 121.630 57.000 ;
        RECT 121.960 56.740 122.190 56.950 ;
        RECT 121.960 55.130 124.860 56.740 ;
        RECT 111.980 54.940 121.600 55.030 ;
        RECT 121.960 54.990 122.190 55.130 ;
        RECT 111.800 54.710 121.800 54.940 ;
        RECT 111.980 53.660 121.600 54.710 ;
        RECT 123.100 53.915 124.850 55.130 ;
        RECT 107.850 52.300 109.710 52.310 ;
        RECT 98.140 51.290 99.120 51.360 ;
        RECT 103.120 51.280 109.710 52.300 ;
        RECT 107.850 51.270 109.710 51.280 ;
        RECT 108.670 45.740 109.710 51.270 ;
        RECT 120.710 51.740 121.520 53.660 ;
        RECT 123.070 52.165 124.880 53.915 ;
        RECT 129.970 51.740 131.150 60.070 ;
        RECT 120.710 50.330 131.150 51.740 ;
        RECT 120.710 50.280 130.660 50.330 ;
        RECT 120.710 48.430 121.520 50.280 ;
        RECT 130.890 50.200 131.120 50.330 ;
        RECT 131.290 50.040 132.950 60.360 ;
        RECT 133.180 60.040 133.410 60.200 ;
        RECT 133.090 51.555 134.240 60.040 ;
        RECT 133.090 50.565 140.620 51.555 ;
        RECT 133.090 50.350 134.240 50.565 ;
        RECT 133.180 50.200 133.410 50.350 ;
        RECT 131.170 49.810 133.130 50.040 ;
        RECT 131.290 49.780 132.950 49.810 ;
        RECT 131.040 48.480 133.190 49.600 ;
        RECT 139.630 49.190 140.620 50.565 ;
        RECT 147.510 49.190 147.990 49.220 ;
        RECT 139.630 48.710 147.990 49.190 ;
        RECT 110.570 46.650 111.350 47.420 ;
        RECT 112.040 47.390 121.710 48.430 ;
        RECT 131.610 47.770 132.610 48.480 ;
        RECT 111.880 47.160 121.880 47.390 ;
        RECT 102.650 44.740 109.710 45.740 ;
        RECT 109.850 45.580 111.350 46.650 ;
        RECT 110.570 44.820 111.350 45.580 ;
        RECT 111.490 45.150 111.720 47.110 ;
        RECT 112.040 47.030 121.710 47.160 ;
        RECT 122.040 46.960 122.270 47.110 ;
        RECT 123.930 46.960 124.690 46.990 ;
        RECT 122.010 45.920 124.690 46.960 ;
        RECT 122.010 45.890 135.380 45.920 ;
        RECT 111.980 45.100 121.770 45.330 ;
        RECT 122.010 45.270 136.060 45.890 ;
        RECT 122.040 45.150 122.270 45.270 ;
        RECT 111.880 44.870 121.880 45.100 ;
        RECT 123.930 45.080 136.060 45.270 ;
        RECT 108.670 43.880 109.710 44.740 ;
        RECT 108.640 42.840 109.740 43.880 ;
        RECT 111.980 43.690 121.770 44.870 ;
        RECT 112.130 42.320 113.110 43.690 ;
        RECT 107.020 41.340 113.110 42.320 ;
        RECT 107.020 40.370 108.000 41.340 ;
        RECT 103.910 39.370 108.000 40.370 ;
        RECT 108.640 39.610 113.100 40.650 ;
        RECT 112.060 39.430 113.100 39.610 ;
        RECT 103.910 37.110 104.910 39.370 ;
        RECT 98.280 33.230 99.140 33.250 ;
        RECT 98.240 32.940 102.340 33.230 ;
        RECT 107.020 33.120 108.000 39.370 ;
        RECT 110.620 37.750 111.350 38.490 ;
        RECT 112.040 38.430 121.810 39.430 ;
        RECT 111.880 38.200 121.880 38.430 ;
        RECT 109.710 36.690 111.350 37.750 ;
        RECT 110.620 35.850 111.350 36.690 ;
        RECT 111.490 36.190 111.720 38.150 ;
        RECT 112.040 38.010 121.810 38.200 ;
        RECT 122.040 38.000 122.270 38.150 ;
        RECT 123.930 38.000 124.690 45.080 ;
        RECT 129.750 43.250 130.030 43.270 ;
        RECT 112.080 36.140 121.760 36.350 ;
        RECT 122.010 36.300 124.690 38.000 ;
        RECT 128.060 43.210 130.030 43.250 ;
        RECT 128.060 42.930 133.270 43.210 ;
        RECT 128.060 42.760 130.030 42.930 ;
        RECT 128.060 37.825 128.640 42.760 ;
        RECT 128.930 41.320 129.410 42.340 ;
        RECT 129.750 41.700 130.030 42.760 ;
        RECT 128.930 40.960 129.450 41.320 ;
        RECT 128.950 40.580 129.450 40.960 ;
        RECT 128.930 40.120 129.450 40.580 ;
        RECT 128.950 39.160 129.450 40.120 ;
        RECT 129.010 39.110 129.450 39.160 ;
        RECT 130.520 38.660 130.860 41.680 ;
        RECT 131.650 39.870 132.130 42.340 ;
        RECT 131.640 39.320 132.130 39.870 ;
        RECT 132.990 39.380 133.270 42.930 ;
        RECT 134.940 42.340 135.410 43.910 ;
        RECT 134.930 40.960 135.410 42.340 ;
        RECT 135.720 41.710 136.050 45.080 ;
        RECT 137.650 41.880 138.130 42.340 ;
        RECT 134.940 40.580 135.410 40.960 ;
        RECT 134.930 40.120 135.410 40.580 ;
        RECT 134.940 40.110 135.410 40.120 ;
        RECT 136.580 39.380 136.860 41.600 ;
        RECT 137.650 40.960 138.140 41.880 ;
        RECT 137.660 40.580 138.140 40.960 ;
        RECT 137.650 40.120 138.140 40.580 ;
        RECT 131.640 39.270 132.120 39.320 ;
        RECT 132.990 39.100 136.860 39.380 ;
        RECT 137.660 39.240 138.140 40.120 ;
        RECT 139.630 41.875 140.620 48.710 ;
        RECT 147.510 48.680 147.990 48.710 ;
        RECT 144.500 47.040 146.070 47.060 ;
        RECT 146.780 47.040 148.350 47.060 ;
        RECT 149.060 47.040 150.630 47.060 ;
        RECT 151.370 47.040 152.940 47.070 ;
        RECT 144.300 46.810 146.260 47.040 ;
        RECT 146.590 46.810 148.550 47.040 ;
        RECT 148.880 46.810 150.840 47.040 ;
        RECT 151.170 46.810 153.130 47.040 ;
        RECT 144.020 46.540 144.250 46.650 ;
        RECT 142.950 41.875 144.320 46.540 ;
        RECT 139.630 40.885 144.320 41.875 ;
        RECT 137.660 39.180 138.130 39.240 ;
        RECT 130.420 38.410 131.000 38.660 ;
        RECT 131.180 38.590 131.650 38.640 ;
        RECT 122.040 36.190 122.270 36.300 ;
        RECT 123.930 36.290 124.690 36.300 ;
        RECT 111.880 35.910 121.880 36.140 ;
        RECT 112.080 34.700 121.760 35.910 ;
        RECT 98.240 32.350 102.585 32.940 ;
        RECT 98.240 32.120 102.340 32.350 ;
        RECT 103.140 32.170 108.010 33.120 ;
        RECT 120.780 32.980 121.760 34.700 ;
        RECT 127.035 33.715 128.785 37.825 ;
        RECT 130.340 37.750 131.000 38.410 ;
        RECT 130.420 37.480 131.000 37.750 ;
        RECT 131.170 37.630 131.650 38.590 ;
        RECT 131.180 37.590 131.650 37.630 ;
        RECT 130.420 37.230 131.040 37.480 ;
        RECT 130.210 36.230 131.210 37.230 ;
        RECT 131.560 35.170 132.480 35.660 ;
        RECT 130.860 33.640 133.180 35.170 ;
        RECT 131.170 33.260 133.130 33.490 ;
        RECT 130.890 32.980 131.120 33.100 ;
        RECT 103.830 30.520 105.270 32.030 ;
        RECT 104.180 30.110 105.030 30.520 ;
        RECT 107.020 24.740 108.000 32.170 ;
        RECT 120.780 32.020 131.180 32.980 ;
        RECT 120.780 30.690 121.760 32.020 ;
        RECT 112.060 30.330 121.760 30.690 ;
        RECT 112.060 29.470 121.730 30.330 ;
        RECT 110.630 28.690 111.330 29.470 ;
        RECT 111.880 29.240 121.880 29.470 ;
        RECT 109.720 27.720 111.330 28.690 ;
        RECT 110.630 26.980 111.330 27.720 ;
        RECT 111.490 27.230 111.720 29.190 ;
        RECT 112.060 29.090 121.730 29.240 ;
        RECT 122.040 29.080 122.270 29.190 ;
        RECT 123.100 29.080 124.850 31.155 ;
        RECT 112.030 27.180 121.740 27.340 ;
        RECT 121.970 27.330 124.850 29.080 ;
        RECT 122.040 27.230 122.270 27.330 ;
        RECT 111.880 26.950 121.880 27.180 ;
        RECT 112.030 25.810 121.740 26.950 ;
        RECT 112.080 24.740 113.060 25.810 ;
        RECT 107.020 23.760 113.060 24.740 ;
        RECT 129.890 23.170 131.180 32.020 ;
        RECT 130.890 23.100 131.120 23.170 ;
        RECT 131.320 22.940 133.020 33.260 ;
        RECT 133.180 32.980 133.410 33.100 ;
        RECT 133.160 32.940 134.270 32.980 ;
        RECT 139.630 32.940 140.620 40.885 ;
        RECT 142.950 36.830 144.320 40.885 ;
        RECT 144.500 46.370 146.070 46.810 ;
        RECT 144.500 36.910 145.870 46.370 ;
        RECT 146.310 46.220 146.540 46.650 ;
        RECT 146.780 46.420 148.350 46.810 ;
        RECT 146.780 46.370 148.060 46.420 ;
        RECT 146.120 42.000 146.740 46.220 ;
        RECT 146.100 40.380 146.740 42.000 ;
        RECT 146.120 37.250 146.740 40.380 ;
        RECT 144.020 36.650 144.250 36.830 ;
        RECT 144.500 36.490 146.070 36.910 ;
        RECT 146.310 36.650 146.540 37.250 ;
        RECT 147.060 36.910 148.060 46.370 ;
        RECT 148.600 46.210 148.830 46.650 ;
        RECT 149.060 46.420 150.630 46.810 ;
        RECT 149.290 46.410 150.630 46.420 ;
        RECT 148.430 44.750 149.010 46.210 ;
        RECT 148.430 42.900 149.020 44.750 ;
        RECT 148.430 37.200 149.010 42.900 ;
        RECT 146.780 36.830 148.060 36.910 ;
        RECT 146.780 36.490 148.350 36.830 ;
        RECT 148.600 36.650 148.830 37.200 ;
        RECT 149.290 36.910 150.310 46.410 ;
        RECT 150.890 46.120 151.120 46.650 ;
        RECT 151.370 46.410 152.940 46.810 ;
        RECT 151.720 46.400 152.940 46.410 ;
        RECT 150.690 42.020 151.350 46.120 ;
        RECT 150.650 40.360 151.350 42.020 ;
        RECT 150.690 37.270 151.350 40.360 ;
        RECT 149.290 36.830 150.630 36.910 ;
        RECT 149.060 36.490 150.630 36.830 ;
        RECT 150.890 36.650 151.120 37.270 ;
        RECT 151.720 36.910 152.740 46.400 ;
        RECT 153.180 46.170 153.410 46.650 ;
        RECT 153.010 37.280 153.480 46.170 ;
        RECT 153.620 40.270 154.250 42.130 ;
        RECT 151.370 36.850 152.740 36.910 ;
        RECT 151.370 36.490 152.940 36.850 ;
        RECT 153.180 36.650 153.410 37.280 ;
        RECT 144.300 36.260 146.260 36.490 ;
        RECT 146.590 36.260 148.550 36.490 ;
        RECT 148.880 36.260 150.840 36.490 ;
        RECT 151.170 36.260 153.130 36.490 ;
        RECT 144.500 35.120 146.070 36.260 ;
        RECT 146.780 35.120 148.350 36.260 ;
        RECT 149.060 35.120 150.630 36.260 ;
        RECT 151.370 35.130 152.940 36.260 ;
        RECT 145.035 34.015 145.745 35.120 ;
        RECT 147.205 34.015 147.915 35.120 ;
        RECT 149.425 34.015 150.135 35.120 ;
        RECT 151.795 34.015 152.505 35.130 ;
        RECT 145.035 33.305 152.505 34.015 ;
        RECT 133.160 31.950 140.620 32.940 ;
        RECT 133.160 23.210 134.270 31.950 ;
        RECT 133.180 23.100 133.410 23.210 ;
        RECT 131.170 22.710 133.130 22.940 ;
        RECT 142.740 22.885 143.450 22.900 ;
        RECT 146.650 22.885 147.150 22.910 ;
        RECT 150.305 22.890 151.015 33.305 ;
        RECT 150.305 22.885 151.020 22.890 ;
        RECT 131.320 22.680 133.020 22.710 ;
        RECT 132.100 21.050 132.880 22.680 ;
        RECT 139.155 22.330 151.020 22.885 ;
        RECT 139.155 22.175 151.015 22.330 ;
        RECT 131.860 20.050 135.170 21.050 ;
        RECT 113.660 19.080 114.700 19.440 ;
        RECT 110.590 17.590 111.550 18.210 ;
        RECT 113.590 17.830 115.020 19.080 ;
        RECT 139.155 17.670 139.865 22.175 ;
        RECT 142.740 21.230 143.450 22.175 ;
        RECT 142.740 20.220 144.210 21.230 ;
        RECT 145.125 21.220 145.835 22.175 ;
        RECT 146.650 22.130 147.150 22.175 ;
        RECT 144.980 20.410 146.630 21.220 ;
        RECT 147.425 21.210 148.135 22.175 ;
        RECT 145.170 20.220 146.630 20.410 ;
        RECT 147.420 20.220 148.730 21.210 ;
        RECT 150.305 21.200 151.015 22.175 ;
        RECT 149.520 20.220 151.230 21.200 ;
        RECT 142.530 19.990 144.490 20.220 ;
        RECT 144.820 19.990 146.780 20.220 ;
        RECT 147.110 19.990 149.070 20.220 ;
        RECT 149.400 19.990 151.360 20.220 ;
        RECT 142.250 19.670 142.480 19.830 ;
        RECT 141.350 17.670 142.550 19.670 ;
        RECT 110.590 17.070 114.990 17.590 ;
        RECT 134.850 17.480 142.550 17.670 ;
        RECT 134.795 17.230 142.550 17.480 ;
        RECT 110.590 16.470 111.550 17.070 ;
        RECT 134.850 17.050 142.550 17.230 ;
        RECT 141.350 14.970 142.550 17.050 ;
        RECT 142.740 19.620 144.210 19.990 ;
        RECT 142.740 15.090 144.200 19.620 ;
        RECT 144.540 19.310 144.770 19.830 ;
        RECT 145.170 19.720 146.630 19.990 ;
        RECT 146.830 19.720 147.060 19.830 ;
        RECT 144.390 15.380 144.920 19.310 ;
        RECT 142.250 14.830 142.480 14.970 ;
        RECT 142.740 14.670 144.370 15.090 ;
        RECT 144.540 14.830 144.770 15.380 ;
        RECT 145.170 15.090 146.480 19.720 ;
        RECT 146.820 19.550 147.070 19.720 ;
        RECT 147.420 19.700 148.730 19.990 ;
        RECT 146.670 15.160 147.110 19.550 ;
        RECT 144.980 14.930 146.480 15.090 ;
        RECT 146.820 15.000 147.070 15.160 ;
        RECT 147.380 15.070 148.730 19.700 ;
        RECT 149.120 19.310 149.350 19.830 ;
        RECT 149.520 19.790 151.230 19.990 ;
        RECT 149.520 19.630 151.020 19.790 ;
        RECT 148.970 17.920 149.540 19.310 ;
        RECT 148.950 16.790 149.540 17.920 ;
        RECT 148.970 15.410 149.540 16.790 ;
        RECT 144.980 14.670 146.630 14.930 ;
        RECT 146.830 14.830 147.060 15.000 ;
        RECT 147.380 14.960 148.910 15.070 ;
        RECT 147.230 14.670 148.910 14.960 ;
        RECT 149.120 14.830 149.350 15.410 ;
        RECT 149.710 15.070 151.020 19.630 ;
        RECT 151.410 19.610 151.640 19.830 ;
        RECT 151.290 15.070 151.730 19.610 ;
        RECT 149.520 14.870 151.020 15.070 ;
        RECT 149.520 14.670 151.230 14.870 ;
        RECT 151.410 14.830 151.640 15.070 ;
        RECT 151.870 14.850 152.480 18.430 ;
        RECT 142.530 14.440 144.490 14.670 ;
        RECT 144.820 14.440 146.780 14.670 ;
        RECT 147.110 14.440 149.070 14.670 ;
        RECT 149.400 14.440 151.360 14.670 ;
        RECT 142.740 14.420 144.370 14.440 ;
        RECT 144.980 14.410 146.630 14.440 ;
        RECT 147.230 14.410 148.910 14.440 ;
        RECT 149.520 14.410 151.230 14.440 ;
        RECT 154.170 11.520 155.170 13.490 ;
        RECT 128.580 7.150 129.580 9.120 ;
      LAYER met2 ;
        RECT 84.950 221.280 85.250 221.290 ;
        RECT 84.915 221.000 85.285 221.280 ;
        RECT 84.950 220.540 85.250 221.000 ;
        RECT 64.250 220.240 85.250 220.540 ;
        RECT 88.630 220.390 88.930 220.400 ;
        RECT 64.250 207.320 64.550 220.240 ;
        RECT 88.595 220.110 88.965 220.390 ;
        RECT 88.630 219.430 88.930 220.110 ;
        RECT 73.890 219.130 88.930 219.430 ;
        RECT 73.890 208.620 74.190 219.130 ;
        RECT 114.390 219.110 114.690 219.120 ;
        RECT 114.355 218.830 114.725 219.110 ;
        RECT 114.390 217.820 114.690 218.830 ;
        RECT 83.600 217.520 114.690 217.820 ;
        RECT 83.600 208.620 83.900 217.520 ;
        RECT 93.220 212.020 93.520 212.030 ;
        RECT 93.185 211.740 93.555 212.020 ;
        RECT 64.260 207.110 64.540 207.320 ;
        RECT 73.890 207.110 74.200 208.620 ;
        RECT 64.260 206.970 67.230 207.110 ;
        RECT 64.260 206.620 64.540 206.970 ;
        RECT 65.355 201.075 66.895 201.445 ;
        RECT 67.090 197.850 67.230 206.970 ;
        RECT 73.530 206.970 74.200 207.110 ;
        RECT 69.610 203.795 71.150 204.165 ;
        RECT 73.530 200.310 73.670 206.970 ;
        RECT 73.890 206.780 74.200 206.970 ;
        RECT 73.920 206.620 74.200 206.780 ;
        RECT 83.580 207.680 83.900 208.620 ;
        RECT 83.580 207.110 83.860 207.680 ;
        RECT 93.220 207.670 93.520 211.740 ;
        RECT 83.580 206.970 84.250 207.110 ;
        RECT 83.580 206.620 83.860 206.970 ;
        RECT 78.120 203.795 79.660 204.165 ;
        RECT 73.865 201.075 75.405 201.445 ;
        RECT 82.375 201.075 83.915 201.445 ;
        RECT 73.530 200.170 74.130 200.310 ;
        RECT 76.230 200.250 76.490 200.570 ;
        RECT 69.610 198.355 71.150 198.725 ;
        RECT 73.990 197.850 74.130 200.170 ;
        RECT 75.770 198.890 76.030 199.210 ;
        RECT 75.830 198.190 75.970 198.890 ;
        RECT 76.290 198.190 76.430 200.250 ;
        RECT 77.610 199.230 77.870 199.550 ;
        RECT 75.770 197.870 76.030 198.190 ;
        RECT 76.230 197.870 76.490 198.190 ;
        RECT 67.030 197.530 67.290 197.850 ;
        RECT 73.930 197.530 74.190 197.850 ;
        RECT 77.670 197.510 77.810 199.230 ;
        RECT 79.910 198.890 80.170 199.210 ;
        RECT 80.830 198.890 81.090 199.210 ;
        RECT 78.120 198.355 79.660 198.725 ;
        RECT 77.610 197.190 77.870 197.510 ;
        RECT 65.355 195.635 66.895 196.005 ;
        RECT 73.865 195.635 75.405 196.005 ;
        RECT 77.670 195.470 77.810 197.190 ;
        RECT 79.970 195.470 80.110 198.890 ;
        RECT 80.890 197.850 81.030 198.890 ;
        RECT 84.110 198.190 84.250 206.970 ;
        RECT 93.240 206.620 93.520 207.670 ;
        RECT 86.630 203.795 88.170 204.165 ;
        RECT 93.310 203.630 93.450 206.620 ;
        RECT 95.140 203.795 96.680 204.165 ;
        RECT 93.250 203.310 93.510 203.630 ;
        RECT 85.890 201.610 86.150 201.930 ;
        RECT 85.430 199.570 85.690 199.890 ;
        RECT 84.050 197.870 84.310 198.190 ;
        RECT 80.830 197.530 81.090 197.850 ;
        RECT 85.490 197.170 85.630 199.570 ;
        RECT 85.950 197.850 86.090 201.610 ;
        RECT 90.885 201.075 92.425 201.445 ;
        RECT 86.630 198.355 88.170 198.725 ;
        RECT 95.140 198.355 96.680 198.725 ;
        RECT 85.890 197.530 86.150 197.850 ;
        RECT 85.430 196.850 85.690 197.170 ;
        RECT 82.375 195.635 83.915 196.005 ;
        RECT 77.610 195.150 77.870 195.470 ;
        RECT 79.910 195.150 80.170 195.470 ;
        RECT 85.950 193.770 86.090 197.530 ;
        RECT 86.350 196.850 86.610 197.170 ;
        RECT 86.410 194.790 86.550 196.850 ;
        RECT 90.885 195.635 92.425 196.005 ;
        RECT 86.350 194.470 86.610 194.790 ;
        RECT 85.890 193.450 86.150 193.770 ;
        RECT 69.610 192.915 71.150 193.285 ;
        RECT 78.120 192.915 79.660 193.285 ;
        RECT 86.630 192.915 88.170 193.285 ;
        RECT 95.140 192.915 96.680 193.285 ;
        RECT 65.355 190.195 66.895 190.565 ;
        RECT 73.865 190.195 75.405 190.565 ;
        RECT 82.375 190.195 83.915 190.565 ;
        RECT 90.885 190.195 92.425 190.565 ;
        RECT 69.610 187.475 71.150 187.845 ;
        RECT 78.120 187.475 79.660 187.845 ;
        RECT 86.630 187.475 88.170 187.845 ;
        RECT 95.140 187.475 96.680 187.845 ;
        RECT 65.355 184.755 66.895 185.125 ;
        RECT 73.865 184.755 75.405 185.125 ;
        RECT 82.375 184.755 83.915 185.125 ;
        RECT 90.885 184.755 92.425 185.125 ;
        RECT 69.610 182.035 71.150 182.405 ;
        RECT 78.120 182.035 79.660 182.405 ;
        RECT 86.630 182.035 88.170 182.405 ;
        RECT 95.140 182.035 96.680 182.405 ;
        RECT 65.355 179.315 66.895 179.685 ;
        RECT 73.865 179.315 75.405 179.685 ;
        RECT 82.375 179.315 83.915 179.685 ;
        RECT 90.885 179.315 92.425 179.685 ;
        RECT 69.610 176.595 71.150 176.965 ;
        RECT 78.120 176.595 79.660 176.965 ;
        RECT 86.630 176.595 88.170 176.965 ;
        RECT 95.140 176.595 96.680 176.965 ;
        RECT 65.355 173.875 66.895 174.245 ;
        RECT 73.865 173.875 75.405 174.245 ;
        RECT 82.375 173.875 83.915 174.245 ;
        RECT 90.885 173.875 92.425 174.245 ;
        RECT 69.610 171.155 71.150 171.525 ;
        RECT 78.120 171.155 79.660 171.525 ;
        RECT 86.630 171.155 88.170 171.525 ;
        RECT 95.140 171.155 96.680 171.525 ;
        RECT 124.975 78.055 125.365 78.070 ;
        RECT 124.975 77.785 126.565 78.055 ;
        RECT 124.975 77.770 125.365 77.785 ;
        RECT 109.220 63.790 110.090 65.460 ;
        RECT 111.460 62.760 112.010 63.310 ;
        RECT 109.850 55.240 110.690 56.480 ;
        RECT 104.140 53.270 104.650 53.750 ;
        RECT 98.090 51.340 99.170 52.320 ;
        RECT 102.680 45.740 103.680 45.770 ;
        RECT 101.465 44.740 103.680 45.740 ;
        RECT 109.800 45.630 110.790 46.600 ;
        RECT 102.680 44.710 103.680 44.740 ;
        RECT 108.670 39.580 109.710 43.910 ;
        RECT 103.910 38.140 104.910 38.185 ;
        RECT 103.880 37.140 104.940 38.140 ;
        RECT 103.910 37.095 104.910 37.140 ;
        RECT 109.660 36.740 110.850 37.700 ;
        RECT 123.100 35.495 124.850 53.945 ;
        RECT 126.295 37.005 126.565 77.785 ;
        RECT 149.630 64.310 151.050 64.980 ;
        RECT 151.760 64.330 152.440 64.980 ;
        RECT 148.440 49.190 149.090 49.230 ;
        RECT 153.040 49.190 153.520 49.230 ;
        RECT 131.560 47.820 132.660 48.880 ;
        RECT 147.480 48.710 153.520 49.190 ;
        RECT 148.440 44.700 149.090 48.710 ;
        RECT 153.040 44.780 153.520 48.710 ;
        RECT 134.890 43.220 135.460 43.860 ;
        RECT 148.390 42.960 149.090 44.700 ;
        RECT 152.980 42.990 153.530 44.780 ;
        RECT 148.390 42.950 149.070 42.960 ;
        RECT 146.050 40.430 146.790 41.950 ;
        RECT 150.600 40.410 151.360 41.970 ;
        RECT 153.520 40.320 154.300 42.080 ;
        RECT 128.960 39.160 129.500 39.790 ;
        RECT 131.590 39.320 132.170 39.820 ;
        RECT 137.610 39.230 138.180 39.760 ;
        RECT 131.130 37.640 131.700 38.590 ;
        RECT 130.585 37.005 130.855 37.055 ;
        RECT 126.295 36.735 130.855 37.005 ;
        RECT 130.585 36.685 130.855 36.735 ;
        RECT 123.100 33.745 128.815 35.495 ;
        RECT 131.510 34.820 132.530 35.610 ;
        RECT 98.230 32.230 99.190 33.200 ;
        RECT 123.100 31.125 124.850 33.745 ;
        RECT 104.130 30.160 105.080 31.020 ;
        RECT 123.070 29.375 124.880 31.125 ;
        RECT 109.670 27.770 110.810 28.640 ;
        RECT 146.640 22.860 147.150 22.900 ;
        RECT 146.600 22.180 147.200 22.860 ;
        RECT 150.490 22.360 151.770 22.860 ;
        RECT 134.140 21.050 135.140 21.080 ;
        RECT 134.140 20.050 136.355 21.050 ;
        RECT 134.140 20.020 135.140 20.050 ;
        RECT 113.610 18.520 114.750 19.390 ;
        RECT 146.640 19.250 147.150 22.180 ;
        RECT 146.620 18.530 147.150 19.250 ;
        RECT 151.270 19.130 151.770 22.360 ;
        RECT 151.240 18.490 151.780 19.130 ;
        RECT 110.540 16.520 111.600 18.160 ;
        RECT 144.360 16.820 144.940 17.850 ;
        RECT 148.900 16.840 149.540 17.870 ;
        RECT 151.840 16.300 152.460 17.010 ;
        RECT 154.170 13.460 155.170 14.605 ;
        RECT 154.140 12.460 155.200 13.460 ;
        RECT 128.580 9.090 129.580 9.975 ;
        RECT 128.550 8.090 129.610 9.090 ;
      LAYER met3 ;
        RECT 84.910 221.760 85.290 222.080 ;
        RECT 84.950 221.305 85.250 221.760 ;
        RECT 88.590 221.490 88.970 221.810 ;
        RECT 84.935 220.975 85.265 221.305 ;
        RECT 88.630 220.415 88.930 221.490 ;
        RECT 149.950 220.900 150.270 220.940 ;
        RECT 93.220 220.600 150.270 220.900 ;
        RECT 88.615 220.085 88.945 220.415 ;
        RECT 93.220 212.045 93.520 220.600 ;
        RECT 149.950 220.560 150.270 220.600 ;
        RECT 114.350 219.760 114.730 220.080 ;
        RECT 114.390 219.135 114.690 219.760 ;
        RECT 114.375 218.805 114.705 219.135 ;
        RECT 93.205 211.715 93.535 212.045 ;
        RECT 118.030 209.370 118.410 209.690 ;
        RECT 118.070 206.830 118.370 209.370 ;
        RECT 118.060 206.450 118.380 206.830 ;
        RECT 69.590 203.815 71.170 204.145 ;
        RECT 78.100 203.815 79.680 204.145 ;
        RECT 86.610 203.815 88.190 204.145 ;
        RECT 95.120 203.815 96.700 204.145 ;
        RECT 65.335 201.095 66.915 201.425 ;
        RECT 73.845 201.095 75.425 201.425 ;
        RECT 82.355 201.095 83.935 201.425 ;
        RECT 90.865 201.095 92.445 201.425 ;
        RECT 69.590 198.375 71.170 198.705 ;
        RECT 78.100 198.375 79.680 198.705 ;
        RECT 86.610 198.375 88.190 198.705 ;
        RECT 95.120 198.375 96.700 198.705 ;
        RECT 65.335 195.655 66.915 195.985 ;
        RECT 73.845 195.655 75.425 195.985 ;
        RECT 82.355 195.655 83.935 195.985 ;
        RECT 90.865 195.655 92.445 195.985 ;
        RECT 69.590 192.935 71.170 193.265 ;
        RECT 78.100 192.935 79.680 193.265 ;
        RECT 86.610 192.935 88.190 193.265 ;
        RECT 95.120 192.935 96.700 193.265 ;
        RECT 65.335 190.215 66.915 190.545 ;
        RECT 73.845 190.215 75.425 190.545 ;
        RECT 82.355 190.215 83.935 190.545 ;
        RECT 90.865 190.215 92.445 190.545 ;
        RECT 69.590 187.495 71.170 187.825 ;
        RECT 78.100 187.495 79.680 187.825 ;
        RECT 86.610 187.495 88.190 187.825 ;
        RECT 95.120 187.495 96.700 187.825 ;
        RECT 65.335 184.775 66.915 185.105 ;
        RECT 73.845 184.775 75.425 185.105 ;
        RECT 82.355 184.775 83.935 185.105 ;
        RECT 90.865 184.775 92.445 185.105 ;
        RECT 69.590 182.055 71.170 182.385 ;
        RECT 78.100 182.055 79.680 182.385 ;
        RECT 86.610 182.055 88.190 182.385 ;
        RECT 95.120 182.055 96.700 182.385 ;
        RECT 65.335 179.335 66.915 179.665 ;
        RECT 73.845 179.335 75.425 179.665 ;
        RECT 82.355 179.335 83.935 179.665 ;
        RECT 90.865 179.335 92.445 179.665 ;
        RECT 69.590 176.615 71.170 176.945 ;
        RECT 78.100 176.615 79.680 176.945 ;
        RECT 86.610 176.615 88.190 176.945 ;
        RECT 95.120 176.615 96.700 176.945 ;
        RECT 65.335 173.895 66.915 174.225 ;
        RECT 73.845 173.895 75.425 174.225 ;
        RECT 82.355 173.895 83.935 174.225 ;
        RECT 90.865 173.895 92.445 174.225 ;
        RECT 69.590 171.175 71.170 171.505 ;
        RECT 78.100 171.175 79.680 171.505 ;
        RECT 86.610 171.175 88.190 171.505 ;
        RECT 95.120 171.175 96.700 171.505 ;
        RECT 52.965 168.440 54.555 168.465 ;
        RECT 45.290 166.840 54.560 168.440 ;
        RECT 52.965 166.815 54.555 166.840 ;
        RECT 118.030 84.160 118.410 84.480 ;
        RECT 118.070 83.140 118.370 84.160 ;
        RECT 118.060 82.760 118.380 83.140 ;
        RECT 123.950 78.070 124.330 78.080 ;
        RECT 124.995 78.070 125.345 78.095 ;
        RECT 123.950 77.770 125.345 78.070 ;
        RECT 123.950 77.760 124.330 77.770 ;
        RECT 124.995 77.745 125.345 77.770 ;
        RECT 109.245 63.740 110.065 65.510 ;
        RECT 149.655 64.260 151.025 65.030 ;
        RECT 151.785 64.280 152.415 65.030 ;
        RECT 111.485 62.710 111.985 63.360 ;
        RECT 109.875 55.190 110.665 56.530 ;
        RECT 104.165 53.220 104.625 53.800 ;
        RECT 98.115 51.290 99.145 52.370 ;
        RECT 131.585 47.770 132.635 48.930 ;
        RECT 101.485 45.740 102.535 45.765 ;
        RECT 95.550 44.740 102.535 45.740 ;
        RECT 109.825 45.580 110.765 46.650 ;
        RECT 42.945 21.390 44.435 21.415 ;
        RECT 42.940 19.890 54.520 21.390 ;
        RECT 42.945 19.865 44.435 19.890 ;
        RECT 95.550 4.650 96.550 44.740 ;
        RECT 101.485 44.715 102.535 44.740 ;
        RECT 134.915 43.170 135.435 43.910 ;
        RECT 146.075 40.380 146.765 42.000 ;
        RECT 150.625 40.360 151.335 42.020 ;
        RECT 153.545 40.270 154.275 42.130 ;
        RECT 128.985 39.110 129.475 39.840 ;
        RECT 131.615 39.270 132.145 39.870 ;
        RECT 137.635 39.180 138.155 39.810 ;
        RECT 103.885 37.115 104.935 38.165 ;
        RECT 103.910 36.610 104.910 37.115 ;
        RECT 109.685 36.690 110.825 37.750 ;
        RECT 131.155 37.590 131.675 38.640 ;
        RECT 101.560 35.610 104.910 36.610 ;
        RECT 98.255 32.180 99.165 33.250 ;
        RECT 101.560 6.440 102.560 35.610 ;
        RECT 131.535 34.770 132.505 35.660 ;
        RECT 104.155 30.110 105.055 31.070 ;
        RECT 109.695 27.720 110.785 28.690 ;
        RECT 135.285 21.050 136.335 21.075 ;
        RECT 135.285 20.050 157.270 21.050 ;
        RECT 135.285 20.025 136.335 20.050 ;
        RECT 113.635 18.470 114.725 19.440 ;
        RECT 110.565 16.470 111.575 18.210 ;
        RECT 144.385 16.770 144.915 17.900 ;
        RECT 148.925 16.790 149.515 17.920 ;
        RECT 151.865 16.250 152.435 17.060 ;
        RECT 154.170 14.585 155.170 15.530 ;
        RECT 154.145 13.535 155.195 14.585 ;
        RECT 128.580 9.955 129.580 10.810 ;
        RECT 128.555 8.905 129.605 9.955 ;
        RECT 101.560 5.780 135.210 6.440 ;
        RECT 101.560 5.440 135.230 5.780 ;
        RECT 95.550 3.650 113.300 4.650 ;
        RECT 134.210 4.370 135.230 5.440 ;
        RECT 112.250 3.440 113.300 3.650 ;
        RECT 112.250 2.665 113.150 3.440 ;
        RECT 134.330 3.225 135.230 4.370 ;
        RECT 112.225 1.775 113.175 2.665 ;
        RECT 134.305 2.335 135.255 3.225 ;
        RECT 156.270 2.720 157.270 20.050 ;
        RECT 134.330 2.330 135.230 2.335 ;
        RECT 112.250 1.770 113.150 1.775 ;
      LAYER met4 ;
        RECT 3.980 224.760 3.990 225.250 ;
        RECT 3.980 223.750 4.280 224.760 ;
        RECT 7.670 223.750 7.970 224.760 ;
        RECT 11.350 223.750 11.650 224.760 ;
        RECT 15.030 223.750 15.330 224.760 ;
        RECT 18.710 223.750 19.010 224.760 ;
        RECT 22.390 223.750 22.690 224.760 ;
        RECT 26.070 223.750 26.370 224.760 ;
        RECT 29.750 223.750 30.050 224.760 ;
        RECT 33.430 223.750 33.730 224.760 ;
        RECT 37.110 223.750 37.410 224.760 ;
        RECT 40.790 223.750 41.090 224.760 ;
        RECT 44.470 223.750 44.770 224.760 ;
        RECT 48.150 223.750 48.450 224.760 ;
        RECT 51.830 223.750 52.130 224.760 ;
        RECT 55.510 223.750 55.810 224.760 ;
        RECT 59.190 223.750 59.490 224.760 ;
        RECT 62.870 223.750 63.170 224.760 ;
        RECT 66.550 223.750 66.850 224.760 ;
        RECT 70.230 223.750 70.530 224.760 ;
        RECT 73.910 223.750 74.210 224.760 ;
        RECT 77.590 223.750 77.890 224.760 ;
        RECT 81.270 223.750 81.570 224.760 ;
        RECT 3.980 223.450 81.900 223.750 ;
        RECT 5.480 223.420 6.980 223.450 ;
        RECT 15.030 223.410 15.330 223.450 ;
        RECT 18.710 223.440 22.710 223.450 ;
        RECT 26.070 223.420 26.370 223.450 ;
        RECT 29.750 223.400 30.050 223.450 ;
        RECT 44.470 223.420 44.770 223.450 ;
        RECT 2.500 219.050 2.520 220.550 ;
        RECT 45.230 220.110 45.530 223.450 ;
        RECT 51.830 223.420 52.130 223.450 ;
        RECT 55.510 223.440 55.810 223.450 ;
        RECT 59.190 223.440 59.490 223.450 ;
        RECT 62.870 223.390 63.170 223.450 ;
        RECT 84.950 222.085 85.250 224.760 ;
        RECT 84.935 221.755 85.265 222.085 ;
        RECT 88.630 221.815 88.930 224.760 ;
        RECT 88.615 221.485 88.945 221.815 ;
        RECT 45.230 219.810 49.000 220.110 ;
        RECT 114.390 220.085 114.690 224.760 ;
        RECT 114.375 219.755 114.705 220.085 ;
        RECT 118.070 209.695 118.370 224.760 ;
        RECT 149.945 220.900 150.275 220.915 ;
        RECT 151.190 220.900 151.490 224.760 ;
        RECT 149.945 220.600 151.490 220.900 ;
        RECT 149.945 220.585 150.275 220.600 ;
        RECT 118.055 209.365 118.385 209.695 ;
        RECT 118.055 206.475 118.385 206.805 ;
        RECT 65.325 171.630 66.925 204.220 ;
        RECT 69.580 171.810 71.180 204.220 ;
        RECT 65.310 171.100 66.925 171.630 ;
        RECT 45.315 168.440 46.925 168.445 ;
        RECT 65.310 168.440 66.910 171.100 ;
        RECT 0.900 166.840 1.000 168.440 ;
        RECT 2.500 166.840 46.925 168.440 ;
        RECT 52.960 166.840 66.910 168.440 ;
        RECT 45.315 166.835 46.925 166.840 ;
        RECT 69.560 163.975 71.230 171.810 ;
        RECT 73.835 171.100 75.435 204.220 ;
        RECT 78.090 171.100 79.690 204.220 ;
        RECT 82.345 171.100 83.945 204.220 ;
        RECT 86.600 171.100 88.200 204.220 ;
        RECT 90.855 171.100 92.455 204.220 ;
        RECT 95.110 171.100 96.710 204.220 ;
        RECT 48.985 162.305 49.000 163.975 ;
        RECT 50.500 162.305 71.230 163.975 ;
        RECT 118.070 84.485 118.370 206.475 ;
        RECT 118.055 84.155 118.385 84.485 ;
        RECT 118.055 82.785 118.385 83.115 ;
        RECT 118.070 78.070 118.370 82.785 ;
        RECT 123.975 78.070 124.305 78.085 ;
        RECT 117.980 77.770 124.305 78.070 ;
        RECT 118.070 77.250 118.370 77.770 ;
        RECT 123.975 77.755 124.305 77.770 ;
        RECT 50.500 71.880 149.390 71.980 ;
        RECT 50.500 70.940 149.400 71.880 ;
        RECT 50.500 70.480 149.390 70.940 ;
        RECT 109.265 65.450 110.045 65.465 ;
        RECT 97.830 63.810 110.045 65.450 ;
        RECT 52.985 21.390 54.495 21.395 ;
        RECT 97.830 21.390 99.470 63.810 ;
        RECT 109.265 63.785 110.045 63.810 ;
        RECT 147.890 65.370 149.390 70.480 ;
        RECT 147.890 63.870 153.360 65.370 ;
        RECT 110.720 60.810 112.220 63.340 ;
        RECT 109.270 60.100 132.930 60.810 ;
        RECT 147.890 60.100 150.680 63.870 ;
        RECT 109.270 59.310 150.680 60.100 ;
        RECT 109.270 54.550 110.770 59.310 ;
        RECT 103.400 53.050 110.770 54.550 ;
        RECT 109.270 37.705 110.770 53.050 ;
        RECT 131.430 58.600 150.680 59.310 ;
        RECT 131.430 48.340 132.930 58.600 ;
        RECT 131.430 46.840 138.710 48.340 ;
        RECT 127.890 42.720 135.990 44.360 ;
        RECT 109.270 36.735 110.805 37.705 ;
        RECT 109.270 31.370 110.770 36.735 ;
        RECT 103.940 29.870 110.770 31.370 ;
        RECT 2.500 19.890 44.440 21.390 ;
        RECT 52.985 19.890 99.470 21.390 ;
        RECT 109.270 21.650 110.770 29.870 ;
        RECT 109.270 20.150 114.800 21.650 ;
        RECT 52.985 19.885 54.495 19.890 ;
        RECT 93.510 19.690 95.010 19.890 ;
        RECT 97.830 18.150 99.470 19.890 ;
        RECT 113.300 18.900 114.800 20.150 ;
        RECT 113.655 18.515 114.705 18.900 ;
        RECT 110.585 18.150 111.555 18.165 ;
        RECT 97.830 16.515 111.555 18.150 ;
        RECT 97.830 16.510 111.420 16.515 ;
        RECT 107.700 12.980 109.340 16.510 ;
        RECT 127.890 12.980 129.530 42.720 ;
        RECT 131.570 39.270 132.590 39.880 ;
        RECT 131.590 38.595 132.590 39.270 ;
        RECT 131.175 37.635 132.590 38.595 ;
        RECT 131.570 36.140 132.590 37.635 ;
        RECT 137.210 36.140 138.710 46.840 ;
        RECT 149.180 41.975 150.680 58.600 ;
        RECT 146.095 41.660 146.745 41.955 ;
        RECT 149.180 41.660 151.315 41.975 ;
        RECT 153.565 41.660 154.255 42.085 ;
        RECT 144.840 40.160 155.170 41.660 ;
        RECT 131.000 34.640 138.710 36.140 ;
        RECT 144.405 17.670 144.895 17.855 ;
        RECT 148.945 17.670 149.495 17.875 ;
        RECT 153.670 17.670 155.170 40.160 ;
        RECT 143.440 16.170 155.170 17.670 ;
        RECT 154.170 15.505 155.170 16.170 ;
        RECT 154.165 14.495 155.175 15.505 ;
        RECT 107.700 12.470 129.530 12.980 ;
        RECT 107.700 11.340 129.580 12.470 ;
        RECT 128.580 10.785 129.580 11.340 ;
        RECT 128.575 9.775 129.585 10.785 ;
        RECT 112.250 1.000 113.150 2.670 ;
        RECT 134.330 1.000 135.230 3.230 ;
        RECT 156.265 2.745 157.275 3.755 ;
        RECT 156.270 1.000 157.270 2.745 ;
        RECT 156.270 0.030 156.410 1.000 ;
  END
END tt_um_brucemack_sb_mixer
END LIBRARY

