VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_lcasimon_tdc
  CLASS BLOCK ;
  FOREIGN tt_um_lcasimon_tdc ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 86.799995 ;
    ANTENNADIFFAREA 3.136000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 107.460 173.520 110.295 173.950 ;
        RECT 107.460 169.170 107.890 173.520 ;
        RECT 108.065 169.370 109.325 173.320 ;
        RECT 107.460 168.740 110.295 169.170 ;
      LAYER nwell ;
        RECT 110.395 168.690 114.355 174.000 ;
        RECT 56.000 113.440 62.890 151.600 ;
      LAYER pwell ;
        RECT 64.305 151.120 67.005 151.550 ;
        RECT 64.305 142.530 64.735 151.120 ;
        RECT 65.275 142.730 66.035 150.920 ;
        RECT 66.575 142.530 67.005 151.120 ;
        RECT 91.785 151.120 94.485 151.550 ;
        RECT 64.305 142.100 67.005 142.530 ;
        RECT 72.460 142.400 77.900 142.830 ;
        RECT 64.305 137.910 67.005 138.340 ;
        RECT 64.305 117.640 64.735 137.910 ;
        RECT 65.275 117.840 66.035 137.710 ;
        RECT 66.575 117.640 67.005 137.910 ;
        RECT 64.305 117.210 67.005 117.640 ;
      LAYER nwell ;
        RECT 68.010 117.160 71.310 138.390 ;
        RECT 56.000 111.570 67.465 113.440 ;
      LAYER pwell ;
        RECT 67.540 112.960 70.375 113.390 ;
      LAYER nwell ;
        RECT 63.505 88.770 67.465 111.570 ;
      LAYER pwell ;
        RECT 68.985 89.450 69.745 112.760 ;
        RECT 69.945 89.250 70.375 112.960 ;
        RECT 72.460 113.090 72.890 142.400 ;
        RECT 73.430 113.250 74.190 142.240 ;
        RECT 76.170 113.650 76.930 141.840 ;
        RECT 77.470 113.090 77.900 142.400 ;
        RECT 72.460 112.660 77.900 113.090 ;
        RECT 80.890 142.400 86.330 142.830 ;
        RECT 80.890 113.090 81.320 142.400 ;
        RECT 81.860 113.650 82.620 141.840 ;
        RECT 84.600 113.250 85.360 142.240 ;
        RECT 85.900 113.090 86.330 142.400 ;
        RECT 91.785 142.530 92.215 151.120 ;
        RECT 92.755 142.730 93.515 150.920 ;
        RECT 94.055 142.530 94.485 151.120 ;
        RECT 91.785 142.100 94.485 142.530 ;
      LAYER nwell ;
        RECT 87.480 117.160 90.780 138.390 ;
      LAYER pwell ;
        RECT 91.785 137.910 94.485 138.340 ;
        RECT 91.785 117.640 92.215 137.910 ;
        RECT 92.755 117.840 93.515 137.710 ;
        RECT 94.055 117.640 94.485 137.910 ;
        RECT 91.785 117.210 94.485 117.640 ;
      LAYER nwell ;
        RECT 95.900 113.440 102.790 151.600 ;
      LAYER pwell ;
        RECT 80.890 112.660 86.330 113.090 ;
        RECT 88.415 112.960 91.250 113.390 ;
        RECT 67.540 88.820 70.375 89.250 ;
        RECT 88.415 89.250 88.845 112.960 ;
        RECT 89.045 89.450 89.805 112.760 ;
      LAYER nwell ;
        RECT 91.325 111.570 102.790 113.440 ;
        RECT 108.455 113.625 114.195 164.850 ;
      LAYER pwell ;
        RECT 121.710 164.330 125.980 164.760 ;
        RECT 114.795 117.970 117.695 118.205 ;
        RECT 121.710 117.970 122.140 164.330 ;
        RECT 114.795 117.775 122.140 117.970 ;
        RECT 114.795 114.365 115.225 117.775 ;
        RECT 115.765 114.525 116.725 117.615 ;
        RECT 117.265 117.540 122.140 117.775 ;
        RECT 117.265 114.365 118.495 117.540 ;
        RECT 114.795 113.935 118.495 114.365 ;
        RECT 88.415 88.820 91.250 89.250 ;
      LAYER nwell ;
        RECT 91.325 88.770 95.285 111.570 ;
        RECT 108.455 109.175 117.745 113.625 ;
      LAYER pwell ;
        RECT 118.065 109.830 118.495 113.935 ;
        RECT 119.035 109.990 120.295 117.380 ;
        RECT 120.835 109.830 122.140 117.540 ;
        RECT 118.065 109.400 122.140 109.830 ;
        RECT 71.345 82.290 74.460 82.720 ;
        RECT 71.345 77.940 71.775 82.290 ;
        RECT 72.315 78.140 73.575 82.090 ;
        RECT 71.345 77.510 74.460 77.940 ;
      LAYER nwell ;
        RECT 74.680 77.460 83.880 82.770 ;
      LAYER pwell ;
        RECT 84.100 82.290 87.215 82.720 ;
        RECT 84.985 78.140 86.245 82.090 ;
        RECT 86.785 77.940 87.215 82.290 ;
        RECT 84.100 77.510 87.215 77.940 ;
        RECT 88.375 82.640 91.210 83.070 ;
        RECT 88.375 78.290 88.805 82.640 ;
        RECT 88.980 78.490 90.240 82.440 ;
        RECT 88.375 77.860 91.210 78.290 ;
      LAYER nwell ;
        RECT 91.310 77.810 95.270 83.120 ;
        RECT 108.455 79.425 114.195 109.175 ;
      LAYER pwell ;
        RECT 114.795 83.770 117.695 84.005 ;
        RECT 121.710 83.770 122.140 109.400 ;
        RECT 114.795 83.575 122.140 83.770 ;
        RECT 114.795 80.165 115.225 83.575 ;
        RECT 115.765 80.325 116.725 83.415 ;
        RECT 117.265 83.340 122.140 83.575 ;
        RECT 117.265 80.165 118.495 83.340 ;
        RECT 114.795 79.735 118.495 80.165 ;
        RECT 64.595 71.980 67.430 72.410 ;
        RECT 64.595 63.330 65.025 71.980 ;
        RECT 65.200 63.530 66.460 71.780 ;
        RECT 64.595 62.900 67.430 63.330 ;
      LAYER nwell ;
        RECT 67.530 62.850 71.490 72.460 ;
      LAYER pwell ;
        RECT 73.615 71.980 76.450 72.410 ;
        RECT 73.615 63.330 74.045 71.980 ;
        RECT 74.220 63.530 75.480 71.780 ;
        RECT 73.615 62.900 76.450 63.330 ;
      LAYER nwell ;
        RECT 76.550 62.850 83.940 72.460 ;
      LAYER pwell ;
        RECT 84.040 71.980 86.875 72.410 ;
        RECT 85.010 63.530 86.270 71.780 ;
        RECT 86.445 63.330 86.875 71.980 ;
        RECT 84.040 62.900 86.875 63.330 ;
        RECT 88.375 71.980 91.210 72.410 ;
        RECT 88.375 63.330 88.805 71.980 ;
        RECT 88.980 63.530 90.240 71.780 ;
        RECT 88.375 62.900 91.210 63.330 ;
      LAYER nwell ;
        RECT 91.310 62.850 95.270 72.460 ;
        RECT 108.455 70.450 117.745 79.425 ;
      LAYER pwell ;
        RECT 118.065 75.630 118.495 79.735 ;
        RECT 119.035 75.790 120.295 83.180 ;
        RECT 120.835 76.860 122.140 83.340 ;
        RECT 122.680 77.020 123.640 164.170 ;
        RECT 124.050 77.020 125.010 164.170 ;
        RECT 125.550 76.860 125.980 164.330 ;
        RECT 120.835 76.430 125.980 76.860 ;
        RECT 120.835 75.630 121.265 76.430 ;
        RECT 118.065 75.200 121.265 75.630 ;
      LAYER nwell ;
        RECT 108.455 65.140 124.005 70.450 ;
      LAYER pwell ;
        RECT 124.325 69.930 127.225 70.360 ;
      LAYER nwell ;
        RECT 108.455 62.660 117.745 65.140 ;
      LAYER pwell ;
        RECT 124.325 65.110 124.755 69.930 ;
      LAYER nwell ;
        RECT 114.590 59.740 117.745 62.660 ;
      LAYER pwell ;
        RECT 118.340 64.680 124.755 65.110 ;
        RECT 118.340 60.410 118.770 64.680 ;
        RECT 119.310 60.570 120.270 64.520 ;
        RECT 122.025 60.570 122.985 64.520 ;
        RECT 123.525 60.500 124.755 64.680 ;
        RECT 125.295 60.660 126.255 69.770 ;
        RECT 126.795 60.500 127.225 69.930 ;
        RECT 123.525 60.410 127.225 60.500 ;
        RECT 118.340 60.070 127.225 60.410 ;
        RECT 118.340 59.980 123.955 60.070 ;
      LAYER li1 ;
        RECT 107.590 173.650 110.165 173.820 ;
        RECT 110.575 173.650 114.175 173.820 ;
        RECT 107.590 169.040 107.760 173.650 ;
        RECT 108.195 172.980 109.195 173.150 ;
        RECT 111.545 172.980 113.545 173.150 ;
        RECT 108.195 172.550 109.195 172.720 ;
        RECT 109.365 172.370 109.695 172.900 ;
        RECT 111.045 172.370 111.375 172.900 ;
        RECT 111.545 172.550 113.545 172.720 ;
        RECT 108.195 172.120 109.195 172.290 ;
        RECT 111.545 172.120 113.545 172.290 ;
        RECT 108.195 171.690 109.195 171.860 ;
        RECT 109.365 171.510 109.695 172.040 ;
        RECT 111.045 171.510 111.375 172.040 ;
        RECT 111.545 171.690 113.545 171.860 ;
        RECT 108.195 171.260 109.195 171.430 ;
        RECT 111.545 171.260 113.545 171.430 ;
        RECT 108.195 170.830 109.195 171.000 ;
        RECT 109.365 170.650 109.695 171.180 ;
        RECT 111.045 170.650 111.375 171.180 ;
        RECT 111.545 170.830 113.545 171.000 ;
        RECT 108.195 170.400 109.195 170.570 ;
        RECT 111.545 170.400 113.545 170.570 ;
        RECT 108.195 169.970 109.195 170.140 ;
        RECT 109.365 169.790 109.695 170.320 ;
        RECT 111.045 169.790 111.375 170.320 ;
        RECT 111.545 169.970 113.545 170.140 ;
        RECT 108.195 169.540 109.195 169.710 ;
        RECT 111.545 169.540 113.545 169.710 ;
        RECT 114.005 169.040 114.175 173.650 ;
        RECT 107.590 168.870 110.165 169.040 ;
        RECT 110.575 168.870 114.175 169.040 ;
        RECT 108.635 164.500 114.015 164.670 ;
        RECT 56.180 151.250 62.710 151.420 ;
        RECT 56.180 111.920 56.350 151.250 ;
        RECT 60.740 150.580 61.740 150.750 ;
        RECT 60.240 149.440 60.570 150.330 ;
        RECT 60.740 149.800 61.740 149.970 ;
        RECT 60.740 149.020 61.740 149.190 ;
        RECT 61.910 147.160 62.240 148.770 ;
        RECT 60.740 146.740 61.740 146.910 ;
        RECT 61.910 144.880 62.240 146.490 ;
        RECT 60.740 144.460 61.740 144.630 ;
        RECT 60.240 143.320 60.570 144.210 ;
        RECT 60.740 143.680 61.740 143.850 ;
        RECT 60.740 142.900 61.740 143.070 ;
        RECT 60.240 141.760 60.570 142.650 ;
        RECT 60.740 142.120 61.740 142.290 ;
        RECT 57.150 141.340 58.150 141.510 ;
        RECT 60.740 141.340 61.740 141.510 ;
        RECT 58.320 139.480 58.650 141.090 ;
        RECT 60.240 139.480 60.570 141.090 ;
        RECT 61.910 139.480 62.240 141.090 ;
        RECT 57.150 139.060 58.150 139.230 ;
        RECT 60.740 139.060 61.740 139.230 ;
        RECT 58.320 137.200 58.650 138.810 ;
        RECT 60.240 137.200 60.570 138.810 ;
        RECT 61.910 137.200 62.240 138.810 ;
        RECT 57.150 136.780 58.150 136.950 ;
        RECT 60.740 136.780 61.740 136.950 ;
        RECT 58.320 134.920 58.650 136.530 ;
        RECT 60.240 134.920 60.570 136.530 ;
        RECT 61.910 134.920 62.240 136.530 ;
        RECT 57.150 134.500 58.150 134.670 ;
        RECT 60.740 134.500 61.740 134.670 ;
        RECT 58.320 132.640 58.650 134.250 ;
        RECT 60.240 132.640 60.570 134.250 ;
        RECT 61.910 132.640 62.240 134.250 ;
        RECT 57.150 132.220 58.150 132.390 ;
        RECT 60.740 132.220 61.740 132.390 ;
        RECT 58.320 130.360 58.650 131.970 ;
        RECT 60.240 130.360 60.570 131.970 ;
        RECT 61.910 130.360 62.240 131.970 ;
        RECT 57.150 129.940 58.150 130.110 ;
        RECT 60.740 129.940 61.740 130.110 ;
        RECT 56.650 128.080 56.980 129.690 ;
        RECT 60.240 128.080 60.570 129.690 ;
        RECT 61.910 128.080 62.240 129.690 ;
        RECT 57.150 127.660 58.150 127.830 ;
        RECT 60.740 127.660 61.740 127.830 ;
        RECT 56.650 125.800 56.980 127.410 ;
        RECT 60.240 125.800 60.570 127.410 ;
        RECT 61.910 125.800 62.240 127.410 ;
        RECT 57.150 125.380 58.150 125.550 ;
        RECT 60.740 125.380 61.740 125.550 ;
        RECT 58.320 123.520 58.650 125.130 ;
        RECT 60.240 123.520 60.570 125.130 ;
        RECT 61.910 123.520 62.240 125.130 ;
        RECT 57.150 123.100 58.150 123.270 ;
        RECT 60.740 123.100 61.740 123.270 ;
        RECT 58.320 121.240 58.650 122.850 ;
        RECT 60.240 121.240 60.570 122.850 ;
        RECT 61.910 121.240 62.240 122.850 ;
        RECT 57.150 120.820 58.150 120.990 ;
        RECT 60.740 120.820 61.740 120.990 ;
        RECT 58.320 118.960 58.650 120.570 ;
        RECT 60.240 118.960 60.570 120.570 ;
        RECT 61.910 118.960 62.240 120.570 ;
        RECT 57.150 118.540 58.150 118.710 ;
        RECT 60.740 118.540 61.740 118.710 ;
        RECT 58.320 116.680 58.650 118.290 ;
        RECT 60.240 116.680 60.570 118.290 ;
        RECT 61.910 116.680 62.240 118.290 ;
        RECT 57.150 116.260 58.150 116.430 ;
        RECT 60.740 116.260 61.740 116.430 ;
        RECT 58.320 114.400 58.650 116.010 ;
        RECT 60.240 114.400 60.570 116.010 ;
        RECT 61.910 114.400 62.240 116.010 ;
        RECT 57.150 113.980 58.150 114.150 ;
        RECT 60.740 113.980 61.740 114.150 ;
        RECT 60.240 112.840 60.570 113.730 ;
        RECT 60.740 113.200 61.740 113.370 ;
        RECT 60.740 112.420 61.740 112.590 ;
        RECT 62.540 111.920 62.710 151.250 ;
        RECT 64.435 151.250 66.875 151.420 ;
        RECT 64.435 142.400 64.605 151.250 ;
        RECT 65.405 150.580 65.905 150.750 ;
        RECT 65.405 149.800 65.905 149.970 ;
        RECT 66.075 149.440 66.405 150.330 ;
        RECT 65.405 149.020 65.905 149.190 ;
        RECT 64.905 147.160 65.235 148.770 ;
        RECT 65.405 146.740 65.905 146.910 ;
        RECT 64.905 144.880 65.235 146.490 ;
        RECT 65.405 144.460 65.905 144.630 ;
        RECT 65.405 143.680 65.905 143.850 ;
        RECT 66.075 143.320 66.405 144.210 ;
        RECT 65.405 142.900 65.905 143.070 ;
        RECT 66.705 142.400 66.875 151.250 ;
        RECT 91.915 151.250 94.355 151.420 ;
        RECT 64.435 142.230 66.875 142.400 ;
        RECT 72.590 142.530 77.770 142.700 ;
        RECT 64.435 138.040 66.875 138.210 ;
        RECT 64.435 117.510 64.605 138.040 ;
        RECT 65.405 137.370 65.905 137.540 ;
        RECT 64.905 135.185 65.235 137.155 ;
        RECT 65.405 136.090 65.905 136.260 ;
        RECT 66.075 135.185 66.405 137.155 ;
        RECT 65.405 134.810 65.905 134.980 ;
        RECT 64.905 132.950 65.235 134.560 ;
        RECT 66.075 132.950 66.405 134.560 ;
        RECT 65.405 132.530 65.905 132.700 ;
        RECT 64.905 130.670 65.235 132.280 ;
        RECT 66.075 130.670 66.405 132.280 ;
        RECT 65.405 130.250 65.905 130.420 ;
        RECT 64.905 128.065 65.235 130.035 ;
        RECT 65.405 128.970 65.905 129.140 ;
        RECT 66.075 128.065 66.405 130.035 ;
        RECT 65.405 127.690 65.905 127.860 ;
        RECT 64.905 125.505 65.235 127.475 ;
        RECT 65.405 126.410 65.905 126.580 ;
        RECT 66.075 125.505 66.405 127.475 ;
        RECT 65.405 125.130 65.905 125.300 ;
        RECT 64.905 123.270 65.235 124.880 ;
        RECT 65.405 122.850 65.905 123.020 ;
        RECT 64.905 120.990 65.235 122.600 ;
        RECT 65.405 120.570 65.905 120.740 ;
        RECT 64.905 118.385 65.235 120.355 ;
        RECT 65.405 119.290 65.905 119.460 ;
        RECT 66.075 118.385 66.405 120.355 ;
        RECT 65.405 118.010 65.905 118.180 ;
        RECT 66.705 117.510 66.875 138.040 ;
        RECT 64.435 117.340 66.875 117.510 ;
        RECT 68.190 138.040 71.130 138.210 ;
        RECT 68.190 117.510 68.360 138.040 ;
        RECT 69.160 137.370 70.160 137.540 ;
        RECT 68.660 135.185 68.990 137.155 ;
        RECT 69.160 136.090 70.160 136.260 ;
        RECT 70.330 135.185 70.660 137.155 ;
        RECT 69.160 134.810 70.160 134.980 ;
        RECT 68.660 132.950 68.990 134.560 ;
        RECT 70.330 132.950 70.660 134.560 ;
        RECT 69.160 132.530 70.160 132.700 ;
        RECT 68.660 130.670 68.990 132.280 ;
        RECT 70.330 130.670 70.660 132.280 ;
        RECT 69.160 130.250 70.160 130.420 ;
        RECT 68.660 128.065 68.990 130.035 ;
        RECT 69.160 128.970 70.160 129.140 ;
        RECT 70.330 128.065 70.660 130.035 ;
        RECT 69.160 127.690 70.160 127.860 ;
        RECT 68.660 125.505 68.990 127.475 ;
        RECT 69.160 126.410 70.160 126.580 ;
        RECT 70.330 125.505 70.660 127.475 ;
        RECT 69.160 125.130 70.160 125.300 ;
        RECT 70.330 123.270 70.660 124.880 ;
        RECT 69.160 122.850 70.160 123.020 ;
        RECT 70.330 120.990 70.660 122.600 ;
        RECT 69.160 120.570 70.160 120.740 ;
        RECT 68.660 118.385 68.990 120.355 ;
        RECT 69.160 119.290 70.160 119.460 ;
        RECT 70.330 118.385 70.660 120.355 ;
        RECT 69.160 118.010 70.160 118.180 ;
        RECT 70.960 117.510 71.130 138.040 ;
        RECT 68.190 117.340 71.130 117.510 ;
        RECT 56.180 111.750 62.710 111.920 ;
        RECT 63.685 113.090 67.285 113.260 ;
        RECT 67.670 113.090 70.245 113.260 ;
        RECT 63.685 89.120 63.855 113.090 ;
        RECT 64.315 112.420 65.315 112.590 ;
        RECT 69.115 112.420 69.615 112.590 ;
        RECT 65.485 110.560 65.815 112.170 ;
        RECT 68.615 110.560 68.945 112.170 ;
        RECT 64.315 110.140 65.315 110.310 ;
        RECT 69.115 110.140 69.615 110.310 ;
        RECT 65.485 108.280 65.815 109.890 ;
        RECT 68.615 108.280 68.945 109.890 ;
        RECT 64.315 107.860 65.315 108.030 ;
        RECT 69.115 107.860 69.615 108.030 ;
        RECT 65.485 106.000 65.815 107.610 ;
        RECT 68.615 106.000 68.945 107.610 ;
        RECT 64.315 105.580 65.315 105.750 ;
        RECT 69.115 105.580 69.615 105.750 ;
        RECT 65.485 103.720 65.815 105.330 ;
        RECT 68.615 103.720 68.945 105.330 ;
        RECT 64.315 103.300 65.315 103.470 ;
        RECT 69.115 103.300 69.615 103.470 ;
        RECT 65.485 101.440 65.815 103.050 ;
        RECT 68.615 101.440 68.945 103.050 ;
        RECT 64.315 101.020 65.315 101.190 ;
        RECT 69.115 101.020 69.615 101.190 ;
        RECT 65.485 99.160 65.815 100.770 ;
        RECT 68.615 99.160 68.945 100.770 ;
        RECT 64.315 98.740 65.315 98.910 ;
        RECT 69.115 98.740 69.615 98.910 ;
        RECT 65.485 96.880 65.815 98.490 ;
        RECT 68.615 96.880 68.945 98.490 ;
        RECT 64.315 96.460 65.315 96.630 ;
        RECT 69.115 96.460 69.615 96.630 ;
        RECT 65.485 94.600 65.815 96.210 ;
        RECT 68.615 94.600 68.945 96.210 ;
        RECT 64.315 94.180 65.315 94.350 ;
        RECT 69.115 94.180 69.615 94.350 ;
        RECT 65.485 92.320 65.815 93.930 ;
        RECT 68.615 92.320 68.945 93.930 ;
        RECT 64.315 91.900 65.315 92.070 ;
        RECT 69.115 91.900 69.615 92.070 ;
        RECT 65.485 90.040 65.815 91.650 ;
        RECT 68.615 90.040 68.945 91.650 ;
        RECT 64.315 89.620 65.315 89.790 ;
        RECT 69.115 89.620 69.615 89.790 ;
        RECT 70.075 89.120 70.245 113.090 ;
        RECT 72.590 112.960 72.760 142.530 ;
        RECT 73.560 141.900 74.060 142.070 ;
        RECT 73.560 140.620 74.060 140.790 ;
        RECT 74.230 139.715 74.560 141.685 ;
        RECT 76.300 141.500 76.800 141.670 ;
        RECT 73.560 139.340 74.060 139.510 ;
        RECT 73.060 137.480 73.390 139.090 ;
        RECT 74.230 137.480 74.560 139.090 ;
        RECT 75.800 138.595 76.130 141.285 ;
        RECT 76.970 138.595 77.300 141.285 ;
        RECT 76.300 138.220 76.800 138.390 ;
        RECT 73.560 137.060 74.060 137.230 ;
        RECT 73.060 135.200 73.390 136.810 ;
        RECT 74.230 135.200 74.560 136.810 ;
        RECT 75.800 135.315 76.130 138.005 ;
        RECT 76.970 135.315 77.300 138.005 ;
        RECT 73.560 134.780 74.060 134.950 ;
        RECT 76.300 134.940 76.800 135.110 ;
        RECT 73.060 132.920 73.390 134.530 ;
        RECT 74.230 132.920 74.560 134.530 ;
        RECT 73.560 132.500 74.060 132.670 ;
        RECT 73.060 130.640 73.390 132.250 ;
        RECT 74.230 130.640 74.560 132.250 ;
        RECT 73.560 130.220 74.060 130.390 ;
        RECT 73.060 128.035 73.390 130.005 ;
        RECT 73.560 128.940 74.060 129.110 ;
        RECT 74.230 128.035 74.560 130.005 ;
        RECT 76.970 128.060 77.300 134.710 ;
        RECT 73.560 127.660 74.060 127.830 ;
        RECT 76.300 127.660 76.800 127.830 ;
        RECT 73.060 125.475 73.390 127.445 ;
        RECT 73.560 126.380 74.060 126.550 ;
        RECT 74.230 125.475 74.560 127.445 ;
        RECT 73.560 125.100 74.060 125.270 ;
        RECT 73.060 123.240 73.390 124.850 ;
        RECT 74.230 123.240 74.560 124.850 ;
        RECT 73.560 122.820 74.060 122.990 ;
        RECT 73.060 120.960 73.390 122.570 ;
        RECT 74.230 120.960 74.560 122.570 ;
        RECT 76.970 120.780 77.300 127.430 ;
        RECT 73.560 120.540 74.060 120.710 ;
        RECT 76.300 120.380 76.800 120.550 ;
        RECT 73.060 118.680 73.390 120.290 ;
        RECT 74.230 118.680 74.560 120.290 ;
        RECT 73.560 118.260 74.060 118.430 ;
        RECT 73.060 116.400 73.390 118.010 ;
        RECT 74.230 116.400 74.560 118.010 ;
        RECT 75.800 117.475 76.130 120.165 ;
        RECT 76.970 117.475 77.300 120.165 ;
        RECT 76.300 117.100 76.800 117.270 ;
        RECT 73.560 115.980 74.060 116.150 ;
        RECT 73.560 114.700 74.060 114.870 ;
        RECT 74.230 113.795 74.560 115.765 ;
        RECT 75.800 114.195 76.130 116.885 ;
        RECT 76.970 114.195 77.300 116.885 ;
        RECT 76.300 113.820 76.800 113.990 ;
        RECT 73.560 113.420 74.060 113.590 ;
        RECT 77.600 112.960 77.770 142.530 ;
        RECT 72.590 112.790 77.770 112.960 ;
        RECT 81.020 142.530 86.200 142.700 ;
        RECT 81.020 112.960 81.190 142.530 ;
        RECT 84.730 141.900 85.230 142.070 ;
        RECT 81.990 141.500 82.490 141.670 ;
        RECT 81.490 138.595 81.820 141.285 ;
        RECT 82.660 138.595 82.990 141.285 ;
        RECT 84.230 139.715 84.560 141.685 ;
        RECT 84.730 140.620 85.230 140.790 ;
        RECT 84.730 139.340 85.230 139.510 ;
        RECT 81.990 138.220 82.490 138.390 ;
        RECT 81.490 135.315 81.820 138.005 ;
        RECT 82.660 135.315 82.990 138.005 ;
        RECT 84.230 137.480 84.560 139.090 ;
        RECT 85.400 137.480 85.730 139.090 ;
        RECT 84.730 137.060 85.230 137.230 ;
        RECT 84.230 135.200 84.560 136.810 ;
        RECT 85.400 135.200 85.730 136.810 ;
        RECT 81.990 134.940 82.490 135.110 ;
        RECT 84.730 134.780 85.230 134.950 ;
        RECT 81.490 128.060 81.820 134.710 ;
        RECT 84.230 132.920 84.560 134.530 ;
        RECT 85.400 132.920 85.730 134.530 ;
        RECT 84.730 132.500 85.230 132.670 ;
        RECT 84.230 130.640 84.560 132.250 ;
        RECT 85.400 130.640 85.730 132.250 ;
        RECT 84.730 130.220 85.230 130.390 ;
        RECT 84.230 128.035 84.560 130.005 ;
        RECT 84.730 128.940 85.230 129.110 ;
        RECT 85.400 128.035 85.730 130.005 ;
        RECT 81.990 127.660 82.490 127.830 ;
        RECT 84.730 127.660 85.230 127.830 ;
        RECT 81.490 120.780 81.820 127.430 ;
        RECT 84.230 125.475 84.560 127.445 ;
        RECT 84.730 126.380 85.230 126.550 ;
        RECT 85.400 125.475 85.730 127.445 ;
        RECT 84.730 125.100 85.230 125.270 ;
        RECT 84.230 123.240 84.560 124.850 ;
        RECT 85.400 123.240 85.730 124.850 ;
        RECT 84.730 122.820 85.230 122.990 ;
        RECT 84.230 120.960 84.560 122.570 ;
        RECT 85.400 120.960 85.730 122.570 ;
        RECT 81.990 120.380 82.490 120.550 ;
        RECT 84.730 120.540 85.230 120.710 ;
        RECT 81.490 117.475 81.820 120.165 ;
        RECT 82.660 117.475 82.990 120.165 ;
        RECT 84.230 118.680 84.560 120.290 ;
        RECT 85.400 118.680 85.730 120.290 ;
        RECT 84.730 118.260 85.230 118.430 ;
        RECT 81.990 117.100 82.490 117.270 ;
        RECT 81.490 114.195 81.820 116.885 ;
        RECT 82.660 114.195 82.990 116.885 ;
        RECT 84.230 116.400 84.560 118.010 ;
        RECT 85.400 116.400 85.730 118.010 ;
        RECT 84.730 115.980 85.230 116.150 ;
        RECT 81.990 113.820 82.490 113.990 ;
        RECT 84.230 113.795 84.560 115.765 ;
        RECT 84.730 114.700 85.230 114.870 ;
        RECT 84.730 113.420 85.230 113.590 ;
        RECT 86.030 112.960 86.200 142.530 ;
        RECT 91.915 142.400 92.085 151.250 ;
        RECT 92.885 150.580 93.385 150.750 ;
        RECT 92.385 149.440 92.715 150.330 ;
        RECT 92.885 149.800 93.385 149.970 ;
        RECT 92.885 149.020 93.385 149.190 ;
        RECT 93.555 147.160 93.885 148.770 ;
        RECT 92.885 146.740 93.385 146.910 ;
        RECT 93.555 144.880 93.885 146.490 ;
        RECT 92.885 144.460 93.385 144.630 ;
        RECT 92.385 143.320 92.715 144.210 ;
        RECT 92.885 143.680 93.385 143.850 ;
        RECT 92.885 142.900 93.385 143.070 ;
        RECT 94.185 142.400 94.355 151.250 ;
        RECT 91.915 142.230 94.355 142.400 ;
        RECT 96.080 151.250 102.610 151.420 ;
        RECT 87.660 138.040 90.600 138.210 ;
        RECT 87.660 117.510 87.830 138.040 ;
        RECT 88.630 137.370 89.630 137.540 ;
        RECT 88.130 135.185 88.460 137.155 ;
        RECT 88.630 136.090 89.630 136.260 ;
        RECT 89.800 135.185 90.130 137.155 ;
        RECT 88.630 134.810 89.630 134.980 ;
        RECT 88.130 132.950 88.460 134.560 ;
        RECT 89.800 132.950 90.130 134.560 ;
        RECT 88.630 132.530 89.630 132.700 ;
        RECT 88.130 130.670 88.460 132.280 ;
        RECT 89.800 130.670 90.130 132.280 ;
        RECT 88.630 130.250 89.630 130.420 ;
        RECT 88.130 128.065 88.460 130.035 ;
        RECT 88.630 128.970 89.630 129.140 ;
        RECT 89.800 128.065 90.130 130.035 ;
        RECT 88.630 127.690 89.630 127.860 ;
        RECT 88.130 125.505 88.460 127.475 ;
        RECT 88.630 126.410 89.630 126.580 ;
        RECT 89.800 125.505 90.130 127.475 ;
        RECT 88.630 125.130 89.630 125.300 ;
        RECT 88.130 123.270 88.460 124.880 ;
        RECT 88.630 122.850 89.630 123.020 ;
        RECT 88.130 120.990 88.460 122.600 ;
        RECT 88.630 120.570 89.630 120.740 ;
        RECT 88.130 118.385 88.460 120.355 ;
        RECT 88.630 119.290 89.630 119.460 ;
        RECT 89.800 118.385 90.130 120.355 ;
        RECT 88.630 118.010 89.630 118.180 ;
        RECT 90.430 117.510 90.600 138.040 ;
        RECT 87.660 117.340 90.600 117.510 ;
        RECT 91.915 138.040 94.355 138.210 ;
        RECT 91.915 117.510 92.085 138.040 ;
        RECT 92.885 137.370 93.385 137.540 ;
        RECT 92.385 135.185 92.715 137.155 ;
        RECT 92.885 136.090 93.385 136.260 ;
        RECT 93.555 135.185 93.885 137.155 ;
        RECT 92.885 134.810 93.385 134.980 ;
        RECT 92.385 132.950 92.715 134.560 ;
        RECT 93.555 132.950 93.885 134.560 ;
        RECT 92.885 132.530 93.385 132.700 ;
        RECT 92.385 130.670 92.715 132.280 ;
        RECT 93.555 130.670 93.885 132.280 ;
        RECT 92.885 130.250 93.385 130.420 ;
        RECT 92.385 128.065 92.715 130.035 ;
        RECT 92.885 128.970 93.385 129.140 ;
        RECT 93.555 128.065 93.885 130.035 ;
        RECT 92.885 127.690 93.385 127.860 ;
        RECT 92.385 125.505 92.715 127.475 ;
        RECT 92.885 126.410 93.385 126.580 ;
        RECT 93.555 125.505 93.885 127.475 ;
        RECT 92.885 125.130 93.385 125.300 ;
        RECT 93.555 123.270 93.885 124.880 ;
        RECT 92.885 122.850 93.385 123.020 ;
        RECT 93.555 120.990 93.885 122.600 ;
        RECT 92.885 120.570 93.385 120.740 ;
        RECT 92.385 118.385 92.715 120.355 ;
        RECT 92.885 119.290 93.385 119.460 ;
        RECT 93.555 118.385 93.885 120.355 ;
        RECT 92.885 118.010 93.385 118.180 ;
        RECT 94.185 117.510 94.355 138.040 ;
        RECT 91.915 117.340 94.355 117.510 ;
        RECT 81.020 112.790 86.200 112.960 ;
        RECT 88.545 113.090 91.120 113.260 ;
        RECT 91.505 113.090 95.105 113.260 ;
        RECT 63.685 88.950 67.285 89.120 ;
        RECT 67.670 88.950 70.245 89.120 ;
        RECT 88.545 89.120 88.715 113.090 ;
        RECT 89.175 112.420 89.675 112.590 ;
        RECT 93.475 112.420 94.475 112.590 ;
        RECT 89.845 110.560 90.175 112.170 ;
        RECT 92.975 110.560 93.305 112.170 ;
        RECT 89.175 110.140 89.675 110.310 ;
        RECT 93.475 110.140 94.475 110.310 ;
        RECT 89.845 108.280 90.175 109.890 ;
        RECT 92.975 108.280 93.305 109.890 ;
        RECT 89.175 107.860 89.675 108.030 ;
        RECT 93.475 107.860 94.475 108.030 ;
        RECT 89.845 106.000 90.175 107.610 ;
        RECT 92.975 106.000 93.305 107.610 ;
        RECT 89.175 105.580 89.675 105.750 ;
        RECT 93.475 105.580 94.475 105.750 ;
        RECT 89.845 103.720 90.175 105.330 ;
        RECT 92.975 103.720 93.305 105.330 ;
        RECT 89.175 103.300 89.675 103.470 ;
        RECT 93.475 103.300 94.475 103.470 ;
        RECT 89.845 101.440 90.175 103.050 ;
        RECT 92.975 101.440 93.305 103.050 ;
        RECT 89.175 101.020 89.675 101.190 ;
        RECT 93.475 101.020 94.475 101.190 ;
        RECT 89.845 99.160 90.175 100.770 ;
        RECT 92.975 99.160 93.305 100.770 ;
        RECT 89.175 98.740 89.675 98.910 ;
        RECT 93.475 98.740 94.475 98.910 ;
        RECT 89.845 96.880 90.175 98.490 ;
        RECT 92.975 96.880 93.305 98.490 ;
        RECT 89.175 96.460 89.675 96.630 ;
        RECT 93.475 96.460 94.475 96.630 ;
        RECT 89.845 94.600 90.175 96.210 ;
        RECT 92.975 94.600 93.305 96.210 ;
        RECT 89.175 94.180 89.675 94.350 ;
        RECT 93.475 94.180 94.475 94.350 ;
        RECT 89.845 92.320 90.175 93.930 ;
        RECT 92.975 92.320 93.305 93.930 ;
        RECT 89.175 91.900 89.675 92.070 ;
        RECT 93.475 91.900 94.475 92.070 ;
        RECT 89.845 90.040 90.175 91.650 ;
        RECT 92.975 90.040 93.305 91.650 ;
        RECT 89.175 89.620 89.675 89.790 ;
        RECT 93.475 89.620 94.475 89.790 ;
        RECT 94.935 89.120 95.105 113.090 ;
        RECT 96.080 111.920 96.250 151.250 ;
        RECT 97.050 150.580 98.050 150.750 ;
        RECT 97.050 149.800 98.050 149.970 ;
        RECT 98.220 149.440 98.550 150.330 ;
        RECT 97.050 149.020 98.050 149.190 ;
        RECT 96.550 147.160 96.880 148.770 ;
        RECT 97.050 146.740 98.050 146.910 ;
        RECT 96.550 144.880 96.880 146.490 ;
        RECT 97.050 144.460 98.050 144.630 ;
        RECT 97.050 143.680 98.050 143.850 ;
        RECT 98.220 143.320 98.550 144.210 ;
        RECT 97.050 142.900 98.050 143.070 ;
        RECT 97.050 142.120 98.050 142.290 ;
        RECT 98.220 141.760 98.550 142.650 ;
        RECT 97.050 141.340 98.050 141.510 ;
        RECT 100.640 141.340 101.640 141.510 ;
        RECT 96.550 139.480 96.880 141.090 ;
        RECT 98.220 139.480 98.550 141.090 ;
        RECT 100.140 139.480 100.470 141.090 ;
        RECT 97.050 139.060 98.050 139.230 ;
        RECT 100.640 139.060 101.640 139.230 ;
        RECT 96.550 137.200 96.880 138.810 ;
        RECT 98.220 137.200 98.550 138.810 ;
        RECT 100.140 137.200 100.470 138.810 ;
        RECT 97.050 136.780 98.050 136.950 ;
        RECT 100.640 136.780 101.640 136.950 ;
        RECT 96.550 134.920 96.880 136.530 ;
        RECT 98.220 134.920 98.550 136.530 ;
        RECT 100.140 134.920 100.470 136.530 ;
        RECT 97.050 134.500 98.050 134.670 ;
        RECT 100.640 134.500 101.640 134.670 ;
        RECT 96.550 132.640 96.880 134.250 ;
        RECT 98.220 132.640 98.550 134.250 ;
        RECT 100.140 132.640 100.470 134.250 ;
        RECT 97.050 132.220 98.050 132.390 ;
        RECT 100.640 132.220 101.640 132.390 ;
        RECT 96.550 130.360 96.880 131.970 ;
        RECT 98.220 130.360 98.550 131.970 ;
        RECT 100.140 130.360 100.470 131.970 ;
        RECT 97.050 129.940 98.050 130.110 ;
        RECT 100.640 129.940 101.640 130.110 ;
        RECT 96.550 128.080 96.880 129.690 ;
        RECT 98.220 128.080 98.550 129.690 ;
        RECT 101.810 128.080 102.140 129.690 ;
        RECT 97.050 127.660 98.050 127.830 ;
        RECT 100.640 127.660 101.640 127.830 ;
        RECT 96.550 125.800 96.880 127.410 ;
        RECT 98.220 125.800 98.550 127.410 ;
        RECT 101.810 125.800 102.140 127.410 ;
        RECT 97.050 125.380 98.050 125.550 ;
        RECT 100.640 125.380 101.640 125.550 ;
        RECT 96.550 123.520 96.880 125.130 ;
        RECT 98.220 123.520 98.550 125.130 ;
        RECT 100.140 123.520 100.470 125.130 ;
        RECT 97.050 123.100 98.050 123.270 ;
        RECT 100.640 123.100 101.640 123.270 ;
        RECT 96.550 121.240 96.880 122.850 ;
        RECT 98.220 121.240 98.550 122.850 ;
        RECT 100.140 121.240 100.470 122.850 ;
        RECT 97.050 120.820 98.050 120.990 ;
        RECT 100.640 120.820 101.640 120.990 ;
        RECT 96.550 118.960 96.880 120.570 ;
        RECT 98.220 118.960 98.550 120.570 ;
        RECT 100.140 118.960 100.470 120.570 ;
        RECT 97.050 118.540 98.050 118.710 ;
        RECT 100.640 118.540 101.640 118.710 ;
        RECT 96.550 116.680 96.880 118.290 ;
        RECT 98.220 116.680 98.550 118.290 ;
        RECT 100.140 116.680 100.470 118.290 ;
        RECT 97.050 116.260 98.050 116.430 ;
        RECT 100.640 116.260 101.640 116.430 ;
        RECT 96.550 114.400 96.880 116.010 ;
        RECT 98.220 114.400 98.550 116.010 ;
        RECT 100.140 114.400 100.470 116.010 ;
        RECT 97.050 113.980 98.050 114.150 ;
        RECT 100.640 113.980 101.640 114.150 ;
        RECT 97.050 113.200 98.050 113.370 ;
        RECT 98.220 112.840 98.550 113.730 ;
        RECT 97.050 112.420 98.050 112.590 ;
        RECT 102.440 111.920 102.610 151.250 ;
        RECT 96.080 111.750 102.610 111.920 ;
        RECT 88.545 88.950 91.120 89.120 ;
        RECT 91.505 88.950 95.105 89.120 ;
        RECT 88.505 82.770 91.080 82.940 ;
        RECT 91.490 82.770 95.090 82.940 ;
        RECT 71.475 82.420 74.330 82.590 ;
        RECT 74.860 82.420 83.700 82.590 ;
        RECT 84.230 82.420 87.085 82.590 ;
        RECT 71.475 77.810 71.645 82.420 ;
        RECT 72.445 81.750 73.445 81.920 ;
        RECT 75.745 81.750 76.745 81.920 ;
        RECT 77.395 81.750 78.395 81.920 ;
        RECT 71.945 81.140 72.275 81.670 ;
        RECT 72.445 81.320 73.445 81.490 ;
        RECT 73.615 81.140 73.945 81.670 ;
        RECT 75.245 81.140 75.575 81.670 ;
        RECT 75.745 81.320 76.745 81.490 ;
        RECT 77.395 81.320 78.395 81.490 ;
        RECT 78.565 81.140 78.895 81.670 ;
        RECT 72.445 80.890 73.445 81.060 ;
        RECT 75.745 80.890 76.745 81.060 ;
        RECT 77.395 80.890 78.395 81.060 ;
        RECT 71.945 80.280 72.275 80.810 ;
        RECT 72.445 80.460 73.445 80.630 ;
        RECT 73.615 80.280 73.945 80.810 ;
        RECT 75.245 80.280 75.575 80.810 ;
        RECT 75.745 80.460 76.745 80.630 ;
        RECT 77.395 80.460 78.395 80.630 ;
        RECT 78.565 80.280 78.895 80.810 ;
        RECT 72.445 80.030 73.445 80.200 ;
        RECT 75.745 80.030 76.745 80.200 ;
        RECT 77.395 80.030 78.395 80.200 ;
        RECT 71.945 79.420 72.275 79.950 ;
        RECT 72.445 79.600 73.445 79.770 ;
        RECT 73.615 79.420 73.945 79.950 ;
        RECT 75.245 79.420 75.575 79.950 ;
        RECT 75.745 79.600 76.745 79.770 ;
        RECT 77.395 79.600 78.395 79.770 ;
        RECT 78.565 79.420 78.895 79.950 ;
        RECT 72.445 79.170 73.445 79.340 ;
        RECT 75.745 79.170 76.745 79.340 ;
        RECT 77.395 79.170 78.395 79.340 ;
        RECT 71.945 78.560 72.275 79.090 ;
        RECT 72.445 78.740 73.445 78.910 ;
        RECT 73.615 78.560 73.945 79.090 ;
        RECT 75.245 78.560 75.575 79.090 ;
        RECT 75.745 78.740 76.745 78.910 ;
        RECT 77.395 78.740 78.395 78.910 ;
        RECT 78.565 78.560 78.895 79.090 ;
        RECT 72.445 78.310 73.445 78.480 ;
        RECT 75.745 78.310 76.745 78.480 ;
        RECT 77.395 78.310 78.395 78.480 ;
        RECT 79.195 77.810 79.365 82.420 ;
        RECT 80.165 81.750 81.165 81.920 ;
        RECT 81.815 81.750 82.815 81.920 ;
        RECT 85.115 81.750 86.115 81.920 ;
        RECT 79.665 81.140 79.995 81.670 ;
        RECT 80.165 81.320 81.165 81.490 ;
        RECT 81.815 81.320 82.815 81.490 ;
        RECT 82.985 81.140 83.315 81.670 ;
        RECT 84.615 81.140 84.945 81.670 ;
        RECT 85.115 81.320 86.115 81.490 ;
        RECT 86.285 81.140 86.615 81.670 ;
        RECT 80.165 80.890 81.165 81.060 ;
        RECT 81.815 80.890 82.815 81.060 ;
        RECT 85.115 80.890 86.115 81.060 ;
        RECT 79.665 80.280 79.995 80.810 ;
        RECT 80.165 80.460 81.165 80.630 ;
        RECT 81.815 80.460 82.815 80.630 ;
        RECT 82.985 80.280 83.315 80.810 ;
        RECT 84.615 80.280 84.945 80.810 ;
        RECT 85.115 80.460 86.115 80.630 ;
        RECT 86.285 80.280 86.615 80.810 ;
        RECT 80.165 80.030 81.165 80.200 ;
        RECT 81.815 80.030 82.815 80.200 ;
        RECT 85.115 80.030 86.115 80.200 ;
        RECT 79.665 79.420 79.995 79.950 ;
        RECT 80.165 79.600 81.165 79.770 ;
        RECT 81.815 79.600 82.815 79.770 ;
        RECT 82.985 79.420 83.315 79.950 ;
        RECT 84.615 79.420 84.945 79.950 ;
        RECT 85.115 79.600 86.115 79.770 ;
        RECT 86.285 79.420 86.615 79.950 ;
        RECT 80.165 79.170 81.165 79.340 ;
        RECT 81.815 79.170 82.815 79.340 ;
        RECT 85.115 79.170 86.115 79.340 ;
        RECT 79.665 78.560 79.995 79.090 ;
        RECT 80.165 78.740 81.165 78.910 ;
        RECT 81.815 78.740 82.815 78.910 ;
        RECT 82.985 78.560 83.315 79.090 ;
        RECT 84.615 78.560 84.945 79.090 ;
        RECT 85.115 78.740 86.115 78.910 ;
        RECT 86.285 78.560 86.615 79.090 ;
        RECT 80.165 78.310 81.165 78.480 ;
        RECT 81.815 78.310 82.815 78.480 ;
        RECT 85.115 78.310 86.115 78.480 ;
        RECT 86.915 77.810 87.085 82.420 ;
        RECT 88.505 78.160 88.675 82.770 ;
        RECT 89.110 82.100 90.110 82.270 ;
        RECT 92.460 82.100 94.460 82.270 ;
        RECT 89.110 81.670 90.110 81.840 ;
        RECT 90.280 81.490 90.610 82.020 ;
        RECT 91.960 81.490 92.290 82.020 ;
        RECT 92.460 81.670 94.460 81.840 ;
        RECT 89.110 81.240 90.110 81.410 ;
        RECT 92.460 81.240 94.460 81.410 ;
        RECT 89.110 80.810 90.110 80.980 ;
        RECT 90.280 80.630 90.610 81.160 ;
        RECT 91.960 80.630 92.290 81.160 ;
        RECT 92.460 80.810 94.460 80.980 ;
        RECT 89.110 80.380 90.110 80.550 ;
        RECT 92.460 80.380 94.460 80.550 ;
        RECT 89.110 79.950 90.110 80.120 ;
        RECT 90.280 79.770 90.610 80.300 ;
        RECT 91.960 79.770 92.290 80.300 ;
        RECT 92.460 79.950 94.460 80.120 ;
        RECT 89.110 79.520 90.110 79.690 ;
        RECT 92.460 79.520 94.460 79.690 ;
        RECT 89.110 79.090 90.110 79.260 ;
        RECT 90.280 78.910 90.610 79.440 ;
        RECT 91.960 78.910 92.290 79.440 ;
        RECT 92.460 79.090 94.460 79.260 ;
        RECT 89.110 78.660 90.110 78.830 ;
        RECT 92.460 78.660 94.460 78.830 ;
        RECT 94.920 78.160 95.090 82.770 ;
        RECT 88.505 77.990 91.080 78.160 ;
        RECT 91.490 77.990 95.090 78.160 ;
        RECT 71.475 77.640 74.330 77.810 ;
        RECT 74.860 77.640 83.700 77.810 ;
        RECT 84.230 77.640 87.085 77.810 ;
        RECT 64.725 72.110 67.300 72.280 ;
        RECT 67.710 72.110 71.310 72.280 ;
        RECT 64.725 63.200 64.895 72.110 ;
        RECT 65.330 71.440 66.330 71.610 ;
        RECT 68.680 71.440 70.680 71.610 ;
        RECT 65.330 71.010 66.330 71.180 ;
        RECT 66.500 70.830 66.830 71.360 ;
        RECT 68.180 70.830 68.510 71.360 ;
        RECT 68.680 71.010 70.680 71.180 ;
        RECT 65.330 70.580 66.330 70.750 ;
        RECT 68.680 70.580 70.680 70.750 ;
        RECT 65.330 70.150 66.330 70.320 ;
        RECT 66.500 69.970 66.830 70.500 ;
        RECT 68.180 69.970 68.510 70.500 ;
        RECT 68.680 70.150 70.680 70.320 ;
        RECT 65.330 69.720 66.330 69.890 ;
        RECT 68.680 69.720 70.680 69.890 ;
        RECT 65.330 69.290 66.330 69.460 ;
        RECT 66.500 69.110 66.830 69.640 ;
        RECT 68.180 69.110 68.510 69.640 ;
        RECT 68.680 69.290 70.680 69.460 ;
        RECT 65.330 68.860 66.330 69.030 ;
        RECT 68.680 68.860 70.680 69.030 ;
        RECT 65.330 68.430 66.330 68.600 ;
        RECT 66.500 68.250 66.830 68.780 ;
        RECT 68.180 68.250 68.510 68.780 ;
        RECT 68.680 68.430 70.680 68.600 ;
        RECT 65.330 68.000 66.330 68.170 ;
        RECT 68.680 68.000 70.680 68.170 ;
        RECT 65.330 67.570 66.330 67.740 ;
        RECT 66.500 67.390 66.830 67.920 ;
        RECT 68.180 67.390 68.510 67.920 ;
        RECT 68.680 67.570 70.680 67.740 ;
        RECT 65.330 67.140 66.330 67.310 ;
        RECT 68.680 67.140 70.680 67.310 ;
        RECT 65.330 66.710 66.330 66.880 ;
        RECT 66.500 66.530 66.830 67.060 ;
        RECT 68.180 66.530 68.510 67.060 ;
        RECT 68.680 66.710 70.680 66.880 ;
        RECT 65.330 66.280 66.330 66.450 ;
        RECT 68.680 66.280 70.680 66.450 ;
        RECT 65.330 65.850 66.330 66.020 ;
        RECT 66.500 65.670 66.830 66.200 ;
        RECT 68.180 65.670 68.510 66.200 ;
        RECT 68.680 65.850 70.680 66.020 ;
        RECT 65.330 65.420 66.330 65.590 ;
        RECT 68.680 65.420 70.680 65.590 ;
        RECT 65.330 64.990 66.330 65.160 ;
        RECT 66.500 64.810 66.830 65.340 ;
        RECT 68.180 64.810 68.510 65.340 ;
        RECT 68.680 64.990 70.680 65.160 ;
        RECT 65.330 64.560 66.330 64.730 ;
        RECT 68.680 64.560 70.680 64.730 ;
        RECT 65.330 64.130 66.330 64.300 ;
        RECT 66.500 63.950 66.830 64.480 ;
        RECT 68.180 63.950 68.510 64.480 ;
        RECT 68.680 64.130 70.680 64.300 ;
        RECT 65.330 63.700 66.330 63.870 ;
        RECT 68.680 63.700 70.680 63.870 ;
        RECT 71.140 63.200 71.310 72.110 ;
        RECT 64.725 63.030 67.300 63.200 ;
        RECT 67.710 63.030 71.310 63.200 ;
        RECT 73.745 72.110 76.320 72.280 ;
        RECT 76.730 72.110 83.760 72.280 ;
        RECT 84.170 72.110 86.745 72.280 ;
        RECT 73.745 63.200 73.915 72.110 ;
        RECT 74.350 71.440 75.350 71.610 ;
        RECT 77.700 71.440 79.700 71.610 ;
        RECT 74.350 71.010 75.350 71.180 ;
        RECT 75.520 70.830 75.850 71.360 ;
        RECT 77.200 70.830 77.530 71.360 ;
        RECT 77.700 71.010 79.700 71.180 ;
        RECT 74.350 70.580 75.350 70.750 ;
        RECT 77.700 70.580 79.700 70.750 ;
        RECT 74.350 70.150 75.350 70.320 ;
        RECT 75.520 69.970 75.850 70.500 ;
        RECT 77.200 69.970 77.530 70.500 ;
        RECT 77.700 70.150 79.700 70.320 ;
        RECT 74.350 69.720 75.350 69.890 ;
        RECT 77.700 69.720 79.700 69.890 ;
        RECT 74.350 69.290 75.350 69.460 ;
        RECT 75.520 69.110 75.850 69.640 ;
        RECT 77.200 69.110 77.530 69.640 ;
        RECT 77.700 69.290 79.700 69.460 ;
        RECT 74.350 68.860 75.350 69.030 ;
        RECT 77.700 68.860 79.700 69.030 ;
        RECT 74.350 68.430 75.350 68.600 ;
        RECT 75.520 68.250 75.850 68.780 ;
        RECT 77.200 68.250 77.530 68.780 ;
        RECT 77.700 68.430 79.700 68.600 ;
        RECT 74.350 68.000 75.350 68.170 ;
        RECT 77.700 68.000 79.700 68.170 ;
        RECT 74.350 67.570 75.350 67.740 ;
        RECT 75.520 67.390 75.850 67.920 ;
        RECT 77.200 67.390 77.530 67.920 ;
        RECT 77.700 67.570 79.700 67.740 ;
        RECT 74.350 67.140 75.350 67.310 ;
        RECT 77.700 67.140 79.700 67.310 ;
        RECT 74.350 66.710 75.350 66.880 ;
        RECT 75.520 66.530 75.850 67.060 ;
        RECT 77.200 66.530 77.530 67.060 ;
        RECT 77.700 66.710 79.700 66.880 ;
        RECT 74.350 66.280 75.350 66.450 ;
        RECT 77.700 66.280 79.700 66.450 ;
        RECT 74.350 65.850 75.350 66.020 ;
        RECT 75.520 65.670 75.850 66.200 ;
        RECT 77.200 65.670 77.530 66.200 ;
        RECT 77.700 65.850 79.700 66.020 ;
        RECT 74.350 65.420 75.350 65.590 ;
        RECT 77.700 65.420 79.700 65.590 ;
        RECT 74.350 64.990 75.350 65.160 ;
        RECT 75.520 64.810 75.850 65.340 ;
        RECT 77.200 64.810 77.530 65.340 ;
        RECT 77.700 64.990 79.700 65.160 ;
        RECT 74.350 64.560 75.350 64.730 ;
        RECT 77.700 64.560 79.700 64.730 ;
        RECT 74.350 64.130 75.350 64.300 ;
        RECT 75.520 63.950 75.850 64.480 ;
        RECT 77.200 63.950 77.530 64.480 ;
        RECT 77.700 64.130 79.700 64.300 ;
        RECT 74.350 63.700 75.350 63.870 ;
        RECT 77.700 63.700 79.700 63.870 ;
        RECT 80.160 63.200 80.330 72.110 ;
        RECT 80.790 71.440 82.790 71.610 ;
        RECT 85.140 71.440 86.140 71.610 ;
        RECT 80.790 71.010 82.790 71.180 ;
        RECT 82.960 70.830 83.290 71.360 ;
        RECT 84.640 70.830 84.970 71.360 ;
        RECT 85.140 71.010 86.140 71.180 ;
        RECT 80.790 70.580 82.790 70.750 ;
        RECT 85.140 70.580 86.140 70.750 ;
        RECT 80.790 70.150 82.790 70.320 ;
        RECT 82.960 69.970 83.290 70.500 ;
        RECT 84.640 69.970 84.970 70.500 ;
        RECT 85.140 70.150 86.140 70.320 ;
        RECT 80.790 69.720 82.790 69.890 ;
        RECT 85.140 69.720 86.140 69.890 ;
        RECT 80.790 69.290 82.790 69.460 ;
        RECT 82.960 69.110 83.290 69.640 ;
        RECT 84.640 69.110 84.970 69.640 ;
        RECT 85.140 69.290 86.140 69.460 ;
        RECT 80.790 68.860 82.790 69.030 ;
        RECT 85.140 68.860 86.140 69.030 ;
        RECT 80.790 68.430 82.790 68.600 ;
        RECT 82.960 68.250 83.290 68.780 ;
        RECT 84.640 68.250 84.970 68.780 ;
        RECT 85.140 68.430 86.140 68.600 ;
        RECT 80.790 68.000 82.790 68.170 ;
        RECT 85.140 68.000 86.140 68.170 ;
        RECT 80.790 67.570 82.790 67.740 ;
        RECT 82.960 67.390 83.290 67.920 ;
        RECT 84.640 67.390 84.970 67.920 ;
        RECT 85.140 67.570 86.140 67.740 ;
        RECT 80.790 67.140 82.790 67.310 ;
        RECT 85.140 67.140 86.140 67.310 ;
        RECT 80.790 66.710 82.790 66.880 ;
        RECT 82.960 66.530 83.290 67.060 ;
        RECT 84.640 66.530 84.970 67.060 ;
        RECT 85.140 66.710 86.140 66.880 ;
        RECT 80.790 66.280 82.790 66.450 ;
        RECT 85.140 66.280 86.140 66.450 ;
        RECT 80.790 65.850 82.790 66.020 ;
        RECT 82.960 65.670 83.290 66.200 ;
        RECT 84.640 65.670 84.970 66.200 ;
        RECT 85.140 65.850 86.140 66.020 ;
        RECT 80.790 65.420 82.790 65.590 ;
        RECT 85.140 65.420 86.140 65.590 ;
        RECT 80.790 64.990 82.790 65.160 ;
        RECT 82.960 64.810 83.290 65.340 ;
        RECT 84.640 64.810 84.970 65.340 ;
        RECT 85.140 64.990 86.140 65.160 ;
        RECT 80.790 64.560 82.790 64.730 ;
        RECT 85.140 64.560 86.140 64.730 ;
        RECT 80.790 64.130 82.790 64.300 ;
        RECT 82.960 63.950 83.290 64.480 ;
        RECT 84.640 63.950 84.970 64.480 ;
        RECT 85.140 64.130 86.140 64.300 ;
        RECT 80.790 63.700 82.790 63.870 ;
        RECT 85.140 63.700 86.140 63.870 ;
        RECT 86.575 63.200 86.745 72.110 ;
        RECT 73.745 63.030 76.320 63.200 ;
        RECT 76.730 63.030 83.760 63.200 ;
        RECT 84.170 63.030 86.745 63.200 ;
        RECT 88.505 72.110 91.080 72.280 ;
        RECT 91.490 72.110 95.090 72.280 ;
        RECT 88.505 63.200 88.675 72.110 ;
        RECT 89.110 71.440 90.110 71.610 ;
        RECT 92.460 71.440 94.460 71.610 ;
        RECT 89.110 71.010 90.110 71.180 ;
        RECT 90.280 70.830 90.610 71.360 ;
        RECT 91.960 70.830 92.290 71.360 ;
        RECT 92.460 71.010 94.460 71.180 ;
        RECT 89.110 70.580 90.110 70.750 ;
        RECT 92.460 70.580 94.460 70.750 ;
        RECT 89.110 70.150 90.110 70.320 ;
        RECT 90.280 69.970 90.610 70.500 ;
        RECT 91.960 69.970 92.290 70.500 ;
        RECT 92.460 70.150 94.460 70.320 ;
        RECT 89.110 69.720 90.110 69.890 ;
        RECT 92.460 69.720 94.460 69.890 ;
        RECT 89.110 69.290 90.110 69.460 ;
        RECT 90.280 69.110 90.610 69.640 ;
        RECT 91.960 69.110 92.290 69.640 ;
        RECT 92.460 69.290 94.460 69.460 ;
        RECT 89.110 68.860 90.110 69.030 ;
        RECT 92.460 68.860 94.460 69.030 ;
        RECT 89.110 68.430 90.110 68.600 ;
        RECT 90.280 68.250 90.610 68.780 ;
        RECT 91.960 68.250 92.290 68.780 ;
        RECT 92.460 68.430 94.460 68.600 ;
        RECT 89.110 68.000 90.110 68.170 ;
        RECT 92.460 68.000 94.460 68.170 ;
        RECT 89.110 67.570 90.110 67.740 ;
        RECT 90.280 67.390 90.610 67.920 ;
        RECT 91.960 67.390 92.290 67.920 ;
        RECT 92.460 67.570 94.460 67.740 ;
        RECT 89.110 67.140 90.110 67.310 ;
        RECT 92.460 67.140 94.460 67.310 ;
        RECT 89.110 66.710 90.110 66.880 ;
        RECT 90.280 66.530 90.610 67.060 ;
        RECT 91.960 66.530 92.290 67.060 ;
        RECT 92.460 66.710 94.460 66.880 ;
        RECT 89.110 66.280 90.110 66.450 ;
        RECT 92.460 66.280 94.460 66.450 ;
        RECT 89.110 65.850 90.110 66.020 ;
        RECT 90.280 65.670 90.610 66.200 ;
        RECT 91.960 65.670 92.290 66.200 ;
        RECT 92.460 65.850 94.460 66.020 ;
        RECT 89.110 65.420 90.110 65.590 ;
        RECT 92.460 65.420 94.460 65.590 ;
        RECT 89.110 64.990 90.110 65.160 ;
        RECT 90.280 64.810 90.610 65.340 ;
        RECT 91.960 64.810 92.290 65.340 ;
        RECT 92.460 64.990 94.460 65.160 ;
        RECT 89.110 64.560 90.110 64.730 ;
        RECT 92.460 64.560 94.460 64.730 ;
        RECT 89.110 64.130 90.110 64.300 ;
        RECT 90.280 63.950 90.610 64.480 ;
        RECT 91.960 63.950 92.290 64.480 ;
        RECT 92.460 64.130 94.460 64.300 ;
        RECT 89.110 63.700 90.110 63.870 ;
        RECT 92.460 63.700 94.460 63.870 ;
        RECT 94.920 63.200 95.090 72.110 ;
        RECT 88.505 63.030 91.080 63.200 ;
        RECT 91.490 63.030 95.090 63.200 ;
        RECT 108.635 63.010 108.805 164.500 ;
        RECT 109.605 163.830 110.305 164.000 ;
        RECT 110.975 163.830 111.675 164.000 ;
        RECT 112.345 163.830 113.045 164.000 ;
        RECT 110.475 161.970 110.805 163.580 ;
        RECT 111.845 161.970 112.175 163.580 ;
        RECT 109.605 161.550 110.305 161.720 ;
        RECT 110.975 161.550 111.675 161.720 ;
        RECT 112.345 161.550 113.045 161.720 ;
        RECT 110.475 159.690 110.805 161.300 ;
        RECT 111.845 159.690 112.175 161.300 ;
        RECT 109.605 159.270 110.305 159.440 ;
        RECT 110.975 159.270 111.675 159.440 ;
        RECT 112.345 159.270 113.045 159.440 ;
        RECT 110.475 157.410 110.805 159.020 ;
        RECT 111.845 157.410 112.175 159.020 ;
        RECT 109.605 156.990 110.305 157.160 ;
        RECT 110.975 156.990 111.675 157.160 ;
        RECT 112.345 156.990 113.045 157.160 ;
        RECT 110.475 155.130 110.805 156.740 ;
        RECT 111.845 155.130 112.175 156.740 ;
        RECT 109.605 154.710 110.305 154.880 ;
        RECT 110.975 154.710 111.675 154.880 ;
        RECT 112.345 154.710 113.045 154.880 ;
        RECT 110.475 152.850 110.805 154.460 ;
        RECT 111.845 152.850 112.175 154.460 ;
        RECT 109.605 152.430 110.305 152.600 ;
        RECT 110.975 152.430 111.675 152.600 ;
        RECT 112.345 152.430 113.045 152.600 ;
        RECT 110.475 150.570 110.805 152.180 ;
        RECT 111.845 150.570 112.175 152.180 ;
        RECT 109.605 150.150 110.305 150.320 ;
        RECT 110.975 150.150 111.675 150.320 ;
        RECT 112.345 150.150 113.045 150.320 ;
        RECT 110.475 148.290 110.805 149.900 ;
        RECT 111.845 148.290 112.175 149.900 ;
        RECT 109.605 147.870 110.305 148.040 ;
        RECT 110.975 147.870 111.675 148.040 ;
        RECT 112.345 147.870 113.045 148.040 ;
        RECT 110.475 146.010 110.805 147.620 ;
        RECT 111.845 146.010 112.175 147.620 ;
        RECT 109.605 145.590 110.305 145.760 ;
        RECT 110.975 145.590 111.675 145.760 ;
        RECT 112.345 145.590 113.045 145.760 ;
        RECT 110.475 143.730 110.805 145.340 ;
        RECT 111.845 143.730 112.175 145.340 ;
        RECT 109.605 143.310 110.305 143.480 ;
        RECT 110.975 143.310 111.675 143.480 ;
        RECT 112.345 143.310 113.045 143.480 ;
        RECT 110.475 141.450 110.805 143.060 ;
        RECT 111.845 141.450 112.175 143.060 ;
        RECT 109.605 141.030 110.305 141.200 ;
        RECT 110.975 141.030 111.675 141.200 ;
        RECT 112.345 141.030 113.045 141.200 ;
        RECT 110.475 139.170 110.805 140.780 ;
        RECT 111.845 139.170 112.175 140.780 ;
        RECT 109.605 138.750 110.305 138.920 ;
        RECT 110.975 138.750 111.675 138.920 ;
        RECT 112.345 138.750 113.045 138.920 ;
        RECT 110.475 136.890 110.805 138.500 ;
        RECT 111.845 136.890 112.175 138.500 ;
        RECT 109.605 136.470 110.305 136.640 ;
        RECT 110.975 136.470 111.675 136.640 ;
        RECT 112.345 136.470 113.045 136.640 ;
        RECT 110.475 134.610 110.805 136.220 ;
        RECT 111.845 134.610 112.175 136.220 ;
        RECT 109.605 134.190 110.305 134.360 ;
        RECT 110.975 134.190 111.675 134.360 ;
        RECT 112.345 134.190 113.045 134.360 ;
        RECT 110.475 132.330 110.805 133.940 ;
        RECT 111.845 132.330 112.175 133.940 ;
        RECT 109.605 131.910 110.305 132.080 ;
        RECT 110.975 131.910 111.675 132.080 ;
        RECT 112.345 131.910 113.045 132.080 ;
        RECT 110.475 130.050 110.805 131.660 ;
        RECT 111.845 130.050 112.175 131.660 ;
        RECT 109.605 129.630 110.305 129.800 ;
        RECT 110.975 129.630 111.675 129.800 ;
        RECT 112.345 129.630 113.045 129.800 ;
        RECT 110.475 127.770 110.805 129.380 ;
        RECT 111.845 127.770 112.175 129.380 ;
        RECT 109.605 127.350 110.305 127.520 ;
        RECT 110.975 127.350 111.675 127.520 ;
        RECT 112.345 127.350 113.045 127.520 ;
        RECT 110.475 125.490 110.805 127.100 ;
        RECT 111.845 125.490 112.175 127.100 ;
        RECT 109.605 125.070 110.305 125.240 ;
        RECT 110.975 125.070 111.675 125.240 ;
        RECT 112.345 125.070 113.045 125.240 ;
        RECT 110.475 123.210 110.805 124.820 ;
        RECT 111.845 123.210 112.175 124.820 ;
        RECT 109.605 122.790 110.305 122.960 ;
        RECT 110.975 122.790 111.675 122.960 ;
        RECT 112.345 122.790 113.045 122.960 ;
        RECT 110.475 120.930 110.805 122.540 ;
        RECT 111.845 120.930 112.175 122.540 ;
        RECT 109.605 120.510 110.305 120.680 ;
        RECT 110.975 120.510 111.675 120.680 ;
        RECT 112.345 120.510 113.045 120.680 ;
        RECT 110.475 118.650 110.805 120.260 ;
        RECT 111.845 118.650 112.175 120.260 ;
        RECT 109.605 118.230 110.305 118.400 ;
        RECT 110.975 118.230 111.675 118.400 ;
        RECT 112.345 118.230 113.045 118.400 ;
        RECT 110.475 116.370 110.805 117.980 ;
        RECT 111.845 116.370 112.175 117.980 ;
        RECT 109.605 115.950 110.305 116.120 ;
        RECT 110.975 115.950 111.675 116.120 ;
        RECT 112.345 115.950 113.045 116.120 ;
        RECT 110.475 114.090 110.805 115.700 ;
        RECT 111.845 114.090 112.175 115.700 ;
        RECT 109.605 113.670 110.305 113.840 ;
        RECT 110.975 113.670 111.675 113.840 ;
        RECT 112.345 113.670 113.045 113.840 ;
        RECT 110.475 111.810 110.805 113.420 ;
        RECT 111.845 111.810 112.175 113.420 ;
        RECT 109.605 111.390 110.305 111.560 ;
        RECT 110.975 111.390 111.675 111.560 ;
        RECT 112.345 111.390 113.045 111.560 ;
        RECT 110.475 109.530 110.805 111.140 ;
        RECT 111.845 109.530 112.175 111.140 ;
        RECT 109.605 109.110 110.305 109.280 ;
        RECT 110.975 109.110 111.675 109.280 ;
        RECT 112.345 109.110 113.045 109.280 ;
        RECT 110.475 107.250 110.805 108.860 ;
        RECT 111.845 107.250 112.175 108.860 ;
        RECT 109.605 106.830 110.305 107.000 ;
        RECT 110.975 106.830 111.675 107.000 ;
        RECT 112.345 106.830 113.045 107.000 ;
        RECT 110.475 104.970 110.805 106.580 ;
        RECT 111.845 104.970 112.175 106.580 ;
        RECT 109.605 104.550 110.305 104.720 ;
        RECT 110.975 104.550 111.675 104.720 ;
        RECT 112.345 104.550 113.045 104.720 ;
        RECT 110.475 102.690 110.805 104.300 ;
        RECT 111.845 102.690 112.175 104.300 ;
        RECT 109.605 102.270 110.305 102.440 ;
        RECT 110.975 102.270 111.675 102.440 ;
        RECT 112.345 102.270 113.045 102.440 ;
        RECT 110.475 100.410 110.805 102.020 ;
        RECT 111.845 100.410 112.175 102.020 ;
        RECT 109.605 99.990 110.305 100.160 ;
        RECT 110.975 99.990 111.675 100.160 ;
        RECT 112.345 99.990 113.045 100.160 ;
        RECT 110.475 98.130 110.805 99.740 ;
        RECT 111.845 98.130 112.175 99.740 ;
        RECT 109.605 97.710 110.305 97.880 ;
        RECT 110.975 97.710 111.675 97.880 ;
        RECT 112.345 97.710 113.045 97.880 ;
        RECT 110.475 95.850 110.805 97.460 ;
        RECT 111.845 95.850 112.175 97.460 ;
        RECT 109.605 95.430 110.305 95.600 ;
        RECT 110.975 95.430 111.675 95.600 ;
        RECT 112.345 95.430 113.045 95.600 ;
        RECT 110.475 93.570 110.805 95.180 ;
        RECT 111.845 93.570 112.175 95.180 ;
        RECT 109.605 93.150 110.305 93.320 ;
        RECT 110.975 93.150 111.675 93.320 ;
        RECT 112.345 93.150 113.045 93.320 ;
        RECT 110.475 91.290 110.805 92.900 ;
        RECT 111.845 91.290 112.175 92.900 ;
        RECT 109.605 90.870 110.305 91.040 ;
        RECT 110.975 90.870 111.675 91.040 ;
        RECT 112.345 90.870 113.045 91.040 ;
        RECT 110.475 89.010 110.805 90.620 ;
        RECT 111.845 89.010 112.175 90.620 ;
        RECT 109.605 88.590 110.305 88.760 ;
        RECT 110.975 88.590 111.675 88.760 ;
        RECT 112.345 88.590 113.045 88.760 ;
        RECT 110.475 86.730 110.805 88.340 ;
        RECT 111.845 86.730 112.175 88.340 ;
        RECT 109.605 86.310 110.305 86.480 ;
        RECT 110.975 86.310 111.675 86.480 ;
        RECT 112.345 86.310 113.045 86.480 ;
        RECT 110.475 84.450 110.805 86.060 ;
        RECT 111.845 84.450 112.175 86.060 ;
        RECT 109.605 84.030 110.305 84.200 ;
        RECT 110.975 84.030 111.675 84.200 ;
        RECT 112.345 84.030 113.045 84.200 ;
        RECT 110.475 82.170 110.805 83.780 ;
        RECT 111.845 82.170 112.175 83.780 ;
        RECT 109.605 81.750 110.305 81.920 ;
        RECT 110.975 81.750 111.675 81.920 ;
        RECT 112.345 81.750 113.045 81.920 ;
        RECT 110.475 79.890 110.805 81.500 ;
        RECT 111.845 79.890 112.175 81.500 ;
        RECT 109.605 79.470 110.305 79.640 ;
        RECT 110.975 79.470 111.675 79.640 ;
        RECT 112.345 79.470 113.045 79.640 ;
        RECT 110.475 77.610 110.805 79.220 ;
        RECT 111.845 77.610 112.175 79.220 ;
        RECT 109.605 77.190 110.305 77.360 ;
        RECT 110.975 77.190 111.675 77.360 ;
        RECT 112.345 77.190 113.045 77.360 ;
        RECT 110.475 75.330 110.805 76.940 ;
        RECT 111.845 75.330 112.175 76.940 ;
        RECT 109.605 74.910 110.305 75.080 ;
        RECT 110.975 74.910 111.675 75.080 ;
        RECT 112.345 74.910 113.045 75.080 ;
        RECT 110.475 73.050 110.805 74.660 ;
        RECT 111.845 73.050 112.175 74.660 ;
        RECT 109.605 72.630 110.305 72.800 ;
        RECT 110.975 72.630 111.675 72.800 ;
        RECT 112.345 72.630 113.045 72.800 ;
        RECT 110.475 70.770 110.805 72.380 ;
        RECT 111.845 70.770 112.175 72.380 ;
        RECT 109.605 70.350 110.305 70.520 ;
        RECT 110.975 70.350 111.675 70.520 ;
        RECT 112.345 70.350 113.045 70.520 ;
        RECT 110.475 68.490 110.805 70.100 ;
        RECT 111.845 68.490 112.175 70.100 ;
        RECT 109.605 68.070 110.305 68.240 ;
        RECT 110.975 68.070 111.675 68.240 ;
        RECT 112.345 68.070 113.045 68.240 ;
        RECT 110.475 66.210 110.805 67.820 ;
        RECT 111.845 66.210 112.175 67.820 ;
        RECT 109.605 65.790 110.305 65.960 ;
        RECT 110.975 65.790 111.675 65.960 ;
        RECT 112.345 65.790 113.045 65.960 ;
        RECT 110.475 63.930 110.805 65.540 ;
        RECT 111.845 63.930 112.175 65.540 ;
        RECT 109.605 63.510 110.305 63.680 ;
        RECT 110.975 63.510 111.675 63.680 ;
        RECT 112.345 63.510 113.045 63.680 ;
        RECT 113.845 63.010 114.015 164.500 ;
        RECT 121.840 164.460 125.850 164.630 ;
        RECT 114.925 117.905 117.565 118.075 ;
        RECT 114.925 114.235 115.095 117.905 ;
        RECT 115.895 117.275 116.595 117.445 ;
        RECT 115.895 116.845 116.595 117.015 ;
        RECT 116.765 116.845 117.095 117.015 ;
        RECT 115.895 116.415 116.595 116.585 ;
        RECT 115.395 115.985 115.725 116.155 ;
        RECT 115.895 115.985 116.595 116.155 ;
        RECT 115.895 115.555 116.595 115.725 ;
        RECT 115.895 115.125 116.595 115.295 ;
        RECT 116.765 115.125 117.095 115.295 ;
        RECT 115.895 114.695 116.595 114.865 ;
        RECT 117.395 114.235 117.565 117.905 ;
        RECT 114.925 114.065 117.565 114.235 ;
        RECT 118.195 117.670 121.135 117.840 ;
        RECT 114.925 113.275 117.565 113.445 ;
        RECT 114.925 109.525 115.095 113.275 ;
        RECT 115.895 112.605 116.595 112.775 ;
        RECT 115.395 112.175 115.725 112.345 ;
        RECT 115.895 112.175 116.595 112.345 ;
        RECT 115.895 111.745 116.595 111.915 ;
        RECT 115.895 111.315 116.595 111.485 ;
        RECT 116.765 111.315 117.095 111.485 ;
        RECT 115.895 110.885 116.595 111.055 ;
        RECT 115.395 110.455 115.725 110.625 ;
        RECT 115.895 110.455 116.595 110.625 ;
        RECT 115.895 110.025 116.595 110.195 ;
        RECT 117.395 109.525 117.565 113.275 ;
        RECT 118.195 109.700 118.365 117.670 ;
        RECT 119.165 117.040 120.165 117.210 ;
        RECT 118.665 116.610 118.995 116.780 ;
        RECT 119.165 116.610 120.165 116.780 ;
        RECT 119.165 116.180 120.165 116.350 ;
        RECT 118.665 115.750 118.995 115.920 ;
        RECT 119.165 115.750 120.165 115.920 ;
        RECT 119.165 115.320 120.165 115.490 ;
        RECT 118.665 114.890 118.995 115.060 ;
        RECT 119.165 114.890 120.165 115.060 ;
        RECT 119.165 114.460 120.165 114.630 ;
        RECT 119.165 114.030 120.165 114.200 ;
        RECT 120.335 114.030 120.665 114.200 ;
        RECT 119.165 113.600 120.165 113.770 ;
        RECT 119.165 113.170 120.165 113.340 ;
        RECT 120.335 113.170 120.665 113.340 ;
        RECT 119.165 112.740 120.165 112.910 ;
        RECT 118.665 112.310 118.995 112.480 ;
        RECT 119.165 112.310 120.165 112.480 ;
        RECT 119.165 111.880 120.165 112.050 ;
        RECT 118.665 111.450 118.995 111.620 ;
        RECT 119.165 111.450 120.165 111.620 ;
        RECT 119.165 111.020 120.165 111.190 ;
        RECT 118.665 110.590 118.995 110.760 ;
        RECT 119.165 110.590 120.165 110.760 ;
        RECT 119.165 110.160 120.165 110.330 ;
        RECT 120.965 109.700 121.135 117.670 ;
        RECT 118.195 109.530 121.135 109.700 ;
        RECT 114.925 109.355 117.565 109.525 ;
        RECT 114.925 83.705 117.565 83.875 ;
        RECT 114.925 80.035 115.095 83.705 ;
        RECT 115.895 83.075 116.595 83.245 ;
        RECT 115.895 82.645 116.595 82.815 ;
        RECT 116.765 82.645 117.095 82.815 ;
        RECT 115.895 82.215 116.595 82.385 ;
        RECT 115.395 81.785 115.725 81.955 ;
        RECT 115.895 81.785 116.595 81.955 ;
        RECT 115.895 81.355 116.595 81.525 ;
        RECT 115.895 80.925 116.595 81.095 ;
        RECT 116.765 80.925 117.095 81.095 ;
        RECT 115.895 80.495 116.595 80.665 ;
        RECT 117.395 80.035 117.565 83.705 ;
        RECT 114.925 79.865 117.565 80.035 ;
        RECT 118.195 83.470 121.135 83.640 ;
        RECT 114.925 79.075 117.565 79.245 ;
        RECT 114.925 75.325 115.095 79.075 ;
        RECT 115.895 78.405 116.595 78.575 ;
        RECT 115.395 77.975 115.725 78.145 ;
        RECT 115.895 77.975 116.595 78.145 ;
        RECT 115.895 77.545 116.595 77.715 ;
        RECT 115.895 77.115 116.595 77.285 ;
        RECT 116.765 77.115 117.095 77.285 ;
        RECT 115.895 76.685 116.595 76.855 ;
        RECT 115.395 76.255 115.725 76.425 ;
        RECT 115.895 76.255 116.595 76.425 ;
        RECT 115.895 75.825 116.595 75.995 ;
        RECT 117.395 75.325 117.565 79.075 ;
        RECT 118.195 75.500 118.365 83.470 ;
        RECT 119.165 82.840 120.165 83.010 ;
        RECT 118.665 82.410 118.995 82.580 ;
        RECT 119.165 82.410 120.165 82.580 ;
        RECT 119.165 81.980 120.165 82.150 ;
        RECT 118.665 81.550 118.995 81.720 ;
        RECT 119.165 81.550 120.165 81.720 ;
        RECT 119.165 81.120 120.165 81.290 ;
        RECT 118.665 80.690 118.995 80.860 ;
        RECT 119.165 80.690 120.165 80.860 ;
        RECT 119.165 80.260 120.165 80.430 ;
        RECT 119.165 79.830 120.165 80.000 ;
        RECT 120.335 79.830 120.665 80.000 ;
        RECT 119.165 79.400 120.165 79.570 ;
        RECT 119.165 78.970 120.165 79.140 ;
        RECT 120.335 78.970 120.665 79.140 ;
        RECT 119.165 78.540 120.165 78.710 ;
        RECT 118.665 78.110 118.995 78.280 ;
        RECT 119.165 78.110 120.165 78.280 ;
        RECT 119.165 77.680 120.165 77.850 ;
        RECT 118.665 77.250 118.995 77.420 ;
        RECT 119.165 77.250 120.165 77.420 ;
        RECT 119.165 76.820 120.165 76.990 ;
        RECT 118.665 76.390 118.995 76.560 ;
        RECT 119.165 76.390 120.165 76.560 ;
        RECT 119.165 75.960 120.165 76.130 ;
        RECT 120.965 75.500 121.135 83.470 ;
        RECT 121.840 76.730 122.010 164.460 ;
        RECT 122.810 163.830 123.510 164.000 ;
        RECT 124.180 163.830 124.880 164.000 ;
        RECT 122.310 161.970 122.640 163.580 ;
        RECT 125.050 161.970 125.380 163.580 ;
        RECT 122.810 161.550 123.510 161.720 ;
        RECT 124.180 161.550 124.880 161.720 ;
        RECT 122.310 159.690 122.640 161.300 ;
        RECT 125.050 159.690 125.380 161.300 ;
        RECT 122.810 159.270 123.510 159.440 ;
        RECT 124.180 159.270 124.880 159.440 ;
        RECT 122.310 157.410 122.640 159.020 ;
        RECT 123.680 157.410 124.010 159.020 ;
        RECT 125.050 157.410 125.380 159.020 ;
        RECT 122.810 156.990 123.510 157.160 ;
        RECT 124.180 156.990 124.880 157.160 ;
        RECT 122.310 155.130 122.640 156.740 ;
        RECT 123.680 155.130 124.010 156.740 ;
        RECT 125.050 155.130 125.380 156.740 ;
        RECT 122.810 154.710 123.510 154.880 ;
        RECT 124.180 154.710 124.880 154.880 ;
        RECT 122.310 152.850 122.640 154.460 ;
        RECT 123.680 152.850 124.010 154.460 ;
        RECT 125.050 152.850 125.380 154.460 ;
        RECT 122.810 152.430 123.510 152.600 ;
        RECT 124.180 152.430 124.880 152.600 ;
        RECT 122.310 150.570 122.640 152.180 ;
        RECT 123.680 150.570 124.010 152.180 ;
        RECT 125.050 150.570 125.380 152.180 ;
        RECT 122.810 150.150 123.510 150.320 ;
        RECT 124.180 150.150 124.880 150.320 ;
        RECT 122.310 148.290 122.640 149.900 ;
        RECT 123.680 148.290 124.010 149.900 ;
        RECT 125.050 148.290 125.380 149.900 ;
        RECT 122.810 147.870 123.510 148.040 ;
        RECT 124.180 147.870 124.880 148.040 ;
        RECT 122.310 146.010 122.640 147.620 ;
        RECT 123.680 146.010 124.010 147.620 ;
        RECT 125.050 146.010 125.380 147.620 ;
        RECT 122.810 145.590 123.510 145.760 ;
        RECT 124.180 145.590 124.880 145.760 ;
        RECT 122.310 143.730 122.640 145.340 ;
        RECT 123.680 143.730 124.010 145.340 ;
        RECT 125.050 143.730 125.380 145.340 ;
        RECT 122.810 143.310 123.510 143.480 ;
        RECT 124.180 143.310 124.880 143.480 ;
        RECT 122.310 141.450 122.640 143.060 ;
        RECT 123.680 141.450 124.010 143.060 ;
        RECT 125.050 141.450 125.380 143.060 ;
        RECT 122.810 141.030 123.510 141.200 ;
        RECT 124.180 141.030 124.880 141.200 ;
        RECT 122.310 139.170 122.640 140.780 ;
        RECT 123.680 139.170 124.010 140.780 ;
        RECT 125.050 139.170 125.380 140.780 ;
        RECT 122.810 138.750 123.510 138.920 ;
        RECT 124.180 138.750 124.880 138.920 ;
        RECT 122.310 136.890 122.640 138.500 ;
        RECT 123.680 136.890 124.010 138.500 ;
        RECT 125.050 136.890 125.380 138.500 ;
        RECT 122.810 136.470 123.510 136.640 ;
        RECT 124.180 136.470 124.880 136.640 ;
        RECT 122.310 134.610 122.640 136.220 ;
        RECT 123.680 134.610 124.010 136.220 ;
        RECT 125.050 134.610 125.380 136.220 ;
        RECT 122.810 134.190 123.510 134.360 ;
        RECT 124.180 134.190 124.880 134.360 ;
        RECT 122.310 132.330 122.640 133.940 ;
        RECT 123.680 132.330 124.010 133.940 ;
        RECT 125.050 132.330 125.380 133.940 ;
        RECT 122.810 131.910 123.510 132.080 ;
        RECT 124.180 131.910 124.880 132.080 ;
        RECT 122.310 130.050 122.640 131.660 ;
        RECT 123.680 130.050 124.010 131.660 ;
        RECT 125.050 130.050 125.380 131.660 ;
        RECT 122.810 129.630 123.510 129.800 ;
        RECT 124.180 129.630 124.880 129.800 ;
        RECT 122.310 127.770 122.640 129.380 ;
        RECT 123.680 127.770 124.010 129.380 ;
        RECT 125.050 127.770 125.380 129.380 ;
        RECT 122.810 127.350 123.510 127.520 ;
        RECT 124.180 127.350 124.880 127.520 ;
        RECT 122.310 125.490 122.640 127.100 ;
        RECT 123.680 125.490 124.010 127.100 ;
        RECT 125.050 125.490 125.380 127.100 ;
        RECT 122.810 125.070 123.510 125.240 ;
        RECT 124.180 125.070 124.880 125.240 ;
        RECT 122.310 123.210 122.640 124.820 ;
        RECT 123.680 123.210 124.010 124.820 ;
        RECT 125.050 123.210 125.380 124.820 ;
        RECT 122.810 122.790 123.510 122.960 ;
        RECT 124.180 122.790 124.880 122.960 ;
        RECT 122.310 120.930 122.640 122.540 ;
        RECT 123.680 120.930 124.010 122.540 ;
        RECT 125.050 120.930 125.380 122.540 ;
        RECT 122.810 120.510 123.510 120.680 ;
        RECT 124.180 120.510 124.880 120.680 ;
        RECT 122.310 118.650 122.640 120.260 ;
        RECT 123.680 118.650 124.010 120.260 ;
        RECT 125.050 118.650 125.380 120.260 ;
        RECT 122.810 118.230 123.510 118.400 ;
        RECT 124.180 118.230 124.880 118.400 ;
        RECT 122.310 116.370 122.640 117.980 ;
        RECT 123.680 116.370 124.010 117.980 ;
        RECT 125.050 116.370 125.380 117.980 ;
        RECT 122.810 115.950 123.510 116.120 ;
        RECT 124.180 115.950 124.880 116.120 ;
        RECT 122.310 114.090 122.640 115.700 ;
        RECT 123.680 114.090 124.010 115.700 ;
        RECT 125.050 114.090 125.380 115.700 ;
        RECT 122.810 113.670 123.510 113.840 ;
        RECT 124.180 113.670 124.880 113.840 ;
        RECT 122.310 111.810 122.640 113.420 ;
        RECT 123.680 111.810 124.010 113.420 ;
        RECT 125.050 111.810 125.380 113.420 ;
        RECT 122.810 111.390 123.510 111.560 ;
        RECT 124.180 111.390 124.880 111.560 ;
        RECT 122.310 109.530 122.640 111.140 ;
        RECT 123.680 109.530 124.010 111.140 ;
        RECT 125.050 109.530 125.380 111.140 ;
        RECT 122.810 109.110 123.510 109.280 ;
        RECT 124.180 109.110 124.880 109.280 ;
        RECT 122.310 107.250 122.640 108.860 ;
        RECT 123.680 107.250 124.010 108.860 ;
        RECT 125.050 107.250 125.380 108.860 ;
        RECT 122.810 106.830 123.510 107.000 ;
        RECT 124.180 106.830 124.880 107.000 ;
        RECT 122.310 104.970 122.640 106.580 ;
        RECT 123.680 104.970 124.010 106.580 ;
        RECT 125.050 104.970 125.380 106.580 ;
        RECT 122.810 104.550 123.510 104.720 ;
        RECT 124.180 104.550 124.880 104.720 ;
        RECT 122.310 102.690 122.640 104.300 ;
        RECT 123.680 102.690 124.010 104.300 ;
        RECT 125.050 102.690 125.380 104.300 ;
        RECT 122.810 102.270 123.510 102.440 ;
        RECT 124.180 102.270 124.880 102.440 ;
        RECT 122.310 100.410 122.640 102.020 ;
        RECT 123.680 100.410 124.010 102.020 ;
        RECT 125.050 100.410 125.380 102.020 ;
        RECT 122.810 99.990 123.510 100.160 ;
        RECT 124.180 99.990 124.880 100.160 ;
        RECT 122.310 98.130 122.640 99.740 ;
        RECT 123.680 98.130 124.010 99.740 ;
        RECT 125.050 98.130 125.380 99.740 ;
        RECT 122.810 97.710 123.510 97.880 ;
        RECT 124.180 97.710 124.880 97.880 ;
        RECT 122.310 95.850 122.640 97.460 ;
        RECT 123.680 95.850 124.010 97.460 ;
        RECT 125.050 95.850 125.380 97.460 ;
        RECT 122.810 95.430 123.510 95.600 ;
        RECT 124.180 95.430 124.880 95.600 ;
        RECT 122.310 93.570 122.640 95.180 ;
        RECT 123.680 93.570 124.010 95.180 ;
        RECT 125.050 93.570 125.380 95.180 ;
        RECT 122.810 93.150 123.510 93.320 ;
        RECT 124.180 93.150 124.880 93.320 ;
        RECT 122.310 91.290 122.640 92.900 ;
        RECT 123.680 91.290 124.010 92.900 ;
        RECT 125.050 91.290 125.380 92.900 ;
        RECT 122.810 90.870 123.510 91.040 ;
        RECT 124.180 90.870 124.880 91.040 ;
        RECT 122.310 89.010 122.640 90.620 ;
        RECT 125.050 89.010 125.380 90.620 ;
        RECT 122.810 88.590 123.510 88.760 ;
        RECT 124.180 88.590 124.880 88.760 ;
        RECT 122.310 86.730 122.640 88.340 ;
        RECT 125.050 86.730 125.380 88.340 ;
        RECT 122.810 86.310 123.510 86.480 ;
        RECT 124.180 86.310 124.880 86.480 ;
        RECT 122.310 84.450 122.640 86.060 ;
        RECT 125.050 84.450 125.380 86.060 ;
        RECT 122.810 84.030 123.510 84.200 ;
        RECT 124.180 84.030 124.880 84.200 ;
        RECT 122.310 82.170 122.640 83.780 ;
        RECT 125.050 82.170 125.380 83.780 ;
        RECT 122.810 81.750 123.510 81.920 ;
        RECT 124.180 81.750 124.880 81.920 ;
        RECT 122.310 79.890 122.640 81.500 ;
        RECT 125.050 79.890 125.380 81.500 ;
        RECT 122.810 79.470 123.510 79.640 ;
        RECT 124.180 79.470 124.880 79.640 ;
        RECT 122.310 77.610 122.640 79.220 ;
        RECT 123.680 77.610 124.010 79.220 ;
        RECT 125.050 77.610 125.380 79.220 ;
        RECT 122.810 77.190 123.510 77.360 ;
        RECT 124.180 77.190 124.880 77.360 ;
        RECT 125.680 76.730 125.850 164.460 ;
        RECT 121.840 76.560 125.850 76.730 ;
        RECT 118.195 75.330 121.135 75.500 ;
        RECT 114.925 75.155 117.565 75.325 ;
        RECT 108.635 62.840 114.015 63.010 ;
        RECT 114.775 70.380 117.415 70.550 ;
        RECT 114.775 60.090 114.945 70.380 ;
        RECT 115.745 69.710 116.445 69.880 ;
        RECT 116.615 67.850 116.945 69.460 ;
        RECT 115.745 67.430 116.445 67.600 ;
        RECT 115.245 65.570 115.575 67.180 ;
        RECT 115.745 65.150 116.445 65.320 ;
        RECT 115.245 63.290 115.575 64.900 ;
        RECT 115.745 62.870 116.445 63.040 ;
        RECT 116.615 61.010 116.945 62.620 ;
        RECT 115.745 60.590 116.445 60.760 ;
        RECT 117.245 60.090 117.415 70.380 ;
        RECT 118.470 70.100 123.825 70.270 ;
        RECT 118.470 65.490 118.640 70.100 ;
        RECT 119.440 69.430 120.140 69.600 ;
        RECT 122.155 69.430 122.855 69.600 ;
        RECT 118.940 69.000 119.270 69.170 ;
        RECT 119.440 69.000 120.140 69.170 ;
        RECT 121.655 69.000 121.985 69.170 ;
        RECT 122.155 69.000 122.855 69.170 ;
        RECT 119.440 68.570 120.140 68.740 ;
        RECT 122.155 68.570 122.855 68.740 ;
        RECT 119.440 68.140 120.140 68.310 ;
        RECT 120.310 68.140 120.640 68.310 ;
        RECT 122.155 68.140 122.855 68.310 ;
        RECT 123.025 68.140 123.355 68.310 ;
        RECT 119.440 67.710 120.140 67.880 ;
        RECT 122.155 67.710 122.855 67.880 ;
        RECT 119.440 67.280 120.140 67.450 ;
        RECT 120.310 67.280 120.640 67.450 ;
        RECT 122.155 67.280 122.855 67.450 ;
        RECT 123.025 67.280 123.355 67.450 ;
        RECT 119.440 66.850 120.140 67.020 ;
        RECT 122.155 66.850 122.855 67.020 ;
        RECT 118.940 66.420 119.270 66.590 ;
        RECT 119.440 66.420 120.140 66.590 ;
        RECT 121.655 66.420 121.985 66.590 ;
        RECT 122.155 66.420 122.855 66.590 ;
        RECT 119.440 65.990 120.140 66.160 ;
        RECT 122.155 65.990 122.855 66.160 ;
        RECT 123.655 65.490 123.825 70.100 ;
        RECT 118.470 65.320 123.825 65.490 ;
        RECT 124.455 70.060 127.095 70.230 ;
        RECT 118.470 64.810 123.825 64.980 ;
        RECT 118.470 60.280 118.640 64.810 ;
        RECT 119.440 64.180 120.140 64.350 ;
        RECT 122.155 64.180 122.855 64.350 ;
        RECT 118.940 63.750 119.270 63.920 ;
        RECT 119.440 63.750 120.140 63.920 ;
        RECT 121.655 63.750 121.985 63.920 ;
        RECT 122.155 63.750 122.855 63.920 ;
        RECT 119.440 63.320 120.140 63.490 ;
        RECT 122.155 63.320 122.855 63.490 ;
        RECT 119.440 62.890 120.140 63.060 ;
        RECT 120.310 62.890 120.640 63.060 ;
        RECT 122.155 62.890 122.855 63.060 ;
        RECT 123.025 62.890 123.355 63.060 ;
        RECT 119.440 62.460 120.140 62.630 ;
        RECT 122.155 62.460 122.855 62.630 ;
        RECT 119.440 62.030 120.140 62.200 ;
        RECT 120.310 62.030 120.640 62.200 ;
        RECT 122.155 62.030 122.855 62.200 ;
        RECT 123.025 62.030 123.355 62.200 ;
        RECT 119.440 61.600 120.140 61.770 ;
        RECT 122.155 61.600 122.855 61.770 ;
        RECT 118.940 61.170 119.270 61.340 ;
        RECT 119.440 61.170 120.140 61.340 ;
        RECT 121.655 61.170 121.985 61.340 ;
        RECT 122.155 61.170 122.855 61.340 ;
        RECT 119.440 60.740 120.140 60.910 ;
        RECT 122.155 60.740 122.855 60.910 ;
        RECT 123.655 60.280 123.825 64.810 ;
        RECT 118.470 60.110 123.825 60.280 ;
        RECT 124.455 60.370 124.625 70.060 ;
        RECT 125.425 69.430 126.125 69.600 ;
        RECT 124.925 69.000 125.255 69.170 ;
        RECT 125.425 69.000 126.125 69.170 ;
        RECT 125.425 68.570 126.125 68.740 ;
        RECT 124.925 68.140 125.255 68.310 ;
        RECT 125.425 68.140 126.125 68.310 ;
        RECT 125.425 67.710 126.125 67.880 ;
        RECT 124.925 67.280 125.255 67.450 ;
        RECT 125.425 67.280 126.125 67.450 ;
        RECT 125.425 66.850 126.125 67.020 ;
        RECT 124.925 66.420 125.255 66.590 ;
        RECT 125.425 66.420 126.125 66.590 ;
        RECT 125.425 65.990 126.125 66.160 ;
        RECT 125.425 65.560 126.125 65.730 ;
        RECT 126.295 65.560 126.625 65.730 ;
        RECT 125.425 65.130 126.125 65.300 ;
        RECT 125.425 64.700 126.125 64.870 ;
        RECT 126.295 64.700 126.625 64.870 ;
        RECT 125.425 64.270 126.125 64.440 ;
        RECT 124.925 63.840 125.255 64.010 ;
        RECT 125.425 63.840 126.125 64.010 ;
        RECT 125.425 63.410 126.125 63.580 ;
        RECT 124.925 62.980 125.255 63.150 ;
        RECT 125.425 62.980 126.125 63.150 ;
        RECT 125.425 62.550 126.125 62.720 ;
        RECT 124.925 62.120 125.255 62.290 ;
        RECT 125.425 62.120 126.125 62.290 ;
        RECT 125.425 61.690 126.125 61.860 ;
        RECT 124.925 61.260 125.255 61.430 ;
        RECT 125.425 61.260 126.125 61.430 ;
        RECT 125.425 60.830 126.125 61.000 ;
        RECT 126.925 60.370 127.095 70.060 ;
        RECT 124.455 60.200 127.095 60.370 ;
        RECT 114.775 59.920 117.415 60.090 ;
      LAYER mcon ;
        RECT 107.890 173.650 108.060 173.820 ;
        RECT 108.250 173.650 108.420 173.820 ;
        RECT 108.610 173.650 108.780 173.820 ;
        RECT 108.970 173.650 109.140 173.820 ;
        RECT 109.330 173.650 109.500 173.820 ;
        RECT 109.690 173.650 109.860 173.820 ;
        RECT 111.185 173.650 111.355 173.820 ;
        RECT 111.545 173.650 111.715 173.820 ;
        RECT 111.905 173.650 112.075 173.820 ;
        RECT 112.265 173.650 112.435 173.820 ;
        RECT 112.625 173.650 112.795 173.820 ;
        RECT 112.985 173.650 113.155 173.820 ;
        RECT 113.345 173.650 113.515 173.820 ;
        RECT 113.705 173.650 113.875 173.820 ;
        RECT 107.590 173.300 107.760 173.470 ;
        RECT 114.005 173.300 114.175 173.470 ;
        RECT 107.590 172.940 107.760 173.110 ;
        RECT 108.430 172.980 108.600 173.150 ;
        RECT 108.790 172.980 108.960 173.150 ;
        RECT 111.740 172.980 111.910 173.150 ;
        RECT 112.100 172.980 112.270 173.150 ;
        RECT 112.460 172.980 112.630 173.150 ;
        RECT 112.820 172.980 112.990 173.150 ;
        RECT 113.180 172.980 113.350 173.150 ;
        RECT 114.005 172.940 114.175 173.110 ;
        RECT 107.590 172.580 107.760 172.750 ;
        RECT 109.445 172.730 109.615 172.900 ;
        RECT 108.430 172.550 108.600 172.720 ;
        RECT 108.790 172.550 108.960 172.720 ;
        RECT 107.590 172.220 107.760 172.390 ;
        RECT 109.445 172.370 109.615 172.540 ;
        RECT 111.125 172.730 111.295 172.900 ;
        RECT 111.740 172.550 111.910 172.720 ;
        RECT 112.100 172.550 112.270 172.720 ;
        RECT 112.460 172.550 112.630 172.720 ;
        RECT 112.820 172.550 112.990 172.720 ;
        RECT 113.180 172.550 113.350 172.720 ;
        RECT 114.005 172.580 114.175 172.750 ;
        RECT 111.125 172.370 111.295 172.540 ;
        RECT 108.430 172.120 108.600 172.290 ;
        RECT 108.790 172.120 108.960 172.290 ;
        RECT 111.740 172.120 111.910 172.290 ;
        RECT 112.100 172.120 112.270 172.290 ;
        RECT 112.460 172.120 112.630 172.290 ;
        RECT 112.820 172.120 112.990 172.290 ;
        RECT 113.180 172.120 113.350 172.290 ;
        RECT 114.005 172.220 114.175 172.390 ;
        RECT 107.590 171.860 107.760 172.030 ;
        RECT 109.445 171.870 109.615 172.040 ;
        RECT 108.430 171.690 108.600 171.860 ;
        RECT 108.790 171.690 108.960 171.860 ;
        RECT 107.590 171.500 107.760 171.670 ;
        RECT 109.445 171.510 109.615 171.680 ;
        RECT 111.125 171.870 111.295 172.040 ;
        RECT 114.005 171.860 114.175 172.030 ;
        RECT 111.740 171.690 111.910 171.860 ;
        RECT 112.100 171.690 112.270 171.860 ;
        RECT 112.460 171.690 112.630 171.860 ;
        RECT 112.820 171.690 112.990 171.860 ;
        RECT 113.180 171.690 113.350 171.860 ;
        RECT 111.125 171.510 111.295 171.680 ;
        RECT 114.005 171.500 114.175 171.670 ;
        RECT 107.590 171.140 107.760 171.310 ;
        RECT 108.430 171.260 108.600 171.430 ;
        RECT 108.790 171.260 108.960 171.430 ;
        RECT 111.740 171.260 111.910 171.430 ;
        RECT 112.100 171.260 112.270 171.430 ;
        RECT 112.460 171.260 112.630 171.430 ;
        RECT 112.820 171.260 112.990 171.430 ;
        RECT 113.180 171.260 113.350 171.430 ;
        RECT 109.445 171.010 109.615 171.180 ;
        RECT 107.590 170.780 107.760 170.950 ;
        RECT 108.430 170.830 108.600 171.000 ;
        RECT 108.790 170.830 108.960 171.000 ;
        RECT 109.445 170.650 109.615 170.820 ;
        RECT 111.125 171.010 111.295 171.180 ;
        RECT 114.005 171.140 114.175 171.310 ;
        RECT 111.740 170.830 111.910 171.000 ;
        RECT 112.100 170.830 112.270 171.000 ;
        RECT 112.460 170.830 112.630 171.000 ;
        RECT 112.820 170.830 112.990 171.000 ;
        RECT 113.180 170.830 113.350 171.000 ;
        RECT 111.125 170.650 111.295 170.820 ;
        RECT 114.005 170.780 114.175 170.950 ;
        RECT 107.590 170.420 107.760 170.590 ;
        RECT 108.430 170.400 108.600 170.570 ;
        RECT 108.790 170.400 108.960 170.570 ;
        RECT 111.740 170.400 111.910 170.570 ;
        RECT 112.100 170.400 112.270 170.570 ;
        RECT 112.460 170.400 112.630 170.570 ;
        RECT 112.820 170.400 112.990 170.570 ;
        RECT 113.180 170.400 113.350 170.570 ;
        RECT 114.005 170.420 114.175 170.590 ;
        RECT 107.590 170.060 107.760 170.230 ;
        RECT 109.445 170.150 109.615 170.320 ;
        RECT 108.430 169.970 108.600 170.140 ;
        RECT 108.790 169.970 108.960 170.140 ;
        RECT 107.590 169.700 107.760 169.870 ;
        RECT 109.445 169.790 109.615 169.960 ;
        RECT 111.125 170.150 111.295 170.320 ;
        RECT 111.740 169.970 111.910 170.140 ;
        RECT 112.100 169.970 112.270 170.140 ;
        RECT 112.460 169.970 112.630 170.140 ;
        RECT 112.820 169.970 112.990 170.140 ;
        RECT 113.180 169.970 113.350 170.140 ;
        RECT 114.005 170.060 114.175 170.230 ;
        RECT 111.125 169.790 111.295 169.960 ;
        RECT 108.430 169.540 108.600 169.710 ;
        RECT 108.790 169.540 108.960 169.710 ;
        RECT 111.740 169.540 111.910 169.710 ;
        RECT 112.100 169.540 112.270 169.710 ;
        RECT 112.460 169.540 112.630 169.710 ;
        RECT 112.820 169.540 112.990 169.710 ;
        RECT 113.180 169.540 113.350 169.710 ;
        RECT 114.005 169.700 114.175 169.870 ;
        RECT 107.590 169.340 107.760 169.510 ;
        RECT 114.005 169.340 114.175 169.510 ;
        RECT 107.890 168.870 108.060 169.040 ;
        RECT 108.250 168.870 108.420 169.040 ;
        RECT 108.610 168.870 108.780 169.040 ;
        RECT 108.970 168.870 109.140 169.040 ;
        RECT 109.330 168.870 109.500 169.040 ;
        RECT 109.690 168.870 109.860 169.040 ;
        RECT 111.185 168.870 111.355 169.040 ;
        RECT 111.545 168.870 111.715 169.040 ;
        RECT 111.905 168.870 112.075 169.040 ;
        RECT 112.265 168.870 112.435 169.040 ;
        RECT 112.625 168.870 112.795 169.040 ;
        RECT 112.985 168.870 113.155 169.040 ;
        RECT 113.345 168.870 113.515 169.040 ;
        RECT 113.705 168.870 113.875 169.040 ;
        RECT 108.635 164.440 108.805 164.610 ;
        RECT 109.105 164.500 109.275 164.670 ;
        RECT 109.465 164.500 109.635 164.670 ;
        RECT 109.825 164.500 109.995 164.670 ;
        RECT 110.185 164.500 110.355 164.670 ;
        RECT 110.545 164.500 110.715 164.670 ;
        RECT 110.905 164.500 111.075 164.670 ;
        RECT 111.265 164.500 111.435 164.670 ;
        RECT 111.625 164.500 111.795 164.670 ;
        RECT 111.985 164.500 112.155 164.670 ;
        RECT 112.345 164.500 112.515 164.670 ;
        RECT 112.705 164.500 112.875 164.670 ;
        RECT 113.065 164.500 113.235 164.670 ;
        RECT 113.425 164.500 113.595 164.670 ;
        RECT 113.785 164.500 113.955 164.670 ;
        RECT 108.635 164.080 108.805 164.250 ;
        RECT 113.845 164.060 114.015 164.230 ;
        RECT 108.635 163.720 108.805 163.890 ;
        RECT 109.690 163.830 109.860 164.000 ;
        RECT 110.050 163.830 110.220 164.000 ;
        RECT 111.060 163.830 111.230 164.000 ;
        RECT 111.420 163.830 111.590 164.000 ;
        RECT 112.430 163.830 112.600 164.000 ;
        RECT 112.790 163.830 112.960 164.000 ;
        RECT 113.845 163.700 114.015 163.870 ;
        RECT 108.635 163.360 108.805 163.530 ;
        RECT 108.635 163.000 108.805 163.170 ;
        RECT 108.635 162.640 108.805 162.810 ;
        RECT 108.635 162.280 108.805 162.450 ;
        RECT 108.635 161.920 108.805 162.090 ;
        RECT 110.555 163.410 110.725 163.580 ;
        RECT 110.555 163.050 110.725 163.220 ;
        RECT 110.555 162.690 110.725 162.860 ;
        RECT 110.555 162.330 110.725 162.500 ;
        RECT 110.555 161.970 110.725 162.140 ;
        RECT 111.925 163.410 112.095 163.580 ;
        RECT 111.925 163.050 112.095 163.220 ;
        RECT 111.925 162.690 112.095 162.860 ;
        RECT 111.925 162.330 112.095 162.500 ;
        RECT 111.925 161.970 112.095 162.140 ;
        RECT 113.845 163.340 114.015 163.510 ;
        RECT 113.845 162.980 114.015 163.150 ;
        RECT 113.845 162.620 114.015 162.790 ;
        RECT 113.845 162.260 114.015 162.430 ;
        RECT 108.635 161.560 108.805 161.730 ;
        RECT 113.845 161.900 114.015 162.070 ;
        RECT 109.690 161.550 109.860 161.720 ;
        RECT 110.050 161.550 110.220 161.720 ;
        RECT 111.060 161.550 111.230 161.720 ;
        RECT 111.420 161.550 111.590 161.720 ;
        RECT 112.430 161.550 112.600 161.720 ;
        RECT 112.790 161.550 112.960 161.720 ;
        RECT 108.635 161.200 108.805 161.370 ;
        RECT 113.845 161.540 114.015 161.710 ;
        RECT 108.635 160.840 108.805 161.010 ;
        RECT 108.635 160.480 108.805 160.650 ;
        RECT 108.635 160.120 108.805 160.290 ;
        RECT 108.635 159.760 108.805 159.930 ;
        RECT 110.555 161.130 110.725 161.300 ;
        RECT 110.555 160.770 110.725 160.940 ;
        RECT 110.555 160.410 110.725 160.580 ;
        RECT 110.555 160.050 110.725 160.220 ;
        RECT 110.555 159.690 110.725 159.860 ;
        RECT 111.925 161.130 112.095 161.300 ;
        RECT 111.925 160.770 112.095 160.940 ;
        RECT 111.925 160.410 112.095 160.580 ;
        RECT 111.925 160.050 112.095 160.220 ;
        RECT 111.925 159.690 112.095 159.860 ;
        RECT 113.845 161.180 114.015 161.350 ;
        RECT 113.845 160.820 114.015 160.990 ;
        RECT 113.845 160.460 114.015 160.630 ;
        RECT 113.845 160.100 114.015 160.270 ;
        RECT 113.845 159.740 114.015 159.910 ;
        RECT 108.635 159.400 108.805 159.570 ;
        RECT 109.690 159.270 109.860 159.440 ;
        RECT 110.050 159.270 110.220 159.440 ;
        RECT 111.060 159.270 111.230 159.440 ;
        RECT 111.420 159.270 111.590 159.440 ;
        RECT 112.430 159.270 112.600 159.440 ;
        RECT 112.790 159.270 112.960 159.440 ;
        RECT 113.845 159.380 114.015 159.550 ;
        RECT 108.635 159.040 108.805 159.210 ;
        RECT 113.845 159.020 114.015 159.190 ;
        RECT 108.635 158.680 108.805 158.850 ;
        RECT 108.635 158.320 108.805 158.490 ;
        RECT 108.635 157.960 108.805 158.130 ;
        RECT 108.635 157.600 108.805 157.770 ;
        RECT 110.555 158.850 110.725 159.020 ;
        RECT 110.555 158.490 110.725 158.660 ;
        RECT 110.555 158.130 110.725 158.300 ;
        RECT 110.555 157.770 110.725 157.940 ;
        RECT 110.555 157.410 110.725 157.580 ;
        RECT 111.925 158.850 112.095 159.020 ;
        RECT 111.925 158.490 112.095 158.660 ;
        RECT 111.925 158.130 112.095 158.300 ;
        RECT 111.925 157.770 112.095 157.940 ;
        RECT 111.925 157.410 112.095 157.580 ;
        RECT 113.845 158.660 114.015 158.830 ;
        RECT 113.845 158.300 114.015 158.470 ;
        RECT 113.845 157.940 114.015 158.110 ;
        RECT 113.845 157.580 114.015 157.750 ;
        RECT 108.635 157.240 108.805 157.410 ;
        RECT 113.845 157.220 114.015 157.390 ;
        RECT 108.635 156.880 108.805 157.050 ;
        RECT 109.690 156.990 109.860 157.160 ;
        RECT 110.050 156.990 110.220 157.160 ;
        RECT 111.060 156.990 111.230 157.160 ;
        RECT 111.420 156.990 111.590 157.160 ;
        RECT 112.430 156.990 112.600 157.160 ;
        RECT 112.790 156.990 112.960 157.160 ;
        RECT 113.845 156.860 114.015 157.030 ;
        RECT 108.635 156.520 108.805 156.690 ;
        RECT 108.635 156.160 108.805 156.330 ;
        RECT 108.635 155.800 108.805 155.970 ;
        RECT 108.635 155.440 108.805 155.610 ;
        RECT 108.635 155.080 108.805 155.250 ;
        RECT 110.555 156.570 110.725 156.740 ;
        RECT 110.555 156.210 110.725 156.380 ;
        RECT 110.555 155.850 110.725 156.020 ;
        RECT 110.555 155.490 110.725 155.660 ;
        RECT 110.555 155.130 110.725 155.300 ;
        RECT 111.925 156.570 112.095 156.740 ;
        RECT 111.925 156.210 112.095 156.380 ;
        RECT 111.925 155.850 112.095 156.020 ;
        RECT 111.925 155.490 112.095 155.660 ;
        RECT 111.925 155.130 112.095 155.300 ;
        RECT 113.845 156.500 114.015 156.670 ;
        RECT 113.845 156.140 114.015 156.310 ;
        RECT 113.845 155.780 114.015 155.950 ;
        RECT 113.845 155.420 114.015 155.590 ;
        RECT 108.635 154.720 108.805 154.890 ;
        RECT 113.845 155.060 114.015 155.230 ;
        RECT 109.690 154.710 109.860 154.880 ;
        RECT 110.050 154.710 110.220 154.880 ;
        RECT 111.060 154.710 111.230 154.880 ;
        RECT 111.420 154.710 111.590 154.880 ;
        RECT 112.430 154.710 112.600 154.880 ;
        RECT 112.790 154.710 112.960 154.880 ;
        RECT 108.635 154.360 108.805 154.530 ;
        RECT 113.845 154.700 114.015 154.870 ;
        RECT 108.635 154.000 108.805 154.170 ;
        RECT 108.635 153.640 108.805 153.810 ;
        RECT 108.635 153.280 108.805 153.450 ;
        RECT 108.635 152.920 108.805 153.090 ;
        RECT 110.555 154.290 110.725 154.460 ;
        RECT 110.555 153.930 110.725 154.100 ;
        RECT 110.555 153.570 110.725 153.740 ;
        RECT 110.555 153.210 110.725 153.380 ;
        RECT 110.555 152.850 110.725 153.020 ;
        RECT 111.925 154.290 112.095 154.460 ;
        RECT 111.925 153.930 112.095 154.100 ;
        RECT 111.925 153.570 112.095 153.740 ;
        RECT 111.925 153.210 112.095 153.380 ;
        RECT 111.925 152.850 112.095 153.020 ;
        RECT 113.845 154.340 114.015 154.510 ;
        RECT 113.845 153.980 114.015 154.150 ;
        RECT 113.845 153.620 114.015 153.790 ;
        RECT 113.845 153.260 114.015 153.430 ;
        RECT 113.845 152.900 114.015 153.070 ;
        RECT 108.635 152.560 108.805 152.730 ;
        RECT 109.690 152.430 109.860 152.600 ;
        RECT 110.050 152.430 110.220 152.600 ;
        RECT 111.060 152.430 111.230 152.600 ;
        RECT 111.420 152.430 111.590 152.600 ;
        RECT 112.430 152.430 112.600 152.600 ;
        RECT 112.790 152.430 112.960 152.600 ;
        RECT 113.845 152.540 114.015 152.710 ;
        RECT 108.635 152.200 108.805 152.370 ;
        RECT 113.845 152.180 114.015 152.350 ;
        RECT 108.635 151.840 108.805 152.010 ;
        RECT 108.635 151.480 108.805 151.650 ;
        RECT 56.480 151.250 56.650 151.420 ;
        RECT 56.840 151.250 57.010 151.420 ;
        RECT 57.200 151.250 57.370 151.420 ;
        RECT 57.560 151.250 57.730 151.420 ;
        RECT 57.920 151.250 58.090 151.420 ;
        RECT 58.280 151.250 58.450 151.420 ;
        RECT 58.640 151.250 58.810 151.420 ;
        RECT 59.000 151.250 59.170 151.420 ;
        RECT 59.360 151.250 59.530 151.420 ;
        RECT 59.720 151.250 59.890 151.420 ;
        RECT 60.080 151.250 60.250 151.420 ;
        RECT 60.440 151.250 60.610 151.420 ;
        RECT 60.800 151.250 60.970 151.420 ;
        RECT 61.160 151.250 61.330 151.420 ;
        RECT 61.520 151.250 61.690 151.420 ;
        RECT 61.880 151.250 62.050 151.420 ;
        RECT 62.240 151.250 62.410 151.420 ;
        RECT 56.180 150.900 56.350 151.070 ;
        RECT 62.540 150.900 62.710 151.070 ;
        RECT 56.180 150.540 56.350 150.710 ;
        RECT 60.975 150.580 61.145 150.750 ;
        RECT 61.335 150.580 61.505 150.750 ;
        RECT 56.180 150.180 56.350 150.350 ;
        RECT 62.540 150.540 62.710 150.710 ;
        RECT 56.180 149.820 56.350 149.990 ;
        RECT 56.180 149.460 56.350 149.630 ;
        RECT 60.320 150.160 60.490 150.330 ;
        RECT 62.540 150.180 62.710 150.350 ;
        RECT 60.320 149.800 60.490 149.970 ;
        RECT 60.975 149.800 61.145 149.970 ;
        RECT 61.335 149.800 61.505 149.970 ;
        RECT 62.540 149.820 62.710 149.990 ;
        RECT 60.320 149.440 60.490 149.610 ;
        RECT 62.540 149.460 62.710 149.630 ;
        RECT 56.180 149.100 56.350 149.270 ;
        RECT 60.975 149.020 61.145 149.190 ;
        RECT 61.335 149.020 61.505 149.190 ;
        RECT 62.540 149.100 62.710 149.270 ;
        RECT 56.180 148.740 56.350 148.910 ;
        RECT 56.180 148.380 56.350 148.550 ;
        RECT 56.180 148.020 56.350 148.190 ;
        RECT 56.180 147.660 56.350 147.830 ;
        RECT 56.180 147.300 56.350 147.470 ;
        RECT 61.990 148.600 62.160 148.770 ;
        RECT 61.990 148.240 62.160 148.410 ;
        RECT 61.990 147.880 62.160 148.050 ;
        RECT 61.990 147.520 62.160 147.690 ;
        RECT 61.990 147.160 62.160 147.330 ;
        RECT 62.540 148.740 62.710 148.910 ;
        RECT 62.540 148.380 62.710 148.550 ;
        RECT 62.540 148.020 62.710 148.190 ;
        RECT 62.540 147.660 62.710 147.830 ;
        RECT 62.540 147.300 62.710 147.470 ;
        RECT 56.180 146.940 56.350 147.110 ;
        RECT 62.540 146.940 62.710 147.110 ;
        RECT 56.180 146.580 56.350 146.750 ;
        RECT 60.975 146.740 61.145 146.910 ;
        RECT 61.335 146.740 61.505 146.910 ;
        RECT 62.540 146.580 62.710 146.750 ;
        RECT 56.180 146.220 56.350 146.390 ;
        RECT 56.180 145.860 56.350 146.030 ;
        RECT 56.180 145.500 56.350 145.670 ;
        RECT 56.180 145.140 56.350 145.310 ;
        RECT 56.180 144.780 56.350 144.950 ;
        RECT 61.990 146.320 62.160 146.490 ;
        RECT 61.990 145.960 62.160 146.130 ;
        RECT 61.990 145.600 62.160 145.770 ;
        RECT 61.990 145.240 62.160 145.410 ;
        RECT 61.990 144.880 62.160 145.050 ;
        RECT 62.540 146.220 62.710 146.390 ;
        RECT 62.540 145.860 62.710 146.030 ;
        RECT 62.540 145.500 62.710 145.670 ;
        RECT 62.540 145.140 62.710 145.310 ;
        RECT 62.540 144.780 62.710 144.950 ;
        RECT 56.180 144.420 56.350 144.590 ;
        RECT 60.975 144.460 61.145 144.630 ;
        RECT 61.335 144.460 61.505 144.630 ;
        RECT 56.180 144.060 56.350 144.230 ;
        RECT 62.540 144.420 62.710 144.590 ;
        RECT 56.180 143.700 56.350 143.870 ;
        RECT 56.180 143.340 56.350 143.510 ;
        RECT 60.320 144.040 60.490 144.210 ;
        RECT 62.540 144.060 62.710 144.230 ;
        RECT 60.320 143.680 60.490 143.850 ;
        RECT 60.975 143.680 61.145 143.850 ;
        RECT 61.335 143.680 61.505 143.850 ;
        RECT 62.540 143.700 62.710 143.870 ;
        RECT 60.320 143.320 60.490 143.490 ;
        RECT 62.540 143.340 62.710 143.510 ;
        RECT 56.180 142.980 56.350 143.150 ;
        RECT 60.975 142.900 61.145 143.070 ;
        RECT 61.335 142.900 61.505 143.070 ;
        RECT 62.540 142.980 62.710 143.150 ;
        RECT 56.180 142.620 56.350 142.790 ;
        RECT 56.180 142.260 56.350 142.430 ;
        RECT 56.180 141.900 56.350 142.070 ;
        RECT 60.320 142.480 60.490 142.650 ;
        RECT 62.540 142.620 62.710 142.790 ;
        RECT 60.320 142.120 60.490 142.290 ;
        RECT 60.975 142.120 61.145 142.290 ;
        RECT 61.335 142.120 61.505 142.290 ;
        RECT 62.540 142.260 62.710 142.430 ;
        RECT 60.320 141.760 60.490 141.930 ;
        RECT 64.965 151.250 65.135 151.420 ;
        RECT 65.325 151.250 65.495 151.420 ;
        RECT 65.685 151.250 65.855 151.420 ;
        RECT 66.045 151.250 66.215 151.420 ;
        RECT 66.405 151.250 66.575 151.420 ;
        RECT 64.435 150.900 64.605 151.070 ;
        RECT 66.705 150.900 66.875 151.070 ;
        RECT 64.435 150.540 64.605 150.710 ;
        RECT 65.570 150.580 65.740 150.750 ;
        RECT 64.435 150.180 64.605 150.350 ;
        RECT 66.705 150.540 66.875 150.710 ;
        RECT 64.435 149.820 64.605 149.990 ;
        RECT 66.155 150.160 66.325 150.330 ;
        RECT 65.570 149.800 65.740 149.970 ;
        RECT 66.155 149.800 66.325 149.970 ;
        RECT 64.435 149.460 64.605 149.630 ;
        RECT 66.155 149.440 66.325 149.610 ;
        RECT 66.705 150.180 66.875 150.350 ;
        RECT 66.705 149.820 66.875 149.990 ;
        RECT 66.705 149.460 66.875 149.630 ;
        RECT 64.435 149.100 64.605 149.270 ;
        RECT 65.570 149.020 65.740 149.190 ;
        RECT 66.705 149.100 66.875 149.270 ;
        RECT 64.435 148.740 64.605 148.910 ;
        RECT 64.435 148.380 64.605 148.550 ;
        RECT 64.435 148.020 64.605 148.190 ;
        RECT 64.435 147.660 64.605 147.830 ;
        RECT 64.435 147.300 64.605 147.470 ;
        RECT 64.985 148.600 65.155 148.770 ;
        RECT 64.985 148.240 65.155 148.410 ;
        RECT 64.985 147.880 65.155 148.050 ;
        RECT 64.985 147.520 65.155 147.690 ;
        RECT 64.985 147.160 65.155 147.330 ;
        RECT 66.705 148.740 66.875 148.910 ;
        RECT 66.705 148.380 66.875 148.550 ;
        RECT 66.705 148.020 66.875 148.190 ;
        RECT 66.705 147.660 66.875 147.830 ;
        RECT 66.705 147.300 66.875 147.470 ;
        RECT 64.435 146.940 64.605 147.110 ;
        RECT 66.705 146.940 66.875 147.110 ;
        RECT 64.435 146.580 64.605 146.750 ;
        RECT 65.570 146.740 65.740 146.910 ;
        RECT 66.705 146.580 66.875 146.750 ;
        RECT 64.435 146.220 64.605 146.390 ;
        RECT 64.435 145.860 64.605 146.030 ;
        RECT 64.435 145.500 64.605 145.670 ;
        RECT 64.435 145.140 64.605 145.310 ;
        RECT 64.435 144.780 64.605 144.950 ;
        RECT 64.985 146.320 65.155 146.490 ;
        RECT 64.985 145.960 65.155 146.130 ;
        RECT 64.985 145.600 65.155 145.770 ;
        RECT 64.985 145.240 65.155 145.410 ;
        RECT 64.985 144.880 65.155 145.050 ;
        RECT 66.705 146.220 66.875 146.390 ;
        RECT 66.705 145.860 66.875 146.030 ;
        RECT 66.705 145.500 66.875 145.670 ;
        RECT 66.705 145.140 66.875 145.310 ;
        RECT 66.705 144.780 66.875 144.950 ;
        RECT 64.435 144.420 64.605 144.590 ;
        RECT 65.570 144.460 65.740 144.630 ;
        RECT 64.435 144.060 64.605 144.230 ;
        RECT 66.705 144.420 66.875 144.590 ;
        RECT 64.435 143.700 64.605 143.870 ;
        RECT 66.155 144.040 66.325 144.210 ;
        RECT 65.570 143.680 65.740 143.850 ;
        RECT 66.155 143.680 66.325 143.850 ;
        RECT 64.435 143.340 64.605 143.510 ;
        RECT 66.155 143.320 66.325 143.490 ;
        RECT 66.705 144.060 66.875 144.230 ;
        RECT 66.705 143.700 66.875 143.870 ;
        RECT 66.705 143.340 66.875 143.510 ;
        RECT 64.435 142.980 64.605 143.150 ;
        RECT 65.570 142.900 65.740 143.070 ;
        RECT 66.705 142.980 66.875 143.150 ;
        RECT 64.435 142.620 64.605 142.790 ;
        RECT 66.705 142.620 66.875 142.790 ;
        RECT 92.215 151.250 92.385 151.420 ;
        RECT 92.575 151.250 92.745 151.420 ;
        RECT 92.935 151.250 93.105 151.420 ;
        RECT 93.295 151.250 93.465 151.420 ;
        RECT 93.655 151.250 93.825 151.420 ;
        RECT 91.915 150.900 92.085 151.070 ;
        RECT 94.185 150.900 94.355 151.070 ;
        RECT 91.915 150.540 92.085 150.710 ;
        RECT 93.050 150.580 93.220 150.750 ;
        RECT 91.915 150.180 92.085 150.350 ;
        RECT 94.185 150.540 94.355 150.710 ;
        RECT 91.915 149.820 92.085 149.990 ;
        RECT 91.915 149.460 92.085 149.630 ;
        RECT 92.465 150.160 92.635 150.330 ;
        RECT 94.185 150.180 94.355 150.350 ;
        RECT 92.465 149.800 92.635 149.970 ;
        RECT 93.050 149.800 93.220 149.970 ;
        RECT 94.185 149.820 94.355 149.990 ;
        RECT 92.465 149.440 92.635 149.610 ;
        RECT 94.185 149.460 94.355 149.630 ;
        RECT 91.915 149.100 92.085 149.270 ;
        RECT 93.050 149.020 93.220 149.190 ;
        RECT 94.185 149.100 94.355 149.270 ;
        RECT 91.915 148.740 92.085 148.910 ;
        RECT 91.915 148.380 92.085 148.550 ;
        RECT 91.915 148.020 92.085 148.190 ;
        RECT 91.915 147.660 92.085 147.830 ;
        RECT 91.915 147.300 92.085 147.470 ;
        RECT 93.635 148.600 93.805 148.770 ;
        RECT 93.635 148.240 93.805 148.410 ;
        RECT 93.635 147.880 93.805 148.050 ;
        RECT 93.635 147.520 93.805 147.690 ;
        RECT 93.635 147.160 93.805 147.330 ;
        RECT 94.185 148.740 94.355 148.910 ;
        RECT 94.185 148.380 94.355 148.550 ;
        RECT 94.185 148.020 94.355 148.190 ;
        RECT 94.185 147.660 94.355 147.830 ;
        RECT 94.185 147.300 94.355 147.470 ;
        RECT 91.915 146.940 92.085 147.110 ;
        RECT 94.185 146.940 94.355 147.110 ;
        RECT 91.915 146.580 92.085 146.750 ;
        RECT 93.050 146.740 93.220 146.910 ;
        RECT 94.185 146.580 94.355 146.750 ;
        RECT 91.915 146.220 92.085 146.390 ;
        RECT 91.915 145.860 92.085 146.030 ;
        RECT 91.915 145.500 92.085 145.670 ;
        RECT 91.915 145.140 92.085 145.310 ;
        RECT 91.915 144.780 92.085 144.950 ;
        RECT 93.635 146.320 93.805 146.490 ;
        RECT 93.635 145.960 93.805 146.130 ;
        RECT 93.635 145.600 93.805 145.770 ;
        RECT 93.635 145.240 93.805 145.410 ;
        RECT 93.635 144.880 93.805 145.050 ;
        RECT 94.185 146.220 94.355 146.390 ;
        RECT 94.185 145.860 94.355 146.030 ;
        RECT 94.185 145.500 94.355 145.670 ;
        RECT 94.185 145.140 94.355 145.310 ;
        RECT 94.185 144.780 94.355 144.950 ;
        RECT 91.915 144.420 92.085 144.590 ;
        RECT 93.050 144.460 93.220 144.630 ;
        RECT 91.915 144.060 92.085 144.230 ;
        RECT 94.185 144.420 94.355 144.590 ;
        RECT 91.915 143.700 92.085 143.870 ;
        RECT 91.915 143.340 92.085 143.510 ;
        RECT 92.465 144.040 92.635 144.210 ;
        RECT 94.185 144.060 94.355 144.230 ;
        RECT 92.465 143.680 92.635 143.850 ;
        RECT 93.050 143.680 93.220 143.850 ;
        RECT 94.185 143.700 94.355 143.870 ;
        RECT 92.465 143.320 92.635 143.490 ;
        RECT 94.185 143.340 94.355 143.510 ;
        RECT 91.915 142.980 92.085 143.150 ;
        RECT 93.050 142.900 93.220 143.070 ;
        RECT 94.185 142.980 94.355 143.150 ;
        RECT 64.965 142.230 65.135 142.400 ;
        RECT 65.325 142.230 65.495 142.400 ;
        RECT 65.685 142.230 65.855 142.400 ;
        RECT 66.045 142.230 66.215 142.400 ;
        RECT 66.405 142.230 66.575 142.400 ;
        RECT 72.980 142.530 73.150 142.700 ;
        RECT 73.340 142.530 73.510 142.700 ;
        RECT 73.700 142.530 73.870 142.700 ;
        RECT 74.060 142.530 74.230 142.700 ;
        RECT 74.420 142.530 74.590 142.700 ;
        RECT 74.780 142.530 74.950 142.700 ;
        RECT 75.140 142.530 75.310 142.700 ;
        RECT 75.500 142.530 75.670 142.700 ;
        RECT 75.860 142.530 76.030 142.700 ;
        RECT 76.220 142.530 76.390 142.700 ;
        RECT 76.580 142.530 76.750 142.700 ;
        RECT 76.940 142.530 77.110 142.700 ;
        RECT 77.300 142.530 77.470 142.700 ;
        RECT 62.540 141.900 62.710 142.070 ;
        RECT 56.180 141.540 56.350 141.710 ;
        RECT 62.540 141.540 62.710 141.710 ;
        RECT 56.180 141.180 56.350 141.350 ;
        RECT 57.385 141.340 57.555 141.510 ;
        RECT 57.745 141.340 57.915 141.510 ;
        RECT 60.975 141.340 61.145 141.510 ;
        RECT 61.335 141.340 61.505 141.510 ;
        RECT 62.540 141.180 62.710 141.350 ;
        RECT 56.180 140.820 56.350 140.990 ;
        RECT 56.180 140.460 56.350 140.630 ;
        RECT 56.180 140.100 56.350 140.270 ;
        RECT 56.180 139.740 56.350 139.910 ;
        RECT 56.180 139.380 56.350 139.550 ;
        RECT 58.400 140.920 58.570 141.090 ;
        RECT 58.400 140.560 58.570 140.730 ;
        RECT 58.400 140.200 58.570 140.370 ;
        RECT 58.400 139.840 58.570 140.010 ;
        RECT 58.400 139.480 58.570 139.650 ;
        RECT 60.320 140.920 60.490 141.090 ;
        RECT 60.320 140.560 60.490 140.730 ;
        RECT 60.320 140.200 60.490 140.370 ;
        RECT 60.320 139.840 60.490 140.010 ;
        RECT 60.320 139.480 60.490 139.650 ;
        RECT 61.990 140.920 62.160 141.090 ;
        RECT 61.990 140.560 62.160 140.730 ;
        RECT 61.990 140.200 62.160 140.370 ;
        RECT 61.990 139.840 62.160 140.010 ;
        RECT 61.990 139.480 62.160 139.650 ;
        RECT 62.540 140.820 62.710 140.990 ;
        RECT 62.540 140.460 62.710 140.630 ;
        RECT 62.540 140.100 62.710 140.270 ;
        RECT 62.540 139.740 62.710 139.910 ;
        RECT 62.540 139.380 62.710 139.550 ;
        RECT 56.180 139.020 56.350 139.190 ;
        RECT 57.385 139.060 57.555 139.230 ;
        RECT 57.745 139.060 57.915 139.230 ;
        RECT 60.975 139.060 61.145 139.230 ;
        RECT 61.335 139.060 61.505 139.230 ;
        RECT 56.180 138.660 56.350 138.830 ;
        RECT 62.540 139.020 62.710 139.190 ;
        RECT 56.180 138.300 56.350 138.470 ;
        RECT 56.180 137.940 56.350 138.110 ;
        RECT 56.180 137.580 56.350 137.750 ;
        RECT 56.180 137.220 56.350 137.390 ;
        RECT 58.400 138.640 58.570 138.810 ;
        RECT 58.400 138.280 58.570 138.450 ;
        RECT 58.400 137.920 58.570 138.090 ;
        RECT 58.400 137.560 58.570 137.730 ;
        RECT 58.400 137.200 58.570 137.370 ;
        RECT 60.320 138.640 60.490 138.810 ;
        RECT 60.320 138.280 60.490 138.450 ;
        RECT 60.320 137.920 60.490 138.090 ;
        RECT 60.320 137.560 60.490 137.730 ;
        RECT 60.320 137.200 60.490 137.370 ;
        RECT 61.990 138.640 62.160 138.810 ;
        RECT 61.990 138.280 62.160 138.450 ;
        RECT 61.990 137.920 62.160 138.090 ;
        RECT 61.990 137.560 62.160 137.730 ;
        RECT 61.990 137.200 62.160 137.370 ;
        RECT 62.540 138.660 62.710 138.830 ;
        RECT 62.540 138.300 62.710 138.470 ;
        RECT 72.590 142.180 72.760 142.350 ;
        RECT 77.600 142.180 77.770 142.350 ;
        RECT 72.590 141.820 72.760 141.990 ;
        RECT 73.725 141.900 73.895 142.070 ;
        RECT 77.600 141.820 77.770 141.990 ;
        RECT 72.590 141.460 72.760 141.630 ;
        RECT 72.590 141.100 72.760 141.270 ;
        RECT 72.590 140.740 72.760 140.910 ;
        RECT 74.310 141.515 74.480 141.685 ;
        RECT 76.465 141.500 76.635 141.670 ;
        RECT 74.310 141.155 74.480 141.325 ;
        RECT 77.600 141.460 77.770 141.630 ;
        RECT 74.310 140.795 74.480 140.965 ;
        RECT 73.725 140.620 73.895 140.790 ;
        RECT 72.590 140.380 72.760 140.550 ;
        RECT 72.590 140.020 72.760 140.190 ;
        RECT 72.590 139.660 72.760 139.830 ;
        RECT 74.310 140.435 74.480 140.605 ;
        RECT 74.310 140.075 74.480 140.245 ;
        RECT 74.310 139.715 74.480 139.885 ;
        RECT 75.880 141.115 76.050 141.285 ;
        RECT 75.880 140.755 76.050 140.925 ;
        RECT 75.880 140.395 76.050 140.565 ;
        RECT 75.880 140.035 76.050 140.205 ;
        RECT 75.880 139.675 76.050 139.845 ;
        RECT 72.590 139.300 72.760 139.470 ;
        RECT 73.725 139.340 73.895 139.510 ;
        RECT 72.590 138.940 72.760 139.110 ;
        RECT 75.880 139.315 76.050 139.485 ;
        RECT 72.590 138.580 72.760 138.750 ;
        RECT 72.590 138.220 72.760 138.390 ;
        RECT 62.540 137.940 62.710 138.110 ;
        RECT 62.540 137.580 62.710 137.750 ;
        RECT 62.540 137.220 62.710 137.390 ;
        RECT 56.180 136.860 56.350 137.030 ;
        RECT 57.385 136.780 57.555 136.950 ;
        RECT 57.745 136.780 57.915 136.950 ;
        RECT 60.975 136.780 61.145 136.950 ;
        RECT 61.335 136.780 61.505 136.950 ;
        RECT 62.540 136.860 62.710 137.030 ;
        RECT 56.180 136.500 56.350 136.670 ;
        RECT 56.180 136.140 56.350 136.310 ;
        RECT 56.180 135.780 56.350 135.950 ;
        RECT 56.180 135.420 56.350 135.590 ;
        RECT 56.180 135.060 56.350 135.230 ;
        RECT 58.400 136.360 58.570 136.530 ;
        RECT 58.400 136.000 58.570 136.170 ;
        RECT 58.400 135.640 58.570 135.810 ;
        RECT 58.400 135.280 58.570 135.450 ;
        RECT 58.400 134.920 58.570 135.090 ;
        RECT 60.320 136.360 60.490 136.530 ;
        RECT 60.320 136.000 60.490 136.170 ;
        RECT 60.320 135.640 60.490 135.810 ;
        RECT 60.320 135.280 60.490 135.450 ;
        RECT 60.320 134.920 60.490 135.090 ;
        RECT 61.990 136.360 62.160 136.530 ;
        RECT 61.990 136.000 62.160 136.170 ;
        RECT 61.990 135.640 62.160 135.810 ;
        RECT 61.990 135.280 62.160 135.450 ;
        RECT 61.990 134.920 62.160 135.090 ;
        RECT 62.540 136.500 62.710 136.670 ;
        RECT 62.540 136.140 62.710 136.310 ;
        RECT 62.540 135.780 62.710 135.950 ;
        RECT 62.540 135.420 62.710 135.590 ;
        RECT 62.540 135.060 62.710 135.230 ;
        RECT 56.180 134.700 56.350 134.870 ;
        RECT 62.540 134.700 62.710 134.870 ;
        RECT 56.180 134.340 56.350 134.510 ;
        RECT 57.385 134.500 57.555 134.670 ;
        RECT 57.745 134.500 57.915 134.670 ;
        RECT 60.975 134.500 61.145 134.670 ;
        RECT 61.335 134.500 61.505 134.670 ;
        RECT 62.540 134.340 62.710 134.510 ;
        RECT 56.180 133.980 56.350 134.150 ;
        RECT 56.180 133.620 56.350 133.790 ;
        RECT 56.180 133.260 56.350 133.430 ;
        RECT 56.180 132.900 56.350 133.070 ;
        RECT 56.180 132.540 56.350 132.710 ;
        RECT 58.400 134.080 58.570 134.250 ;
        RECT 58.400 133.720 58.570 133.890 ;
        RECT 58.400 133.360 58.570 133.530 ;
        RECT 58.400 133.000 58.570 133.170 ;
        RECT 58.400 132.640 58.570 132.810 ;
        RECT 60.320 134.080 60.490 134.250 ;
        RECT 60.320 133.720 60.490 133.890 ;
        RECT 60.320 133.360 60.490 133.530 ;
        RECT 60.320 133.000 60.490 133.170 ;
        RECT 60.320 132.640 60.490 132.810 ;
        RECT 61.990 134.080 62.160 134.250 ;
        RECT 61.990 133.720 62.160 133.890 ;
        RECT 61.990 133.360 62.160 133.530 ;
        RECT 61.990 133.000 62.160 133.170 ;
        RECT 61.990 132.640 62.160 132.810 ;
        RECT 62.540 133.980 62.710 134.150 ;
        RECT 62.540 133.620 62.710 133.790 ;
        RECT 62.540 133.260 62.710 133.430 ;
        RECT 62.540 132.900 62.710 133.070 ;
        RECT 62.540 132.540 62.710 132.710 ;
        RECT 56.180 132.180 56.350 132.350 ;
        RECT 57.385 132.220 57.555 132.390 ;
        RECT 57.745 132.220 57.915 132.390 ;
        RECT 60.975 132.220 61.145 132.390 ;
        RECT 61.335 132.220 61.505 132.390 ;
        RECT 56.180 131.820 56.350 131.990 ;
        RECT 62.540 132.180 62.710 132.350 ;
        RECT 56.180 131.460 56.350 131.630 ;
        RECT 56.180 131.100 56.350 131.270 ;
        RECT 56.180 130.740 56.350 130.910 ;
        RECT 56.180 130.380 56.350 130.550 ;
        RECT 58.400 131.800 58.570 131.970 ;
        RECT 58.400 131.440 58.570 131.610 ;
        RECT 58.400 131.080 58.570 131.250 ;
        RECT 58.400 130.720 58.570 130.890 ;
        RECT 58.400 130.360 58.570 130.530 ;
        RECT 60.320 131.800 60.490 131.970 ;
        RECT 60.320 131.440 60.490 131.610 ;
        RECT 60.320 131.080 60.490 131.250 ;
        RECT 60.320 130.720 60.490 130.890 ;
        RECT 60.320 130.360 60.490 130.530 ;
        RECT 61.990 131.800 62.160 131.970 ;
        RECT 61.990 131.440 62.160 131.610 ;
        RECT 61.990 131.080 62.160 131.250 ;
        RECT 61.990 130.720 62.160 130.890 ;
        RECT 61.990 130.360 62.160 130.530 ;
        RECT 62.540 131.820 62.710 131.990 ;
        RECT 62.540 131.460 62.710 131.630 ;
        RECT 62.540 131.100 62.710 131.270 ;
        RECT 62.540 130.740 62.710 130.910 ;
        RECT 62.540 130.380 62.710 130.550 ;
        RECT 56.180 130.020 56.350 130.190 ;
        RECT 57.385 129.940 57.555 130.110 ;
        RECT 57.745 129.940 57.915 130.110 ;
        RECT 60.975 129.940 61.145 130.110 ;
        RECT 61.335 129.940 61.505 130.110 ;
        RECT 62.540 130.020 62.710 130.190 ;
        RECT 56.180 129.660 56.350 129.830 ;
        RECT 56.180 129.300 56.350 129.470 ;
        RECT 56.180 128.940 56.350 129.110 ;
        RECT 56.180 128.580 56.350 128.750 ;
        RECT 56.180 128.220 56.350 128.390 ;
        RECT 56.730 129.520 56.900 129.690 ;
        RECT 56.730 129.160 56.900 129.330 ;
        RECT 56.730 128.800 56.900 128.970 ;
        RECT 56.730 128.440 56.900 128.610 ;
        RECT 56.730 128.080 56.900 128.250 ;
        RECT 60.320 129.520 60.490 129.690 ;
        RECT 60.320 129.160 60.490 129.330 ;
        RECT 60.320 128.800 60.490 128.970 ;
        RECT 60.320 128.440 60.490 128.610 ;
        RECT 60.320 128.080 60.490 128.250 ;
        RECT 61.990 129.520 62.160 129.690 ;
        RECT 61.990 129.160 62.160 129.330 ;
        RECT 61.990 128.800 62.160 128.970 ;
        RECT 61.990 128.440 62.160 128.610 ;
        RECT 61.990 128.080 62.160 128.250 ;
        RECT 62.540 129.660 62.710 129.830 ;
        RECT 62.540 129.300 62.710 129.470 ;
        RECT 62.540 128.940 62.710 129.110 ;
        RECT 62.540 128.580 62.710 128.750 ;
        RECT 62.540 128.220 62.710 128.390 ;
        RECT 56.180 127.860 56.350 128.030 ;
        RECT 62.540 127.860 62.710 128.030 ;
        RECT 56.180 127.500 56.350 127.670 ;
        RECT 57.385 127.660 57.555 127.830 ;
        RECT 57.745 127.660 57.915 127.830 ;
        RECT 60.975 127.660 61.145 127.830 ;
        RECT 61.335 127.660 61.505 127.830 ;
        RECT 62.540 127.500 62.710 127.670 ;
        RECT 56.180 127.140 56.350 127.310 ;
        RECT 56.180 126.780 56.350 126.950 ;
        RECT 56.180 126.420 56.350 126.590 ;
        RECT 56.180 126.060 56.350 126.230 ;
        RECT 56.180 125.700 56.350 125.870 ;
        RECT 56.730 127.240 56.900 127.410 ;
        RECT 56.730 126.880 56.900 127.050 ;
        RECT 56.730 126.520 56.900 126.690 ;
        RECT 56.730 126.160 56.900 126.330 ;
        RECT 56.730 125.800 56.900 125.970 ;
        RECT 60.320 127.240 60.490 127.410 ;
        RECT 60.320 126.880 60.490 127.050 ;
        RECT 60.320 126.520 60.490 126.690 ;
        RECT 60.320 126.160 60.490 126.330 ;
        RECT 60.320 125.800 60.490 125.970 ;
        RECT 61.990 127.240 62.160 127.410 ;
        RECT 61.990 126.880 62.160 127.050 ;
        RECT 61.990 126.520 62.160 126.690 ;
        RECT 61.990 126.160 62.160 126.330 ;
        RECT 61.990 125.800 62.160 125.970 ;
        RECT 62.540 127.140 62.710 127.310 ;
        RECT 62.540 126.780 62.710 126.950 ;
        RECT 62.540 126.420 62.710 126.590 ;
        RECT 62.540 126.060 62.710 126.230 ;
        RECT 62.540 125.700 62.710 125.870 ;
        RECT 56.180 125.340 56.350 125.510 ;
        RECT 57.385 125.380 57.555 125.550 ;
        RECT 57.745 125.380 57.915 125.550 ;
        RECT 60.975 125.380 61.145 125.550 ;
        RECT 61.335 125.380 61.505 125.550 ;
        RECT 56.180 124.980 56.350 125.150 ;
        RECT 62.540 125.340 62.710 125.510 ;
        RECT 56.180 124.620 56.350 124.790 ;
        RECT 56.180 124.260 56.350 124.430 ;
        RECT 56.180 123.900 56.350 124.070 ;
        RECT 56.180 123.540 56.350 123.710 ;
        RECT 58.400 124.960 58.570 125.130 ;
        RECT 58.400 124.600 58.570 124.770 ;
        RECT 58.400 124.240 58.570 124.410 ;
        RECT 58.400 123.880 58.570 124.050 ;
        RECT 58.400 123.520 58.570 123.690 ;
        RECT 60.320 124.960 60.490 125.130 ;
        RECT 60.320 124.600 60.490 124.770 ;
        RECT 60.320 124.240 60.490 124.410 ;
        RECT 60.320 123.880 60.490 124.050 ;
        RECT 60.320 123.520 60.490 123.690 ;
        RECT 61.990 124.960 62.160 125.130 ;
        RECT 61.990 124.600 62.160 124.770 ;
        RECT 61.990 124.240 62.160 124.410 ;
        RECT 61.990 123.880 62.160 124.050 ;
        RECT 61.990 123.520 62.160 123.690 ;
        RECT 62.540 124.980 62.710 125.150 ;
        RECT 62.540 124.620 62.710 124.790 ;
        RECT 62.540 124.260 62.710 124.430 ;
        RECT 62.540 123.900 62.710 124.070 ;
        RECT 62.540 123.540 62.710 123.710 ;
        RECT 56.180 123.180 56.350 123.350 ;
        RECT 57.385 123.100 57.555 123.270 ;
        RECT 57.745 123.100 57.915 123.270 ;
        RECT 60.975 123.100 61.145 123.270 ;
        RECT 61.335 123.100 61.505 123.270 ;
        RECT 62.540 123.180 62.710 123.350 ;
        RECT 56.180 122.820 56.350 122.990 ;
        RECT 56.180 122.460 56.350 122.630 ;
        RECT 56.180 122.100 56.350 122.270 ;
        RECT 56.180 121.740 56.350 121.910 ;
        RECT 56.180 121.380 56.350 121.550 ;
        RECT 58.400 122.680 58.570 122.850 ;
        RECT 58.400 122.320 58.570 122.490 ;
        RECT 58.400 121.960 58.570 122.130 ;
        RECT 58.400 121.600 58.570 121.770 ;
        RECT 58.400 121.240 58.570 121.410 ;
        RECT 60.320 122.680 60.490 122.850 ;
        RECT 60.320 122.320 60.490 122.490 ;
        RECT 60.320 121.960 60.490 122.130 ;
        RECT 60.320 121.600 60.490 121.770 ;
        RECT 60.320 121.240 60.490 121.410 ;
        RECT 61.990 122.680 62.160 122.850 ;
        RECT 61.990 122.320 62.160 122.490 ;
        RECT 61.990 121.960 62.160 122.130 ;
        RECT 61.990 121.600 62.160 121.770 ;
        RECT 61.990 121.240 62.160 121.410 ;
        RECT 62.540 122.820 62.710 122.990 ;
        RECT 62.540 122.460 62.710 122.630 ;
        RECT 62.540 122.100 62.710 122.270 ;
        RECT 62.540 121.740 62.710 121.910 ;
        RECT 62.540 121.380 62.710 121.550 ;
        RECT 56.180 121.020 56.350 121.190 ;
        RECT 62.540 121.020 62.710 121.190 ;
        RECT 56.180 120.660 56.350 120.830 ;
        RECT 57.385 120.820 57.555 120.990 ;
        RECT 57.745 120.820 57.915 120.990 ;
        RECT 60.975 120.820 61.145 120.990 ;
        RECT 61.335 120.820 61.505 120.990 ;
        RECT 62.540 120.660 62.710 120.830 ;
        RECT 56.180 120.300 56.350 120.470 ;
        RECT 56.180 119.940 56.350 120.110 ;
        RECT 56.180 119.580 56.350 119.750 ;
        RECT 56.180 119.220 56.350 119.390 ;
        RECT 56.180 118.860 56.350 119.030 ;
        RECT 58.400 120.400 58.570 120.570 ;
        RECT 58.400 120.040 58.570 120.210 ;
        RECT 58.400 119.680 58.570 119.850 ;
        RECT 58.400 119.320 58.570 119.490 ;
        RECT 58.400 118.960 58.570 119.130 ;
        RECT 60.320 120.400 60.490 120.570 ;
        RECT 60.320 120.040 60.490 120.210 ;
        RECT 60.320 119.680 60.490 119.850 ;
        RECT 60.320 119.320 60.490 119.490 ;
        RECT 60.320 118.960 60.490 119.130 ;
        RECT 61.990 120.400 62.160 120.570 ;
        RECT 61.990 120.040 62.160 120.210 ;
        RECT 61.990 119.680 62.160 119.850 ;
        RECT 61.990 119.320 62.160 119.490 ;
        RECT 61.990 118.960 62.160 119.130 ;
        RECT 62.540 120.300 62.710 120.470 ;
        RECT 62.540 119.940 62.710 120.110 ;
        RECT 62.540 119.580 62.710 119.750 ;
        RECT 62.540 119.220 62.710 119.390 ;
        RECT 62.540 118.860 62.710 119.030 ;
        RECT 56.180 118.500 56.350 118.670 ;
        RECT 57.385 118.540 57.555 118.710 ;
        RECT 57.745 118.540 57.915 118.710 ;
        RECT 60.975 118.540 61.145 118.710 ;
        RECT 61.335 118.540 61.505 118.710 ;
        RECT 56.180 118.140 56.350 118.310 ;
        RECT 62.540 118.500 62.710 118.670 ;
        RECT 56.180 117.780 56.350 117.950 ;
        RECT 56.180 117.420 56.350 117.590 ;
        RECT 56.180 117.060 56.350 117.230 ;
        RECT 56.180 116.700 56.350 116.870 ;
        RECT 58.400 118.120 58.570 118.290 ;
        RECT 58.400 117.760 58.570 117.930 ;
        RECT 58.400 117.400 58.570 117.570 ;
        RECT 58.400 117.040 58.570 117.210 ;
        RECT 58.400 116.680 58.570 116.850 ;
        RECT 60.320 118.120 60.490 118.290 ;
        RECT 60.320 117.760 60.490 117.930 ;
        RECT 60.320 117.400 60.490 117.570 ;
        RECT 60.320 117.040 60.490 117.210 ;
        RECT 60.320 116.680 60.490 116.850 ;
        RECT 61.990 118.120 62.160 118.290 ;
        RECT 61.990 117.760 62.160 117.930 ;
        RECT 61.990 117.400 62.160 117.570 ;
        RECT 61.990 117.040 62.160 117.210 ;
        RECT 61.990 116.680 62.160 116.850 ;
        RECT 62.540 118.140 62.710 118.310 ;
        RECT 62.540 117.780 62.710 117.950 ;
        RECT 62.540 117.420 62.710 117.590 ;
        RECT 64.965 138.040 65.135 138.210 ;
        RECT 65.325 138.040 65.495 138.210 ;
        RECT 65.685 138.040 65.855 138.210 ;
        RECT 66.045 138.040 66.215 138.210 ;
        RECT 66.405 138.040 66.575 138.210 ;
        RECT 64.435 137.690 64.605 137.860 ;
        RECT 66.705 137.690 66.875 137.860 ;
        RECT 64.435 137.330 64.605 137.500 ;
        RECT 65.570 137.370 65.740 137.540 ;
        RECT 66.705 137.330 66.875 137.500 ;
        RECT 64.435 136.970 64.605 137.140 ;
        RECT 64.435 136.610 64.605 136.780 ;
        RECT 64.435 136.250 64.605 136.420 ;
        RECT 64.435 135.890 64.605 136.060 ;
        RECT 64.435 135.530 64.605 135.700 ;
        RECT 64.435 135.170 64.605 135.340 ;
        RECT 64.985 136.985 65.155 137.155 ;
        RECT 64.985 136.625 65.155 136.795 ;
        RECT 64.985 136.265 65.155 136.435 ;
        RECT 66.155 136.985 66.325 137.155 ;
        RECT 66.155 136.625 66.325 136.795 ;
        RECT 66.155 136.265 66.325 136.435 ;
        RECT 65.570 136.090 65.740 136.260 ;
        RECT 64.985 135.905 65.155 136.075 ;
        RECT 64.985 135.545 65.155 135.715 ;
        RECT 64.985 135.185 65.155 135.355 ;
        RECT 66.155 135.905 66.325 136.075 ;
        RECT 66.155 135.545 66.325 135.715 ;
        RECT 66.155 135.185 66.325 135.355 ;
        RECT 66.705 136.970 66.875 137.140 ;
        RECT 66.705 136.610 66.875 136.780 ;
        RECT 66.705 136.250 66.875 136.420 ;
        RECT 66.705 135.890 66.875 136.060 ;
        RECT 66.705 135.530 66.875 135.700 ;
        RECT 66.705 135.170 66.875 135.340 ;
        RECT 64.435 134.810 64.605 134.980 ;
        RECT 65.570 134.810 65.740 134.980 ;
        RECT 66.705 134.810 66.875 134.980 ;
        RECT 64.435 134.450 64.605 134.620 ;
        RECT 64.435 134.090 64.605 134.260 ;
        RECT 64.435 133.730 64.605 133.900 ;
        RECT 64.435 133.370 64.605 133.540 ;
        RECT 64.435 133.010 64.605 133.180 ;
        RECT 64.985 134.390 65.155 134.560 ;
        RECT 64.985 134.030 65.155 134.200 ;
        RECT 64.985 133.670 65.155 133.840 ;
        RECT 64.985 133.310 65.155 133.480 ;
        RECT 64.985 132.950 65.155 133.120 ;
        RECT 66.155 134.390 66.325 134.560 ;
        RECT 66.155 134.030 66.325 134.200 ;
        RECT 66.155 133.670 66.325 133.840 ;
        RECT 66.155 133.310 66.325 133.480 ;
        RECT 66.155 132.950 66.325 133.120 ;
        RECT 66.705 134.450 66.875 134.620 ;
        RECT 66.705 134.090 66.875 134.260 ;
        RECT 66.705 133.730 66.875 133.900 ;
        RECT 66.705 133.370 66.875 133.540 ;
        RECT 66.705 133.010 66.875 133.180 ;
        RECT 64.435 132.650 64.605 132.820 ;
        RECT 65.570 132.530 65.740 132.700 ;
        RECT 66.705 132.650 66.875 132.820 ;
        RECT 64.435 132.290 64.605 132.460 ;
        RECT 66.705 132.290 66.875 132.460 ;
        RECT 64.435 131.930 64.605 132.100 ;
        RECT 64.435 131.570 64.605 131.740 ;
        RECT 64.435 131.210 64.605 131.380 ;
        RECT 64.435 130.850 64.605 131.020 ;
        RECT 64.985 132.110 65.155 132.280 ;
        RECT 64.985 131.750 65.155 131.920 ;
        RECT 64.985 131.390 65.155 131.560 ;
        RECT 64.985 131.030 65.155 131.200 ;
        RECT 64.985 130.670 65.155 130.840 ;
        RECT 66.155 132.110 66.325 132.280 ;
        RECT 66.155 131.750 66.325 131.920 ;
        RECT 66.155 131.390 66.325 131.560 ;
        RECT 66.155 131.030 66.325 131.200 ;
        RECT 66.155 130.670 66.325 130.840 ;
        RECT 66.705 131.930 66.875 132.100 ;
        RECT 66.705 131.570 66.875 131.740 ;
        RECT 66.705 131.210 66.875 131.380 ;
        RECT 66.705 130.850 66.875 131.020 ;
        RECT 64.435 130.490 64.605 130.660 ;
        RECT 66.705 130.490 66.875 130.660 ;
        RECT 64.435 130.130 64.605 130.300 ;
        RECT 65.570 130.250 65.740 130.420 ;
        RECT 66.705 130.130 66.875 130.300 ;
        RECT 64.435 129.770 64.605 129.940 ;
        RECT 64.435 129.410 64.605 129.580 ;
        RECT 64.435 129.050 64.605 129.220 ;
        RECT 64.435 128.690 64.605 128.860 ;
        RECT 64.435 128.330 64.605 128.500 ;
        RECT 64.435 127.970 64.605 128.140 ;
        RECT 64.985 129.865 65.155 130.035 ;
        RECT 64.985 129.505 65.155 129.675 ;
        RECT 64.985 129.145 65.155 129.315 ;
        RECT 66.155 129.865 66.325 130.035 ;
        RECT 66.155 129.505 66.325 129.675 ;
        RECT 66.155 129.145 66.325 129.315 ;
        RECT 65.570 128.970 65.740 129.140 ;
        RECT 64.985 128.785 65.155 128.955 ;
        RECT 64.985 128.425 65.155 128.595 ;
        RECT 64.985 128.065 65.155 128.235 ;
        RECT 66.155 128.785 66.325 128.955 ;
        RECT 66.155 128.425 66.325 128.595 ;
        RECT 66.155 128.065 66.325 128.235 ;
        RECT 66.705 129.770 66.875 129.940 ;
        RECT 66.705 129.410 66.875 129.580 ;
        RECT 66.705 129.050 66.875 129.220 ;
        RECT 66.705 128.690 66.875 128.860 ;
        RECT 66.705 128.330 66.875 128.500 ;
        RECT 66.705 127.970 66.875 128.140 ;
        RECT 64.435 127.610 64.605 127.780 ;
        RECT 65.570 127.690 65.740 127.860 ;
        RECT 66.705 127.610 66.875 127.780 ;
        RECT 64.435 127.250 64.605 127.420 ;
        RECT 64.435 126.890 64.605 127.060 ;
        RECT 64.435 126.530 64.605 126.700 ;
        RECT 64.435 126.170 64.605 126.340 ;
        RECT 64.435 125.810 64.605 125.980 ;
        RECT 64.435 125.450 64.605 125.620 ;
        RECT 64.985 127.305 65.155 127.475 ;
        RECT 64.985 126.945 65.155 127.115 ;
        RECT 64.985 126.585 65.155 126.755 ;
        RECT 66.155 127.305 66.325 127.475 ;
        RECT 66.155 126.945 66.325 127.115 ;
        RECT 66.155 126.585 66.325 126.755 ;
        RECT 65.570 126.410 65.740 126.580 ;
        RECT 64.985 126.225 65.155 126.395 ;
        RECT 64.985 125.865 65.155 126.035 ;
        RECT 64.985 125.505 65.155 125.675 ;
        RECT 66.155 126.225 66.325 126.395 ;
        RECT 66.155 125.865 66.325 126.035 ;
        RECT 66.155 125.505 66.325 125.675 ;
        RECT 66.705 127.250 66.875 127.420 ;
        RECT 66.705 126.890 66.875 127.060 ;
        RECT 66.705 126.530 66.875 126.700 ;
        RECT 66.705 126.170 66.875 126.340 ;
        RECT 66.705 125.810 66.875 125.980 ;
        RECT 66.705 125.450 66.875 125.620 ;
        RECT 64.435 125.090 64.605 125.260 ;
        RECT 65.570 125.130 65.740 125.300 ;
        RECT 64.435 124.730 64.605 124.900 ;
        RECT 66.705 125.090 66.875 125.260 ;
        RECT 64.435 124.370 64.605 124.540 ;
        RECT 64.435 124.010 64.605 124.180 ;
        RECT 64.435 123.650 64.605 123.820 ;
        RECT 64.435 123.290 64.605 123.460 ;
        RECT 64.985 124.710 65.155 124.880 ;
        RECT 64.985 124.350 65.155 124.520 ;
        RECT 64.985 123.990 65.155 124.160 ;
        RECT 64.985 123.630 65.155 123.800 ;
        RECT 64.985 123.270 65.155 123.440 ;
        RECT 66.705 124.730 66.875 124.900 ;
        RECT 66.705 124.370 66.875 124.540 ;
        RECT 66.705 124.010 66.875 124.180 ;
        RECT 66.705 123.650 66.875 123.820 ;
        RECT 66.705 123.290 66.875 123.460 ;
        RECT 64.435 122.930 64.605 123.100 ;
        RECT 65.570 122.850 65.740 123.020 ;
        RECT 66.705 122.930 66.875 123.100 ;
        RECT 64.435 122.570 64.605 122.740 ;
        RECT 64.435 122.210 64.605 122.380 ;
        RECT 64.435 121.850 64.605 122.020 ;
        RECT 64.435 121.490 64.605 121.660 ;
        RECT 64.435 121.130 64.605 121.300 ;
        RECT 64.985 122.430 65.155 122.600 ;
        RECT 64.985 122.070 65.155 122.240 ;
        RECT 64.985 121.710 65.155 121.880 ;
        RECT 64.985 121.350 65.155 121.520 ;
        RECT 64.985 120.990 65.155 121.160 ;
        RECT 66.705 122.570 66.875 122.740 ;
        RECT 66.705 122.210 66.875 122.380 ;
        RECT 66.705 121.850 66.875 122.020 ;
        RECT 66.705 121.490 66.875 121.660 ;
        RECT 66.705 121.130 66.875 121.300 ;
        RECT 64.435 120.770 64.605 120.940 ;
        RECT 66.705 120.770 66.875 120.940 ;
        RECT 64.435 120.410 64.605 120.580 ;
        RECT 65.570 120.570 65.740 120.740 ;
        RECT 66.705 120.410 66.875 120.580 ;
        RECT 64.435 120.050 64.605 120.220 ;
        RECT 64.435 119.690 64.605 119.860 ;
        RECT 64.435 119.330 64.605 119.500 ;
        RECT 64.435 118.970 64.605 119.140 ;
        RECT 64.435 118.610 64.605 118.780 ;
        RECT 64.435 118.250 64.605 118.420 ;
        RECT 64.985 120.185 65.155 120.355 ;
        RECT 64.985 119.825 65.155 119.995 ;
        RECT 64.985 119.465 65.155 119.635 ;
        RECT 66.155 120.185 66.325 120.355 ;
        RECT 66.155 119.825 66.325 119.995 ;
        RECT 66.155 119.465 66.325 119.635 ;
        RECT 65.570 119.290 65.740 119.460 ;
        RECT 64.985 119.105 65.155 119.275 ;
        RECT 64.985 118.745 65.155 118.915 ;
        RECT 64.985 118.385 65.155 118.555 ;
        RECT 66.155 119.105 66.325 119.275 ;
        RECT 66.155 118.745 66.325 118.915 ;
        RECT 66.155 118.385 66.325 118.555 ;
        RECT 66.705 120.050 66.875 120.220 ;
        RECT 66.705 119.690 66.875 119.860 ;
        RECT 66.705 119.330 66.875 119.500 ;
        RECT 66.705 118.970 66.875 119.140 ;
        RECT 66.705 118.610 66.875 118.780 ;
        RECT 66.705 118.250 66.875 118.420 ;
        RECT 64.435 117.890 64.605 118.060 ;
        RECT 65.570 118.010 65.740 118.180 ;
        RECT 66.705 117.890 66.875 118.060 ;
        RECT 64.965 117.340 65.135 117.510 ;
        RECT 65.325 117.340 65.495 117.510 ;
        RECT 65.685 117.340 65.855 117.510 ;
        RECT 66.045 117.340 66.215 117.510 ;
        RECT 66.405 117.340 66.575 117.510 ;
        RECT 68.500 138.040 68.670 138.210 ;
        RECT 68.860 138.040 69.030 138.210 ;
        RECT 69.220 138.040 69.390 138.210 ;
        RECT 69.580 138.040 69.750 138.210 ;
        RECT 69.940 138.040 70.110 138.210 ;
        RECT 70.300 138.040 70.470 138.210 ;
        RECT 70.660 138.040 70.830 138.210 ;
        RECT 68.190 137.690 68.360 137.860 ;
        RECT 70.960 137.690 71.130 137.860 ;
        RECT 68.190 137.330 68.360 137.500 ;
        RECT 69.395 137.370 69.565 137.540 ;
        RECT 69.755 137.370 69.925 137.540 ;
        RECT 70.960 137.330 71.130 137.500 ;
        RECT 68.190 136.970 68.360 137.140 ;
        RECT 68.190 136.610 68.360 136.780 ;
        RECT 68.190 136.250 68.360 136.420 ;
        RECT 68.190 135.890 68.360 136.060 ;
        RECT 68.190 135.530 68.360 135.700 ;
        RECT 68.190 135.170 68.360 135.340 ;
        RECT 68.740 136.985 68.910 137.155 ;
        RECT 68.740 136.625 68.910 136.795 ;
        RECT 68.740 136.265 68.910 136.435 ;
        RECT 70.410 136.985 70.580 137.155 ;
        RECT 70.410 136.625 70.580 136.795 ;
        RECT 70.410 136.265 70.580 136.435 ;
        RECT 69.395 136.090 69.565 136.260 ;
        RECT 69.755 136.090 69.925 136.260 ;
        RECT 68.740 135.905 68.910 136.075 ;
        RECT 68.740 135.545 68.910 135.715 ;
        RECT 68.740 135.185 68.910 135.355 ;
        RECT 70.410 135.905 70.580 136.075 ;
        RECT 70.410 135.545 70.580 135.715 ;
        RECT 70.410 135.185 70.580 135.355 ;
        RECT 70.960 136.970 71.130 137.140 ;
        RECT 70.960 136.610 71.130 136.780 ;
        RECT 70.960 136.250 71.130 136.420 ;
        RECT 70.960 135.890 71.130 136.060 ;
        RECT 70.960 135.530 71.130 135.700 ;
        RECT 70.960 135.170 71.130 135.340 ;
        RECT 68.190 134.810 68.360 134.980 ;
        RECT 69.395 134.810 69.565 134.980 ;
        RECT 69.755 134.810 69.925 134.980 ;
        RECT 70.960 134.810 71.130 134.980 ;
        RECT 68.190 134.450 68.360 134.620 ;
        RECT 68.190 134.090 68.360 134.260 ;
        RECT 68.190 133.730 68.360 133.900 ;
        RECT 68.190 133.370 68.360 133.540 ;
        RECT 68.190 133.010 68.360 133.180 ;
        RECT 68.740 134.390 68.910 134.560 ;
        RECT 68.740 134.030 68.910 134.200 ;
        RECT 68.740 133.670 68.910 133.840 ;
        RECT 68.740 133.310 68.910 133.480 ;
        RECT 68.740 132.950 68.910 133.120 ;
        RECT 70.410 134.390 70.580 134.560 ;
        RECT 70.410 134.030 70.580 134.200 ;
        RECT 70.410 133.670 70.580 133.840 ;
        RECT 70.410 133.310 70.580 133.480 ;
        RECT 70.410 132.950 70.580 133.120 ;
        RECT 70.960 134.450 71.130 134.620 ;
        RECT 70.960 134.090 71.130 134.260 ;
        RECT 70.960 133.730 71.130 133.900 ;
        RECT 70.960 133.370 71.130 133.540 ;
        RECT 70.960 133.010 71.130 133.180 ;
        RECT 68.190 132.650 68.360 132.820 ;
        RECT 69.395 132.530 69.565 132.700 ;
        RECT 69.755 132.530 69.925 132.700 ;
        RECT 70.960 132.650 71.130 132.820 ;
        RECT 68.190 132.290 68.360 132.460 ;
        RECT 70.960 132.290 71.130 132.460 ;
        RECT 68.190 131.930 68.360 132.100 ;
        RECT 68.190 131.570 68.360 131.740 ;
        RECT 68.190 131.210 68.360 131.380 ;
        RECT 68.190 130.850 68.360 131.020 ;
        RECT 68.740 132.110 68.910 132.280 ;
        RECT 68.740 131.750 68.910 131.920 ;
        RECT 68.740 131.390 68.910 131.560 ;
        RECT 68.740 131.030 68.910 131.200 ;
        RECT 68.740 130.670 68.910 130.840 ;
        RECT 70.410 132.110 70.580 132.280 ;
        RECT 70.410 131.750 70.580 131.920 ;
        RECT 70.410 131.390 70.580 131.560 ;
        RECT 70.410 131.030 70.580 131.200 ;
        RECT 70.410 130.670 70.580 130.840 ;
        RECT 70.960 131.930 71.130 132.100 ;
        RECT 70.960 131.570 71.130 131.740 ;
        RECT 70.960 131.210 71.130 131.380 ;
        RECT 70.960 130.850 71.130 131.020 ;
        RECT 68.190 130.490 68.360 130.660 ;
        RECT 70.960 130.490 71.130 130.660 ;
        RECT 68.190 130.130 68.360 130.300 ;
        RECT 69.395 130.250 69.565 130.420 ;
        RECT 69.755 130.250 69.925 130.420 ;
        RECT 70.960 130.130 71.130 130.300 ;
        RECT 68.190 129.770 68.360 129.940 ;
        RECT 68.190 129.410 68.360 129.580 ;
        RECT 68.190 129.050 68.360 129.220 ;
        RECT 68.190 128.690 68.360 128.860 ;
        RECT 68.190 128.330 68.360 128.500 ;
        RECT 68.190 127.970 68.360 128.140 ;
        RECT 68.740 129.865 68.910 130.035 ;
        RECT 68.740 129.505 68.910 129.675 ;
        RECT 68.740 129.145 68.910 129.315 ;
        RECT 70.410 129.865 70.580 130.035 ;
        RECT 70.410 129.505 70.580 129.675 ;
        RECT 70.410 129.145 70.580 129.315 ;
        RECT 69.395 128.970 69.565 129.140 ;
        RECT 69.755 128.970 69.925 129.140 ;
        RECT 68.740 128.785 68.910 128.955 ;
        RECT 68.740 128.425 68.910 128.595 ;
        RECT 68.740 128.065 68.910 128.235 ;
        RECT 70.410 128.785 70.580 128.955 ;
        RECT 70.410 128.425 70.580 128.595 ;
        RECT 70.410 128.065 70.580 128.235 ;
        RECT 70.960 129.770 71.130 129.940 ;
        RECT 70.960 129.410 71.130 129.580 ;
        RECT 70.960 129.050 71.130 129.220 ;
        RECT 70.960 128.690 71.130 128.860 ;
        RECT 70.960 128.330 71.130 128.500 ;
        RECT 70.960 127.970 71.130 128.140 ;
        RECT 68.190 127.610 68.360 127.780 ;
        RECT 69.395 127.690 69.565 127.860 ;
        RECT 69.755 127.690 69.925 127.860 ;
        RECT 70.960 127.610 71.130 127.780 ;
        RECT 68.190 127.250 68.360 127.420 ;
        RECT 68.190 126.890 68.360 127.060 ;
        RECT 68.190 126.530 68.360 126.700 ;
        RECT 68.190 126.170 68.360 126.340 ;
        RECT 68.190 125.810 68.360 125.980 ;
        RECT 68.190 125.450 68.360 125.620 ;
        RECT 68.740 127.305 68.910 127.475 ;
        RECT 68.740 126.945 68.910 127.115 ;
        RECT 68.740 126.585 68.910 126.755 ;
        RECT 70.410 127.305 70.580 127.475 ;
        RECT 70.410 126.945 70.580 127.115 ;
        RECT 70.410 126.585 70.580 126.755 ;
        RECT 69.395 126.410 69.565 126.580 ;
        RECT 69.755 126.410 69.925 126.580 ;
        RECT 68.740 126.225 68.910 126.395 ;
        RECT 68.740 125.865 68.910 126.035 ;
        RECT 68.740 125.505 68.910 125.675 ;
        RECT 70.410 126.225 70.580 126.395 ;
        RECT 70.410 125.865 70.580 126.035 ;
        RECT 70.410 125.505 70.580 125.675 ;
        RECT 70.960 127.250 71.130 127.420 ;
        RECT 70.960 126.890 71.130 127.060 ;
        RECT 70.960 126.530 71.130 126.700 ;
        RECT 70.960 126.170 71.130 126.340 ;
        RECT 70.960 125.810 71.130 125.980 ;
        RECT 70.960 125.450 71.130 125.620 ;
        RECT 68.190 125.090 68.360 125.260 ;
        RECT 69.395 125.130 69.565 125.300 ;
        RECT 69.755 125.130 69.925 125.300 ;
        RECT 68.190 124.730 68.360 124.900 ;
        RECT 70.960 125.090 71.130 125.260 ;
        RECT 68.190 124.370 68.360 124.540 ;
        RECT 68.190 124.010 68.360 124.180 ;
        RECT 68.190 123.650 68.360 123.820 ;
        RECT 68.190 123.290 68.360 123.460 ;
        RECT 70.410 124.710 70.580 124.880 ;
        RECT 70.410 124.350 70.580 124.520 ;
        RECT 70.410 123.990 70.580 124.160 ;
        RECT 70.410 123.630 70.580 123.800 ;
        RECT 70.410 123.270 70.580 123.440 ;
        RECT 70.960 124.730 71.130 124.900 ;
        RECT 70.960 124.370 71.130 124.540 ;
        RECT 70.960 124.010 71.130 124.180 ;
        RECT 70.960 123.650 71.130 123.820 ;
        RECT 70.960 123.290 71.130 123.460 ;
        RECT 68.190 122.930 68.360 123.100 ;
        RECT 69.395 122.850 69.565 123.020 ;
        RECT 69.755 122.850 69.925 123.020 ;
        RECT 70.960 122.930 71.130 123.100 ;
        RECT 68.190 122.570 68.360 122.740 ;
        RECT 68.190 122.210 68.360 122.380 ;
        RECT 68.190 121.850 68.360 122.020 ;
        RECT 68.190 121.490 68.360 121.660 ;
        RECT 68.190 121.130 68.360 121.300 ;
        RECT 70.410 122.430 70.580 122.600 ;
        RECT 70.410 122.070 70.580 122.240 ;
        RECT 70.410 121.710 70.580 121.880 ;
        RECT 70.410 121.350 70.580 121.520 ;
        RECT 70.410 120.990 70.580 121.160 ;
        RECT 70.960 122.570 71.130 122.740 ;
        RECT 70.960 122.210 71.130 122.380 ;
        RECT 70.960 121.850 71.130 122.020 ;
        RECT 70.960 121.490 71.130 121.660 ;
        RECT 70.960 121.130 71.130 121.300 ;
        RECT 68.190 120.770 68.360 120.940 ;
        RECT 70.960 120.770 71.130 120.940 ;
        RECT 68.190 120.410 68.360 120.580 ;
        RECT 69.395 120.570 69.565 120.740 ;
        RECT 69.755 120.570 69.925 120.740 ;
        RECT 70.960 120.410 71.130 120.580 ;
        RECT 68.190 120.050 68.360 120.220 ;
        RECT 68.190 119.690 68.360 119.860 ;
        RECT 68.190 119.330 68.360 119.500 ;
        RECT 68.190 118.970 68.360 119.140 ;
        RECT 68.190 118.610 68.360 118.780 ;
        RECT 68.190 118.250 68.360 118.420 ;
        RECT 68.740 120.185 68.910 120.355 ;
        RECT 68.740 119.825 68.910 119.995 ;
        RECT 68.740 119.465 68.910 119.635 ;
        RECT 70.410 120.185 70.580 120.355 ;
        RECT 70.410 119.825 70.580 119.995 ;
        RECT 70.410 119.465 70.580 119.635 ;
        RECT 69.395 119.290 69.565 119.460 ;
        RECT 69.755 119.290 69.925 119.460 ;
        RECT 68.740 119.105 68.910 119.275 ;
        RECT 68.740 118.745 68.910 118.915 ;
        RECT 68.740 118.385 68.910 118.555 ;
        RECT 70.410 119.105 70.580 119.275 ;
        RECT 70.410 118.745 70.580 118.915 ;
        RECT 70.410 118.385 70.580 118.555 ;
        RECT 70.960 120.050 71.130 120.220 ;
        RECT 70.960 119.690 71.130 119.860 ;
        RECT 70.960 119.330 71.130 119.500 ;
        RECT 70.960 118.970 71.130 119.140 ;
        RECT 70.960 118.610 71.130 118.780 ;
        RECT 70.960 118.250 71.130 118.420 ;
        RECT 68.190 117.890 68.360 118.060 ;
        RECT 69.395 118.010 69.565 118.180 ;
        RECT 69.755 118.010 69.925 118.180 ;
        RECT 70.960 117.890 71.130 118.060 ;
        RECT 68.500 117.340 68.670 117.510 ;
        RECT 68.860 117.340 69.030 117.510 ;
        RECT 69.220 117.340 69.390 117.510 ;
        RECT 69.580 117.340 69.750 117.510 ;
        RECT 69.940 117.340 70.110 117.510 ;
        RECT 70.300 117.340 70.470 117.510 ;
        RECT 70.660 117.340 70.830 117.510 ;
        RECT 72.590 137.860 72.760 138.030 ;
        RECT 72.590 137.500 72.760 137.670 ;
        RECT 73.140 138.920 73.310 139.090 ;
        RECT 73.140 138.560 73.310 138.730 ;
        RECT 73.140 138.200 73.310 138.370 ;
        RECT 73.140 137.840 73.310 138.010 ;
        RECT 73.140 137.480 73.310 137.650 ;
        RECT 74.310 138.920 74.480 139.090 ;
        RECT 74.310 138.560 74.480 138.730 ;
        RECT 75.880 138.955 76.050 139.125 ;
        RECT 75.880 138.595 76.050 138.765 ;
        RECT 77.050 141.115 77.220 141.285 ;
        RECT 77.050 140.755 77.220 140.925 ;
        RECT 77.050 140.395 77.220 140.565 ;
        RECT 77.050 140.035 77.220 140.205 ;
        RECT 77.050 139.675 77.220 139.845 ;
        RECT 77.050 139.315 77.220 139.485 ;
        RECT 77.050 138.955 77.220 139.125 ;
        RECT 77.050 138.595 77.220 138.765 ;
        RECT 77.600 141.100 77.770 141.270 ;
        RECT 77.600 140.740 77.770 140.910 ;
        RECT 77.600 140.380 77.770 140.550 ;
        RECT 77.600 140.020 77.770 140.190 ;
        RECT 77.600 139.660 77.770 139.830 ;
        RECT 77.600 139.300 77.770 139.470 ;
        RECT 77.600 138.940 77.770 139.110 ;
        RECT 77.600 138.580 77.770 138.750 ;
        RECT 74.310 138.200 74.480 138.370 ;
        RECT 76.465 138.220 76.635 138.390 ;
        RECT 77.600 138.220 77.770 138.390 ;
        RECT 74.310 137.840 74.480 138.010 ;
        RECT 74.310 137.480 74.480 137.650 ;
        RECT 75.880 137.835 76.050 138.005 ;
        RECT 72.590 137.140 72.760 137.310 ;
        RECT 75.880 137.475 76.050 137.645 ;
        RECT 73.725 137.060 73.895 137.230 ;
        RECT 75.880 137.115 76.050 137.285 ;
        RECT 72.590 136.780 72.760 136.950 ;
        RECT 72.590 136.420 72.760 136.590 ;
        RECT 72.590 136.060 72.760 136.230 ;
        RECT 72.590 135.700 72.760 135.870 ;
        RECT 72.590 135.340 72.760 135.510 ;
        RECT 73.140 136.640 73.310 136.810 ;
        RECT 73.140 136.280 73.310 136.450 ;
        RECT 73.140 135.920 73.310 136.090 ;
        RECT 73.140 135.560 73.310 135.730 ;
        RECT 73.140 135.200 73.310 135.370 ;
        RECT 74.310 136.640 74.480 136.810 ;
        RECT 74.310 136.280 74.480 136.450 ;
        RECT 74.310 135.920 74.480 136.090 ;
        RECT 74.310 135.560 74.480 135.730 ;
        RECT 74.310 135.200 74.480 135.370 ;
        RECT 75.880 136.755 76.050 136.925 ;
        RECT 75.880 136.395 76.050 136.565 ;
        RECT 75.880 136.035 76.050 136.205 ;
        RECT 75.880 135.675 76.050 135.845 ;
        RECT 75.880 135.315 76.050 135.485 ;
        RECT 77.050 137.835 77.220 138.005 ;
        RECT 77.050 137.475 77.220 137.645 ;
        RECT 77.050 137.115 77.220 137.285 ;
        RECT 77.050 136.755 77.220 136.925 ;
        RECT 77.050 136.395 77.220 136.565 ;
        RECT 77.050 136.035 77.220 136.205 ;
        RECT 77.050 135.675 77.220 135.845 ;
        RECT 77.050 135.315 77.220 135.485 ;
        RECT 77.600 137.860 77.770 138.030 ;
        RECT 77.600 137.500 77.770 137.670 ;
        RECT 77.600 137.140 77.770 137.310 ;
        RECT 77.600 136.780 77.770 136.950 ;
        RECT 77.600 136.420 77.770 136.590 ;
        RECT 77.600 136.060 77.770 136.230 ;
        RECT 77.600 135.700 77.770 135.870 ;
        RECT 77.600 135.340 77.770 135.510 ;
        RECT 72.590 134.980 72.760 135.150 ;
        RECT 72.590 134.620 72.760 134.790 ;
        RECT 73.725 134.780 73.895 134.950 ;
        RECT 76.465 134.940 76.635 135.110 ;
        RECT 77.600 134.980 77.770 135.150 ;
        RECT 77.050 134.540 77.220 134.710 ;
        RECT 72.590 134.260 72.760 134.430 ;
        RECT 72.590 133.900 72.760 134.070 ;
        RECT 72.590 133.540 72.760 133.710 ;
        RECT 72.590 133.180 72.760 133.350 ;
        RECT 72.590 132.820 72.760 132.990 ;
        RECT 73.140 134.360 73.310 134.530 ;
        RECT 73.140 134.000 73.310 134.170 ;
        RECT 73.140 133.640 73.310 133.810 ;
        RECT 73.140 133.280 73.310 133.450 ;
        RECT 73.140 132.920 73.310 133.090 ;
        RECT 74.310 134.360 74.480 134.530 ;
        RECT 74.310 134.000 74.480 134.170 ;
        RECT 74.310 133.640 74.480 133.810 ;
        RECT 74.310 133.280 74.480 133.450 ;
        RECT 74.310 132.920 74.480 133.090 ;
        RECT 77.050 134.180 77.220 134.350 ;
        RECT 77.050 133.820 77.220 133.990 ;
        RECT 77.050 133.460 77.220 133.630 ;
        RECT 77.050 133.100 77.220 133.270 ;
        RECT 77.050 132.740 77.220 132.910 ;
        RECT 72.590 132.460 72.760 132.630 ;
        RECT 73.725 132.500 73.895 132.670 ;
        RECT 72.590 132.100 72.760 132.270 ;
        RECT 77.050 132.380 77.220 132.550 ;
        RECT 72.590 131.740 72.760 131.910 ;
        RECT 72.590 131.380 72.760 131.550 ;
        RECT 72.590 131.020 72.760 131.190 ;
        RECT 72.590 130.660 72.760 130.830 ;
        RECT 73.140 132.080 73.310 132.250 ;
        RECT 73.140 131.720 73.310 131.890 ;
        RECT 73.140 131.360 73.310 131.530 ;
        RECT 73.140 131.000 73.310 131.170 ;
        RECT 73.140 130.640 73.310 130.810 ;
        RECT 74.310 132.080 74.480 132.250 ;
        RECT 74.310 131.720 74.480 131.890 ;
        RECT 74.310 131.360 74.480 131.530 ;
        RECT 74.310 131.000 74.480 131.170 ;
        RECT 74.310 130.640 74.480 130.810 ;
        RECT 77.050 132.020 77.220 132.190 ;
        RECT 77.050 131.660 77.220 131.830 ;
        RECT 77.050 131.300 77.220 131.470 ;
        RECT 77.050 130.940 77.220 131.110 ;
        RECT 72.590 130.300 72.760 130.470 ;
        RECT 77.050 130.580 77.220 130.750 ;
        RECT 73.725 130.220 73.895 130.390 ;
        RECT 77.050 130.220 77.220 130.390 ;
        RECT 72.590 129.940 72.760 130.110 ;
        RECT 72.590 129.580 72.760 129.750 ;
        RECT 72.590 129.220 72.760 129.390 ;
        RECT 72.590 128.860 72.760 129.030 ;
        RECT 72.590 128.500 72.760 128.670 ;
        RECT 72.590 128.140 72.760 128.310 ;
        RECT 73.140 129.835 73.310 130.005 ;
        RECT 73.140 129.475 73.310 129.645 ;
        RECT 73.140 129.115 73.310 129.285 ;
        RECT 74.310 129.835 74.480 130.005 ;
        RECT 74.310 129.475 74.480 129.645 ;
        RECT 74.310 129.115 74.480 129.285 ;
        RECT 73.725 128.940 73.895 129.110 ;
        RECT 73.140 128.755 73.310 128.925 ;
        RECT 73.140 128.395 73.310 128.565 ;
        RECT 73.140 128.035 73.310 128.205 ;
        RECT 74.310 128.755 74.480 128.925 ;
        RECT 74.310 128.395 74.480 128.565 ;
        RECT 74.310 128.035 74.480 128.205 ;
        RECT 77.050 129.860 77.220 130.030 ;
        RECT 77.050 129.500 77.220 129.670 ;
        RECT 77.050 129.140 77.220 129.310 ;
        RECT 77.050 128.780 77.220 128.950 ;
        RECT 77.050 128.420 77.220 128.590 ;
        RECT 77.050 128.060 77.220 128.230 ;
        RECT 77.600 134.620 77.770 134.790 ;
        RECT 77.600 134.260 77.770 134.430 ;
        RECT 77.600 133.900 77.770 134.070 ;
        RECT 77.600 133.540 77.770 133.710 ;
        RECT 77.600 133.180 77.770 133.350 ;
        RECT 77.600 132.820 77.770 132.990 ;
        RECT 77.600 132.460 77.770 132.630 ;
        RECT 77.600 132.100 77.770 132.270 ;
        RECT 77.600 131.740 77.770 131.910 ;
        RECT 77.600 131.380 77.770 131.550 ;
        RECT 77.600 131.020 77.770 131.190 ;
        RECT 77.600 130.660 77.770 130.830 ;
        RECT 77.600 130.300 77.770 130.470 ;
        RECT 77.600 129.940 77.770 130.110 ;
        RECT 77.600 129.580 77.770 129.750 ;
        RECT 77.600 129.220 77.770 129.390 ;
        RECT 77.600 128.860 77.770 129.030 ;
        RECT 77.600 128.500 77.770 128.670 ;
        RECT 77.600 128.140 77.770 128.310 ;
        RECT 72.590 127.780 72.760 127.950 ;
        RECT 73.725 127.660 73.895 127.830 ;
        RECT 76.465 127.660 76.635 127.830 ;
        RECT 77.600 127.780 77.770 127.950 ;
        RECT 72.590 127.420 72.760 127.590 ;
        RECT 72.590 127.060 72.760 127.230 ;
        RECT 72.590 126.700 72.760 126.870 ;
        RECT 72.590 126.340 72.760 126.510 ;
        RECT 72.590 125.980 72.760 126.150 ;
        RECT 72.590 125.620 72.760 125.790 ;
        RECT 73.140 127.275 73.310 127.445 ;
        RECT 73.140 126.915 73.310 127.085 ;
        RECT 73.140 126.555 73.310 126.725 ;
        RECT 74.310 127.275 74.480 127.445 ;
        RECT 74.310 126.915 74.480 127.085 ;
        RECT 74.310 126.555 74.480 126.725 ;
        RECT 73.725 126.380 73.895 126.550 ;
        RECT 73.140 126.195 73.310 126.365 ;
        RECT 73.140 125.835 73.310 126.005 ;
        RECT 73.140 125.475 73.310 125.645 ;
        RECT 74.310 126.195 74.480 126.365 ;
        RECT 74.310 125.835 74.480 126.005 ;
        RECT 74.310 125.475 74.480 125.645 ;
        RECT 77.050 127.260 77.220 127.430 ;
        RECT 77.050 126.900 77.220 127.070 ;
        RECT 77.050 126.540 77.220 126.710 ;
        RECT 77.050 126.180 77.220 126.350 ;
        RECT 77.050 125.820 77.220 125.990 ;
        RECT 72.590 125.260 72.760 125.430 ;
        RECT 77.050 125.460 77.220 125.630 ;
        RECT 73.725 125.100 73.895 125.270 ;
        RECT 77.050 125.100 77.220 125.270 ;
        RECT 72.590 124.900 72.760 125.070 ;
        RECT 72.590 124.540 72.760 124.710 ;
        RECT 72.590 124.180 72.760 124.350 ;
        RECT 72.590 123.820 72.760 123.990 ;
        RECT 72.590 123.460 72.760 123.630 ;
        RECT 72.590 123.100 72.760 123.270 ;
        RECT 73.140 124.680 73.310 124.850 ;
        RECT 73.140 124.320 73.310 124.490 ;
        RECT 73.140 123.960 73.310 124.130 ;
        RECT 73.140 123.600 73.310 123.770 ;
        RECT 73.140 123.240 73.310 123.410 ;
        RECT 74.310 124.680 74.480 124.850 ;
        RECT 74.310 124.320 74.480 124.490 ;
        RECT 74.310 123.960 74.480 124.130 ;
        RECT 74.310 123.600 74.480 123.770 ;
        RECT 74.310 123.240 74.480 123.410 ;
        RECT 77.050 124.740 77.220 124.910 ;
        RECT 77.050 124.380 77.220 124.550 ;
        RECT 77.050 124.020 77.220 124.190 ;
        RECT 77.050 123.660 77.220 123.830 ;
        RECT 77.050 123.300 77.220 123.470 ;
        RECT 72.590 122.740 72.760 122.910 ;
        RECT 73.725 122.820 73.895 122.990 ;
        RECT 77.050 122.940 77.220 123.110 ;
        RECT 77.050 122.580 77.220 122.750 ;
        RECT 72.590 122.380 72.760 122.550 ;
        RECT 72.590 122.020 72.760 122.190 ;
        RECT 72.590 121.660 72.760 121.830 ;
        RECT 72.590 121.300 72.760 121.470 ;
        RECT 72.590 120.940 72.760 121.110 ;
        RECT 73.140 122.400 73.310 122.570 ;
        RECT 73.140 122.040 73.310 122.210 ;
        RECT 73.140 121.680 73.310 121.850 ;
        RECT 73.140 121.320 73.310 121.490 ;
        RECT 73.140 120.960 73.310 121.130 ;
        RECT 74.310 122.400 74.480 122.570 ;
        RECT 74.310 122.040 74.480 122.210 ;
        RECT 74.310 121.680 74.480 121.850 ;
        RECT 74.310 121.320 74.480 121.490 ;
        RECT 74.310 120.960 74.480 121.130 ;
        RECT 77.050 122.220 77.220 122.390 ;
        RECT 77.050 121.860 77.220 122.030 ;
        RECT 77.050 121.500 77.220 121.670 ;
        RECT 77.050 121.140 77.220 121.310 ;
        RECT 77.050 120.780 77.220 120.950 ;
        RECT 77.600 127.420 77.770 127.590 ;
        RECT 77.600 127.060 77.770 127.230 ;
        RECT 77.600 126.700 77.770 126.870 ;
        RECT 77.600 126.340 77.770 126.510 ;
        RECT 77.600 125.980 77.770 126.150 ;
        RECT 77.600 125.620 77.770 125.790 ;
        RECT 77.600 125.260 77.770 125.430 ;
        RECT 77.600 124.900 77.770 125.070 ;
        RECT 77.600 124.540 77.770 124.710 ;
        RECT 77.600 124.180 77.770 124.350 ;
        RECT 77.600 123.820 77.770 123.990 ;
        RECT 77.600 123.460 77.770 123.630 ;
        RECT 77.600 123.100 77.770 123.270 ;
        RECT 77.600 122.740 77.770 122.910 ;
        RECT 77.600 122.380 77.770 122.550 ;
        RECT 77.600 122.020 77.770 122.190 ;
        RECT 77.600 121.660 77.770 121.830 ;
        RECT 77.600 121.300 77.770 121.470 ;
        RECT 77.600 120.940 77.770 121.110 ;
        RECT 72.590 120.580 72.760 120.750 ;
        RECT 73.725 120.540 73.895 120.710 ;
        RECT 77.600 120.580 77.770 120.750 ;
        RECT 72.590 120.220 72.760 120.390 ;
        RECT 76.465 120.380 76.635 120.550 ;
        RECT 72.590 119.860 72.760 120.030 ;
        RECT 72.590 119.500 72.760 119.670 ;
        RECT 72.590 119.140 72.760 119.310 ;
        RECT 72.590 118.780 72.760 118.950 ;
        RECT 73.140 120.120 73.310 120.290 ;
        RECT 73.140 119.760 73.310 119.930 ;
        RECT 73.140 119.400 73.310 119.570 ;
        RECT 73.140 119.040 73.310 119.210 ;
        RECT 73.140 118.680 73.310 118.850 ;
        RECT 74.310 120.120 74.480 120.290 ;
        RECT 77.600 120.220 77.770 120.390 ;
        RECT 74.310 119.760 74.480 119.930 ;
        RECT 74.310 119.400 74.480 119.570 ;
        RECT 74.310 119.040 74.480 119.210 ;
        RECT 74.310 118.680 74.480 118.850 ;
        RECT 75.880 119.995 76.050 120.165 ;
        RECT 75.880 119.635 76.050 119.805 ;
        RECT 75.880 119.275 76.050 119.445 ;
        RECT 75.880 118.915 76.050 119.085 ;
        RECT 72.590 118.420 72.760 118.590 ;
        RECT 75.880 118.555 76.050 118.725 ;
        RECT 73.725 118.260 73.895 118.430 ;
        RECT 72.590 118.060 72.760 118.230 ;
        RECT 75.880 118.195 76.050 118.365 ;
        RECT 72.590 117.700 72.760 117.870 ;
        RECT 72.590 117.340 72.760 117.510 ;
        RECT 62.540 117.060 62.710 117.230 ;
        RECT 62.540 116.700 62.710 116.870 ;
        RECT 56.180 116.340 56.350 116.510 ;
        RECT 57.385 116.260 57.555 116.430 ;
        RECT 57.745 116.260 57.915 116.430 ;
        RECT 60.975 116.260 61.145 116.430 ;
        RECT 61.335 116.260 61.505 116.430 ;
        RECT 62.540 116.340 62.710 116.510 ;
        RECT 56.180 115.980 56.350 116.150 ;
        RECT 56.180 115.620 56.350 115.790 ;
        RECT 56.180 115.260 56.350 115.430 ;
        RECT 56.180 114.900 56.350 115.070 ;
        RECT 56.180 114.540 56.350 114.710 ;
        RECT 58.400 115.840 58.570 116.010 ;
        RECT 58.400 115.480 58.570 115.650 ;
        RECT 58.400 115.120 58.570 115.290 ;
        RECT 58.400 114.760 58.570 114.930 ;
        RECT 58.400 114.400 58.570 114.570 ;
        RECT 60.320 115.840 60.490 116.010 ;
        RECT 60.320 115.480 60.490 115.650 ;
        RECT 60.320 115.120 60.490 115.290 ;
        RECT 60.320 114.760 60.490 114.930 ;
        RECT 60.320 114.400 60.490 114.570 ;
        RECT 61.990 115.840 62.160 116.010 ;
        RECT 61.990 115.480 62.160 115.650 ;
        RECT 61.990 115.120 62.160 115.290 ;
        RECT 61.990 114.760 62.160 114.930 ;
        RECT 61.990 114.400 62.160 114.570 ;
        RECT 62.540 115.980 62.710 116.150 ;
        RECT 62.540 115.620 62.710 115.790 ;
        RECT 62.540 115.260 62.710 115.430 ;
        RECT 62.540 114.900 62.710 115.070 ;
        RECT 62.540 114.540 62.710 114.710 ;
        RECT 56.180 114.180 56.350 114.350 ;
        RECT 62.540 114.180 62.710 114.350 ;
        RECT 56.180 113.820 56.350 113.990 ;
        RECT 57.385 113.980 57.555 114.150 ;
        RECT 57.745 113.980 57.915 114.150 ;
        RECT 60.975 113.980 61.145 114.150 ;
        RECT 61.335 113.980 61.505 114.150 ;
        RECT 62.540 113.820 62.710 113.990 ;
        RECT 56.180 113.460 56.350 113.630 ;
        RECT 56.180 113.100 56.350 113.270 ;
        RECT 56.180 112.740 56.350 112.910 ;
        RECT 60.320 113.560 60.490 113.730 ;
        RECT 62.540 113.460 62.710 113.630 ;
        RECT 60.320 113.200 60.490 113.370 ;
        RECT 60.975 113.200 61.145 113.370 ;
        RECT 61.335 113.200 61.505 113.370 ;
        RECT 60.320 112.840 60.490 113.010 ;
        RECT 62.540 113.100 62.710 113.270 ;
        RECT 72.590 116.980 72.760 117.150 ;
        RECT 72.590 116.620 72.760 116.790 ;
        RECT 72.590 116.260 72.760 116.430 ;
        RECT 73.140 117.840 73.310 118.010 ;
        RECT 73.140 117.480 73.310 117.650 ;
        RECT 73.140 117.120 73.310 117.290 ;
        RECT 73.140 116.760 73.310 116.930 ;
        RECT 73.140 116.400 73.310 116.570 ;
        RECT 74.310 117.840 74.480 118.010 ;
        RECT 74.310 117.480 74.480 117.650 ;
        RECT 75.880 117.835 76.050 118.005 ;
        RECT 75.880 117.475 76.050 117.645 ;
        RECT 77.050 119.995 77.220 120.165 ;
        RECT 77.050 119.635 77.220 119.805 ;
        RECT 77.050 119.275 77.220 119.445 ;
        RECT 77.050 118.915 77.220 119.085 ;
        RECT 77.050 118.555 77.220 118.725 ;
        RECT 77.050 118.195 77.220 118.365 ;
        RECT 77.050 117.835 77.220 118.005 ;
        RECT 77.050 117.475 77.220 117.645 ;
        RECT 77.600 119.860 77.770 120.030 ;
        RECT 77.600 119.500 77.770 119.670 ;
        RECT 77.600 119.140 77.770 119.310 ;
        RECT 77.600 118.780 77.770 118.950 ;
        RECT 77.600 118.420 77.770 118.590 ;
        RECT 77.600 118.060 77.770 118.230 ;
        RECT 77.600 117.700 77.770 117.870 ;
        RECT 74.310 117.120 74.480 117.290 ;
        RECT 77.600 117.340 77.770 117.510 ;
        RECT 76.465 117.100 76.635 117.270 ;
        RECT 74.310 116.760 74.480 116.930 ;
        RECT 77.600 116.980 77.770 117.150 ;
        RECT 74.310 116.400 74.480 116.570 ;
        RECT 75.880 116.715 76.050 116.885 ;
        RECT 75.880 116.355 76.050 116.525 ;
        RECT 72.590 115.900 72.760 116.070 ;
        RECT 73.725 115.980 73.895 116.150 ;
        RECT 75.880 115.995 76.050 116.165 ;
        RECT 72.590 115.540 72.760 115.710 ;
        RECT 72.590 115.180 72.760 115.350 ;
        RECT 72.590 114.820 72.760 114.990 ;
        RECT 74.310 115.595 74.480 115.765 ;
        RECT 74.310 115.235 74.480 115.405 ;
        RECT 74.310 114.875 74.480 115.045 ;
        RECT 73.725 114.700 73.895 114.870 ;
        RECT 72.590 114.460 72.760 114.630 ;
        RECT 72.590 114.100 72.760 114.270 ;
        RECT 72.590 113.740 72.760 113.910 ;
        RECT 74.310 114.515 74.480 114.685 ;
        RECT 74.310 114.155 74.480 114.325 ;
        RECT 75.880 115.635 76.050 115.805 ;
        RECT 75.880 115.275 76.050 115.445 ;
        RECT 75.880 114.915 76.050 115.085 ;
        RECT 75.880 114.555 76.050 114.725 ;
        RECT 75.880 114.195 76.050 114.365 ;
        RECT 77.050 116.715 77.220 116.885 ;
        RECT 77.050 116.355 77.220 116.525 ;
        RECT 77.050 115.995 77.220 116.165 ;
        RECT 77.050 115.635 77.220 115.805 ;
        RECT 77.050 115.275 77.220 115.445 ;
        RECT 77.050 114.915 77.220 115.085 ;
        RECT 77.050 114.555 77.220 114.725 ;
        RECT 77.050 114.195 77.220 114.365 ;
        RECT 77.600 116.620 77.770 116.790 ;
        RECT 77.600 116.260 77.770 116.430 ;
        RECT 77.600 115.900 77.770 116.070 ;
        RECT 77.600 115.540 77.770 115.710 ;
        RECT 77.600 115.180 77.770 115.350 ;
        RECT 77.600 114.820 77.770 114.990 ;
        RECT 77.600 114.460 77.770 114.630 ;
        RECT 77.600 114.100 77.770 114.270 ;
        RECT 74.310 113.795 74.480 113.965 ;
        RECT 76.465 113.820 76.635 113.990 ;
        RECT 77.600 113.740 77.770 113.910 ;
        RECT 72.590 113.380 72.760 113.550 ;
        RECT 73.725 113.420 73.895 113.590 ;
        RECT 62.540 112.740 62.710 112.910 ;
        RECT 56.180 112.380 56.350 112.550 ;
        RECT 60.975 112.420 61.145 112.590 ;
        RECT 61.335 112.420 61.505 112.590 ;
        RECT 62.540 112.380 62.710 112.550 ;
        RECT 56.480 111.750 56.650 111.920 ;
        RECT 56.840 111.750 57.010 111.920 ;
        RECT 57.200 111.750 57.370 111.920 ;
        RECT 57.560 111.750 57.730 111.920 ;
        RECT 57.920 111.750 58.090 111.920 ;
        RECT 58.280 111.750 58.450 111.920 ;
        RECT 58.640 111.750 58.810 111.920 ;
        RECT 59.000 111.750 59.170 111.920 ;
        RECT 59.360 111.750 59.530 111.920 ;
        RECT 59.720 111.750 59.890 111.920 ;
        RECT 60.080 111.750 60.250 111.920 ;
        RECT 60.440 111.750 60.610 111.920 ;
        RECT 60.800 111.750 60.970 111.920 ;
        RECT 61.160 111.750 61.330 111.920 ;
        RECT 61.520 111.750 61.690 111.920 ;
        RECT 61.880 111.750 62.050 111.920 ;
        RECT 62.240 111.750 62.410 111.920 ;
        RECT 63.985 113.090 64.155 113.260 ;
        RECT 64.345 113.090 64.515 113.260 ;
        RECT 64.705 113.090 64.875 113.260 ;
        RECT 65.065 113.090 65.235 113.260 ;
        RECT 65.425 113.090 65.595 113.260 ;
        RECT 65.785 113.090 65.955 113.260 ;
        RECT 66.145 113.090 66.315 113.260 ;
        RECT 66.505 113.090 66.675 113.260 ;
        RECT 67.975 113.090 68.145 113.260 ;
        RECT 68.335 113.090 68.505 113.260 ;
        RECT 68.695 113.090 68.865 113.260 ;
        RECT 69.055 113.090 69.225 113.260 ;
        RECT 69.415 113.090 69.585 113.260 ;
        RECT 69.775 113.090 69.945 113.260 ;
        RECT 63.685 112.740 63.855 112.910 ;
        RECT 70.075 112.740 70.245 112.910 ;
        RECT 77.600 113.380 77.770 113.550 ;
        RECT 72.980 112.790 73.150 112.960 ;
        RECT 73.340 112.790 73.510 112.960 ;
        RECT 73.700 112.790 73.870 112.960 ;
        RECT 74.060 112.790 74.230 112.960 ;
        RECT 74.420 112.790 74.590 112.960 ;
        RECT 74.780 112.790 74.950 112.960 ;
        RECT 75.140 112.790 75.310 112.960 ;
        RECT 75.500 112.790 75.670 112.960 ;
        RECT 75.860 112.790 76.030 112.960 ;
        RECT 76.220 112.790 76.390 112.960 ;
        RECT 76.580 112.790 76.750 112.960 ;
        RECT 76.940 112.790 77.110 112.960 ;
        RECT 77.300 112.790 77.470 112.960 ;
        RECT 81.320 142.530 81.490 142.700 ;
        RECT 81.680 142.530 81.850 142.700 ;
        RECT 82.040 142.530 82.210 142.700 ;
        RECT 82.400 142.530 82.570 142.700 ;
        RECT 82.760 142.530 82.930 142.700 ;
        RECT 83.120 142.530 83.290 142.700 ;
        RECT 83.480 142.530 83.650 142.700 ;
        RECT 83.840 142.530 84.010 142.700 ;
        RECT 84.200 142.530 84.370 142.700 ;
        RECT 84.560 142.530 84.730 142.700 ;
        RECT 84.920 142.530 85.090 142.700 ;
        RECT 85.280 142.530 85.450 142.700 ;
        RECT 85.640 142.530 85.810 142.700 ;
        RECT 81.020 142.180 81.190 142.350 ;
        RECT 86.030 142.180 86.200 142.350 ;
        RECT 91.915 142.620 92.085 142.790 ;
        RECT 94.185 142.620 94.355 142.790 ;
        RECT 92.215 142.230 92.385 142.400 ;
        RECT 92.575 142.230 92.745 142.400 ;
        RECT 92.935 142.230 93.105 142.400 ;
        RECT 93.295 142.230 93.465 142.400 ;
        RECT 93.655 142.230 93.825 142.400 ;
        RECT 96.380 151.250 96.550 151.420 ;
        RECT 96.740 151.250 96.910 151.420 ;
        RECT 97.100 151.250 97.270 151.420 ;
        RECT 97.460 151.250 97.630 151.420 ;
        RECT 97.820 151.250 97.990 151.420 ;
        RECT 98.180 151.250 98.350 151.420 ;
        RECT 98.540 151.250 98.710 151.420 ;
        RECT 98.900 151.250 99.070 151.420 ;
        RECT 99.260 151.250 99.430 151.420 ;
        RECT 99.620 151.250 99.790 151.420 ;
        RECT 99.980 151.250 100.150 151.420 ;
        RECT 100.340 151.250 100.510 151.420 ;
        RECT 100.700 151.250 100.870 151.420 ;
        RECT 101.060 151.250 101.230 151.420 ;
        RECT 101.420 151.250 101.590 151.420 ;
        RECT 101.780 151.250 101.950 151.420 ;
        RECT 102.140 151.250 102.310 151.420 ;
        RECT 96.080 150.900 96.250 151.070 ;
        RECT 102.440 150.900 102.610 151.070 ;
        RECT 96.080 150.540 96.250 150.710 ;
        RECT 97.285 150.580 97.455 150.750 ;
        RECT 97.645 150.580 97.815 150.750 ;
        RECT 96.080 150.180 96.250 150.350 ;
        RECT 102.440 150.540 102.610 150.710 ;
        RECT 96.080 149.820 96.250 149.990 ;
        RECT 98.300 150.160 98.470 150.330 ;
        RECT 97.285 149.800 97.455 149.970 ;
        RECT 97.645 149.800 97.815 149.970 ;
        RECT 98.300 149.800 98.470 149.970 ;
        RECT 96.080 149.460 96.250 149.630 ;
        RECT 98.300 149.440 98.470 149.610 ;
        RECT 102.440 150.180 102.610 150.350 ;
        RECT 102.440 149.820 102.610 149.990 ;
        RECT 102.440 149.460 102.610 149.630 ;
        RECT 96.080 149.100 96.250 149.270 ;
        RECT 97.285 149.020 97.455 149.190 ;
        RECT 97.645 149.020 97.815 149.190 ;
        RECT 102.440 149.100 102.610 149.270 ;
        RECT 96.080 148.740 96.250 148.910 ;
        RECT 96.080 148.380 96.250 148.550 ;
        RECT 96.080 148.020 96.250 148.190 ;
        RECT 96.080 147.660 96.250 147.830 ;
        RECT 96.080 147.300 96.250 147.470 ;
        RECT 96.630 148.600 96.800 148.770 ;
        RECT 96.630 148.240 96.800 148.410 ;
        RECT 96.630 147.880 96.800 148.050 ;
        RECT 96.630 147.520 96.800 147.690 ;
        RECT 96.630 147.160 96.800 147.330 ;
        RECT 102.440 148.740 102.610 148.910 ;
        RECT 102.440 148.380 102.610 148.550 ;
        RECT 102.440 148.020 102.610 148.190 ;
        RECT 102.440 147.660 102.610 147.830 ;
        RECT 102.440 147.300 102.610 147.470 ;
        RECT 96.080 146.940 96.250 147.110 ;
        RECT 102.440 146.940 102.610 147.110 ;
        RECT 96.080 146.580 96.250 146.750 ;
        RECT 97.285 146.740 97.455 146.910 ;
        RECT 97.645 146.740 97.815 146.910 ;
        RECT 102.440 146.580 102.610 146.750 ;
        RECT 96.080 146.220 96.250 146.390 ;
        RECT 96.080 145.860 96.250 146.030 ;
        RECT 96.080 145.500 96.250 145.670 ;
        RECT 96.080 145.140 96.250 145.310 ;
        RECT 96.080 144.780 96.250 144.950 ;
        RECT 96.630 146.320 96.800 146.490 ;
        RECT 96.630 145.960 96.800 146.130 ;
        RECT 96.630 145.600 96.800 145.770 ;
        RECT 96.630 145.240 96.800 145.410 ;
        RECT 96.630 144.880 96.800 145.050 ;
        RECT 102.440 146.220 102.610 146.390 ;
        RECT 102.440 145.860 102.610 146.030 ;
        RECT 102.440 145.500 102.610 145.670 ;
        RECT 102.440 145.140 102.610 145.310 ;
        RECT 102.440 144.780 102.610 144.950 ;
        RECT 96.080 144.420 96.250 144.590 ;
        RECT 97.285 144.460 97.455 144.630 ;
        RECT 97.645 144.460 97.815 144.630 ;
        RECT 96.080 144.060 96.250 144.230 ;
        RECT 102.440 144.420 102.610 144.590 ;
        RECT 96.080 143.700 96.250 143.870 ;
        RECT 98.300 144.040 98.470 144.210 ;
        RECT 97.285 143.680 97.455 143.850 ;
        RECT 97.645 143.680 97.815 143.850 ;
        RECT 98.300 143.680 98.470 143.850 ;
        RECT 96.080 143.340 96.250 143.510 ;
        RECT 98.300 143.320 98.470 143.490 ;
        RECT 102.440 144.060 102.610 144.230 ;
        RECT 102.440 143.700 102.610 143.870 ;
        RECT 102.440 143.340 102.610 143.510 ;
        RECT 96.080 142.980 96.250 143.150 ;
        RECT 97.285 142.900 97.455 143.070 ;
        RECT 97.645 142.900 97.815 143.070 ;
        RECT 102.440 142.980 102.610 143.150 ;
        RECT 96.080 142.620 96.250 142.790 ;
        RECT 96.080 142.260 96.250 142.430 ;
        RECT 98.300 142.480 98.470 142.650 ;
        RECT 81.020 141.820 81.190 141.990 ;
        RECT 84.895 141.900 85.065 142.070 ;
        RECT 86.030 141.820 86.200 141.990 ;
        RECT 81.020 141.460 81.190 141.630 ;
        RECT 82.155 141.500 82.325 141.670 ;
        RECT 84.310 141.515 84.480 141.685 ;
        RECT 81.020 141.100 81.190 141.270 ;
        RECT 81.020 140.740 81.190 140.910 ;
        RECT 81.020 140.380 81.190 140.550 ;
        RECT 81.020 140.020 81.190 140.190 ;
        RECT 81.020 139.660 81.190 139.830 ;
        RECT 81.020 139.300 81.190 139.470 ;
        RECT 81.020 138.940 81.190 139.110 ;
        RECT 81.020 138.580 81.190 138.750 ;
        RECT 81.570 141.115 81.740 141.285 ;
        RECT 81.570 140.755 81.740 140.925 ;
        RECT 81.570 140.395 81.740 140.565 ;
        RECT 81.570 140.035 81.740 140.205 ;
        RECT 81.570 139.675 81.740 139.845 ;
        RECT 81.570 139.315 81.740 139.485 ;
        RECT 81.570 138.955 81.740 139.125 ;
        RECT 81.570 138.595 81.740 138.765 ;
        RECT 82.740 141.115 82.910 141.285 ;
        RECT 82.740 140.755 82.910 140.925 ;
        RECT 82.740 140.395 82.910 140.565 ;
        RECT 82.740 140.035 82.910 140.205 ;
        RECT 82.740 139.675 82.910 139.845 ;
        RECT 84.310 141.155 84.480 141.325 ;
        RECT 84.310 140.795 84.480 140.965 ;
        RECT 86.030 141.460 86.200 141.630 ;
        RECT 86.030 141.100 86.200 141.270 ;
        RECT 84.895 140.620 85.065 140.790 ;
        RECT 86.030 140.740 86.200 140.910 ;
        RECT 84.310 140.435 84.480 140.605 ;
        RECT 84.310 140.075 84.480 140.245 ;
        RECT 84.310 139.715 84.480 139.885 ;
        RECT 86.030 140.380 86.200 140.550 ;
        RECT 86.030 140.020 86.200 140.190 ;
        RECT 86.030 139.660 86.200 139.830 ;
        RECT 82.740 139.315 82.910 139.485 ;
        RECT 84.895 139.340 85.065 139.510 ;
        RECT 82.740 138.955 82.910 139.125 ;
        RECT 86.030 139.300 86.200 139.470 ;
        RECT 82.740 138.595 82.910 138.765 ;
        RECT 84.310 138.920 84.480 139.090 ;
        RECT 84.310 138.560 84.480 138.730 ;
        RECT 81.020 138.220 81.190 138.390 ;
        RECT 82.155 138.220 82.325 138.390 ;
        RECT 81.020 137.860 81.190 138.030 ;
        RECT 84.310 138.200 84.480 138.370 ;
        RECT 81.020 137.500 81.190 137.670 ;
        RECT 81.020 137.140 81.190 137.310 ;
        RECT 81.020 136.780 81.190 136.950 ;
        RECT 81.020 136.420 81.190 136.590 ;
        RECT 81.020 136.060 81.190 136.230 ;
        RECT 81.020 135.700 81.190 135.870 ;
        RECT 81.020 135.340 81.190 135.510 ;
        RECT 81.570 137.835 81.740 138.005 ;
        RECT 81.570 137.475 81.740 137.645 ;
        RECT 81.570 137.115 81.740 137.285 ;
        RECT 81.570 136.755 81.740 136.925 ;
        RECT 81.570 136.395 81.740 136.565 ;
        RECT 81.570 136.035 81.740 136.205 ;
        RECT 81.570 135.675 81.740 135.845 ;
        RECT 81.570 135.315 81.740 135.485 ;
        RECT 82.740 137.835 82.910 138.005 ;
        RECT 82.740 137.475 82.910 137.645 ;
        RECT 84.310 137.840 84.480 138.010 ;
        RECT 84.310 137.480 84.480 137.650 ;
        RECT 85.480 138.920 85.650 139.090 ;
        RECT 85.480 138.560 85.650 138.730 ;
        RECT 85.480 138.200 85.650 138.370 ;
        RECT 85.480 137.840 85.650 138.010 ;
        RECT 85.480 137.480 85.650 137.650 ;
        RECT 86.030 138.940 86.200 139.110 ;
        RECT 86.030 138.580 86.200 138.750 ;
        RECT 86.030 138.220 86.200 138.390 ;
        RECT 97.285 142.120 97.455 142.290 ;
        RECT 97.645 142.120 97.815 142.290 ;
        RECT 98.300 142.120 98.470 142.290 ;
        RECT 96.080 141.900 96.250 142.070 ;
        RECT 98.300 141.760 98.470 141.930 ;
        RECT 102.440 142.620 102.610 142.790 ;
        RECT 102.440 142.260 102.610 142.430 ;
        RECT 102.440 141.900 102.610 142.070 ;
        RECT 96.080 141.540 96.250 141.710 ;
        RECT 102.440 141.540 102.610 141.710 ;
        RECT 96.080 141.180 96.250 141.350 ;
        RECT 97.285 141.340 97.455 141.510 ;
        RECT 97.645 141.340 97.815 141.510 ;
        RECT 100.875 141.340 101.045 141.510 ;
        RECT 101.235 141.340 101.405 141.510 ;
        RECT 102.440 141.180 102.610 141.350 ;
        RECT 96.080 140.820 96.250 140.990 ;
        RECT 96.080 140.460 96.250 140.630 ;
        RECT 96.080 140.100 96.250 140.270 ;
        RECT 96.080 139.740 96.250 139.910 ;
        RECT 96.080 139.380 96.250 139.550 ;
        RECT 96.630 140.920 96.800 141.090 ;
        RECT 96.630 140.560 96.800 140.730 ;
        RECT 96.630 140.200 96.800 140.370 ;
        RECT 96.630 139.840 96.800 140.010 ;
        RECT 96.630 139.480 96.800 139.650 ;
        RECT 98.300 140.920 98.470 141.090 ;
        RECT 98.300 140.560 98.470 140.730 ;
        RECT 98.300 140.200 98.470 140.370 ;
        RECT 98.300 139.840 98.470 140.010 ;
        RECT 98.300 139.480 98.470 139.650 ;
        RECT 100.220 140.920 100.390 141.090 ;
        RECT 100.220 140.560 100.390 140.730 ;
        RECT 100.220 140.200 100.390 140.370 ;
        RECT 100.220 139.840 100.390 140.010 ;
        RECT 100.220 139.480 100.390 139.650 ;
        RECT 102.440 140.820 102.610 140.990 ;
        RECT 102.440 140.460 102.610 140.630 ;
        RECT 102.440 140.100 102.610 140.270 ;
        RECT 102.440 139.740 102.610 139.910 ;
        RECT 102.440 139.380 102.610 139.550 ;
        RECT 96.080 139.020 96.250 139.190 ;
        RECT 97.285 139.060 97.455 139.230 ;
        RECT 97.645 139.060 97.815 139.230 ;
        RECT 100.875 139.060 101.045 139.230 ;
        RECT 101.235 139.060 101.405 139.230 ;
        RECT 96.080 138.660 96.250 138.830 ;
        RECT 102.440 139.020 102.610 139.190 ;
        RECT 96.080 138.300 96.250 138.470 ;
        RECT 86.030 137.860 86.200 138.030 ;
        RECT 86.030 137.500 86.200 137.670 ;
        RECT 82.740 137.115 82.910 137.285 ;
        RECT 84.895 137.060 85.065 137.230 ;
        RECT 86.030 137.140 86.200 137.310 ;
        RECT 82.740 136.755 82.910 136.925 ;
        RECT 82.740 136.395 82.910 136.565 ;
        RECT 82.740 136.035 82.910 136.205 ;
        RECT 82.740 135.675 82.910 135.845 ;
        RECT 82.740 135.315 82.910 135.485 ;
        RECT 84.310 136.640 84.480 136.810 ;
        RECT 84.310 136.280 84.480 136.450 ;
        RECT 84.310 135.920 84.480 136.090 ;
        RECT 84.310 135.560 84.480 135.730 ;
        RECT 84.310 135.200 84.480 135.370 ;
        RECT 85.480 136.640 85.650 136.810 ;
        RECT 85.480 136.280 85.650 136.450 ;
        RECT 85.480 135.920 85.650 136.090 ;
        RECT 85.480 135.560 85.650 135.730 ;
        RECT 85.480 135.200 85.650 135.370 ;
        RECT 86.030 136.780 86.200 136.950 ;
        RECT 86.030 136.420 86.200 136.590 ;
        RECT 86.030 136.060 86.200 136.230 ;
        RECT 86.030 135.700 86.200 135.870 ;
        RECT 86.030 135.340 86.200 135.510 ;
        RECT 81.020 134.980 81.190 135.150 ;
        RECT 82.155 134.940 82.325 135.110 ;
        RECT 86.030 134.980 86.200 135.150 ;
        RECT 81.020 134.620 81.190 134.790 ;
        RECT 84.895 134.780 85.065 134.950 ;
        RECT 81.020 134.260 81.190 134.430 ;
        RECT 81.020 133.900 81.190 134.070 ;
        RECT 81.020 133.540 81.190 133.710 ;
        RECT 81.020 133.180 81.190 133.350 ;
        RECT 81.020 132.820 81.190 132.990 ;
        RECT 81.020 132.460 81.190 132.630 ;
        RECT 81.020 132.100 81.190 132.270 ;
        RECT 81.020 131.740 81.190 131.910 ;
        RECT 81.020 131.380 81.190 131.550 ;
        RECT 81.020 131.020 81.190 131.190 ;
        RECT 81.020 130.660 81.190 130.830 ;
        RECT 81.020 130.300 81.190 130.470 ;
        RECT 81.020 129.940 81.190 130.110 ;
        RECT 81.020 129.580 81.190 129.750 ;
        RECT 81.020 129.220 81.190 129.390 ;
        RECT 81.020 128.860 81.190 129.030 ;
        RECT 81.020 128.500 81.190 128.670 ;
        RECT 81.020 128.140 81.190 128.310 ;
        RECT 81.570 134.540 81.740 134.710 ;
        RECT 86.030 134.620 86.200 134.790 ;
        RECT 81.570 134.180 81.740 134.350 ;
        RECT 81.570 133.820 81.740 133.990 ;
        RECT 81.570 133.460 81.740 133.630 ;
        RECT 81.570 133.100 81.740 133.270 ;
        RECT 84.310 134.360 84.480 134.530 ;
        RECT 84.310 134.000 84.480 134.170 ;
        RECT 84.310 133.640 84.480 133.810 ;
        RECT 84.310 133.280 84.480 133.450 ;
        RECT 84.310 132.920 84.480 133.090 ;
        RECT 85.480 134.360 85.650 134.530 ;
        RECT 85.480 134.000 85.650 134.170 ;
        RECT 85.480 133.640 85.650 133.810 ;
        RECT 85.480 133.280 85.650 133.450 ;
        RECT 85.480 132.920 85.650 133.090 ;
        RECT 86.030 134.260 86.200 134.430 ;
        RECT 86.030 133.900 86.200 134.070 ;
        RECT 86.030 133.540 86.200 133.710 ;
        RECT 86.030 133.180 86.200 133.350 ;
        RECT 81.570 132.740 81.740 132.910 ;
        RECT 86.030 132.820 86.200 132.990 ;
        RECT 81.570 132.380 81.740 132.550 ;
        RECT 84.895 132.500 85.065 132.670 ;
        RECT 86.030 132.460 86.200 132.630 ;
        RECT 81.570 132.020 81.740 132.190 ;
        RECT 81.570 131.660 81.740 131.830 ;
        RECT 81.570 131.300 81.740 131.470 ;
        RECT 81.570 130.940 81.740 131.110 ;
        RECT 81.570 130.580 81.740 130.750 ;
        RECT 84.310 132.080 84.480 132.250 ;
        RECT 84.310 131.720 84.480 131.890 ;
        RECT 84.310 131.360 84.480 131.530 ;
        RECT 84.310 131.000 84.480 131.170 ;
        RECT 84.310 130.640 84.480 130.810 ;
        RECT 85.480 132.080 85.650 132.250 ;
        RECT 85.480 131.720 85.650 131.890 ;
        RECT 85.480 131.360 85.650 131.530 ;
        RECT 85.480 131.000 85.650 131.170 ;
        RECT 85.480 130.640 85.650 130.810 ;
        RECT 86.030 132.100 86.200 132.270 ;
        RECT 86.030 131.740 86.200 131.910 ;
        RECT 86.030 131.380 86.200 131.550 ;
        RECT 86.030 131.020 86.200 131.190 ;
        RECT 86.030 130.660 86.200 130.830 ;
        RECT 81.570 130.220 81.740 130.390 ;
        RECT 84.895 130.220 85.065 130.390 ;
        RECT 86.030 130.300 86.200 130.470 ;
        RECT 81.570 129.860 81.740 130.030 ;
        RECT 81.570 129.500 81.740 129.670 ;
        RECT 81.570 129.140 81.740 129.310 ;
        RECT 81.570 128.780 81.740 128.950 ;
        RECT 81.570 128.420 81.740 128.590 ;
        RECT 81.570 128.060 81.740 128.230 ;
        RECT 84.310 129.835 84.480 130.005 ;
        RECT 84.310 129.475 84.480 129.645 ;
        RECT 84.310 129.115 84.480 129.285 ;
        RECT 85.480 129.835 85.650 130.005 ;
        RECT 85.480 129.475 85.650 129.645 ;
        RECT 85.480 129.115 85.650 129.285 ;
        RECT 84.895 128.940 85.065 129.110 ;
        RECT 84.310 128.755 84.480 128.925 ;
        RECT 84.310 128.395 84.480 128.565 ;
        RECT 84.310 128.035 84.480 128.205 ;
        RECT 85.480 128.755 85.650 128.925 ;
        RECT 85.480 128.395 85.650 128.565 ;
        RECT 85.480 128.035 85.650 128.205 ;
        RECT 86.030 129.940 86.200 130.110 ;
        RECT 86.030 129.580 86.200 129.750 ;
        RECT 86.030 129.220 86.200 129.390 ;
        RECT 86.030 128.860 86.200 129.030 ;
        RECT 86.030 128.500 86.200 128.670 ;
        RECT 86.030 128.140 86.200 128.310 ;
        RECT 81.020 127.780 81.190 127.950 ;
        RECT 82.155 127.660 82.325 127.830 ;
        RECT 84.895 127.660 85.065 127.830 ;
        RECT 86.030 127.780 86.200 127.950 ;
        RECT 81.020 127.420 81.190 127.590 ;
        RECT 81.020 127.060 81.190 127.230 ;
        RECT 81.020 126.700 81.190 126.870 ;
        RECT 81.020 126.340 81.190 126.510 ;
        RECT 81.020 125.980 81.190 126.150 ;
        RECT 81.020 125.620 81.190 125.790 ;
        RECT 81.020 125.260 81.190 125.430 ;
        RECT 81.020 124.900 81.190 125.070 ;
        RECT 81.020 124.540 81.190 124.710 ;
        RECT 81.020 124.180 81.190 124.350 ;
        RECT 81.020 123.820 81.190 123.990 ;
        RECT 81.020 123.460 81.190 123.630 ;
        RECT 81.020 123.100 81.190 123.270 ;
        RECT 81.020 122.740 81.190 122.910 ;
        RECT 81.020 122.380 81.190 122.550 ;
        RECT 81.020 122.020 81.190 122.190 ;
        RECT 81.020 121.660 81.190 121.830 ;
        RECT 81.020 121.300 81.190 121.470 ;
        RECT 81.020 120.940 81.190 121.110 ;
        RECT 81.570 127.260 81.740 127.430 ;
        RECT 81.570 126.900 81.740 127.070 ;
        RECT 81.570 126.540 81.740 126.710 ;
        RECT 81.570 126.180 81.740 126.350 ;
        RECT 81.570 125.820 81.740 125.990 ;
        RECT 81.570 125.460 81.740 125.630 ;
        RECT 84.310 127.275 84.480 127.445 ;
        RECT 84.310 126.915 84.480 127.085 ;
        RECT 84.310 126.555 84.480 126.725 ;
        RECT 85.480 127.275 85.650 127.445 ;
        RECT 85.480 126.915 85.650 127.085 ;
        RECT 85.480 126.555 85.650 126.725 ;
        RECT 84.895 126.380 85.065 126.550 ;
        RECT 84.310 126.195 84.480 126.365 ;
        RECT 84.310 125.835 84.480 126.005 ;
        RECT 84.310 125.475 84.480 125.645 ;
        RECT 85.480 126.195 85.650 126.365 ;
        RECT 85.480 125.835 85.650 126.005 ;
        RECT 85.480 125.475 85.650 125.645 ;
        RECT 86.030 127.420 86.200 127.590 ;
        RECT 86.030 127.060 86.200 127.230 ;
        RECT 86.030 126.700 86.200 126.870 ;
        RECT 86.030 126.340 86.200 126.510 ;
        RECT 86.030 125.980 86.200 126.150 ;
        RECT 86.030 125.620 86.200 125.790 ;
        RECT 81.570 125.100 81.740 125.270 ;
        RECT 84.895 125.100 85.065 125.270 ;
        RECT 86.030 125.260 86.200 125.430 ;
        RECT 81.570 124.740 81.740 124.910 ;
        RECT 86.030 124.900 86.200 125.070 ;
        RECT 81.570 124.380 81.740 124.550 ;
        RECT 81.570 124.020 81.740 124.190 ;
        RECT 81.570 123.660 81.740 123.830 ;
        RECT 81.570 123.300 81.740 123.470 ;
        RECT 84.310 124.680 84.480 124.850 ;
        RECT 84.310 124.320 84.480 124.490 ;
        RECT 84.310 123.960 84.480 124.130 ;
        RECT 84.310 123.600 84.480 123.770 ;
        RECT 84.310 123.240 84.480 123.410 ;
        RECT 85.480 124.680 85.650 124.850 ;
        RECT 85.480 124.320 85.650 124.490 ;
        RECT 85.480 123.960 85.650 124.130 ;
        RECT 85.480 123.600 85.650 123.770 ;
        RECT 85.480 123.240 85.650 123.410 ;
        RECT 86.030 124.540 86.200 124.710 ;
        RECT 86.030 124.180 86.200 124.350 ;
        RECT 86.030 123.820 86.200 123.990 ;
        RECT 86.030 123.460 86.200 123.630 ;
        RECT 81.570 122.940 81.740 123.110 ;
        RECT 86.030 123.100 86.200 123.270 ;
        RECT 84.895 122.820 85.065 122.990 ;
        RECT 81.570 122.580 81.740 122.750 ;
        RECT 86.030 122.740 86.200 122.910 ;
        RECT 81.570 122.220 81.740 122.390 ;
        RECT 81.570 121.860 81.740 122.030 ;
        RECT 81.570 121.500 81.740 121.670 ;
        RECT 81.570 121.140 81.740 121.310 ;
        RECT 84.310 122.400 84.480 122.570 ;
        RECT 84.310 122.040 84.480 122.210 ;
        RECT 84.310 121.680 84.480 121.850 ;
        RECT 84.310 121.320 84.480 121.490 ;
        RECT 84.310 120.960 84.480 121.130 ;
        RECT 85.480 122.400 85.650 122.570 ;
        RECT 85.480 122.040 85.650 122.210 ;
        RECT 85.480 121.680 85.650 121.850 ;
        RECT 85.480 121.320 85.650 121.490 ;
        RECT 85.480 120.960 85.650 121.130 ;
        RECT 86.030 122.380 86.200 122.550 ;
        RECT 86.030 122.020 86.200 122.190 ;
        RECT 86.030 121.660 86.200 121.830 ;
        RECT 86.030 121.300 86.200 121.470 ;
        RECT 81.570 120.780 81.740 120.950 ;
        RECT 86.030 120.940 86.200 121.110 ;
        RECT 81.020 120.580 81.190 120.750 ;
        RECT 81.020 120.220 81.190 120.390 ;
        RECT 82.155 120.380 82.325 120.550 ;
        RECT 84.895 120.540 85.065 120.710 ;
        RECT 86.030 120.580 86.200 120.750 ;
        RECT 81.020 119.860 81.190 120.030 ;
        RECT 81.020 119.500 81.190 119.670 ;
        RECT 81.020 119.140 81.190 119.310 ;
        RECT 81.020 118.780 81.190 118.950 ;
        RECT 81.020 118.420 81.190 118.590 ;
        RECT 81.020 118.060 81.190 118.230 ;
        RECT 81.020 117.700 81.190 117.870 ;
        RECT 81.020 117.340 81.190 117.510 ;
        RECT 81.570 119.995 81.740 120.165 ;
        RECT 81.570 119.635 81.740 119.805 ;
        RECT 81.570 119.275 81.740 119.445 ;
        RECT 81.570 118.915 81.740 119.085 ;
        RECT 81.570 118.555 81.740 118.725 ;
        RECT 81.570 118.195 81.740 118.365 ;
        RECT 81.570 117.835 81.740 118.005 ;
        RECT 81.570 117.475 81.740 117.645 ;
        RECT 82.740 119.995 82.910 120.165 ;
        RECT 82.740 119.635 82.910 119.805 ;
        RECT 82.740 119.275 82.910 119.445 ;
        RECT 82.740 118.915 82.910 119.085 ;
        RECT 82.740 118.555 82.910 118.725 ;
        RECT 84.310 120.120 84.480 120.290 ;
        RECT 84.310 119.760 84.480 119.930 ;
        RECT 84.310 119.400 84.480 119.570 ;
        RECT 84.310 119.040 84.480 119.210 ;
        RECT 84.310 118.680 84.480 118.850 ;
        RECT 85.480 120.120 85.650 120.290 ;
        RECT 85.480 119.760 85.650 119.930 ;
        RECT 85.480 119.400 85.650 119.570 ;
        RECT 85.480 119.040 85.650 119.210 ;
        RECT 85.480 118.680 85.650 118.850 ;
        RECT 86.030 120.220 86.200 120.390 ;
        RECT 86.030 119.860 86.200 120.030 ;
        RECT 86.030 119.500 86.200 119.670 ;
        RECT 86.030 119.140 86.200 119.310 ;
        RECT 86.030 118.780 86.200 118.950 ;
        RECT 82.740 118.195 82.910 118.365 ;
        RECT 84.895 118.260 85.065 118.430 ;
        RECT 86.030 118.420 86.200 118.590 ;
        RECT 86.030 118.060 86.200 118.230 ;
        RECT 82.740 117.835 82.910 118.005 ;
        RECT 82.740 117.475 82.910 117.645 ;
        RECT 84.310 117.840 84.480 118.010 ;
        RECT 84.310 117.480 84.480 117.650 ;
        RECT 81.020 116.980 81.190 117.150 ;
        RECT 82.155 117.100 82.325 117.270 ;
        RECT 84.310 117.120 84.480 117.290 ;
        RECT 81.020 116.620 81.190 116.790 ;
        RECT 81.020 116.260 81.190 116.430 ;
        RECT 81.020 115.900 81.190 116.070 ;
        RECT 81.020 115.540 81.190 115.710 ;
        RECT 81.020 115.180 81.190 115.350 ;
        RECT 81.020 114.820 81.190 114.990 ;
        RECT 81.020 114.460 81.190 114.630 ;
        RECT 81.020 114.100 81.190 114.270 ;
        RECT 81.570 116.715 81.740 116.885 ;
        RECT 81.570 116.355 81.740 116.525 ;
        RECT 81.570 115.995 81.740 116.165 ;
        RECT 81.570 115.635 81.740 115.805 ;
        RECT 81.570 115.275 81.740 115.445 ;
        RECT 81.570 114.915 81.740 115.085 ;
        RECT 81.570 114.555 81.740 114.725 ;
        RECT 81.570 114.195 81.740 114.365 ;
        RECT 82.740 116.715 82.910 116.885 ;
        RECT 82.740 116.355 82.910 116.525 ;
        RECT 84.310 116.760 84.480 116.930 ;
        RECT 84.310 116.400 84.480 116.570 ;
        RECT 85.480 117.840 85.650 118.010 ;
        RECT 85.480 117.480 85.650 117.650 ;
        RECT 85.480 117.120 85.650 117.290 ;
        RECT 85.480 116.760 85.650 116.930 ;
        RECT 85.480 116.400 85.650 116.570 ;
        RECT 86.030 117.700 86.200 117.870 ;
        RECT 86.030 117.340 86.200 117.510 ;
        RECT 87.960 138.040 88.130 138.210 ;
        RECT 88.320 138.040 88.490 138.210 ;
        RECT 88.680 138.040 88.850 138.210 ;
        RECT 89.040 138.040 89.210 138.210 ;
        RECT 89.400 138.040 89.570 138.210 ;
        RECT 89.760 138.040 89.930 138.210 ;
        RECT 90.120 138.040 90.290 138.210 ;
        RECT 87.660 137.690 87.830 137.860 ;
        RECT 90.430 137.690 90.600 137.860 ;
        RECT 87.660 137.330 87.830 137.500 ;
        RECT 88.865 137.370 89.035 137.540 ;
        RECT 89.225 137.370 89.395 137.540 ;
        RECT 90.430 137.330 90.600 137.500 ;
        RECT 87.660 136.970 87.830 137.140 ;
        RECT 87.660 136.610 87.830 136.780 ;
        RECT 87.660 136.250 87.830 136.420 ;
        RECT 87.660 135.890 87.830 136.060 ;
        RECT 87.660 135.530 87.830 135.700 ;
        RECT 87.660 135.170 87.830 135.340 ;
        RECT 88.210 136.985 88.380 137.155 ;
        RECT 88.210 136.625 88.380 136.795 ;
        RECT 88.210 136.265 88.380 136.435 ;
        RECT 89.880 136.985 90.050 137.155 ;
        RECT 89.880 136.625 90.050 136.795 ;
        RECT 89.880 136.265 90.050 136.435 ;
        RECT 88.865 136.090 89.035 136.260 ;
        RECT 89.225 136.090 89.395 136.260 ;
        RECT 88.210 135.905 88.380 136.075 ;
        RECT 88.210 135.545 88.380 135.715 ;
        RECT 88.210 135.185 88.380 135.355 ;
        RECT 89.880 135.905 90.050 136.075 ;
        RECT 89.880 135.545 90.050 135.715 ;
        RECT 89.880 135.185 90.050 135.355 ;
        RECT 90.430 136.970 90.600 137.140 ;
        RECT 90.430 136.610 90.600 136.780 ;
        RECT 90.430 136.250 90.600 136.420 ;
        RECT 90.430 135.890 90.600 136.060 ;
        RECT 90.430 135.530 90.600 135.700 ;
        RECT 90.430 135.170 90.600 135.340 ;
        RECT 87.660 134.810 87.830 134.980 ;
        RECT 88.865 134.810 89.035 134.980 ;
        RECT 89.225 134.810 89.395 134.980 ;
        RECT 90.430 134.810 90.600 134.980 ;
        RECT 87.660 134.450 87.830 134.620 ;
        RECT 87.660 134.090 87.830 134.260 ;
        RECT 87.660 133.730 87.830 133.900 ;
        RECT 87.660 133.370 87.830 133.540 ;
        RECT 87.660 133.010 87.830 133.180 ;
        RECT 88.210 134.390 88.380 134.560 ;
        RECT 88.210 134.030 88.380 134.200 ;
        RECT 88.210 133.670 88.380 133.840 ;
        RECT 88.210 133.310 88.380 133.480 ;
        RECT 88.210 132.950 88.380 133.120 ;
        RECT 89.880 134.390 90.050 134.560 ;
        RECT 89.880 134.030 90.050 134.200 ;
        RECT 89.880 133.670 90.050 133.840 ;
        RECT 89.880 133.310 90.050 133.480 ;
        RECT 89.880 132.950 90.050 133.120 ;
        RECT 90.430 134.450 90.600 134.620 ;
        RECT 90.430 134.090 90.600 134.260 ;
        RECT 90.430 133.730 90.600 133.900 ;
        RECT 90.430 133.370 90.600 133.540 ;
        RECT 90.430 133.010 90.600 133.180 ;
        RECT 87.660 132.650 87.830 132.820 ;
        RECT 88.865 132.530 89.035 132.700 ;
        RECT 89.225 132.530 89.395 132.700 ;
        RECT 90.430 132.650 90.600 132.820 ;
        RECT 87.660 132.290 87.830 132.460 ;
        RECT 90.430 132.290 90.600 132.460 ;
        RECT 87.660 131.930 87.830 132.100 ;
        RECT 87.660 131.570 87.830 131.740 ;
        RECT 87.660 131.210 87.830 131.380 ;
        RECT 87.660 130.850 87.830 131.020 ;
        RECT 88.210 132.110 88.380 132.280 ;
        RECT 88.210 131.750 88.380 131.920 ;
        RECT 88.210 131.390 88.380 131.560 ;
        RECT 88.210 131.030 88.380 131.200 ;
        RECT 88.210 130.670 88.380 130.840 ;
        RECT 89.880 132.110 90.050 132.280 ;
        RECT 89.880 131.750 90.050 131.920 ;
        RECT 89.880 131.390 90.050 131.560 ;
        RECT 89.880 131.030 90.050 131.200 ;
        RECT 89.880 130.670 90.050 130.840 ;
        RECT 90.430 131.930 90.600 132.100 ;
        RECT 90.430 131.570 90.600 131.740 ;
        RECT 90.430 131.210 90.600 131.380 ;
        RECT 90.430 130.850 90.600 131.020 ;
        RECT 87.660 130.490 87.830 130.660 ;
        RECT 90.430 130.490 90.600 130.660 ;
        RECT 87.660 130.130 87.830 130.300 ;
        RECT 88.865 130.250 89.035 130.420 ;
        RECT 89.225 130.250 89.395 130.420 ;
        RECT 90.430 130.130 90.600 130.300 ;
        RECT 87.660 129.770 87.830 129.940 ;
        RECT 87.660 129.410 87.830 129.580 ;
        RECT 87.660 129.050 87.830 129.220 ;
        RECT 87.660 128.690 87.830 128.860 ;
        RECT 87.660 128.330 87.830 128.500 ;
        RECT 87.660 127.970 87.830 128.140 ;
        RECT 88.210 129.865 88.380 130.035 ;
        RECT 88.210 129.505 88.380 129.675 ;
        RECT 88.210 129.145 88.380 129.315 ;
        RECT 89.880 129.865 90.050 130.035 ;
        RECT 89.880 129.505 90.050 129.675 ;
        RECT 89.880 129.145 90.050 129.315 ;
        RECT 88.865 128.970 89.035 129.140 ;
        RECT 89.225 128.970 89.395 129.140 ;
        RECT 88.210 128.785 88.380 128.955 ;
        RECT 88.210 128.425 88.380 128.595 ;
        RECT 88.210 128.065 88.380 128.235 ;
        RECT 89.880 128.785 90.050 128.955 ;
        RECT 89.880 128.425 90.050 128.595 ;
        RECT 89.880 128.065 90.050 128.235 ;
        RECT 90.430 129.770 90.600 129.940 ;
        RECT 90.430 129.410 90.600 129.580 ;
        RECT 90.430 129.050 90.600 129.220 ;
        RECT 90.430 128.690 90.600 128.860 ;
        RECT 90.430 128.330 90.600 128.500 ;
        RECT 90.430 127.970 90.600 128.140 ;
        RECT 87.660 127.610 87.830 127.780 ;
        RECT 88.865 127.690 89.035 127.860 ;
        RECT 89.225 127.690 89.395 127.860 ;
        RECT 90.430 127.610 90.600 127.780 ;
        RECT 87.660 127.250 87.830 127.420 ;
        RECT 87.660 126.890 87.830 127.060 ;
        RECT 87.660 126.530 87.830 126.700 ;
        RECT 87.660 126.170 87.830 126.340 ;
        RECT 87.660 125.810 87.830 125.980 ;
        RECT 87.660 125.450 87.830 125.620 ;
        RECT 88.210 127.305 88.380 127.475 ;
        RECT 88.210 126.945 88.380 127.115 ;
        RECT 88.210 126.585 88.380 126.755 ;
        RECT 89.880 127.305 90.050 127.475 ;
        RECT 89.880 126.945 90.050 127.115 ;
        RECT 89.880 126.585 90.050 126.755 ;
        RECT 88.865 126.410 89.035 126.580 ;
        RECT 89.225 126.410 89.395 126.580 ;
        RECT 88.210 126.225 88.380 126.395 ;
        RECT 88.210 125.865 88.380 126.035 ;
        RECT 88.210 125.505 88.380 125.675 ;
        RECT 89.880 126.225 90.050 126.395 ;
        RECT 89.880 125.865 90.050 126.035 ;
        RECT 89.880 125.505 90.050 125.675 ;
        RECT 90.430 127.250 90.600 127.420 ;
        RECT 90.430 126.890 90.600 127.060 ;
        RECT 90.430 126.530 90.600 126.700 ;
        RECT 90.430 126.170 90.600 126.340 ;
        RECT 90.430 125.810 90.600 125.980 ;
        RECT 90.430 125.450 90.600 125.620 ;
        RECT 87.660 125.090 87.830 125.260 ;
        RECT 88.865 125.130 89.035 125.300 ;
        RECT 89.225 125.130 89.395 125.300 ;
        RECT 87.660 124.730 87.830 124.900 ;
        RECT 90.430 125.090 90.600 125.260 ;
        RECT 87.660 124.370 87.830 124.540 ;
        RECT 87.660 124.010 87.830 124.180 ;
        RECT 87.660 123.650 87.830 123.820 ;
        RECT 87.660 123.290 87.830 123.460 ;
        RECT 88.210 124.710 88.380 124.880 ;
        RECT 88.210 124.350 88.380 124.520 ;
        RECT 88.210 123.990 88.380 124.160 ;
        RECT 88.210 123.630 88.380 123.800 ;
        RECT 88.210 123.270 88.380 123.440 ;
        RECT 90.430 124.730 90.600 124.900 ;
        RECT 90.430 124.370 90.600 124.540 ;
        RECT 90.430 124.010 90.600 124.180 ;
        RECT 90.430 123.650 90.600 123.820 ;
        RECT 90.430 123.290 90.600 123.460 ;
        RECT 87.660 122.930 87.830 123.100 ;
        RECT 88.865 122.850 89.035 123.020 ;
        RECT 89.225 122.850 89.395 123.020 ;
        RECT 90.430 122.930 90.600 123.100 ;
        RECT 87.660 122.570 87.830 122.740 ;
        RECT 87.660 122.210 87.830 122.380 ;
        RECT 87.660 121.850 87.830 122.020 ;
        RECT 87.660 121.490 87.830 121.660 ;
        RECT 87.660 121.130 87.830 121.300 ;
        RECT 88.210 122.430 88.380 122.600 ;
        RECT 88.210 122.070 88.380 122.240 ;
        RECT 88.210 121.710 88.380 121.880 ;
        RECT 88.210 121.350 88.380 121.520 ;
        RECT 88.210 120.990 88.380 121.160 ;
        RECT 90.430 122.570 90.600 122.740 ;
        RECT 90.430 122.210 90.600 122.380 ;
        RECT 90.430 121.850 90.600 122.020 ;
        RECT 90.430 121.490 90.600 121.660 ;
        RECT 90.430 121.130 90.600 121.300 ;
        RECT 87.660 120.770 87.830 120.940 ;
        RECT 90.430 120.770 90.600 120.940 ;
        RECT 87.660 120.410 87.830 120.580 ;
        RECT 88.865 120.570 89.035 120.740 ;
        RECT 89.225 120.570 89.395 120.740 ;
        RECT 90.430 120.410 90.600 120.580 ;
        RECT 87.660 120.050 87.830 120.220 ;
        RECT 87.660 119.690 87.830 119.860 ;
        RECT 87.660 119.330 87.830 119.500 ;
        RECT 87.660 118.970 87.830 119.140 ;
        RECT 87.660 118.610 87.830 118.780 ;
        RECT 87.660 118.250 87.830 118.420 ;
        RECT 88.210 120.185 88.380 120.355 ;
        RECT 88.210 119.825 88.380 119.995 ;
        RECT 88.210 119.465 88.380 119.635 ;
        RECT 89.880 120.185 90.050 120.355 ;
        RECT 89.880 119.825 90.050 119.995 ;
        RECT 89.880 119.465 90.050 119.635 ;
        RECT 88.865 119.290 89.035 119.460 ;
        RECT 89.225 119.290 89.395 119.460 ;
        RECT 88.210 119.105 88.380 119.275 ;
        RECT 88.210 118.745 88.380 118.915 ;
        RECT 88.210 118.385 88.380 118.555 ;
        RECT 89.880 119.105 90.050 119.275 ;
        RECT 89.880 118.745 90.050 118.915 ;
        RECT 89.880 118.385 90.050 118.555 ;
        RECT 90.430 120.050 90.600 120.220 ;
        RECT 90.430 119.690 90.600 119.860 ;
        RECT 90.430 119.330 90.600 119.500 ;
        RECT 90.430 118.970 90.600 119.140 ;
        RECT 90.430 118.610 90.600 118.780 ;
        RECT 90.430 118.250 90.600 118.420 ;
        RECT 87.660 117.890 87.830 118.060 ;
        RECT 88.865 118.010 89.035 118.180 ;
        RECT 89.225 118.010 89.395 118.180 ;
        RECT 90.430 117.890 90.600 118.060 ;
        RECT 87.960 117.340 88.130 117.510 ;
        RECT 88.320 117.340 88.490 117.510 ;
        RECT 88.680 117.340 88.850 117.510 ;
        RECT 89.040 117.340 89.210 117.510 ;
        RECT 89.400 117.340 89.570 117.510 ;
        RECT 89.760 117.340 89.930 117.510 ;
        RECT 90.120 117.340 90.290 117.510 ;
        RECT 92.215 138.040 92.385 138.210 ;
        RECT 92.575 138.040 92.745 138.210 ;
        RECT 92.935 138.040 93.105 138.210 ;
        RECT 93.295 138.040 93.465 138.210 ;
        RECT 93.655 138.040 93.825 138.210 ;
        RECT 91.915 137.690 92.085 137.860 ;
        RECT 94.185 137.690 94.355 137.860 ;
        RECT 91.915 137.330 92.085 137.500 ;
        RECT 93.050 137.370 93.220 137.540 ;
        RECT 94.185 137.330 94.355 137.500 ;
        RECT 91.915 136.970 92.085 137.140 ;
        RECT 91.915 136.610 92.085 136.780 ;
        RECT 91.915 136.250 92.085 136.420 ;
        RECT 91.915 135.890 92.085 136.060 ;
        RECT 91.915 135.530 92.085 135.700 ;
        RECT 91.915 135.170 92.085 135.340 ;
        RECT 92.465 136.985 92.635 137.155 ;
        RECT 92.465 136.625 92.635 136.795 ;
        RECT 92.465 136.265 92.635 136.435 ;
        RECT 93.635 136.985 93.805 137.155 ;
        RECT 93.635 136.625 93.805 136.795 ;
        RECT 93.635 136.265 93.805 136.435 ;
        RECT 93.050 136.090 93.220 136.260 ;
        RECT 92.465 135.905 92.635 136.075 ;
        RECT 92.465 135.545 92.635 135.715 ;
        RECT 92.465 135.185 92.635 135.355 ;
        RECT 93.635 135.905 93.805 136.075 ;
        RECT 93.635 135.545 93.805 135.715 ;
        RECT 93.635 135.185 93.805 135.355 ;
        RECT 94.185 136.970 94.355 137.140 ;
        RECT 94.185 136.610 94.355 136.780 ;
        RECT 94.185 136.250 94.355 136.420 ;
        RECT 94.185 135.890 94.355 136.060 ;
        RECT 94.185 135.530 94.355 135.700 ;
        RECT 94.185 135.170 94.355 135.340 ;
        RECT 91.915 134.810 92.085 134.980 ;
        RECT 93.050 134.810 93.220 134.980 ;
        RECT 94.185 134.810 94.355 134.980 ;
        RECT 91.915 134.450 92.085 134.620 ;
        RECT 91.915 134.090 92.085 134.260 ;
        RECT 91.915 133.730 92.085 133.900 ;
        RECT 91.915 133.370 92.085 133.540 ;
        RECT 91.915 133.010 92.085 133.180 ;
        RECT 92.465 134.390 92.635 134.560 ;
        RECT 92.465 134.030 92.635 134.200 ;
        RECT 92.465 133.670 92.635 133.840 ;
        RECT 92.465 133.310 92.635 133.480 ;
        RECT 92.465 132.950 92.635 133.120 ;
        RECT 93.635 134.390 93.805 134.560 ;
        RECT 93.635 134.030 93.805 134.200 ;
        RECT 93.635 133.670 93.805 133.840 ;
        RECT 93.635 133.310 93.805 133.480 ;
        RECT 93.635 132.950 93.805 133.120 ;
        RECT 94.185 134.450 94.355 134.620 ;
        RECT 94.185 134.090 94.355 134.260 ;
        RECT 94.185 133.730 94.355 133.900 ;
        RECT 94.185 133.370 94.355 133.540 ;
        RECT 94.185 133.010 94.355 133.180 ;
        RECT 91.915 132.650 92.085 132.820 ;
        RECT 93.050 132.530 93.220 132.700 ;
        RECT 94.185 132.650 94.355 132.820 ;
        RECT 91.915 132.290 92.085 132.460 ;
        RECT 94.185 132.290 94.355 132.460 ;
        RECT 91.915 131.930 92.085 132.100 ;
        RECT 91.915 131.570 92.085 131.740 ;
        RECT 91.915 131.210 92.085 131.380 ;
        RECT 91.915 130.850 92.085 131.020 ;
        RECT 92.465 132.110 92.635 132.280 ;
        RECT 92.465 131.750 92.635 131.920 ;
        RECT 92.465 131.390 92.635 131.560 ;
        RECT 92.465 131.030 92.635 131.200 ;
        RECT 92.465 130.670 92.635 130.840 ;
        RECT 93.635 132.110 93.805 132.280 ;
        RECT 93.635 131.750 93.805 131.920 ;
        RECT 93.635 131.390 93.805 131.560 ;
        RECT 93.635 131.030 93.805 131.200 ;
        RECT 93.635 130.670 93.805 130.840 ;
        RECT 94.185 131.930 94.355 132.100 ;
        RECT 94.185 131.570 94.355 131.740 ;
        RECT 94.185 131.210 94.355 131.380 ;
        RECT 94.185 130.850 94.355 131.020 ;
        RECT 91.915 130.490 92.085 130.660 ;
        RECT 94.185 130.490 94.355 130.660 ;
        RECT 91.915 130.130 92.085 130.300 ;
        RECT 93.050 130.250 93.220 130.420 ;
        RECT 94.185 130.130 94.355 130.300 ;
        RECT 91.915 129.770 92.085 129.940 ;
        RECT 91.915 129.410 92.085 129.580 ;
        RECT 91.915 129.050 92.085 129.220 ;
        RECT 91.915 128.690 92.085 128.860 ;
        RECT 91.915 128.330 92.085 128.500 ;
        RECT 91.915 127.970 92.085 128.140 ;
        RECT 92.465 129.865 92.635 130.035 ;
        RECT 92.465 129.505 92.635 129.675 ;
        RECT 92.465 129.145 92.635 129.315 ;
        RECT 93.635 129.865 93.805 130.035 ;
        RECT 93.635 129.505 93.805 129.675 ;
        RECT 93.635 129.145 93.805 129.315 ;
        RECT 93.050 128.970 93.220 129.140 ;
        RECT 92.465 128.785 92.635 128.955 ;
        RECT 92.465 128.425 92.635 128.595 ;
        RECT 92.465 128.065 92.635 128.235 ;
        RECT 93.635 128.785 93.805 128.955 ;
        RECT 93.635 128.425 93.805 128.595 ;
        RECT 93.635 128.065 93.805 128.235 ;
        RECT 94.185 129.770 94.355 129.940 ;
        RECT 94.185 129.410 94.355 129.580 ;
        RECT 94.185 129.050 94.355 129.220 ;
        RECT 94.185 128.690 94.355 128.860 ;
        RECT 94.185 128.330 94.355 128.500 ;
        RECT 94.185 127.970 94.355 128.140 ;
        RECT 91.915 127.610 92.085 127.780 ;
        RECT 93.050 127.690 93.220 127.860 ;
        RECT 94.185 127.610 94.355 127.780 ;
        RECT 91.915 127.250 92.085 127.420 ;
        RECT 91.915 126.890 92.085 127.060 ;
        RECT 91.915 126.530 92.085 126.700 ;
        RECT 91.915 126.170 92.085 126.340 ;
        RECT 91.915 125.810 92.085 125.980 ;
        RECT 91.915 125.450 92.085 125.620 ;
        RECT 92.465 127.305 92.635 127.475 ;
        RECT 92.465 126.945 92.635 127.115 ;
        RECT 92.465 126.585 92.635 126.755 ;
        RECT 93.635 127.305 93.805 127.475 ;
        RECT 93.635 126.945 93.805 127.115 ;
        RECT 93.635 126.585 93.805 126.755 ;
        RECT 93.050 126.410 93.220 126.580 ;
        RECT 92.465 126.225 92.635 126.395 ;
        RECT 92.465 125.865 92.635 126.035 ;
        RECT 92.465 125.505 92.635 125.675 ;
        RECT 93.635 126.225 93.805 126.395 ;
        RECT 93.635 125.865 93.805 126.035 ;
        RECT 93.635 125.505 93.805 125.675 ;
        RECT 94.185 127.250 94.355 127.420 ;
        RECT 94.185 126.890 94.355 127.060 ;
        RECT 94.185 126.530 94.355 126.700 ;
        RECT 94.185 126.170 94.355 126.340 ;
        RECT 94.185 125.810 94.355 125.980 ;
        RECT 94.185 125.450 94.355 125.620 ;
        RECT 91.915 125.090 92.085 125.260 ;
        RECT 93.050 125.130 93.220 125.300 ;
        RECT 91.915 124.730 92.085 124.900 ;
        RECT 94.185 125.090 94.355 125.260 ;
        RECT 91.915 124.370 92.085 124.540 ;
        RECT 91.915 124.010 92.085 124.180 ;
        RECT 91.915 123.650 92.085 123.820 ;
        RECT 91.915 123.290 92.085 123.460 ;
        RECT 93.635 124.710 93.805 124.880 ;
        RECT 93.635 124.350 93.805 124.520 ;
        RECT 93.635 123.990 93.805 124.160 ;
        RECT 93.635 123.630 93.805 123.800 ;
        RECT 93.635 123.270 93.805 123.440 ;
        RECT 94.185 124.730 94.355 124.900 ;
        RECT 94.185 124.370 94.355 124.540 ;
        RECT 94.185 124.010 94.355 124.180 ;
        RECT 94.185 123.650 94.355 123.820 ;
        RECT 94.185 123.290 94.355 123.460 ;
        RECT 91.915 122.930 92.085 123.100 ;
        RECT 93.050 122.850 93.220 123.020 ;
        RECT 94.185 122.930 94.355 123.100 ;
        RECT 91.915 122.570 92.085 122.740 ;
        RECT 91.915 122.210 92.085 122.380 ;
        RECT 91.915 121.850 92.085 122.020 ;
        RECT 91.915 121.490 92.085 121.660 ;
        RECT 91.915 121.130 92.085 121.300 ;
        RECT 93.635 122.430 93.805 122.600 ;
        RECT 93.635 122.070 93.805 122.240 ;
        RECT 93.635 121.710 93.805 121.880 ;
        RECT 93.635 121.350 93.805 121.520 ;
        RECT 93.635 120.990 93.805 121.160 ;
        RECT 94.185 122.570 94.355 122.740 ;
        RECT 94.185 122.210 94.355 122.380 ;
        RECT 94.185 121.850 94.355 122.020 ;
        RECT 94.185 121.490 94.355 121.660 ;
        RECT 94.185 121.130 94.355 121.300 ;
        RECT 91.915 120.770 92.085 120.940 ;
        RECT 94.185 120.770 94.355 120.940 ;
        RECT 91.915 120.410 92.085 120.580 ;
        RECT 93.050 120.570 93.220 120.740 ;
        RECT 94.185 120.410 94.355 120.580 ;
        RECT 91.915 120.050 92.085 120.220 ;
        RECT 91.915 119.690 92.085 119.860 ;
        RECT 91.915 119.330 92.085 119.500 ;
        RECT 91.915 118.970 92.085 119.140 ;
        RECT 91.915 118.610 92.085 118.780 ;
        RECT 91.915 118.250 92.085 118.420 ;
        RECT 92.465 120.185 92.635 120.355 ;
        RECT 92.465 119.825 92.635 119.995 ;
        RECT 92.465 119.465 92.635 119.635 ;
        RECT 93.635 120.185 93.805 120.355 ;
        RECT 93.635 119.825 93.805 119.995 ;
        RECT 93.635 119.465 93.805 119.635 ;
        RECT 93.050 119.290 93.220 119.460 ;
        RECT 92.465 119.105 92.635 119.275 ;
        RECT 92.465 118.745 92.635 118.915 ;
        RECT 92.465 118.385 92.635 118.555 ;
        RECT 93.635 119.105 93.805 119.275 ;
        RECT 93.635 118.745 93.805 118.915 ;
        RECT 93.635 118.385 93.805 118.555 ;
        RECT 94.185 120.050 94.355 120.220 ;
        RECT 94.185 119.690 94.355 119.860 ;
        RECT 94.185 119.330 94.355 119.500 ;
        RECT 94.185 118.970 94.355 119.140 ;
        RECT 94.185 118.610 94.355 118.780 ;
        RECT 94.185 118.250 94.355 118.420 ;
        RECT 91.915 117.890 92.085 118.060 ;
        RECT 93.050 118.010 93.220 118.180 ;
        RECT 94.185 117.890 94.355 118.060 ;
        RECT 92.215 117.340 92.385 117.510 ;
        RECT 92.575 117.340 92.745 117.510 ;
        RECT 92.935 117.340 93.105 117.510 ;
        RECT 93.295 117.340 93.465 117.510 ;
        RECT 93.655 117.340 93.825 117.510 ;
        RECT 96.080 137.940 96.250 138.110 ;
        RECT 96.080 137.580 96.250 137.750 ;
        RECT 96.080 137.220 96.250 137.390 ;
        RECT 96.630 138.640 96.800 138.810 ;
        RECT 96.630 138.280 96.800 138.450 ;
        RECT 96.630 137.920 96.800 138.090 ;
        RECT 96.630 137.560 96.800 137.730 ;
        RECT 96.630 137.200 96.800 137.370 ;
        RECT 98.300 138.640 98.470 138.810 ;
        RECT 98.300 138.280 98.470 138.450 ;
        RECT 98.300 137.920 98.470 138.090 ;
        RECT 98.300 137.560 98.470 137.730 ;
        RECT 98.300 137.200 98.470 137.370 ;
        RECT 100.220 138.640 100.390 138.810 ;
        RECT 100.220 138.280 100.390 138.450 ;
        RECT 100.220 137.920 100.390 138.090 ;
        RECT 100.220 137.560 100.390 137.730 ;
        RECT 100.220 137.200 100.390 137.370 ;
        RECT 102.440 138.660 102.610 138.830 ;
        RECT 102.440 138.300 102.610 138.470 ;
        RECT 102.440 137.940 102.610 138.110 ;
        RECT 102.440 137.580 102.610 137.750 ;
        RECT 102.440 137.220 102.610 137.390 ;
        RECT 96.080 136.860 96.250 137.030 ;
        RECT 97.285 136.780 97.455 136.950 ;
        RECT 97.645 136.780 97.815 136.950 ;
        RECT 100.875 136.780 101.045 136.950 ;
        RECT 101.235 136.780 101.405 136.950 ;
        RECT 102.440 136.860 102.610 137.030 ;
        RECT 96.080 136.500 96.250 136.670 ;
        RECT 96.080 136.140 96.250 136.310 ;
        RECT 96.080 135.780 96.250 135.950 ;
        RECT 96.080 135.420 96.250 135.590 ;
        RECT 96.080 135.060 96.250 135.230 ;
        RECT 96.630 136.360 96.800 136.530 ;
        RECT 96.630 136.000 96.800 136.170 ;
        RECT 96.630 135.640 96.800 135.810 ;
        RECT 96.630 135.280 96.800 135.450 ;
        RECT 96.630 134.920 96.800 135.090 ;
        RECT 98.300 136.360 98.470 136.530 ;
        RECT 98.300 136.000 98.470 136.170 ;
        RECT 98.300 135.640 98.470 135.810 ;
        RECT 98.300 135.280 98.470 135.450 ;
        RECT 98.300 134.920 98.470 135.090 ;
        RECT 100.220 136.360 100.390 136.530 ;
        RECT 100.220 136.000 100.390 136.170 ;
        RECT 100.220 135.640 100.390 135.810 ;
        RECT 100.220 135.280 100.390 135.450 ;
        RECT 100.220 134.920 100.390 135.090 ;
        RECT 102.440 136.500 102.610 136.670 ;
        RECT 102.440 136.140 102.610 136.310 ;
        RECT 102.440 135.780 102.610 135.950 ;
        RECT 102.440 135.420 102.610 135.590 ;
        RECT 102.440 135.060 102.610 135.230 ;
        RECT 96.080 134.700 96.250 134.870 ;
        RECT 102.440 134.700 102.610 134.870 ;
        RECT 96.080 134.340 96.250 134.510 ;
        RECT 97.285 134.500 97.455 134.670 ;
        RECT 97.645 134.500 97.815 134.670 ;
        RECT 100.875 134.500 101.045 134.670 ;
        RECT 101.235 134.500 101.405 134.670 ;
        RECT 102.440 134.340 102.610 134.510 ;
        RECT 96.080 133.980 96.250 134.150 ;
        RECT 96.080 133.620 96.250 133.790 ;
        RECT 96.080 133.260 96.250 133.430 ;
        RECT 96.080 132.900 96.250 133.070 ;
        RECT 96.080 132.540 96.250 132.710 ;
        RECT 96.630 134.080 96.800 134.250 ;
        RECT 96.630 133.720 96.800 133.890 ;
        RECT 96.630 133.360 96.800 133.530 ;
        RECT 96.630 133.000 96.800 133.170 ;
        RECT 96.630 132.640 96.800 132.810 ;
        RECT 98.300 134.080 98.470 134.250 ;
        RECT 98.300 133.720 98.470 133.890 ;
        RECT 98.300 133.360 98.470 133.530 ;
        RECT 98.300 133.000 98.470 133.170 ;
        RECT 98.300 132.640 98.470 132.810 ;
        RECT 100.220 134.080 100.390 134.250 ;
        RECT 100.220 133.720 100.390 133.890 ;
        RECT 100.220 133.360 100.390 133.530 ;
        RECT 100.220 133.000 100.390 133.170 ;
        RECT 100.220 132.640 100.390 132.810 ;
        RECT 102.440 133.980 102.610 134.150 ;
        RECT 102.440 133.620 102.610 133.790 ;
        RECT 102.440 133.260 102.610 133.430 ;
        RECT 102.440 132.900 102.610 133.070 ;
        RECT 102.440 132.540 102.610 132.710 ;
        RECT 96.080 132.180 96.250 132.350 ;
        RECT 97.285 132.220 97.455 132.390 ;
        RECT 97.645 132.220 97.815 132.390 ;
        RECT 100.875 132.220 101.045 132.390 ;
        RECT 101.235 132.220 101.405 132.390 ;
        RECT 96.080 131.820 96.250 131.990 ;
        RECT 102.440 132.180 102.610 132.350 ;
        RECT 96.080 131.460 96.250 131.630 ;
        RECT 96.080 131.100 96.250 131.270 ;
        RECT 96.080 130.740 96.250 130.910 ;
        RECT 96.080 130.380 96.250 130.550 ;
        RECT 96.630 131.800 96.800 131.970 ;
        RECT 96.630 131.440 96.800 131.610 ;
        RECT 96.630 131.080 96.800 131.250 ;
        RECT 96.630 130.720 96.800 130.890 ;
        RECT 96.630 130.360 96.800 130.530 ;
        RECT 98.300 131.800 98.470 131.970 ;
        RECT 98.300 131.440 98.470 131.610 ;
        RECT 98.300 131.080 98.470 131.250 ;
        RECT 98.300 130.720 98.470 130.890 ;
        RECT 98.300 130.360 98.470 130.530 ;
        RECT 100.220 131.800 100.390 131.970 ;
        RECT 100.220 131.440 100.390 131.610 ;
        RECT 100.220 131.080 100.390 131.250 ;
        RECT 100.220 130.720 100.390 130.890 ;
        RECT 100.220 130.360 100.390 130.530 ;
        RECT 102.440 131.820 102.610 131.990 ;
        RECT 102.440 131.460 102.610 131.630 ;
        RECT 102.440 131.100 102.610 131.270 ;
        RECT 102.440 130.740 102.610 130.910 ;
        RECT 102.440 130.380 102.610 130.550 ;
        RECT 96.080 130.020 96.250 130.190 ;
        RECT 97.285 129.940 97.455 130.110 ;
        RECT 97.645 129.940 97.815 130.110 ;
        RECT 100.875 129.940 101.045 130.110 ;
        RECT 101.235 129.940 101.405 130.110 ;
        RECT 102.440 130.020 102.610 130.190 ;
        RECT 96.080 129.660 96.250 129.830 ;
        RECT 96.080 129.300 96.250 129.470 ;
        RECT 96.080 128.940 96.250 129.110 ;
        RECT 96.080 128.580 96.250 128.750 ;
        RECT 96.080 128.220 96.250 128.390 ;
        RECT 96.630 129.520 96.800 129.690 ;
        RECT 96.630 129.160 96.800 129.330 ;
        RECT 96.630 128.800 96.800 128.970 ;
        RECT 96.630 128.440 96.800 128.610 ;
        RECT 96.630 128.080 96.800 128.250 ;
        RECT 98.300 129.520 98.470 129.690 ;
        RECT 98.300 129.160 98.470 129.330 ;
        RECT 98.300 128.800 98.470 128.970 ;
        RECT 98.300 128.440 98.470 128.610 ;
        RECT 98.300 128.080 98.470 128.250 ;
        RECT 101.890 129.520 102.060 129.690 ;
        RECT 101.890 129.160 102.060 129.330 ;
        RECT 101.890 128.800 102.060 128.970 ;
        RECT 101.890 128.440 102.060 128.610 ;
        RECT 101.890 128.080 102.060 128.250 ;
        RECT 102.440 129.660 102.610 129.830 ;
        RECT 102.440 129.300 102.610 129.470 ;
        RECT 102.440 128.940 102.610 129.110 ;
        RECT 102.440 128.580 102.610 128.750 ;
        RECT 102.440 128.220 102.610 128.390 ;
        RECT 96.080 127.860 96.250 128.030 ;
        RECT 102.440 127.860 102.610 128.030 ;
        RECT 96.080 127.500 96.250 127.670 ;
        RECT 97.285 127.660 97.455 127.830 ;
        RECT 97.645 127.660 97.815 127.830 ;
        RECT 100.875 127.660 101.045 127.830 ;
        RECT 101.235 127.660 101.405 127.830 ;
        RECT 102.440 127.500 102.610 127.670 ;
        RECT 96.080 127.140 96.250 127.310 ;
        RECT 96.080 126.780 96.250 126.950 ;
        RECT 96.080 126.420 96.250 126.590 ;
        RECT 96.080 126.060 96.250 126.230 ;
        RECT 96.080 125.700 96.250 125.870 ;
        RECT 96.630 127.240 96.800 127.410 ;
        RECT 96.630 126.880 96.800 127.050 ;
        RECT 96.630 126.520 96.800 126.690 ;
        RECT 96.630 126.160 96.800 126.330 ;
        RECT 96.630 125.800 96.800 125.970 ;
        RECT 98.300 127.240 98.470 127.410 ;
        RECT 98.300 126.880 98.470 127.050 ;
        RECT 98.300 126.520 98.470 126.690 ;
        RECT 98.300 126.160 98.470 126.330 ;
        RECT 98.300 125.800 98.470 125.970 ;
        RECT 101.890 127.240 102.060 127.410 ;
        RECT 101.890 126.880 102.060 127.050 ;
        RECT 101.890 126.520 102.060 126.690 ;
        RECT 101.890 126.160 102.060 126.330 ;
        RECT 101.890 125.800 102.060 125.970 ;
        RECT 102.440 127.140 102.610 127.310 ;
        RECT 102.440 126.780 102.610 126.950 ;
        RECT 102.440 126.420 102.610 126.590 ;
        RECT 102.440 126.060 102.610 126.230 ;
        RECT 102.440 125.700 102.610 125.870 ;
        RECT 96.080 125.340 96.250 125.510 ;
        RECT 97.285 125.380 97.455 125.550 ;
        RECT 97.645 125.380 97.815 125.550 ;
        RECT 100.875 125.380 101.045 125.550 ;
        RECT 101.235 125.380 101.405 125.550 ;
        RECT 96.080 124.980 96.250 125.150 ;
        RECT 102.440 125.340 102.610 125.510 ;
        RECT 96.080 124.620 96.250 124.790 ;
        RECT 96.080 124.260 96.250 124.430 ;
        RECT 96.080 123.900 96.250 124.070 ;
        RECT 96.080 123.540 96.250 123.710 ;
        RECT 96.630 124.960 96.800 125.130 ;
        RECT 96.630 124.600 96.800 124.770 ;
        RECT 96.630 124.240 96.800 124.410 ;
        RECT 96.630 123.880 96.800 124.050 ;
        RECT 96.630 123.520 96.800 123.690 ;
        RECT 98.300 124.960 98.470 125.130 ;
        RECT 98.300 124.600 98.470 124.770 ;
        RECT 98.300 124.240 98.470 124.410 ;
        RECT 98.300 123.880 98.470 124.050 ;
        RECT 98.300 123.520 98.470 123.690 ;
        RECT 100.220 124.960 100.390 125.130 ;
        RECT 100.220 124.600 100.390 124.770 ;
        RECT 100.220 124.240 100.390 124.410 ;
        RECT 100.220 123.880 100.390 124.050 ;
        RECT 100.220 123.520 100.390 123.690 ;
        RECT 102.440 124.980 102.610 125.150 ;
        RECT 102.440 124.620 102.610 124.790 ;
        RECT 102.440 124.260 102.610 124.430 ;
        RECT 102.440 123.900 102.610 124.070 ;
        RECT 102.440 123.540 102.610 123.710 ;
        RECT 96.080 123.180 96.250 123.350 ;
        RECT 97.285 123.100 97.455 123.270 ;
        RECT 97.645 123.100 97.815 123.270 ;
        RECT 100.875 123.100 101.045 123.270 ;
        RECT 101.235 123.100 101.405 123.270 ;
        RECT 102.440 123.180 102.610 123.350 ;
        RECT 96.080 122.820 96.250 122.990 ;
        RECT 96.080 122.460 96.250 122.630 ;
        RECT 96.080 122.100 96.250 122.270 ;
        RECT 96.080 121.740 96.250 121.910 ;
        RECT 96.080 121.380 96.250 121.550 ;
        RECT 96.630 122.680 96.800 122.850 ;
        RECT 96.630 122.320 96.800 122.490 ;
        RECT 96.630 121.960 96.800 122.130 ;
        RECT 96.630 121.600 96.800 121.770 ;
        RECT 96.630 121.240 96.800 121.410 ;
        RECT 98.300 122.680 98.470 122.850 ;
        RECT 98.300 122.320 98.470 122.490 ;
        RECT 98.300 121.960 98.470 122.130 ;
        RECT 98.300 121.600 98.470 121.770 ;
        RECT 98.300 121.240 98.470 121.410 ;
        RECT 100.220 122.680 100.390 122.850 ;
        RECT 100.220 122.320 100.390 122.490 ;
        RECT 100.220 121.960 100.390 122.130 ;
        RECT 100.220 121.600 100.390 121.770 ;
        RECT 100.220 121.240 100.390 121.410 ;
        RECT 102.440 122.820 102.610 122.990 ;
        RECT 102.440 122.460 102.610 122.630 ;
        RECT 102.440 122.100 102.610 122.270 ;
        RECT 102.440 121.740 102.610 121.910 ;
        RECT 102.440 121.380 102.610 121.550 ;
        RECT 96.080 121.020 96.250 121.190 ;
        RECT 102.440 121.020 102.610 121.190 ;
        RECT 96.080 120.660 96.250 120.830 ;
        RECT 97.285 120.820 97.455 120.990 ;
        RECT 97.645 120.820 97.815 120.990 ;
        RECT 100.875 120.820 101.045 120.990 ;
        RECT 101.235 120.820 101.405 120.990 ;
        RECT 102.440 120.660 102.610 120.830 ;
        RECT 96.080 120.300 96.250 120.470 ;
        RECT 96.080 119.940 96.250 120.110 ;
        RECT 96.080 119.580 96.250 119.750 ;
        RECT 96.080 119.220 96.250 119.390 ;
        RECT 96.080 118.860 96.250 119.030 ;
        RECT 96.630 120.400 96.800 120.570 ;
        RECT 96.630 120.040 96.800 120.210 ;
        RECT 96.630 119.680 96.800 119.850 ;
        RECT 96.630 119.320 96.800 119.490 ;
        RECT 96.630 118.960 96.800 119.130 ;
        RECT 98.300 120.400 98.470 120.570 ;
        RECT 98.300 120.040 98.470 120.210 ;
        RECT 98.300 119.680 98.470 119.850 ;
        RECT 98.300 119.320 98.470 119.490 ;
        RECT 98.300 118.960 98.470 119.130 ;
        RECT 100.220 120.400 100.390 120.570 ;
        RECT 100.220 120.040 100.390 120.210 ;
        RECT 100.220 119.680 100.390 119.850 ;
        RECT 100.220 119.320 100.390 119.490 ;
        RECT 100.220 118.960 100.390 119.130 ;
        RECT 102.440 120.300 102.610 120.470 ;
        RECT 102.440 119.940 102.610 120.110 ;
        RECT 102.440 119.580 102.610 119.750 ;
        RECT 102.440 119.220 102.610 119.390 ;
        RECT 102.440 118.860 102.610 119.030 ;
        RECT 96.080 118.500 96.250 118.670 ;
        RECT 97.285 118.540 97.455 118.710 ;
        RECT 97.645 118.540 97.815 118.710 ;
        RECT 100.875 118.540 101.045 118.710 ;
        RECT 101.235 118.540 101.405 118.710 ;
        RECT 96.080 118.140 96.250 118.310 ;
        RECT 102.440 118.500 102.610 118.670 ;
        RECT 96.080 117.780 96.250 117.950 ;
        RECT 96.080 117.420 96.250 117.590 ;
        RECT 86.030 116.980 86.200 117.150 ;
        RECT 86.030 116.620 86.200 116.790 ;
        RECT 82.740 115.995 82.910 116.165 ;
        RECT 86.030 116.260 86.200 116.430 ;
        RECT 84.895 115.980 85.065 116.150 ;
        RECT 82.740 115.635 82.910 115.805 ;
        RECT 86.030 115.900 86.200 116.070 ;
        RECT 82.740 115.275 82.910 115.445 ;
        RECT 82.740 114.915 82.910 115.085 ;
        RECT 82.740 114.555 82.910 114.725 ;
        RECT 82.740 114.195 82.910 114.365 ;
        RECT 84.310 115.595 84.480 115.765 ;
        RECT 84.310 115.235 84.480 115.405 ;
        RECT 84.310 114.875 84.480 115.045 ;
        RECT 86.030 115.540 86.200 115.710 ;
        RECT 86.030 115.180 86.200 115.350 ;
        RECT 84.895 114.700 85.065 114.870 ;
        RECT 86.030 114.820 86.200 114.990 ;
        RECT 84.310 114.515 84.480 114.685 ;
        RECT 84.310 114.155 84.480 114.325 ;
        RECT 81.020 113.740 81.190 113.910 ;
        RECT 82.155 113.820 82.325 113.990 ;
        RECT 84.310 113.795 84.480 113.965 ;
        RECT 86.030 114.460 86.200 114.630 ;
        RECT 86.030 114.100 86.200 114.270 ;
        RECT 86.030 113.740 86.200 113.910 ;
        RECT 81.020 113.380 81.190 113.550 ;
        RECT 84.895 113.420 85.065 113.590 ;
        RECT 86.030 113.380 86.200 113.550 ;
        RECT 96.080 117.060 96.250 117.230 ;
        RECT 96.080 116.700 96.250 116.870 ;
        RECT 96.630 118.120 96.800 118.290 ;
        RECT 96.630 117.760 96.800 117.930 ;
        RECT 96.630 117.400 96.800 117.570 ;
        RECT 96.630 117.040 96.800 117.210 ;
        RECT 96.630 116.680 96.800 116.850 ;
        RECT 98.300 118.120 98.470 118.290 ;
        RECT 98.300 117.760 98.470 117.930 ;
        RECT 98.300 117.400 98.470 117.570 ;
        RECT 98.300 117.040 98.470 117.210 ;
        RECT 98.300 116.680 98.470 116.850 ;
        RECT 100.220 118.120 100.390 118.290 ;
        RECT 100.220 117.760 100.390 117.930 ;
        RECT 100.220 117.400 100.390 117.570 ;
        RECT 100.220 117.040 100.390 117.210 ;
        RECT 100.220 116.680 100.390 116.850 ;
        RECT 102.440 118.140 102.610 118.310 ;
        RECT 102.440 117.780 102.610 117.950 ;
        RECT 102.440 117.420 102.610 117.590 ;
        RECT 102.440 117.060 102.610 117.230 ;
        RECT 102.440 116.700 102.610 116.870 ;
        RECT 96.080 116.340 96.250 116.510 ;
        RECT 97.285 116.260 97.455 116.430 ;
        RECT 97.645 116.260 97.815 116.430 ;
        RECT 100.875 116.260 101.045 116.430 ;
        RECT 101.235 116.260 101.405 116.430 ;
        RECT 102.440 116.340 102.610 116.510 ;
        RECT 96.080 115.980 96.250 116.150 ;
        RECT 96.080 115.620 96.250 115.790 ;
        RECT 96.080 115.260 96.250 115.430 ;
        RECT 96.080 114.900 96.250 115.070 ;
        RECT 96.080 114.540 96.250 114.710 ;
        RECT 96.630 115.840 96.800 116.010 ;
        RECT 96.630 115.480 96.800 115.650 ;
        RECT 96.630 115.120 96.800 115.290 ;
        RECT 96.630 114.760 96.800 114.930 ;
        RECT 96.630 114.400 96.800 114.570 ;
        RECT 98.300 115.840 98.470 116.010 ;
        RECT 98.300 115.480 98.470 115.650 ;
        RECT 98.300 115.120 98.470 115.290 ;
        RECT 98.300 114.760 98.470 114.930 ;
        RECT 98.300 114.400 98.470 114.570 ;
        RECT 100.220 115.840 100.390 116.010 ;
        RECT 100.220 115.480 100.390 115.650 ;
        RECT 100.220 115.120 100.390 115.290 ;
        RECT 100.220 114.760 100.390 114.930 ;
        RECT 100.220 114.400 100.390 114.570 ;
        RECT 102.440 115.980 102.610 116.150 ;
        RECT 102.440 115.620 102.610 115.790 ;
        RECT 102.440 115.260 102.610 115.430 ;
        RECT 102.440 114.900 102.610 115.070 ;
        RECT 102.440 114.540 102.610 114.710 ;
        RECT 96.080 114.180 96.250 114.350 ;
        RECT 102.440 114.180 102.610 114.350 ;
        RECT 96.080 113.820 96.250 113.990 ;
        RECT 97.285 113.980 97.455 114.150 ;
        RECT 97.645 113.980 97.815 114.150 ;
        RECT 100.875 113.980 101.045 114.150 ;
        RECT 101.235 113.980 101.405 114.150 ;
        RECT 102.440 113.820 102.610 113.990 ;
        RECT 96.080 113.460 96.250 113.630 ;
        RECT 98.300 113.560 98.470 113.730 ;
        RECT 81.320 112.790 81.490 112.960 ;
        RECT 81.680 112.790 81.850 112.960 ;
        RECT 82.040 112.790 82.210 112.960 ;
        RECT 82.400 112.790 82.570 112.960 ;
        RECT 82.760 112.790 82.930 112.960 ;
        RECT 83.120 112.790 83.290 112.960 ;
        RECT 83.480 112.790 83.650 112.960 ;
        RECT 83.840 112.790 84.010 112.960 ;
        RECT 84.200 112.790 84.370 112.960 ;
        RECT 84.560 112.790 84.730 112.960 ;
        RECT 84.920 112.790 85.090 112.960 ;
        RECT 85.280 112.790 85.450 112.960 ;
        RECT 85.640 112.790 85.810 112.960 ;
        RECT 88.845 113.090 89.015 113.260 ;
        RECT 89.205 113.090 89.375 113.260 ;
        RECT 89.565 113.090 89.735 113.260 ;
        RECT 89.925 113.090 90.095 113.260 ;
        RECT 90.285 113.090 90.455 113.260 ;
        RECT 90.645 113.090 90.815 113.260 ;
        RECT 92.115 113.090 92.285 113.260 ;
        RECT 92.475 113.090 92.645 113.260 ;
        RECT 92.835 113.090 93.005 113.260 ;
        RECT 93.195 113.090 93.365 113.260 ;
        RECT 93.555 113.090 93.725 113.260 ;
        RECT 93.915 113.090 94.085 113.260 ;
        RECT 94.275 113.090 94.445 113.260 ;
        RECT 94.635 113.090 94.805 113.260 ;
        RECT 63.685 112.380 63.855 112.550 ;
        RECT 64.550 112.420 64.720 112.590 ;
        RECT 64.910 112.420 65.080 112.590 ;
        RECT 69.280 112.420 69.450 112.590 ;
        RECT 63.685 112.020 63.855 112.190 ;
        RECT 70.075 112.380 70.245 112.550 ;
        RECT 63.685 111.660 63.855 111.830 ;
        RECT 63.685 111.300 63.855 111.470 ;
        RECT 63.685 110.940 63.855 111.110 ;
        RECT 63.685 110.580 63.855 110.750 ;
        RECT 65.565 112.000 65.735 112.170 ;
        RECT 65.565 111.640 65.735 111.810 ;
        RECT 65.565 111.280 65.735 111.450 ;
        RECT 65.565 110.920 65.735 111.090 ;
        RECT 65.565 110.560 65.735 110.730 ;
        RECT 68.695 112.000 68.865 112.170 ;
        RECT 68.695 111.640 68.865 111.810 ;
        RECT 68.695 111.280 68.865 111.450 ;
        RECT 68.695 110.920 68.865 111.090 ;
        RECT 68.695 110.560 68.865 110.730 ;
        RECT 70.075 112.020 70.245 112.190 ;
        RECT 70.075 111.660 70.245 111.830 ;
        RECT 70.075 111.300 70.245 111.470 ;
        RECT 70.075 110.940 70.245 111.110 ;
        RECT 70.075 110.580 70.245 110.750 ;
        RECT 63.685 110.220 63.855 110.390 ;
        RECT 64.550 110.140 64.720 110.310 ;
        RECT 64.910 110.140 65.080 110.310 ;
        RECT 69.280 110.140 69.450 110.310 ;
        RECT 70.075 110.220 70.245 110.390 ;
        RECT 63.685 109.860 63.855 110.030 ;
        RECT 63.685 109.500 63.855 109.670 ;
        RECT 63.685 109.140 63.855 109.310 ;
        RECT 63.685 108.780 63.855 108.950 ;
        RECT 63.685 108.420 63.855 108.590 ;
        RECT 65.565 109.720 65.735 109.890 ;
        RECT 65.565 109.360 65.735 109.530 ;
        RECT 65.565 109.000 65.735 109.170 ;
        RECT 65.565 108.640 65.735 108.810 ;
        RECT 65.565 108.280 65.735 108.450 ;
        RECT 68.695 109.720 68.865 109.890 ;
        RECT 68.695 109.360 68.865 109.530 ;
        RECT 68.695 109.000 68.865 109.170 ;
        RECT 68.695 108.640 68.865 108.810 ;
        RECT 68.695 108.280 68.865 108.450 ;
        RECT 70.075 109.860 70.245 110.030 ;
        RECT 70.075 109.500 70.245 109.670 ;
        RECT 70.075 109.140 70.245 109.310 ;
        RECT 70.075 108.780 70.245 108.950 ;
        RECT 70.075 108.420 70.245 108.590 ;
        RECT 63.685 108.060 63.855 108.230 ;
        RECT 70.075 108.060 70.245 108.230 ;
        RECT 63.685 107.700 63.855 107.870 ;
        RECT 64.550 107.860 64.720 108.030 ;
        RECT 64.910 107.860 65.080 108.030 ;
        RECT 69.280 107.860 69.450 108.030 ;
        RECT 70.075 107.700 70.245 107.870 ;
        RECT 63.685 107.340 63.855 107.510 ;
        RECT 63.685 106.980 63.855 107.150 ;
        RECT 63.685 106.620 63.855 106.790 ;
        RECT 63.685 106.260 63.855 106.430 ;
        RECT 63.685 105.900 63.855 106.070 ;
        RECT 65.565 107.440 65.735 107.610 ;
        RECT 65.565 107.080 65.735 107.250 ;
        RECT 65.565 106.720 65.735 106.890 ;
        RECT 65.565 106.360 65.735 106.530 ;
        RECT 65.565 106.000 65.735 106.170 ;
        RECT 68.695 107.440 68.865 107.610 ;
        RECT 68.695 107.080 68.865 107.250 ;
        RECT 68.695 106.720 68.865 106.890 ;
        RECT 68.695 106.360 68.865 106.530 ;
        RECT 68.695 106.000 68.865 106.170 ;
        RECT 70.075 107.340 70.245 107.510 ;
        RECT 70.075 106.980 70.245 107.150 ;
        RECT 70.075 106.620 70.245 106.790 ;
        RECT 70.075 106.260 70.245 106.430 ;
        RECT 70.075 105.900 70.245 106.070 ;
        RECT 63.685 105.540 63.855 105.710 ;
        RECT 64.550 105.580 64.720 105.750 ;
        RECT 64.910 105.580 65.080 105.750 ;
        RECT 69.280 105.580 69.450 105.750 ;
        RECT 63.685 105.180 63.855 105.350 ;
        RECT 70.075 105.540 70.245 105.710 ;
        RECT 63.685 104.820 63.855 104.990 ;
        RECT 63.685 104.460 63.855 104.630 ;
        RECT 63.685 104.100 63.855 104.270 ;
        RECT 63.685 103.740 63.855 103.910 ;
        RECT 65.565 105.160 65.735 105.330 ;
        RECT 65.565 104.800 65.735 104.970 ;
        RECT 65.565 104.440 65.735 104.610 ;
        RECT 65.565 104.080 65.735 104.250 ;
        RECT 65.565 103.720 65.735 103.890 ;
        RECT 68.695 105.160 68.865 105.330 ;
        RECT 68.695 104.800 68.865 104.970 ;
        RECT 68.695 104.440 68.865 104.610 ;
        RECT 68.695 104.080 68.865 104.250 ;
        RECT 68.695 103.720 68.865 103.890 ;
        RECT 70.075 105.180 70.245 105.350 ;
        RECT 70.075 104.820 70.245 104.990 ;
        RECT 70.075 104.460 70.245 104.630 ;
        RECT 70.075 104.100 70.245 104.270 ;
        RECT 70.075 103.740 70.245 103.910 ;
        RECT 63.685 103.380 63.855 103.550 ;
        RECT 64.550 103.300 64.720 103.470 ;
        RECT 64.910 103.300 65.080 103.470 ;
        RECT 69.280 103.300 69.450 103.470 ;
        RECT 70.075 103.380 70.245 103.550 ;
        RECT 63.685 103.020 63.855 103.190 ;
        RECT 63.685 102.660 63.855 102.830 ;
        RECT 63.685 102.300 63.855 102.470 ;
        RECT 63.685 101.940 63.855 102.110 ;
        RECT 63.685 101.580 63.855 101.750 ;
        RECT 65.565 102.880 65.735 103.050 ;
        RECT 65.565 102.520 65.735 102.690 ;
        RECT 65.565 102.160 65.735 102.330 ;
        RECT 65.565 101.800 65.735 101.970 ;
        RECT 65.565 101.440 65.735 101.610 ;
        RECT 68.695 102.880 68.865 103.050 ;
        RECT 68.695 102.520 68.865 102.690 ;
        RECT 68.695 102.160 68.865 102.330 ;
        RECT 68.695 101.800 68.865 101.970 ;
        RECT 68.695 101.440 68.865 101.610 ;
        RECT 70.075 103.020 70.245 103.190 ;
        RECT 70.075 102.660 70.245 102.830 ;
        RECT 70.075 102.300 70.245 102.470 ;
        RECT 70.075 101.940 70.245 102.110 ;
        RECT 70.075 101.580 70.245 101.750 ;
        RECT 63.685 101.220 63.855 101.390 ;
        RECT 70.075 101.220 70.245 101.390 ;
        RECT 63.685 100.860 63.855 101.030 ;
        RECT 64.550 101.020 64.720 101.190 ;
        RECT 64.910 101.020 65.080 101.190 ;
        RECT 69.280 101.020 69.450 101.190 ;
        RECT 70.075 100.860 70.245 101.030 ;
        RECT 63.685 100.500 63.855 100.670 ;
        RECT 63.685 100.140 63.855 100.310 ;
        RECT 63.685 99.780 63.855 99.950 ;
        RECT 63.685 99.420 63.855 99.590 ;
        RECT 63.685 99.060 63.855 99.230 ;
        RECT 65.565 100.600 65.735 100.770 ;
        RECT 65.565 100.240 65.735 100.410 ;
        RECT 65.565 99.880 65.735 100.050 ;
        RECT 65.565 99.520 65.735 99.690 ;
        RECT 65.565 99.160 65.735 99.330 ;
        RECT 68.695 100.600 68.865 100.770 ;
        RECT 68.695 100.240 68.865 100.410 ;
        RECT 68.695 99.880 68.865 100.050 ;
        RECT 68.695 99.520 68.865 99.690 ;
        RECT 68.695 99.160 68.865 99.330 ;
        RECT 70.075 100.500 70.245 100.670 ;
        RECT 70.075 100.140 70.245 100.310 ;
        RECT 70.075 99.780 70.245 99.950 ;
        RECT 70.075 99.420 70.245 99.590 ;
        RECT 70.075 99.060 70.245 99.230 ;
        RECT 63.685 98.700 63.855 98.870 ;
        RECT 64.550 98.740 64.720 98.910 ;
        RECT 64.910 98.740 65.080 98.910 ;
        RECT 69.280 98.740 69.450 98.910 ;
        RECT 63.685 98.340 63.855 98.510 ;
        RECT 70.075 98.700 70.245 98.870 ;
        RECT 63.685 97.980 63.855 98.150 ;
        RECT 63.685 97.620 63.855 97.790 ;
        RECT 63.685 97.260 63.855 97.430 ;
        RECT 63.685 96.900 63.855 97.070 ;
        RECT 65.565 98.320 65.735 98.490 ;
        RECT 65.565 97.960 65.735 98.130 ;
        RECT 65.565 97.600 65.735 97.770 ;
        RECT 65.565 97.240 65.735 97.410 ;
        RECT 65.565 96.880 65.735 97.050 ;
        RECT 68.695 98.320 68.865 98.490 ;
        RECT 68.695 97.960 68.865 98.130 ;
        RECT 68.695 97.600 68.865 97.770 ;
        RECT 68.695 97.240 68.865 97.410 ;
        RECT 68.695 96.880 68.865 97.050 ;
        RECT 70.075 98.340 70.245 98.510 ;
        RECT 70.075 97.980 70.245 98.150 ;
        RECT 70.075 97.620 70.245 97.790 ;
        RECT 70.075 97.260 70.245 97.430 ;
        RECT 70.075 96.900 70.245 97.070 ;
        RECT 63.685 96.540 63.855 96.710 ;
        RECT 64.550 96.460 64.720 96.630 ;
        RECT 64.910 96.460 65.080 96.630 ;
        RECT 69.280 96.460 69.450 96.630 ;
        RECT 70.075 96.540 70.245 96.710 ;
        RECT 63.685 96.180 63.855 96.350 ;
        RECT 63.685 95.820 63.855 95.990 ;
        RECT 63.685 95.460 63.855 95.630 ;
        RECT 63.685 95.100 63.855 95.270 ;
        RECT 63.685 94.740 63.855 94.910 ;
        RECT 65.565 96.040 65.735 96.210 ;
        RECT 65.565 95.680 65.735 95.850 ;
        RECT 65.565 95.320 65.735 95.490 ;
        RECT 65.565 94.960 65.735 95.130 ;
        RECT 65.565 94.600 65.735 94.770 ;
        RECT 68.695 96.040 68.865 96.210 ;
        RECT 68.695 95.680 68.865 95.850 ;
        RECT 68.695 95.320 68.865 95.490 ;
        RECT 68.695 94.960 68.865 95.130 ;
        RECT 68.695 94.600 68.865 94.770 ;
        RECT 70.075 96.180 70.245 96.350 ;
        RECT 70.075 95.820 70.245 95.990 ;
        RECT 70.075 95.460 70.245 95.630 ;
        RECT 70.075 95.100 70.245 95.270 ;
        RECT 70.075 94.740 70.245 94.910 ;
        RECT 63.685 94.380 63.855 94.550 ;
        RECT 70.075 94.380 70.245 94.550 ;
        RECT 63.685 94.020 63.855 94.190 ;
        RECT 64.550 94.180 64.720 94.350 ;
        RECT 64.910 94.180 65.080 94.350 ;
        RECT 69.280 94.180 69.450 94.350 ;
        RECT 70.075 94.020 70.245 94.190 ;
        RECT 63.685 93.660 63.855 93.830 ;
        RECT 63.685 93.300 63.855 93.470 ;
        RECT 63.685 92.940 63.855 93.110 ;
        RECT 63.685 92.580 63.855 92.750 ;
        RECT 63.685 92.220 63.855 92.390 ;
        RECT 65.565 93.760 65.735 93.930 ;
        RECT 65.565 93.400 65.735 93.570 ;
        RECT 65.565 93.040 65.735 93.210 ;
        RECT 65.565 92.680 65.735 92.850 ;
        RECT 65.565 92.320 65.735 92.490 ;
        RECT 68.695 93.760 68.865 93.930 ;
        RECT 68.695 93.400 68.865 93.570 ;
        RECT 68.695 93.040 68.865 93.210 ;
        RECT 68.695 92.680 68.865 92.850 ;
        RECT 68.695 92.320 68.865 92.490 ;
        RECT 70.075 93.660 70.245 93.830 ;
        RECT 70.075 93.300 70.245 93.470 ;
        RECT 70.075 92.940 70.245 93.110 ;
        RECT 70.075 92.580 70.245 92.750 ;
        RECT 70.075 92.220 70.245 92.390 ;
        RECT 63.685 91.860 63.855 92.030 ;
        RECT 64.550 91.900 64.720 92.070 ;
        RECT 64.910 91.900 65.080 92.070 ;
        RECT 69.280 91.900 69.450 92.070 ;
        RECT 63.685 91.500 63.855 91.670 ;
        RECT 70.075 91.860 70.245 92.030 ;
        RECT 63.685 91.140 63.855 91.310 ;
        RECT 63.685 90.780 63.855 90.950 ;
        RECT 63.685 90.420 63.855 90.590 ;
        RECT 63.685 90.060 63.855 90.230 ;
        RECT 65.565 91.480 65.735 91.650 ;
        RECT 65.565 91.120 65.735 91.290 ;
        RECT 65.565 90.760 65.735 90.930 ;
        RECT 65.565 90.400 65.735 90.570 ;
        RECT 65.565 90.040 65.735 90.210 ;
        RECT 68.695 91.480 68.865 91.650 ;
        RECT 68.695 91.120 68.865 91.290 ;
        RECT 68.695 90.760 68.865 90.930 ;
        RECT 68.695 90.400 68.865 90.570 ;
        RECT 68.695 90.040 68.865 90.210 ;
        RECT 70.075 91.500 70.245 91.670 ;
        RECT 70.075 91.140 70.245 91.310 ;
        RECT 70.075 90.780 70.245 90.950 ;
        RECT 70.075 90.420 70.245 90.590 ;
        RECT 70.075 90.060 70.245 90.230 ;
        RECT 63.685 89.700 63.855 89.870 ;
        RECT 64.550 89.620 64.720 89.790 ;
        RECT 64.910 89.620 65.080 89.790 ;
        RECT 69.280 89.620 69.450 89.790 ;
        RECT 70.075 89.700 70.245 89.870 ;
        RECT 63.685 89.340 63.855 89.510 ;
        RECT 70.075 89.340 70.245 89.510 ;
        RECT 63.985 88.950 64.155 89.120 ;
        RECT 64.345 88.950 64.515 89.120 ;
        RECT 64.705 88.950 64.875 89.120 ;
        RECT 65.065 88.950 65.235 89.120 ;
        RECT 65.425 88.950 65.595 89.120 ;
        RECT 65.785 88.950 65.955 89.120 ;
        RECT 66.145 88.950 66.315 89.120 ;
        RECT 66.505 88.950 66.675 89.120 ;
        RECT 67.975 88.950 68.145 89.120 ;
        RECT 68.335 88.950 68.505 89.120 ;
        RECT 68.695 88.950 68.865 89.120 ;
        RECT 69.055 88.950 69.225 89.120 ;
        RECT 69.415 88.950 69.585 89.120 ;
        RECT 69.775 88.950 69.945 89.120 ;
        RECT 88.545 112.740 88.715 112.910 ;
        RECT 94.935 112.740 95.105 112.910 ;
        RECT 88.545 112.380 88.715 112.550 ;
        RECT 89.340 112.420 89.510 112.590 ;
        RECT 93.710 112.420 93.880 112.590 ;
        RECT 94.070 112.420 94.240 112.590 ;
        RECT 88.545 112.020 88.715 112.190 ;
        RECT 94.935 112.380 95.105 112.550 ;
        RECT 88.545 111.660 88.715 111.830 ;
        RECT 88.545 111.300 88.715 111.470 ;
        RECT 88.545 110.940 88.715 111.110 ;
        RECT 88.545 110.580 88.715 110.750 ;
        RECT 89.925 112.000 90.095 112.170 ;
        RECT 89.925 111.640 90.095 111.810 ;
        RECT 89.925 111.280 90.095 111.450 ;
        RECT 89.925 110.920 90.095 111.090 ;
        RECT 89.925 110.560 90.095 110.730 ;
        RECT 93.055 112.000 93.225 112.170 ;
        RECT 93.055 111.640 93.225 111.810 ;
        RECT 93.055 111.280 93.225 111.450 ;
        RECT 93.055 110.920 93.225 111.090 ;
        RECT 93.055 110.560 93.225 110.730 ;
        RECT 94.935 112.020 95.105 112.190 ;
        RECT 94.935 111.660 95.105 111.830 ;
        RECT 96.080 113.100 96.250 113.270 ;
        RECT 97.285 113.200 97.455 113.370 ;
        RECT 97.645 113.200 97.815 113.370 ;
        RECT 98.300 113.200 98.470 113.370 ;
        RECT 96.080 112.740 96.250 112.910 ;
        RECT 98.300 112.840 98.470 113.010 ;
        RECT 102.440 113.460 102.610 113.630 ;
        RECT 102.440 113.100 102.610 113.270 ;
        RECT 102.440 112.740 102.610 112.910 ;
        RECT 96.080 112.380 96.250 112.550 ;
        RECT 97.285 112.420 97.455 112.590 ;
        RECT 97.645 112.420 97.815 112.590 ;
        RECT 102.440 112.380 102.610 112.550 ;
        RECT 96.380 111.750 96.550 111.920 ;
        RECT 96.740 111.750 96.910 111.920 ;
        RECT 97.100 111.750 97.270 111.920 ;
        RECT 97.460 111.750 97.630 111.920 ;
        RECT 97.820 111.750 97.990 111.920 ;
        RECT 98.180 111.750 98.350 111.920 ;
        RECT 98.540 111.750 98.710 111.920 ;
        RECT 98.900 111.750 99.070 111.920 ;
        RECT 99.260 111.750 99.430 111.920 ;
        RECT 99.620 111.750 99.790 111.920 ;
        RECT 99.980 111.750 100.150 111.920 ;
        RECT 100.340 111.750 100.510 111.920 ;
        RECT 100.700 111.750 100.870 111.920 ;
        RECT 101.060 111.750 101.230 111.920 ;
        RECT 101.420 111.750 101.590 111.920 ;
        RECT 101.780 111.750 101.950 111.920 ;
        RECT 102.140 111.750 102.310 111.920 ;
        RECT 108.635 151.120 108.805 151.290 ;
        RECT 108.635 150.760 108.805 150.930 ;
        RECT 110.555 152.010 110.725 152.180 ;
        RECT 110.555 151.650 110.725 151.820 ;
        RECT 110.555 151.290 110.725 151.460 ;
        RECT 110.555 150.930 110.725 151.100 ;
        RECT 110.555 150.570 110.725 150.740 ;
        RECT 111.925 152.010 112.095 152.180 ;
        RECT 111.925 151.650 112.095 151.820 ;
        RECT 111.925 151.290 112.095 151.460 ;
        RECT 111.925 150.930 112.095 151.100 ;
        RECT 111.925 150.570 112.095 150.740 ;
        RECT 113.845 151.820 114.015 151.990 ;
        RECT 113.845 151.460 114.015 151.630 ;
        RECT 113.845 151.100 114.015 151.270 ;
        RECT 113.845 150.740 114.015 150.910 ;
        RECT 108.635 150.400 108.805 150.570 ;
        RECT 113.845 150.380 114.015 150.550 ;
        RECT 108.635 150.040 108.805 150.210 ;
        RECT 109.690 150.150 109.860 150.320 ;
        RECT 110.050 150.150 110.220 150.320 ;
        RECT 111.060 150.150 111.230 150.320 ;
        RECT 111.420 150.150 111.590 150.320 ;
        RECT 112.430 150.150 112.600 150.320 ;
        RECT 112.790 150.150 112.960 150.320 ;
        RECT 113.845 150.020 114.015 150.190 ;
        RECT 108.635 149.680 108.805 149.850 ;
        RECT 108.635 149.320 108.805 149.490 ;
        RECT 108.635 148.960 108.805 149.130 ;
        RECT 108.635 148.600 108.805 148.770 ;
        RECT 108.635 148.240 108.805 148.410 ;
        RECT 110.555 149.730 110.725 149.900 ;
        RECT 110.555 149.370 110.725 149.540 ;
        RECT 110.555 149.010 110.725 149.180 ;
        RECT 110.555 148.650 110.725 148.820 ;
        RECT 110.555 148.290 110.725 148.460 ;
        RECT 111.925 149.730 112.095 149.900 ;
        RECT 111.925 149.370 112.095 149.540 ;
        RECT 111.925 149.010 112.095 149.180 ;
        RECT 111.925 148.650 112.095 148.820 ;
        RECT 111.925 148.290 112.095 148.460 ;
        RECT 113.845 149.660 114.015 149.830 ;
        RECT 113.845 149.300 114.015 149.470 ;
        RECT 113.845 148.940 114.015 149.110 ;
        RECT 113.845 148.580 114.015 148.750 ;
        RECT 108.635 147.880 108.805 148.050 ;
        RECT 113.845 148.220 114.015 148.390 ;
        RECT 109.690 147.870 109.860 148.040 ;
        RECT 110.050 147.870 110.220 148.040 ;
        RECT 111.060 147.870 111.230 148.040 ;
        RECT 111.420 147.870 111.590 148.040 ;
        RECT 112.430 147.870 112.600 148.040 ;
        RECT 112.790 147.870 112.960 148.040 ;
        RECT 108.635 147.520 108.805 147.690 ;
        RECT 113.845 147.860 114.015 148.030 ;
        RECT 108.635 147.160 108.805 147.330 ;
        RECT 108.635 146.800 108.805 146.970 ;
        RECT 108.635 146.440 108.805 146.610 ;
        RECT 108.635 146.080 108.805 146.250 ;
        RECT 110.555 147.450 110.725 147.620 ;
        RECT 110.555 147.090 110.725 147.260 ;
        RECT 110.555 146.730 110.725 146.900 ;
        RECT 110.555 146.370 110.725 146.540 ;
        RECT 110.555 146.010 110.725 146.180 ;
        RECT 111.925 147.450 112.095 147.620 ;
        RECT 111.925 147.090 112.095 147.260 ;
        RECT 111.925 146.730 112.095 146.900 ;
        RECT 111.925 146.370 112.095 146.540 ;
        RECT 111.925 146.010 112.095 146.180 ;
        RECT 113.845 147.500 114.015 147.670 ;
        RECT 113.845 147.140 114.015 147.310 ;
        RECT 113.845 146.780 114.015 146.950 ;
        RECT 113.845 146.420 114.015 146.590 ;
        RECT 113.845 146.060 114.015 146.230 ;
        RECT 108.635 145.720 108.805 145.890 ;
        RECT 109.690 145.590 109.860 145.760 ;
        RECT 110.050 145.590 110.220 145.760 ;
        RECT 111.060 145.590 111.230 145.760 ;
        RECT 111.420 145.590 111.590 145.760 ;
        RECT 112.430 145.590 112.600 145.760 ;
        RECT 112.790 145.590 112.960 145.760 ;
        RECT 113.845 145.700 114.015 145.870 ;
        RECT 108.635 145.360 108.805 145.530 ;
        RECT 113.845 145.340 114.015 145.510 ;
        RECT 108.635 145.000 108.805 145.170 ;
        RECT 108.635 144.640 108.805 144.810 ;
        RECT 108.635 144.280 108.805 144.450 ;
        RECT 108.635 143.920 108.805 144.090 ;
        RECT 110.555 145.170 110.725 145.340 ;
        RECT 110.555 144.810 110.725 144.980 ;
        RECT 110.555 144.450 110.725 144.620 ;
        RECT 110.555 144.090 110.725 144.260 ;
        RECT 110.555 143.730 110.725 143.900 ;
        RECT 111.925 145.170 112.095 145.340 ;
        RECT 111.925 144.810 112.095 144.980 ;
        RECT 111.925 144.450 112.095 144.620 ;
        RECT 111.925 144.090 112.095 144.260 ;
        RECT 111.925 143.730 112.095 143.900 ;
        RECT 113.845 144.980 114.015 145.150 ;
        RECT 113.845 144.620 114.015 144.790 ;
        RECT 113.845 144.260 114.015 144.430 ;
        RECT 113.845 143.900 114.015 144.070 ;
        RECT 108.635 143.560 108.805 143.730 ;
        RECT 113.845 143.540 114.015 143.710 ;
        RECT 108.635 143.200 108.805 143.370 ;
        RECT 109.690 143.310 109.860 143.480 ;
        RECT 110.050 143.310 110.220 143.480 ;
        RECT 111.060 143.310 111.230 143.480 ;
        RECT 111.420 143.310 111.590 143.480 ;
        RECT 112.430 143.310 112.600 143.480 ;
        RECT 112.790 143.310 112.960 143.480 ;
        RECT 113.845 143.180 114.015 143.350 ;
        RECT 108.635 142.840 108.805 143.010 ;
        RECT 108.635 142.480 108.805 142.650 ;
        RECT 108.635 142.120 108.805 142.290 ;
        RECT 108.635 141.760 108.805 141.930 ;
        RECT 108.635 141.400 108.805 141.570 ;
        RECT 110.555 142.890 110.725 143.060 ;
        RECT 110.555 142.530 110.725 142.700 ;
        RECT 110.555 142.170 110.725 142.340 ;
        RECT 110.555 141.810 110.725 141.980 ;
        RECT 110.555 141.450 110.725 141.620 ;
        RECT 111.925 142.890 112.095 143.060 ;
        RECT 111.925 142.530 112.095 142.700 ;
        RECT 111.925 142.170 112.095 142.340 ;
        RECT 111.925 141.810 112.095 141.980 ;
        RECT 111.925 141.450 112.095 141.620 ;
        RECT 113.845 142.820 114.015 142.990 ;
        RECT 113.845 142.460 114.015 142.630 ;
        RECT 113.845 142.100 114.015 142.270 ;
        RECT 113.845 141.740 114.015 141.910 ;
        RECT 108.635 141.040 108.805 141.210 ;
        RECT 113.845 141.380 114.015 141.550 ;
        RECT 109.690 141.030 109.860 141.200 ;
        RECT 110.050 141.030 110.220 141.200 ;
        RECT 111.060 141.030 111.230 141.200 ;
        RECT 111.420 141.030 111.590 141.200 ;
        RECT 112.430 141.030 112.600 141.200 ;
        RECT 112.790 141.030 112.960 141.200 ;
        RECT 108.635 140.680 108.805 140.850 ;
        RECT 113.845 141.020 114.015 141.190 ;
        RECT 108.635 140.320 108.805 140.490 ;
        RECT 108.635 139.960 108.805 140.130 ;
        RECT 108.635 139.600 108.805 139.770 ;
        RECT 108.635 139.240 108.805 139.410 ;
        RECT 110.555 140.610 110.725 140.780 ;
        RECT 110.555 140.250 110.725 140.420 ;
        RECT 110.555 139.890 110.725 140.060 ;
        RECT 110.555 139.530 110.725 139.700 ;
        RECT 110.555 139.170 110.725 139.340 ;
        RECT 111.925 140.610 112.095 140.780 ;
        RECT 111.925 140.250 112.095 140.420 ;
        RECT 111.925 139.890 112.095 140.060 ;
        RECT 111.925 139.530 112.095 139.700 ;
        RECT 111.925 139.170 112.095 139.340 ;
        RECT 113.845 140.660 114.015 140.830 ;
        RECT 113.845 140.300 114.015 140.470 ;
        RECT 113.845 139.940 114.015 140.110 ;
        RECT 113.845 139.580 114.015 139.750 ;
        RECT 113.845 139.220 114.015 139.390 ;
        RECT 108.635 138.880 108.805 139.050 ;
        RECT 109.690 138.750 109.860 138.920 ;
        RECT 110.050 138.750 110.220 138.920 ;
        RECT 111.060 138.750 111.230 138.920 ;
        RECT 111.420 138.750 111.590 138.920 ;
        RECT 112.430 138.750 112.600 138.920 ;
        RECT 112.790 138.750 112.960 138.920 ;
        RECT 113.845 138.860 114.015 139.030 ;
        RECT 108.635 138.520 108.805 138.690 ;
        RECT 113.845 138.500 114.015 138.670 ;
        RECT 108.635 138.160 108.805 138.330 ;
        RECT 108.635 137.800 108.805 137.970 ;
        RECT 108.635 137.440 108.805 137.610 ;
        RECT 108.635 137.080 108.805 137.250 ;
        RECT 110.555 138.330 110.725 138.500 ;
        RECT 110.555 137.970 110.725 138.140 ;
        RECT 110.555 137.610 110.725 137.780 ;
        RECT 110.555 137.250 110.725 137.420 ;
        RECT 110.555 136.890 110.725 137.060 ;
        RECT 111.925 138.330 112.095 138.500 ;
        RECT 111.925 137.970 112.095 138.140 ;
        RECT 111.925 137.610 112.095 137.780 ;
        RECT 111.925 137.250 112.095 137.420 ;
        RECT 111.925 136.890 112.095 137.060 ;
        RECT 113.845 138.140 114.015 138.310 ;
        RECT 113.845 137.780 114.015 137.950 ;
        RECT 113.845 137.420 114.015 137.590 ;
        RECT 113.845 137.060 114.015 137.230 ;
        RECT 108.635 136.720 108.805 136.890 ;
        RECT 113.845 136.700 114.015 136.870 ;
        RECT 108.635 136.360 108.805 136.530 ;
        RECT 109.690 136.470 109.860 136.640 ;
        RECT 110.050 136.470 110.220 136.640 ;
        RECT 111.060 136.470 111.230 136.640 ;
        RECT 111.420 136.470 111.590 136.640 ;
        RECT 112.430 136.470 112.600 136.640 ;
        RECT 112.790 136.470 112.960 136.640 ;
        RECT 113.845 136.340 114.015 136.510 ;
        RECT 108.635 136.000 108.805 136.170 ;
        RECT 108.635 135.640 108.805 135.810 ;
        RECT 108.635 135.280 108.805 135.450 ;
        RECT 108.635 134.920 108.805 135.090 ;
        RECT 108.635 134.560 108.805 134.730 ;
        RECT 110.555 136.050 110.725 136.220 ;
        RECT 110.555 135.690 110.725 135.860 ;
        RECT 110.555 135.330 110.725 135.500 ;
        RECT 110.555 134.970 110.725 135.140 ;
        RECT 110.555 134.610 110.725 134.780 ;
        RECT 111.925 136.050 112.095 136.220 ;
        RECT 111.925 135.690 112.095 135.860 ;
        RECT 111.925 135.330 112.095 135.500 ;
        RECT 111.925 134.970 112.095 135.140 ;
        RECT 111.925 134.610 112.095 134.780 ;
        RECT 113.845 135.980 114.015 136.150 ;
        RECT 113.845 135.620 114.015 135.790 ;
        RECT 113.845 135.260 114.015 135.430 ;
        RECT 113.845 134.900 114.015 135.070 ;
        RECT 108.635 134.200 108.805 134.370 ;
        RECT 113.845 134.540 114.015 134.710 ;
        RECT 109.690 134.190 109.860 134.360 ;
        RECT 110.050 134.190 110.220 134.360 ;
        RECT 111.060 134.190 111.230 134.360 ;
        RECT 111.420 134.190 111.590 134.360 ;
        RECT 112.430 134.190 112.600 134.360 ;
        RECT 112.790 134.190 112.960 134.360 ;
        RECT 108.635 133.840 108.805 134.010 ;
        RECT 113.845 134.180 114.015 134.350 ;
        RECT 108.635 133.480 108.805 133.650 ;
        RECT 108.635 133.120 108.805 133.290 ;
        RECT 108.635 132.760 108.805 132.930 ;
        RECT 108.635 132.400 108.805 132.570 ;
        RECT 110.555 133.770 110.725 133.940 ;
        RECT 110.555 133.410 110.725 133.580 ;
        RECT 110.555 133.050 110.725 133.220 ;
        RECT 110.555 132.690 110.725 132.860 ;
        RECT 110.555 132.330 110.725 132.500 ;
        RECT 111.925 133.770 112.095 133.940 ;
        RECT 111.925 133.410 112.095 133.580 ;
        RECT 111.925 133.050 112.095 133.220 ;
        RECT 111.925 132.690 112.095 132.860 ;
        RECT 111.925 132.330 112.095 132.500 ;
        RECT 113.845 133.820 114.015 133.990 ;
        RECT 113.845 133.460 114.015 133.630 ;
        RECT 113.845 133.100 114.015 133.270 ;
        RECT 113.845 132.740 114.015 132.910 ;
        RECT 113.845 132.380 114.015 132.550 ;
        RECT 108.635 132.040 108.805 132.210 ;
        RECT 109.690 131.910 109.860 132.080 ;
        RECT 110.050 131.910 110.220 132.080 ;
        RECT 111.060 131.910 111.230 132.080 ;
        RECT 111.420 131.910 111.590 132.080 ;
        RECT 112.430 131.910 112.600 132.080 ;
        RECT 112.790 131.910 112.960 132.080 ;
        RECT 113.845 132.020 114.015 132.190 ;
        RECT 108.635 131.680 108.805 131.850 ;
        RECT 113.845 131.660 114.015 131.830 ;
        RECT 108.635 131.320 108.805 131.490 ;
        RECT 108.635 130.960 108.805 131.130 ;
        RECT 108.635 130.600 108.805 130.770 ;
        RECT 108.635 130.240 108.805 130.410 ;
        RECT 110.555 131.490 110.725 131.660 ;
        RECT 110.555 131.130 110.725 131.300 ;
        RECT 110.555 130.770 110.725 130.940 ;
        RECT 110.555 130.410 110.725 130.580 ;
        RECT 110.555 130.050 110.725 130.220 ;
        RECT 111.925 131.490 112.095 131.660 ;
        RECT 111.925 131.130 112.095 131.300 ;
        RECT 111.925 130.770 112.095 130.940 ;
        RECT 111.925 130.410 112.095 130.580 ;
        RECT 111.925 130.050 112.095 130.220 ;
        RECT 113.845 131.300 114.015 131.470 ;
        RECT 113.845 130.940 114.015 131.110 ;
        RECT 113.845 130.580 114.015 130.750 ;
        RECT 113.845 130.220 114.015 130.390 ;
        RECT 108.635 129.880 108.805 130.050 ;
        RECT 113.845 129.860 114.015 130.030 ;
        RECT 108.635 129.520 108.805 129.690 ;
        RECT 109.690 129.630 109.860 129.800 ;
        RECT 110.050 129.630 110.220 129.800 ;
        RECT 111.060 129.630 111.230 129.800 ;
        RECT 111.420 129.630 111.590 129.800 ;
        RECT 112.430 129.630 112.600 129.800 ;
        RECT 112.790 129.630 112.960 129.800 ;
        RECT 113.845 129.500 114.015 129.670 ;
        RECT 108.635 129.160 108.805 129.330 ;
        RECT 108.635 128.800 108.805 128.970 ;
        RECT 108.635 128.440 108.805 128.610 ;
        RECT 108.635 128.080 108.805 128.250 ;
        RECT 108.635 127.720 108.805 127.890 ;
        RECT 110.555 129.210 110.725 129.380 ;
        RECT 110.555 128.850 110.725 129.020 ;
        RECT 110.555 128.490 110.725 128.660 ;
        RECT 110.555 128.130 110.725 128.300 ;
        RECT 110.555 127.770 110.725 127.940 ;
        RECT 111.925 129.210 112.095 129.380 ;
        RECT 111.925 128.850 112.095 129.020 ;
        RECT 111.925 128.490 112.095 128.660 ;
        RECT 111.925 128.130 112.095 128.300 ;
        RECT 111.925 127.770 112.095 127.940 ;
        RECT 113.845 129.140 114.015 129.310 ;
        RECT 113.845 128.780 114.015 128.950 ;
        RECT 113.845 128.420 114.015 128.590 ;
        RECT 113.845 128.060 114.015 128.230 ;
        RECT 108.635 127.360 108.805 127.530 ;
        RECT 113.845 127.700 114.015 127.870 ;
        RECT 109.690 127.350 109.860 127.520 ;
        RECT 110.050 127.350 110.220 127.520 ;
        RECT 111.060 127.350 111.230 127.520 ;
        RECT 111.420 127.350 111.590 127.520 ;
        RECT 112.430 127.350 112.600 127.520 ;
        RECT 112.790 127.350 112.960 127.520 ;
        RECT 108.635 127.000 108.805 127.170 ;
        RECT 113.845 127.340 114.015 127.510 ;
        RECT 108.635 126.640 108.805 126.810 ;
        RECT 108.635 126.280 108.805 126.450 ;
        RECT 108.635 125.920 108.805 126.090 ;
        RECT 108.635 125.560 108.805 125.730 ;
        RECT 110.555 126.930 110.725 127.100 ;
        RECT 110.555 126.570 110.725 126.740 ;
        RECT 110.555 126.210 110.725 126.380 ;
        RECT 110.555 125.850 110.725 126.020 ;
        RECT 110.555 125.490 110.725 125.660 ;
        RECT 111.925 126.930 112.095 127.100 ;
        RECT 111.925 126.570 112.095 126.740 ;
        RECT 111.925 126.210 112.095 126.380 ;
        RECT 111.925 125.850 112.095 126.020 ;
        RECT 111.925 125.490 112.095 125.660 ;
        RECT 113.845 126.980 114.015 127.150 ;
        RECT 113.845 126.620 114.015 126.790 ;
        RECT 113.845 126.260 114.015 126.430 ;
        RECT 113.845 125.900 114.015 126.070 ;
        RECT 113.845 125.540 114.015 125.710 ;
        RECT 108.635 125.200 108.805 125.370 ;
        RECT 109.690 125.070 109.860 125.240 ;
        RECT 110.050 125.070 110.220 125.240 ;
        RECT 111.060 125.070 111.230 125.240 ;
        RECT 111.420 125.070 111.590 125.240 ;
        RECT 112.430 125.070 112.600 125.240 ;
        RECT 112.790 125.070 112.960 125.240 ;
        RECT 113.845 125.180 114.015 125.350 ;
        RECT 108.635 124.840 108.805 125.010 ;
        RECT 113.845 124.820 114.015 124.990 ;
        RECT 108.635 124.480 108.805 124.650 ;
        RECT 108.635 124.120 108.805 124.290 ;
        RECT 108.635 123.760 108.805 123.930 ;
        RECT 108.635 123.400 108.805 123.570 ;
        RECT 110.555 124.650 110.725 124.820 ;
        RECT 110.555 124.290 110.725 124.460 ;
        RECT 110.555 123.930 110.725 124.100 ;
        RECT 110.555 123.570 110.725 123.740 ;
        RECT 110.555 123.210 110.725 123.380 ;
        RECT 111.925 124.650 112.095 124.820 ;
        RECT 111.925 124.290 112.095 124.460 ;
        RECT 111.925 123.930 112.095 124.100 ;
        RECT 111.925 123.570 112.095 123.740 ;
        RECT 111.925 123.210 112.095 123.380 ;
        RECT 113.845 124.460 114.015 124.630 ;
        RECT 113.845 124.100 114.015 124.270 ;
        RECT 113.845 123.740 114.015 123.910 ;
        RECT 113.845 123.380 114.015 123.550 ;
        RECT 108.635 123.040 108.805 123.210 ;
        RECT 113.845 123.020 114.015 123.190 ;
        RECT 108.635 122.680 108.805 122.850 ;
        RECT 109.690 122.790 109.860 122.960 ;
        RECT 110.050 122.790 110.220 122.960 ;
        RECT 111.060 122.790 111.230 122.960 ;
        RECT 111.420 122.790 111.590 122.960 ;
        RECT 112.430 122.790 112.600 122.960 ;
        RECT 112.790 122.790 112.960 122.960 ;
        RECT 113.845 122.660 114.015 122.830 ;
        RECT 108.635 122.320 108.805 122.490 ;
        RECT 108.635 121.960 108.805 122.130 ;
        RECT 108.635 121.600 108.805 121.770 ;
        RECT 108.635 121.240 108.805 121.410 ;
        RECT 108.635 120.880 108.805 121.050 ;
        RECT 110.555 122.370 110.725 122.540 ;
        RECT 110.555 122.010 110.725 122.180 ;
        RECT 110.555 121.650 110.725 121.820 ;
        RECT 110.555 121.290 110.725 121.460 ;
        RECT 110.555 120.930 110.725 121.100 ;
        RECT 111.925 122.370 112.095 122.540 ;
        RECT 111.925 122.010 112.095 122.180 ;
        RECT 111.925 121.650 112.095 121.820 ;
        RECT 111.925 121.290 112.095 121.460 ;
        RECT 111.925 120.930 112.095 121.100 ;
        RECT 113.845 122.300 114.015 122.470 ;
        RECT 113.845 121.940 114.015 122.110 ;
        RECT 113.845 121.580 114.015 121.750 ;
        RECT 113.845 121.220 114.015 121.390 ;
        RECT 108.635 120.520 108.805 120.690 ;
        RECT 113.845 120.860 114.015 121.030 ;
        RECT 109.690 120.510 109.860 120.680 ;
        RECT 110.050 120.510 110.220 120.680 ;
        RECT 111.060 120.510 111.230 120.680 ;
        RECT 111.420 120.510 111.590 120.680 ;
        RECT 112.430 120.510 112.600 120.680 ;
        RECT 112.790 120.510 112.960 120.680 ;
        RECT 108.635 120.160 108.805 120.330 ;
        RECT 113.845 120.500 114.015 120.670 ;
        RECT 108.635 119.800 108.805 119.970 ;
        RECT 108.635 119.440 108.805 119.610 ;
        RECT 108.635 119.080 108.805 119.250 ;
        RECT 108.635 118.720 108.805 118.890 ;
        RECT 110.555 120.090 110.725 120.260 ;
        RECT 110.555 119.730 110.725 119.900 ;
        RECT 110.555 119.370 110.725 119.540 ;
        RECT 110.555 119.010 110.725 119.180 ;
        RECT 110.555 118.650 110.725 118.820 ;
        RECT 111.925 120.090 112.095 120.260 ;
        RECT 111.925 119.730 112.095 119.900 ;
        RECT 111.925 119.370 112.095 119.540 ;
        RECT 111.925 119.010 112.095 119.180 ;
        RECT 111.925 118.650 112.095 118.820 ;
        RECT 113.845 120.140 114.015 120.310 ;
        RECT 113.845 119.780 114.015 119.950 ;
        RECT 113.845 119.420 114.015 119.590 ;
        RECT 113.845 119.060 114.015 119.230 ;
        RECT 113.845 118.700 114.015 118.870 ;
        RECT 108.635 118.360 108.805 118.530 ;
        RECT 109.690 118.230 109.860 118.400 ;
        RECT 110.050 118.230 110.220 118.400 ;
        RECT 111.060 118.230 111.230 118.400 ;
        RECT 111.420 118.230 111.590 118.400 ;
        RECT 112.430 118.230 112.600 118.400 ;
        RECT 112.790 118.230 112.960 118.400 ;
        RECT 113.845 118.340 114.015 118.510 ;
        RECT 108.635 118.000 108.805 118.170 ;
        RECT 113.845 117.980 114.015 118.150 ;
        RECT 121.840 164.400 122.010 164.570 ;
        RECT 122.380 164.460 122.550 164.630 ;
        RECT 122.740 164.460 122.910 164.630 ;
        RECT 123.100 164.460 123.270 164.630 ;
        RECT 123.460 164.460 123.630 164.630 ;
        RECT 123.820 164.460 123.990 164.630 ;
        RECT 124.180 164.460 124.350 164.630 ;
        RECT 124.540 164.460 124.710 164.630 ;
        RECT 124.900 164.460 125.070 164.630 ;
        RECT 125.260 164.460 125.430 164.630 ;
        RECT 125.620 164.460 125.790 164.630 ;
        RECT 121.840 164.040 122.010 164.210 ;
        RECT 125.680 164.100 125.850 164.270 ;
        RECT 121.840 163.680 122.010 163.850 ;
        RECT 122.895 163.830 123.065 164.000 ;
        RECT 123.255 163.830 123.425 164.000 ;
        RECT 124.265 163.830 124.435 164.000 ;
        RECT 124.625 163.830 124.795 164.000 ;
        RECT 125.680 163.740 125.850 163.910 ;
        RECT 121.840 163.320 122.010 163.490 ;
        RECT 121.840 162.960 122.010 163.130 ;
        RECT 121.840 162.600 122.010 162.770 ;
        RECT 121.840 162.240 122.010 162.410 ;
        RECT 121.840 161.880 122.010 162.050 ;
        RECT 122.390 163.410 122.560 163.580 ;
        RECT 122.390 163.050 122.560 163.220 ;
        RECT 122.390 162.690 122.560 162.860 ;
        RECT 122.390 162.330 122.560 162.500 ;
        RECT 122.390 161.970 122.560 162.140 ;
        RECT 125.130 163.410 125.300 163.580 ;
        RECT 125.130 163.050 125.300 163.220 ;
        RECT 125.130 162.690 125.300 162.860 ;
        RECT 125.130 162.330 125.300 162.500 ;
        RECT 125.130 161.970 125.300 162.140 ;
        RECT 125.680 163.380 125.850 163.550 ;
        RECT 125.680 163.020 125.850 163.190 ;
        RECT 125.680 162.660 125.850 162.830 ;
        RECT 125.680 162.300 125.850 162.470 ;
        RECT 125.680 161.940 125.850 162.110 ;
        RECT 121.840 161.520 122.010 161.690 ;
        RECT 122.895 161.550 123.065 161.720 ;
        RECT 123.255 161.550 123.425 161.720 ;
        RECT 124.265 161.550 124.435 161.720 ;
        RECT 124.625 161.550 124.795 161.720 ;
        RECT 125.680 161.580 125.850 161.750 ;
        RECT 121.840 161.160 122.010 161.330 ;
        RECT 121.840 160.800 122.010 160.970 ;
        RECT 121.840 160.440 122.010 160.610 ;
        RECT 121.840 160.080 122.010 160.250 ;
        RECT 121.840 159.720 122.010 159.890 ;
        RECT 122.390 161.130 122.560 161.300 ;
        RECT 122.390 160.770 122.560 160.940 ;
        RECT 122.390 160.410 122.560 160.580 ;
        RECT 122.390 160.050 122.560 160.220 ;
        RECT 122.390 159.690 122.560 159.860 ;
        RECT 125.130 161.130 125.300 161.300 ;
        RECT 125.130 160.770 125.300 160.940 ;
        RECT 125.130 160.410 125.300 160.580 ;
        RECT 125.130 160.050 125.300 160.220 ;
        RECT 125.130 159.690 125.300 159.860 ;
        RECT 125.680 161.220 125.850 161.390 ;
        RECT 125.680 160.860 125.850 161.030 ;
        RECT 125.680 160.500 125.850 160.670 ;
        RECT 125.680 160.140 125.850 160.310 ;
        RECT 125.680 159.780 125.850 159.950 ;
        RECT 121.840 159.360 122.010 159.530 ;
        RECT 122.895 159.270 123.065 159.440 ;
        RECT 123.255 159.270 123.425 159.440 ;
        RECT 124.265 159.270 124.435 159.440 ;
        RECT 124.625 159.270 124.795 159.440 ;
        RECT 125.680 159.420 125.850 159.590 ;
        RECT 121.840 159.000 122.010 159.170 ;
        RECT 125.680 159.060 125.850 159.230 ;
        RECT 121.840 158.640 122.010 158.810 ;
        RECT 121.840 158.280 122.010 158.450 ;
        RECT 121.840 157.920 122.010 158.090 ;
        RECT 121.840 157.560 122.010 157.730 ;
        RECT 122.390 158.850 122.560 159.020 ;
        RECT 122.390 158.490 122.560 158.660 ;
        RECT 122.390 158.130 122.560 158.300 ;
        RECT 122.390 157.770 122.560 157.940 ;
        RECT 122.390 157.410 122.560 157.580 ;
        RECT 123.760 158.850 123.930 159.020 ;
        RECT 123.760 158.490 123.930 158.660 ;
        RECT 123.760 158.130 123.930 158.300 ;
        RECT 123.760 157.770 123.930 157.940 ;
        RECT 123.760 157.410 123.930 157.580 ;
        RECT 125.130 158.850 125.300 159.020 ;
        RECT 125.130 158.490 125.300 158.660 ;
        RECT 125.130 158.130 125.300 158.300 ;
        RECT 125.130 157.770 125.300 157.940 ;
        RECT 125.130 157.410 125.300 157.580 ;
        RECT 125.680 158.700 125.850 158.870 ;
        RECT 125.680 158.340 125.850 158.510 ;
        RECT 125.680 157.980 125.850 158.150 ;
        RECT 125.680 157.620 125.850 157.790 ;
        RECT 121.840 157.200 122.010 157.370 ;
        RECT 125.680 157.260 125.850 157.430 ;
        RECT 121.840 156.840 122.010 157.010 ;
        RECT 122.895 156.990 123.065 157.160 ;
        RECT 123.255 156.990 123.425 157.160 ;
        RECT 124.265 156.990 124.435 157.160 ;
        RECT 124.625 156.990 124.795 157.160 ;
        RECT 125.680 156.900 125.850 157.070 ;
        RECT 121.840 156.480 122.010 156.650 ;
        RECT 121.840 156.120 122.010 156.290 ;
        RECT 121.840 155.760 122.010 155.930 ;
        RECT 121.840 155.400 122.010 155.570 ;
        RECT 121.840 155.040 122.010 155.210 ;
        RECT 122.390 156.570 122.560 156.740 ;
        RECT 122.390 156.210 122.560 156.380 ;
        RECT 122.390 155.850 122.560 156.020 ;
        RECT 122.390 155.490 122.560 155.660 ;
        RECT 122.390 155.130 122.560 155.300 ;
        RECT 123.760 156.570 123.930 156.740 ;
        RECT 123.760 156.210 123.930 156.380 ;
        RECT 123.760 155.850 123.930 156.020 ;
        RECT 123.760 155.490 123.930 155.660 ;
        RECT 123.760 155.130 123.930 155.300 ;
        RECT 125.130 156.570 125.300 156.740 ;
        RECT 125.130 156.210 125.300 156.380 ;
        RECT 125.130 155.850 125.300 156.020 ;
        RECT 125.130 155.490 125.300 155.660 ;
        RECT 125.130 155.130 125.300 155.300 ;
        RECT 125.680 156.540 125.850 156.710 ;
        RECT 125.680 156.180 125.850 156.350 ;
        RECT 125.680 155.820 125.850 155.990 ;
        RECT 125.680 155.460 125.850 155.630 ;
        RECT 125.680 155.100 125.850 155.270 ;
        RECT 121.840 154.680 122.010 154.850 ;
        RECT 122.895 154.710 123.065 154.880 ;
        RECT 123.255 154.710 123.425 154.880 ;
        RECT 124.265 154.710 124.435 154.880 ;
        RECT 124.625 154.710 124.795 154.880 ;
        RECT 125.680 154.740 125.850 154.910 ;
        RECT 121.840 154.320 122.010 154.490 ;
        RECT 121.840 153.960 122.010 154.130 ;
        RECT 121.840 153.600 122.010 153.770 ;
        RECT 121.840 153.240 122.010 153.410 ;
        RECT 121.840 152.880 122.010 153.050 ;
        RECT 122.390 154.290 122.560 154.460 ;
        RECT 122.390 153.930 122.560 154.100 ;
        RECT 122.390 153.570 122.560 153.740 ;
        RECT 122.390 153.210 122.560 153.380 ;
        RECT 122.390 152.850 122.560 153.020 ;
        RECT 123.760 154.290 123.930 154.460 ;
        RECT 123.760 153.930 123.930 154.100 ;
        RECT 123.760 153.570 123.930 153.740 ;
        RECT 123.760 153.210 123.930 153.380 ;
        RECT 123.760 152.850 123.930 153.020 ;
        RECT 125.130 154.290 125.300 154.460 ;
        RECT 125.130 153.930 125.300 154.100 ;
        RECT 125.130 153.570 125.300 153.740 ;
        RECT 125.130 153.210 125.300 153.380 ;
        RECT 125.130 152.850 125.300 153.020 ;
        RECT 125.680 154.380 125.850 154.550 ;
        RECT 125.680 154.020 125.850 154.190 ;
        RECT 125.680 153.660 125.850 153.830 ;
        RECT 125.680 153.300 125.850 153.470 ;
        RECT 125.680 152.940 125.850 153.110 ;
        RECT 121.840 152.520 122.010 152.690 ;
        RECT 122.895 152.430 123.065 152.600 ;
        RECT 123.255 152.430 123.425 152.600 ;
        RECT 124.265 152.430 124.435 152.600 ;
        RECT 124.625 152.430 124.795 152.600 ;
        RECT 125.680 152.580 125.850 152.750 ;
        RECT 121.840 152.160 122.010 152.330 ;
        RECT 125.680 152.220 125.850 152.390 ;
        RECT 121.840 151.800 122.010 151.970 ;
        RECT 121.840 151.440 122.010 151.610 ;
        RECT 121.840 151.080 122.010 151.250 ;
        RECT 121.840 150.720 122.010 150.890 ;
        RECT 122.390 152.010 122.560 152.180 ;
        RECT 122.390 151.650 122.560 151.820 ;
        RECT 122.390 151.290 122.560 151.460 ;
        RECT 122.390 150.930 122.560 151.100 ;
        RECT 122.390 150.570 122.560 150.740 ;
        RECT 123.760 152.010 123.930 152.180 ;
        RECT 123.760 151.650 123.930 151.820 ;
        RECT 123.760 151.290 123.930 151.460 ;
        RECT 123.760 150.930 123.930 151.100 ;
        RECT 123.760 150.570 123.930 150.740 ;
        RECT 125.130 152.010 125.300 152.180 ;
        RECT 125.130 151.650 125.300 151.820 ;
        RECT 125.130 151.290 125.300 151.460 ;
        RECT 125.130 150.930 125.300 151.100 ;
        RECT 125.130 150.570 125.300 150.740 ;
        RECT 125.680 151.860 125.850 152.030 ;
        RECT 125.680 151.500 125.850 151.670 ;
        RECT 125.680 151.140 125.850 151.310 ;
        RECT 125.680 150.780 125.850 150.950 ;
        RECT 121.840 150.360 122.010 150.530 ;
        RECT 125.680 150.420 125.850 150.590 ;
        RECT 121.840 150.000 122.010 150.170 ;
        RECT 122.895 150.150 123.065 150.320 ;
        RECT 123.255 150.150 123.425 150.320 ;
        RECT 124.265 150.150 124.435 150.320 ;
        RECT 124.625 150.150 124.795 150.320 ;
        RECT 125.680 150.060 125.850 150.230 ;
        RECT 121.840 149.640 122.010 149.810 ;
        RECT 121.840 149.280 122.010 149.450 ;
        RECT 121.840 148.920 122.010 149.090 ;
        RECT 121.840 148.560 122.010 148.730 ;
        RECT 121.840 148.200 122.010 148.370 ;
        RECT 122.390 149.730 122.560 149.900 ;
        RECT 122.390 149.370 122.560 149.540 ;
        RECT 122.390 149.010 122.560 149.180 ;
        RECT 122.390 148.650 122.560 148.820 ;
        RECT 122.390 148.290 122.560 148.460 ;
        RECT 123.760 149.730 123.930 149.900 ;
        RECT 123.760 149.370 123.930 149.540 ;
        RECT 123.760 149.010 123.930 149.180 ;
        RECT 123.760 148.650 123.930 148.820 ;
        RECT 123.760 148.290 123.930 148.460 ;
        RECT 125.130 149.730 125.300 149.900 ;
        RECT 125.130 149.370 125.300 149.540 ;
        RECT 125.130 149.010 125.300 149.180 ;
        RECT 125.130 148.650 125.300 148.820 ;
        RECT 125.130 148.290 125.300 148.460 ;
        RECT 125.680 149.700 125.850 149.870 ;
        RECT 125.680 149.340 125.850 149.510 ;
        RECT 125.680 148.980 125.850 149.150 ;
        RECT 125.680 148.620 125.850 148.790 ;
        RECT 125.680 148.260 125.850 148.430 ;
        RECT 121.840 147.840 122.010 148.010 ;
        RECT 122.895 147.870 123.065 148.040 ;
        RECT 123.255 147.870 123.425 148.040 ;
        RECT 124.265 147.870 124.435 148.040 ;
        RECT 124.625 147.870 124.795 148.040 ;
        RECT 125.680 147.900 125.850 148.070 ;
        RECT 121.840 147.480 122.010 147.650 ;
        RECT 121.840 147.120 122.010 147.290 ;
        RECT 121.840 146.760 122.010 146.930 ;
        RECT 121.840 146.400 122.010 146.570 ;
        RECT 121.840 146.040 122.010 146.210 ;
        RECT 122.390 147.450 122.560 147.620 ;
        RECT 122.390 147.090 122.560 147.260 ;
        RECT 122.390 146.730 122.560 146.900 ;
        RECT 122.390 146.370 122.560 146.540 ;
        RECT 122.390 146.010 122.560 146.180 ;
        RECT 123.760 147.450 123.930 147.620 ;
        RECT 123.760 147.090 123.930 147.260 ;
        RECT 123.760 146.730 123.930 146.900 ;
        RECT 123.760 146.370 123.930 146.540 ;
        RECT 123.760 146.010 123.930 146.180 ;
        RECT 125.130 147.450 125.300 147.620 ;
        RECT 125.130 147.090 125.300 147.260 ;
        RECT 125.130 146.730 125.300 146.900 ;
        RECT 125.130 146.370 125.300 146.540 ;
        RECT 125.130 146.010 125.300 146.180 ;
        RECT 125.680 147.540 125.850 147.710 ;
        RECT 125.680 147.180 125.850 147.350 ;
        RECT 125.680 146.820 125.850 146.990 ;
        RECT 125.680 146.460 125.850 146.630 ;
        RECT 125.680 146.100 125.850 146.270 ;
        RECT 121.840 145.680 122.010 145.850 ;
        RECT 122.895 145.590 123.065 145.760 ;
        RECT 123.255 145.590 123.425 145.760 ;
        RECT 124.265 145.590 124.435 145.760 ;
        RECT 124.625 145.590 124.795 145.760 ;
        RECT 125.680 145.740 125.850 145.910 ;
        RECT 121.840 145.320 122.010 145.490 ;
        RECT 125.680 145.380 125.850 145.550 ;
        RECT 121.840 144.960 122.010 145.130 ;
        RECT 121.840 144.600 122.010 144.770 ;
        RECT 121.840 144.240 122.010 144.410 ;
        RECT 121.840 143.880 122.010 144.050 ;
        RECT 122.390 145.170 122.560 145.340 ;
        RECT 122.390 144.810 122.560 144.980 ;
        RECT 122.390 144.450 122.560 144.620 ;
        RECT 122.390 144.090 122.560 144.260 ;
        RECT 122.390 143.730 122.560 143.900 ;
        RECT 123.760 145.170 123.930 145.340 ;
        RECT 123.760 144.810 123.930 144.980 ;
        RECT 123.760 144.450 123.930 144.620 ;
        RECT 123.760 144.090 123.930 144.260 ;
        RECT 123.760 143.730 123.930 143.900 ;
        RECT 125.130 145.170 125.300 145.340 ;
        RECT 125.130 144.810 125.300 144.980 ;
        RECT 125.130 144.450 125.300 144.620 ;
        RECT 125.130 144.090 125.300 144.260 ;
        RECT 125.130 143.730 125.300 143.900 ;
        RECT 125.680 145.020 125.850 145.190 ;
        RECT 125.680 144.660 125.850 144.830 ;
        RECT 125.680 144.300 125.850 144.470 ;
        RECT 125.680 143.940 125.850 144.110 ;
        RECT 121.840 143.520 122.010 143.690 ;
        RECT 125.680 143.580 125.850 143.750 ;
        RECT 121.840 143.160 122.010 143.330 ;
        RECT 122.895 143.310 123.065 143.480 ;
        RECT 123.255 143.310 123.425 143.480 ;
        RECT 124.265 143.310 124.435 143.480 ;
        RECT 124.625 143.310 124.795 143.480 ;
        RECT 125.680 143.220 125.850 143.390 ;
        RECT 121.840 142.800 122.010 142.970 ;
        RECT 121.840 142.440 122.010 142.610 ;
        RECT 121.840 142.080 122.010 142.250 ;
        RECT 121.840 141.720 122.010 141.890 ;
        RECT 121.840 141.360 122.010 141.530 ;
        RECT 122.390 142.890 122.560 143.060 ;
        RECT 122.390 142.530 122.560 142.700 ;
        RECT 122.390 142.170 122.560 142.340 ;
        RECT 122.390 141.810 122.560 141.980 ;
        RECT 122.390 141.450 122.560 141.620 ;
        RECT 123.760 142.890 123.930 143.060 ;
        RECT 123.760 142.530 123.930 142.700 ;
        RECT 123.760 142.170 123.930 142.340 ;
        RECT 123.760 141.810 123.930 141.980 ;
        RECT 123.760 141.450 123.930 141.620 ;
        RECT 125.130 142.890 125.300 143.060 ;
        RECT 125.130 142.530 125.300 142.700 ;
        RECT 125.130 142.170 125.300 142.340 ;
        RECT 125.130 141.810 125.300 141.980 ;
        RECT 125.130 141.450 125.300 141.620 ;
        RECT 125.680 142.860 125.850 143.030 ;
        RECT 125.680 142.500 125.850 142.670 ;
        RECT 125.680 142.140 125.850 142.310 ;
        RECT 125.680 141.780 125.850 141.950 ;
        RECT 125.680 141.420 125.850 141.590 ;
        RECT 121.840 141.000 122.010 141.170 ;
        RECT 122.895 141.030 123.065 141.200 ;
        RECT 123.255 141.030 123.425 141.200 ;
        RECT 124.265 141.030 124.435 141.200 ;
        RECT 124.625 141.030 124.795 141.200 ;
        RECT 125.680 141.060 125.850 141.230 ;
        RECT 121.840 140.640 122.010 140.810 ;
        RECT 121.840 140.280 122.010 140.450 ;
        RECT 121.840 139.920 122.010 140.090 ;
        RECT 121.840 139.560 122.010 139.730 ;
        RECT 121.840 139.200 122.010 139.370 ;
        RECT 122.390 140.610 122.560 140.780 ;
        RECT 122.390 140.250 122.560 140.420 ;
        RECT 122.390 139.890 122.560 140.060 ;
        RECT 122.390 139.530 122.560 139.700 ;
        RECT 122.390 139.170 122.560 139.340 ;
        RECT 123.760 140.610 123.930 140.780 ;
        RECT 123.760 140.250 123.930 140.420 ;
        RECT 123.760 139.890 123.930 140.060 ;
        RECT 123.760 139.530 123.930 139.700 ;
        RECT 123.760 139.170 123.930 139.340 ;
        RECT 125.130 140.610 125.300 140.780 ;
        RECT 125.130 140.250 125.300 140.420 ;
        RECT 125.130 139.890 125.300 140.060 ;
        RECT 125.130 139.530 125.300 139.700 ;
        RECT 125.130 139.170 125.300 139.340 ;
        RECT 125.680 140.700 125.850 140.870 ;
        RECT 125.680 140.340 125.850 140.510 ;
        RECT 125.680 139.980 125.850 140.150 ;
        RECT 125.680 139.620 125.850 139.790 ;
        RECT 125.680 139.260 125.850 139.430 ;
        RECT 121.840 138.840 122.010 139.010 ;
        RECT 122.895 138.750 123.065 138.920 ;
        RECT 123.255 138.750 123.425 138.920 ;
        RECT 124.265 138.750 124.435 138.920 ;
        RECT 124.625 138.750 124.795 138.920 ;
        RECT 125.680 138.900 125.850 139.070 ;
        RECT 121.840 138.480 122.010 138.650 ;
        RECT 125.680 138.540 125.850 138.710 ;
        RECT 121.840 138.120 122.010 138.290 ;
        RECT 121.840 137.760 122.010 137.930 ;
        RECT 121.840 137.400 122.010 137.570 ;
        RECT 121.840 137.040 122.010 137.210 ;
        RECT 122.390 138.330 122.560 138.500 ;
        RECT 122.390 137.970 122.560 138.140 ;
        RECT 122.390 137.610 122.560 137.780 ;
        RECT 122.390 137.250 122.560 137.420 ;
        RECT 122.390 136.890 122.560 137.060 ;
        RECT 123.760 138.330 123.930 138.500 ;
        RECT 123.760 137.970 123.930 138.140 ;
        RECT 123.760 137.610 123.930 137.780 ;
        RECT 123.760 137.250 123.930 137.420 ;
        RECT 123.760 136.890 123.930 137.060 ;
        RECT 125.130 138.330 125.300 138.500 ;
        RECT 125.130 137.970 125.300 138.140 ;
        RECT 125.130 137.610 125.300 137.780 ;
        RECT 125.130 137.250 125.300 137.420 ;
        RECT 125.130 136.890 125.300 137.060 ;
        RECT 125.680 138.180 125.850 138.350 ;
        RECT 125.680 137.820 125.850 137.990 ;
        RECT 125.680 137.460 125.850 137.630 ;
        RECT 125.680 137.100 125.850 137.270 ;
        RECT 121.840 136.680 122.010 136.850 ;
        RECT 125.680 136.740 125.850 136.910 ;
        RECT 121.840 136.320 122.010 136.490 ;
        RECT 122.895 136.470 123.065 136.640 ;
        RECT 123.255 136.470 123.425 136.640 ;
        RECT 124.265 136.470 124.435 136.640 ;
        RECT 124.625 136.470 124.795 136.640 ;
        RECT 125.680 136.380 125.850 136.550 ;
        RECT 121.840 135.960 122.010 136.130 ;
        RECT 121.840 135.600 122.010 135.770 ;
        RECT 121.840 135.240 122.010 135.410 ;
        RECT 121.840 134.880 122.010 135.050 ;
        RECT 121.840 134.520 122.010 134.690 ;
        RECT 122.390 136.050 122.560 136.220 ;
        RECT 122.390 135.690 122.560 135.860 ;
        RECT 122.390 135.330 122.560 135.500 ;
        RECT 122.390 134.970 122.560 135.140 ;
        RECT 122.390 134.610 122.560 134.780 ;
        RECT 123.760 136.050 123.930 136.220 ;
        RECT 123.760 135.690 123.930 135.860 ;
        RECT 123.760 135.330 123.930 135.500 ;
        RECT 123.760 134.970 123.930 135.140 ;
        RECT 123.760 134.610 123.930 134.780 ;
        RECT 125.130 136.050 125.300 136.220 ;
        RECT 125.130 135.690 125.300 135.860 ;
        RECT 125.130 135.330 125.300 135.500 ;
        RECT 125.130 134.970 125.300 135.140 ;
        RECT 125.130 134.610 125.300 134.780 ;
        RECT 125.680 136.020 125.850 136.190 ;
        RECT 125.680 135.660 125.850 135.830 ;
        RECT 125.680 135.300 125.850 135.470 ;
        RECT 125.680 134.940 125.850 135.110 ;
        RECT 125.680 134.580 125.850 134.750 ;
        RECT 121.840 134.160 122.010 134.330 ;
        RECT 122.895 134.190 123.065 134.360 ;
        RECT 123.255 134.190 123.425 134.360 ;
        RECT 124.265 134.190 124.435 134.360 ;
        RECT 124.625 134.190 124.795 134.360 ;
        RECT 125.680 134.220 125.850 134.390 ;
        RECT 121.840 133.800 122.010 133.970 ;
        RECT 121.840 133.440 122.010 133.610 ;
        RECT 121.840 133.080 122.010 133.250 ;
        RECT 121.840 132.720 122.010 132.890 ;
        RECT 121.840 132.360 122.010 132.530 ;
        RECT 122.390 133.770 122.560 133.940 ;
        RECT 122.390 133.410 122.560 133.580 ;
        RECT 122.390 133.050 122.560 133.220 ;
        RECT 122.390 132.690 122.560 132.860 ;
        RECT 122.390 132.330 122.560 132.500 ;
        RECT 123.760 133.770 123.930 133.940 ;
        RECT 123.760 133.410 123.930 133.580 ;
        RECT 123.760 133.050 123.930 133.220 ;
        RECT 123.760 132.690 123.930 132.860 ;
        RECT 123.760 132.330 123.930 132.500 ;
        RECT 125.130 133.770 125.300 133.940 ;
        RECT 125.130 133.410 125.300 133.580 ;
        RECT 125.130 133.050 125.300 133.220 ;
        RECT 125.130 132.690 125.300 132.860 ;
        RECT 125.130 132.330 125.300 132.500 ;
        RECT 125.680 133.860 125.850 134.030 ;
        RECT 125.680 133.500 125.850 133.670 ;
        RECT 125.680 133.140 125.850 133.310 ;
        RECT 125.680 132.780 125.850 132.950 ;
        RECT 125.680 132.420 125.850 132.590 ;
        RECT 121.840 132.000 122.010 132.170 ;
        RECT 122.895 131.910 123.065 132.080 ;
        RECT 123.255 131.910 123.425 132.080 ;
        RECT 124.265 131.910 124.435 132.080 ;
        RECT 124.625 131.910 124.795 132.080 ;
        RECT 125.680 132.060 125.850 132.230 ;
        RECT 121.840 131.640 122.010 131.810 ;
        RECT 125.680 131.700 125.850 131.870 ;
        RECT 121.840 131.280 122.010 131.450 ;
        RECT 121.840 130.920 122.010 131.090 ;
        RECT 121.840 130.560 122.010 130.730 ;
        RECT 121.840 130.200 122.010 130.370 ;
        RECT 122.390 131.490 122.560 131.660 ;
        RECT 122.390 131.130 122.560 131.300 ;
        RECT 122.390 130.770 122.560 130.940 ;
        RECT 122.390 130.410 122.560 130.580 ;
        RECT 122.390 130.050 122.560 130.220 ;
        RECT 123.760 131.490 123.930 131.660 ;
        RECT 123.760 131.130 123.930 131.300 ;
        RECT 123.760 130.770 123.930 130.940 ;
        RECT 123.760 130.410 123.930 130.580 ;
        RECT 123.760 130.050 123.930 130.220 ;
        RECT 125.130 131.490 125.300 131.660 ;
        RECT 125.130 131.130 125.300 131.300 ;
        RECT 125.130 130.770 125.300 130.940 ;
        RECT 125.130 130.410 125.300 130.580 ;
        RECT 125.130 130.050 125.300 130.220 ;
        RECT 125.680 131.340 125.850 131.510 ;
        RECT 125.680 130.980 125.850 131.150 ;
        RECT 125.680 130.620 125.850 130.790 ;
        RECT 125.680 130.260 125.850 130.430 ;
        RECT 121.840 129.840 122.010 130.010 ;
        RECT 125.680 129.900 125.850 130.070 ;
        RECT 121.840 129.480 122.010 129.650 ;
        RECT 122.895 129.630 123.065 129.800 ;
        RECT 123.255 129.630 123.425 129.800 ;
        RECT 124.265 129.630 124.435 129.800 ;
        RECT 124.625 129.630 124.795 129.800 ;
        RECT 125.680 129.540 125.850 129.710 ;
        RECT 121.840 129.120 122.010 129.290 ;
        RECT 121.840 128.760 122.010 128.930 ;
        RECT 121.840 128.400 122.010 128.570 ;
        RECT 121.840 128.040 122.010 128.210 ;
        RECT 121.840 127.680 122.010 127.850 ;
        RECT 122.390 129.210 122.560 129.380 ;
        RECT 122.390 128.850 122.560 129.020 ;
        RECT 122.390 128.490 122.560 128.660 ;
        RECT 122.390 128.130 122.560 128.300 ;
        RECT 122.390 127.770 122.560 127.940 ;
        RECT 123.760 129.210 123.930 129.380 ;
        RECT 123.760 128.850 123.930 129.020 ;
        RECT 123.760 128.490 123.930 128.660 ;
        RECT 123.760 128.130 123.930 128.300 ;
        RECT 123.760 127.770 123.930 127.940 ;
        RECT 125.130 129.210 125.300 129.380 ;
        RECT 125.130 128.850 125.300 129.020 ;
        RECT 125.130 128.490 125.300 128.660 ;
        RECT 125.130 128.130 125.300 128.300 ;
        RECT 125.130 127.770 125.300 127.940 ;
        RECT 125.680 129.180 125.850 129.350 ;
        RECT 125.680 128.820 125.850 128.990 ;
        RECT 125.680 128.460 125.850 128.630 ;
        RECT 125.680 128.100 125.850 128.270 ;
        RECT 125.680 127.740 125.850 127.910 ;
        RECT 121.840 127.320 122.010 127.490 ;
        RECT 122.895 127.350 123.065 127.520 ;
        RECT 123.255 127.350 123.425 127.520 ;
        RECT 124.265 127.350 124.435 127.520 ;
        RECT 124.625 127.350 124.795 127.520 ;
        RECT 125.680 127.380 125.850 127.550 ;
        RECT 121.840 126.960 122.010 127.130 ;
        RECT 121.840 126.600 122.010 126.770 ;
        RECT 121.840 126.240 122.010 126.410 ;
        RECT 121.840 125.880 122.010 126.050 ;
        RECT 121.840 125.520 122.010 125.690 ;
        RECT 122.390 126.930 122.560 127.100 ;
        RECT 122.390 126.570 122.560 126.740 ;
        RECT 122.390 126.210 122.560 126.380 ;
        RECT 122.390 125.850 122.560 126.020 ;
        RECT 122.390 125.490 122.560 125.660 ;
        RECT 123.760 126.930 123.930 127.100 ;
        RECT 123.760 126.570 123.930 126.740 ;
        RECT 123.760 126.210 123.930 126.380 ;
        RECT 123.760 125.850 123.930 126.020 ;
        RECT 123.760 125.490 123.930 125.660 ;
        RECT 125.130 126.930 125.300 127.100 ;
        RECT 125.130 126.570 125.300 126.740 ;
        RECT 125.130 126.210 125.300 126.380 ;
        RECT 125.130 125.850 125.300 126.020 ;
        RECT 125.130 125.490 125.300 125.660 ;
        RECT 125.680 127.020 125.850 127.190 ;
        RECT 125.680 126.660 125.850 126.830 ;
        RECT 125.680 126.300 125.850 126.470 ;
        RECT 125.680 125.940 125.850 126.110 ;
        RECT 125.680 125.580 125.850 125.750 ;
        RECT 121.840 125.160 122.010 125.330 ;
        RECT 122.895 125.070 123.065 125.240 ;
        RECT 123.255 125.070 123.425 125.240 ;
        RECT 124.265 125.070 124.435 125.240 ;
        RECT 124.625 125.070 124.795 125.240 ;
        RECT 125.680 125.220 125.850 125.390 ;
        RECT 121.840 124.800 122.010 124.970 ;
        RECT 125.680 124.860 125.850 125.030 ;
        RECT 121.840 124.440 122.010 124.610 ;
        RECT 121.840 124.080 122.010 124.250 ;
        RECT 121.840 123.720 122.010 123.890 ;
        RECT 121.840 123.360 122.010 123.530 ;
        RECT 122.390 124.650 122.560 124.820 ;
        RECT 122.390 124.290 122.560 124.460 ;
        RECT 122.390 123.930 122.560 124.100 ;
        RECT 122.390 123.570 122.560 123.740 ;
        RECT 122.390 123.210 122.560 123.380 ;
        RECT 123.760 124.650 123.930 124.820 ;
        RECT 123.760 124.290 123.930 124.460 ;
        RECT 123.760 123.930 123.930 124.100 ;
        RECT 123.760 123.570 123.930 123.740 ;
        RECT 123.760 123.210 123.930 123.380 ;
        RECT 125.130 124.650 125.300 124.820 ;
        RECT 125.130 124.290 125.300 124.460 ;
        RECT 125.130 123.930 125.300 124.100 ;
        RECT 125.130 123.570 125.300 123.740 ;
        RECT 125.130 123.210 125.300 123.380 ;
        RECT 125.680 124.500 125.850 124.670 ;
        RECT 125.680 124.140 125.850 124.310 ;
        RECT 125.680 123.780 125.850 123.950 ;
        RECT 125.680 123.420 125.850 123.590 ;
        RECT 121.840 123.000 122.010 123.170 ;
        RECT 125.680 123.060 125.850 123.230 ;
        RECT 121.840 122.640 122.010 122.810 ;
        RECT 122.895 122.790 123.065 122.960 ;
        RECT 123.255 122.790 123.425 122.960 ;
        RECT 124.265 122.790 124.435 122.960 ;
        RECT 124.625 122.790 124.795 122.960 ;
        RECT 125.680 122.700 125.850 122.870 ;
        RECT 121.840 122.280 122.010 122.450 ;
        RECT 121.840 121.920 122.010 122.090 ;
        RECT 121.840 121.560 122.010 121.730 ;
        RECT 121.840 121.200 122.010 121.370 ;
        RECT 121.840 120.840 122.010 121.010 ;
        RECT 122.390 122.370 122.560 122.540 ;
        RECT 122.390 122.010 122.560 122.180 ;
        RECT 122.390 121.650 122.560 121.820 ;
        RECT 122.390 121.290 122.560 121.460 ;
        RECT 122.390 120.930 122.560 121.100 ;
        RECT 123.760 122.370 123.930 122.540 ;
        RECT 123.760 122.010 123.930 122.180 ;
        RECT 123.760 121.650 123.930 121.820 ;
        RECT 123.760 121.290 123.930 121.460 ;
        RECT 123.760 120.930 123.930 121.100 ;
        RECT 125.130 122.370 125.300 122.540 ;
        RECT 125.130 122.010 125.300 122.180 ;
        RECT 125.130 121.650 125.300 121.820 ;
        RECT 125.130 121.290 125.300 121.460 ;
        RECT 125.130 120.930 125.300 121.100 ;
        RECT 125.680 122.340 125.850 122.510 ;
        RECT 125.680 121.980 125.850 122.150 ;
        RECT 125.680 121.620 125.850 121.790 ;
        RECT 125.680 121.260 125.850 121.430 ;
        RECT 125.680 120.900 125.850 121.070 ;
        RECT 122.895 120.510 123.065 120.680 ;
        RECT 123.255 120.510 123.425 120.680 ;
        RECT 124.265 120.510 124.435 120.680 ;
        RECT 124.625 120.510 124.795 120.680 ;
        RECT 125.680 120.540 125.850 120.710 ;
        RECT 121.840 120.330 122.010 120.500 ;
        RECT 121.840 119.970 122.010 120.140 ;
        RECT 121.840 119.610 122.010 119.780 ;
        RECT 121.840 119.250 122.010 119.420 ;
        RECT 121.840 118.890 122.010 119.060 ;
        RECT 121.840 118.530 122.010 118.700 ;
        RECT 122.390 120.090 122.560 120.260 ;
        RECT 122.390 119.730 122.560 119.900 ;
        RECT 122.390 119.370 122.560 119.540 ;
        RECT 122.390 119.010 122.560 119.180 ;
        RECT 122.390 118.650 122.560 118.820 ;
        RECT 123.760 120.090 123.930 120.260 ;
        RECT 123.760 119.730 123.930 119.900 ;
        RECT 123.760 119.370 123.930 119.540 ;
        RECT 123.760 119.010 123.930 119.180 ;
        RECT 123.760 118.650 123.930 118.820 ;
        RECT 125.130 120.090 125.300 120.260 ;
        RECT 125.130 119.730 125.300 119.900 ;
        RECT 125.130 119.370 125.300 119.540 ;
        RECT 125.130 119.010 125.300 119.180 ;
        RECT 125.130 118.650 125.300 118.820 ;
        RECT 125.680 120.180 125.850 120.350 ;
        RECT 125.680 119.820 125.850 119.990 ;
        RECT 125.680 119.460 125.850 119.630 ;
        RECT 125.680 119.100 125.850 119.270 ;
        RECT 125.680 118.740 125.850 118.910 ;
        RECT 121.840 118.170 122.010 118.340 ;
        RECT 122.895 118.230 123.065 118.400 ;
        RECT 123.255 118.230 123.425 118.400 ;
        RECT 124.265 118.230 124.435 118.400 ;
        RECT 124.625 118.230 124.795 118.400 ;
        RECT 125.680 118.380 125.850 118.550 ;
        RECT 108.635 117.640 108.805 117.810 ;
        RECT 108.635 117.280 108.805 117.450 ;
        RECT 108.635 116.920 108.805 117.090 ;
        RECT 108.635 116.560 108.805 116.730 ;
        RECT 110.555 117.810 110.725 117.980 ;
        RECT 110.555 117.450 110.725 117.620 ;
        RECT 110.555 117.090 110.725 117.260 ;
        RECT 110.555 116.730 110.725 116.900 ;
        RECT 110.555 116.370 110.725 116.540 ;
        RECT 111.925 117.810 112.095 117.980 ;
        RECT 111.925 117.450 112.095 117.620 ;
        RECT 111.925 117.090 112.095 117.260 ;
        RECT 111.925 116.730 112.095 116.900 ;
        RECT 111.925 116.370 112.095 116.540 ;
        RECT 113.845 117.620 114.015 117.790 ;
        RECT 113.845 117.260 114.015 117.430 ;
        RECT 113.845 116.900 114.015 117.070 ;
        RECT 113.845 116.540 114.015 116.710 ;
        RECT 108.635 116.200 108.805 116.370 ;
        RECT 113.845 116.180 114.015 116.350 ;
        RECT 108.635 115.840 108.805 116.010 ;
        RECT 109.690 115.950 109.860 116.120 ;
        RECT 110.050 115.950 110.220 116.120 ;
        RECT 111.060 115.950 111.230 116.120 ;
        RECT 111.420 115.950 111.590 116.120 ;
        RECT 112.430 115.950 112.600 116.120 ;
        RECT 112.790 115.950 112.960 116.120 ;
        RECT 113.845 115.820 114.015 115.990 ;
        RECT 108.635 115.480 108.805 115.650 ;
        RECT 108.635 115.120 108.805 115.290 ;
        RECT 108.635 114.760 108.805 114.930 ;
        RECT 108.635 114.400 108.805 114.570 ;
        RECT 108.635 114.040 108.805 114.210 ;
        RECT 110.555 115.530 110.725 115.700 ;
        RECT 110.555 115.170 110.725 115.340 ;
        RECT 110.555 114.810 110.725 114.980 ;
        RECT 110.555 114.450 110.725 114.620 ;
        RECT 110.555 114.090 110.725 114.260 ;
        RECT 111.925 115.530 112.095 115.700 ;
        RECT 111.925 115.170 112.095 115.340 ;
        RECT 111.925 114.810 112.095 114.980 ;
        RECT 111.925 114.450 112.095 114.620 ;
        RECT 111.925 114.090 112.095 114.260 ;
        RECT 113.845 115.460 114.015 115.630 ;
        RECT 113.845 115.100 114.015 115.270 ;
        RECT 113.845 114.740 114.015 114.910 ;
        RECT 113.845 114.380 114.015 114.550 ;
        RECT 113.845 114.020 114.015 114.190 ;
        RECT 114.925 117.845 115.095 118.015 ;
        RECT 115.535 117.905 115.705 118.075 ;
        RECT 115.895 117.905 116.065 118.075 ;
        RECT 116.255 117.905 116.425 118.075 ;
        RECT 116.615 117.905 116.785 118.075 ;
        RECT 116.975 117.905 117.145 118.075 ;
        RECT 117.335 117.905 117.505 118.075 ;
        RECT 114.925 117.485 115.095 117.655 ;
        RECT 125.680 118.020 125.850 118.190 ;
        RECT 114.925 117.125 115.095 117.295 ;
        RECT 115.980 117.275 116.150 117.445 ;
        RECT 116.340 117.275 116.510 117.445 ;
        RECT 117.395 117.365 117.565 117.535 ;
        RECT 114.925 116.765 115.095 116.935 ;
        RECT 115.980 116.845 116.150 117.015 ;
        RECT 116.340 116.845 116.510 117.015 ;
        RECT 116.845 116.845 117.015 117.015 ;
        RECT 117.395 117.005 117.565 117.175 ;
        RECT 117.395 116.645 117.565 116.815 ;
        RECT 114.925 116.405 115.095 116.575 ;
        RECT 115.980 116.415 116.150 116.585 ;
        RECT 116.340 116.415 116.510 116.585 ;
        RECT 117.395 116.285 117.565 116.455 ;
        RECT 115.475 115.985 115.645 116.155 ;
        RECT 115.980 115.985 116.150 116.155 ;
        RECT 116.340 115.985 116.510 116.155 ;
        RECT 114.925 115.805 115.095 115.975 ;
        RECT 117.395 115.925 117.565 116.095 ;
        RECT 114.925 115.445 115.095 115.615 ;
        RECT 115.980 115.555 116.150 115.725 ;
        RECT 116.340 115.555 116.510 115.725 ;
        RECT 117.395 115.565 117.565 115.735 ;
        RECT 114.925 115.085 115.095 115.255 ;
        RECT 115.980 115.125 116.150 115.295 ;
        RECT 116.340 115.125 116.510 115.295 ;
        RECT 116.845 115.125 117.015 115.295 ;
        RECT 117.395 115.205 117.565 115.375 ;
        RECT 114.925 114.725 115.095 114.895 ;
        RECT 115.980 114.695 116.150 114.865 ;
        RECT 116.340 114.695 116.510 114.865 ;
        RECT 117.395 114.845 117.565 115.015 ;
        RECT 117.395 114.485 117.565 114.655 ;
        RECT 114.985 114.065 115.155 114.235 ;
        RECT 115.345 114.065 115.515 114.235 ;
        RECT 115.705 114.065 115.875 114.235 ;
        RECT 116.065 114.065 116.235 114.235 ;
        RECT 116.425 114.065 116.595 114.235 ;
        RECT 116.785 114.065 116.955 114.235 ;
        RECT 117.395 114.125 117.565 114.295 ;
        RECT 118.195 117.610 118.365 117.780 ;
        RECT 118.745 117.670 118.915 117.840 ;
        RECT 119.105 117.670 119.275 117.840 ;
        RECT 119.465 117.670 119.635 117.840 ;
        RECT 119.825 117.670 119.995 117.840 ;
        RECT 120.185 117.670 120.355 117.840 ;
        RECT 120.545 117.670 120.715 117.840 ;
        RECT 120.905 117.670 121.075 117.840 ;
        RECT 118.195 117.250 118.365 117.420 ;
        RECT 118.195 116.890 118.365 117.060 ;
        RECT 119.400 117.040 119.570 117.210 ;
        RECT 119.760 117.040 119.930 117.210 ;
        RECT 120.965 117.150 121.135 117.320 ;
        RECT 120.965 116.790 121.135 116.960 ;
        RECT 118.195 116.530 118.365 116.700 ;
        RECT 118.745 116.610 118.915 116.780 ;
        RECT 119.400 116.610 119.570 116.780 ;
        RECT 119.760 116.610 119.930 116.780 ;
        RECT 120.965 116.430 121.135 116.600 ;
        RECT 118.195 116.170 118.365 116.340 ;
        RECT 119.400 116.180 119.570 116.350 ;
        RECT 119.760 116.180 119.930 116.350 ;
        RECT 118.195 115.810 118.365 115.980 ;
        RECT 120.965 116.070 121.135 116.240 ;
        RECT 118.745 115.750 118.915 115.920 ;
        RECT 119.400 115.750 119.570 115.920 ;
        RECT 119.760 115.750 119.930 115.920 ;
        RECT 118.195 115.450 118.365 115.620 ;
        RECT 120.965 115.710 121.135 115.880 ;
        RECT 119.400 115.320 119.570 115.490 ;
        RECT 119.760 115.320 119.930 115.490 ;
        RECT 120.965 115.350 121.135 115.520 ;
        RECT 118.195 115.090 118.365 115.260 ;
        RECT 118.195 114.730 118.365 114.900 ;
        RECT 118.745 114.890 118.915 115.060 ;
        RECT 119.400 114.890 119.570 115.060 ;
        RECT 119.760 114.890 119.930 115.060 ;
        RECT 120.965 114.990 121.135 115.160 ;
        RECT 120.965 114.630 121.135 114.800 ;
        RECT 118.195 114.370 118.365 114.540 ;
        RECT 119.400 114.460 119.570 114.630 ;
        RECT 119.760 114.460 119.930 114.630 ;
        RECT 120.965 114.270 121.135 114.440 ;
        RECT 109.690 113.670 109.860 113.840 ;
        RECT 110.050 113.670 110.220 113.840 ;
        RECT 111.060 113.670 111.230 113.840 ;
        RECT 111.420 113.670 111.590 113.840 ;
        RECT 112.430 113.670 112.600 113.840 ;
        RECT 112.790 113.670 112.960 113.840 ;
        RECT 108.635 113.490 108.805 113.660 ;
        RECT 113.845 113.660 114.015 113.830 ;
        RECT 108.635 113.130 108.805 113.300 ;
        RECT 108.635 112.770 108.805 112.940 ;
        RECT 108.635 112.410 108.805 112.580 ;
        RECT 108.635 112.050 108.805 112.220 ;
        RECT 94.935 111.300 95.105 111.470 ;
        RECT 94.935 110.940 95.105 111.110 ;
        RECT 94.935 110.580 95.105 110.750 ;
        RECT 88.545 110.220 88.715 110.390 ;
        RECT 89.340 110.140 89.510 110.310 ;
        RECT 93.710 110.140 93.880 110.310 ;
        RECT 94.070 110.140 94.240 110.310 ;
        RECT 94.935 110.220 95.105 110.390 ;
        RECT 88.545 109.860 88.715 110.030 ;
        RECT 88.545 109.500 88.715 109.670 ;
        RECT 88.545 109.140 88.715 109.310 ;
        RECT 88.545 108.780 88.715 108.950 ;
        RECT 88.545 108.420 88.715 108.590 ;
        RECT 89.925 109.720 90.095 109.890 ;
        RECT 89.925 109.360 90.095 109.530 ;
        RECT 89.925 109.000 90.095 109.170 ;
        RECT 89.925 108.640 90.095 108.810 ;
        RECT 89.925 108.280 90.095 108.450 ;
        RECT 93.055 109.720 93.225 109.890 ;
        RECT 93.055 109.360 93.225 109.530 ;
        RECT 93.055 109.000 93.225 109.170 ;
        RECT 93.055 108.640 93.225 108.810 ;
        RECT 93.055 108.280 93.225 108.450 ;
        RECT 94.935 109.860 95.105 110.030 ;
        RECT 94.935 109.500 95.105 109.670 ;
        RECT 94.935 109.140 95.105 109.310 ;
        RECT 94.935 108.780 95.105 108.950 ;
        RECT 94.935 108.420 95.105 108.590 ;
        RECT 88.545 108.060 88.715 108.230 ;
        RECT 94.935 108.060 95.105 108.230 ;
        RECT 88.545 107.700 88.715 107.870 ;
        RECT 89.340 107.860 89.510 108.030 ;
        RECT 93.710 107.860 93.880 108.030 ;
        RECT 94.070 107.860 94.240 108.030 ;
        RECT 94.935 107.700 95.105 107.870 ;
        RECT 88.545 107.340 88.715 107.510 ;
        RECT 88.545 106.980 88.715 107.150 ;
        RECT 88.545 106.620 88.715 106.790 ;
        RECT 88.545 106.260 88.715 106.430 ;
        RECT 88.545 105.900 88.715 106.070 ;
        RECT 89.925 107.440 90.095 107.610 ;
        RECT 89.925 107.080 90.095 107.250 ;
        RECT 89.925 106.720 90.095 106.890 ;
        RECT 89.925 106.360 90.095 106.530 ;
        RECT 89.925 106.000 90.095 106.170 ;
        RECT 93.055 107.440 93.225 107.610 ;
        RECT 93.055 107.080 93.225 107.250 ;
        RECT 93.055 106.720 93.225 106.890 ;
        RECT 93.055 106.360 93.225 106.530 ;
        RECT 93.055 106.000 93.225 106.170 ;
        RECT 94.935 107.340 95.105 107.510 ;
        RECT 94.935 106.980 95.105 107.150 ;
        RECT 94.935 106.620 95.105 106.790 ;
        RECT 94.935 106.260 95.105 106.430 ;
        RECT 94.935 105.900 95.105 106.070 ;
        RECT 88.545 105.540 88.715 105.710 ;
        RECT 89.340 105.580 89.510 105.750 ;
        RECT 93.710 105.580 93.880 105.750 ;
        RECT 94.070 105.580 94.240 105.750 ;
        RECT 88.545 105.180 88.715 105.350 ;
        RECT 94.935 105.540 95.105 105.710 ;
        RECT 88.545 104.820 88.715 104.990 ;
        RECT 88.545 104.460 88.715 104.630 ;
        RECT 88.545 104.100 88.715 104.270 ;
        RECT 88.545 103.740 88.715 103.910 ;
        RECT 89.925 105.160 90.095 105.330 ;
        RECT 89.925 104.800 90.095 104.970 ;
        RECT 89.925 104.440 90.095 104.610 ;
        RECT 89.925 104.080 90.095 104.250 ;
        RECT 89.925 103.720 90.095 103.890 ;
        RECT 93.055 105.160 93.225 105.330 ;
        RECT 93.055 104.800 93.225 104.970 ;
        RECT 93.055 104.440 93.225 104.610 ;
        RECT 93.055 104.080 93.225 104.250 ;
        RECT 93.055 103.720 93.225 103.890 ;
        RECT 94.935 105.180 95.105 105.350 ;
        RECT 94.935 104.820 95.105 104.990 ;
        RECT 94.935 104.460 95.105 104.630 ;
        RECT 94.935 104.100 95.105 104.270 ;
        RECT 94.935 103.740 95.105 103.910 ;
        RECT 88.545 103.380 88.715 103.550 ;
        RECT 89.340 103.300 89.510 103.470 ;
        RECT 93.710 103.300 93.880 103.470 ;
        RECT 94.070 103.300 94.240 103.470 ;
        RECT 94.935 103.380 95.105 103.550 ;
        RECT 88.545 103.020 88.715 103.190 ;
        RECT 88.545 102.660 88.715 102.830 ;
        RECT 88.545 102.300 88.715 102.470 ;
        RECT 88.545 101.940 88.715 102.110 ;
        RECT 88.545 101.580 88.715 101.750 ;
        RECT 89.925 102.880 90.095 103.050 ;
        RECT 89.925 102.520 90.095 102.690 ;
        RECT 89.925 102.160 90.095 102.330 ;
        RECT 89.925 101.800 90.095 101.970 ;
        RECT 89.925 101.440 90.095 101.610 ;
        RECT 93.055 102.880 93.225 103.050 ;
        RECT 93.055 102.520 93.225 102.690 ;
        RECT 93.055 102.160 93.225 102.330 ;
        RECT 93.055 101.800 93.225 101.970 ;
        RECT 93.055 101.440 93.225 101.610 ;
        RECT 94.935 103.020 95.105 103.190 ;
        RECT 94.935 102.660 95.105 102.830 ;
        RECT 94.935 102.300 95.105 102.470 ;
        RECT 94.935 101.940 95.105 102.110 ;
        RECT 94.935 101.580 95.105 101.750 ;
        RECT 88.545 101.220 88.715 101.390 ;
        RECT 94.935 101.220 95.105 101.390 ;
        RECT 88.545 100.860 88.715 101.030 ;
        RECT 89.340 101.020 89.510 101.190 ;
        RECT 93.710 101.020 93.880 101.190 ;
        RECT 94.070 101.020 94.240 101.190 ;
        RECT 94.935 100.860 95.105 101.030 ;
        RECT 88.545 100.500 88.715 100.670 ;
        RECT 88.545 100.140 88.715 100.310 ;
        RECT 88.545 99.780 88.715 99.950 ;
        RECT 88.545 99.420 88.715 99.590 ;
        RECT 88.545 99.060 88.715 99.230 ;
        RECT 89.925 100.600 90.095 100.770 ;
        RECT 89.925 100.240 90.095 100.410 ;
        RECT 89.925 99.880 90.095 100.050 ;
        RECT 89.925 99.520 90.095 99.690 ;
        RECT 89.925 99.160 90.095 99.330 ;
        RECT 93.055 100.600 93.225 100.770 ;
        RECT 93.055 100.240 93.225 100.410 ;
        RECT 93.055 99.880 93.225 100.050 ;
        RECT 93.055 99.520 93.225 99.690 ;
        RECT 93.055 99.160 93.225 99.330 ;
        RECT 94.935 100.500 95.105 100.670 ;
        RECT 94.935 100.140 95.105 100.310 ;
        RECT 94.935 99.780 95.105 99.950 ;
        RECT 94.935 99.420 95.105 99.590 ;
        RECT 94.935 99.060 95.105 99.230 ;
        RECT 88.545 98.700 88.715 98.870 ;
        RECT 89.340 98.740 89.510 98.910 ;
        RECT 93.710 98.740 93.880 98.910 ;
        RECT 94.070 98.740 94.240 98.910 ;
        RECT 88.545 98.340 88.715 98.510 ;
        RECT 94.935 98.700 95.105 98.870 ;
        RECT 88.545 97.980 88.715 98.150 ;
        RECT 88.545 97.620 88.715 97.790 ;
        RECT 88.545 97.260 88.715 97.430 ;
        RECT 88.545 96.900 88.715 97.070 ;
        RECT 89.925 98.320 90.095 98.490 ;
        RECT 89.925 97.960 90.095 98.130 ;
        RECT 89.925 97.600 90.095 97.770 ;
        RECT 89.925 97.240 90.095 97.410 ;
        RECT 89.925 96.880 90.095 97.050 ;
        RECT 93.055 98.320 93.225 98.490 ;
        RECT 93.055 97.960 93.225 98.130 ;
        RECT 93.055 97.600 93.225 97.770 ;
        RECT 93.055 97.240 93.225 97.410 ;
        RECT 93.055 96.880 93.225 97.050 ;
        RECT 94.935 98.340 95.105 98.510 ;
        RECT 94.935 97.980 95.105 98.150 ;
        RECT 94.935 97.620 95.105 97.790 ;
        RECT 94.935 97.260 95.105 97.430 ;
        RECT 94.935 96.900 95.105 97.070 ;
        RECT 88.545 96.540 88.715 96.710 ;
        RECT 89.340 96.460 89.510 96.630 ;
        RECT 93.710 96.460 93.880 96.630 ;
        RECT 94.070 96.460 94.240 96.630 ;
        RECT 94.935 96.540 95.105 96.710 ;
        RECT 88.545 96.180 88.715 96.350 ;
        RECT 88.545 95.820 88.715 95.990 ;
        RECT 88.545 95.460 88.715 95.630 ;
        RECT 88.545 95.100 88.715 95.270 ;
        RECT 88.545 94.740 88.715 94.910 ;
        RECT 89.925 96.040 90.095 96.210 ;
        RECT 89.925 95.680 90.095 95.850 ;
        RECT 89.925 95.320 90.095 95.490 ;
        RECT 89.925 94.960 90.095 95.130 ;
        RECT 89.925 94.600 90.095 94.770 ;
        RECT 93.055 96.040 93.225 96.210 ;
        RECT 93.055 95.680 93.225 95.850 ;
        RECT 93.055 95.320 93.225 95.490 ;
        RECT 93.055 94.960 93.225 95.130 ;
        RECT 93.055 94.600 93.225 94.770 ;
        RECT 94.935 96.180 95.105 96.350 ;
        RECT 94.935 95.820 95.105 95.990 ;
        RECT 94.935 95.460 95.105 95.630 ;
        RECT 94.935 95.100 95.105 95.270 ;
        RECT 94.935 94.740 95.105 94.910 ;
        RECT 88.545 94.380 88.715 94.550 ;
        RECT 94.935 94.380 95.105 94.550 ;
        RECT 88.545 94.020 88.715 94.190 ;
        RECT 89.340 94.180 89.510 94.350 ;
        RECT 93.710 94.180 93.880 94.350 ;
        RECT 94.070 94.180 94.240 94.350 ;
        RECT 94.935 94.020 95.105 94.190 ;
        RECT 88.545 93.660 88.715 93.830 ;
        RECT 88.545 93.300 88.715 93.470 ;
        RECT 88.545 92.940 88.715 93.110 ;
        RECT 88.545 92.580 88.715 92.750 ;
        RECT 88.545 92.220 88.715 92.390 ;
        RECT 89.925 93.760 90.095 93.930 ;
        RECT 89.925 93.400 90.095 93.570 ;
        RECT 89.925 93.040 90.095 93.210 ;
        RECT 89.925 92.680 90.095 92.850 ;
        RECT 89.925 92.320 90.095 92.490 ;
        RECT 93.055 93.760 93.225 93.930 ;
        RECT 93.055 93.400 93.225 93.570 ;
        RECT 93.055 93.040 93.225 93.210 ;
        RECT 93.055 92.680 93.225 92.850 ;
        RECT 93.055 92.320 93.225 92.490 ;
        RECT 94.935 93.660 95.105 93.830 ;
        RECT 94.935 93.300 95.105 93.470 ;
        RECT 94.935 92.940 95.105 93.110 ;
        RECT 94.935 92.580 95.105 92.750 ;
        RECT 94.935 92.220 95.105 92.390 ;
        RECT 88.545 91.860 88.715 92.030 ;
        RECT 89.340 91.900 89.510 92.070 ;
        RECT 93.710 91.900 93.880 92.070 ;
        RECT 94.070 91.900 94.240 92.070 ;
        RECT 88.545 91.500 88.715 91.670 ;
        RECT 94.935 91.860 95.105 92.030 ;
        RECT 88.545 91.140 88.715 91.310 ;
        RECT 88.545 90.780 88.715 90.950 ;
        RECT 88.545 90.420 88.715 90.590 ;
        RECT 88.545 90.060 88.715 90.230 ;
        RECT 89.925 91.480 90.095 91.650 ;
        RECT 89.925 91.120 90.095 91.290 ;
        RECT 89.925 90.760 90.095 90.930 ;
        RECT 89.925 90.400 90.095 90.570 ;
        RECT 89.925 90.040 90.095 90.210 ;
        RECT 93.055 91.480 93.225 91.650 ;
        RECT 93.055 91.120 93.225 91.290 ;
        RECT 93.055 90.760 93.225 90.930 ;
        RECT 93.055 90.400 93.225 90.570 ;
        RECT 93.055 90.040 93.225 90.210 ;
        RECT 94.935 91.500 95.105 91.670 ;
        RECT 94.935 91.140 95.105 91.310 ;
        RECT 94.935 90.780 95.105 90.950 ;
        RECT 94.935 90.420 95.105 90.590 ;
        RECT 94.935 90.060 95.105 90.230 ;
        RECT 88.545 89.700 88.715 89.870 ;
        RECT 89.340 89.620 89.510 89.790 ;
        RECT 93.710 89.620 93.880 89.790 ;
        RECT 94.070 89.620 94.240 89.790 ;
        RECT 94.935 89.700 95.105 89.870 ;
        RECT 88.545 89.340 88.715 89.510 ;
        RECT 94.935 89.340 95.105 89.510 ;
        RECT 88.845 88.950 89.015 89.120 ;
        RECT 89.205 88.950 89.375 89.120 ;
        RECT 89.565 88.950 89.735 89.120 ;
        RECT 89.925 88.950 90.095 89.120 ;
        RECT 90.285 88.950 90.455 89.120 ;
        RECT 90.645 88.950 90.815 89.120 ;
        RECT 92.115 88.950 92.285 89.120 ;
        RECT 92.475 88.950 92.645 89.120 ;
        RECT 92.835 88.950 93.005 89.120 ;
        RECT 93.195 88.950 93.365 89.120 ;
        RECT 93.555 88.950 93.725 89.120 ;
        RECT 93.915 88.950 94.085 89.120 ;
        RECT 94.275 88.950 94.445 89.120 ;
        RECT 94.635 88.950 94.805 89.120 ;
        RECT 108.635 111.690 108.805 111.860 ;
        RECT 110.555 113.250 110.725 113.420 ;
        RECT 110.555 112.890 110.725 113.060 ;
        RECT 110.555 112.530 110.725 112.700 ;
        RECT 110.555 112.170 110.725 112.340 ;
        RECT 110.555 111.810 110.725 111.980 ;
        RECT 111.925 113.250 112.095 113.420 ;
        RECT 111.925 112.890 112.095 113.060 ;
        RECT 111.925 112.530 112.095 112.700 ;
        RECT 111.925 112.170 112.095 112.340 ;
        RECT 111.925 111.810 112.095 111.980 ;
        RECT 113.845 113.300 114.015 113.470 ;
        RECT 118.195 114.010 118.365 114.180 ;
        RECT 119.400 114.030 119.570 114.200 ;
        RECT 119.760 114.030 119.930 114.200 ;
        RECT 120.415 114.030 120.585 114.200 ;
        RECT 120.965 113.910 121.135 114.080 ;
        RECT 119.400 113.600 119.570 113.770 ;
        RECT 119.760 113.600 119.930 113.770 ;
        RECT 113.845 112.940 114.015 113.110 ;
        RECT 113.845 112.580 114.015 112.750 ;
        RECT 113.845 112.220 114.015 112.390 ;
        RECT 113.845 111.860 114.015 112.030 ;
        RECT 108.635 111.330 108.805 111.500 ;
        RECT 109.690 111.390 109.860 111.560 ;
        RECT 110.050 111.390 110.220 111.560 ;
        RECT 111.060 111.390 111.230 111.560 ;
        RECT 111.420 111.390 111.590 111.560 ;
        RECT 112.430 111.390 112.600 111.560 ;
        RECT 112.790 111.390 112.960 111.560 ;
        RECT 113.845 111.500 114.015 111.670 ;
        RECT 113.845 111.140 114.015 111.310 ;
        RECT 108.635 110.970 108.805 111.140 ;
        RECT 108.635 110.610 108.805 110.780 ;
        RECT 108.635 110.250 108.805 110.420 ;
        RECT 108.635 109.890 108.805 110.060 ;
        RECT 108.635 109.530 108.805 109.700 ;
        RECT 110.555 110.970 110.725 111.140 ;
        RECT 110.555 110.610 110.725 110.780 ;
        RECT 110.555 110.250 110.725 110.420 ;
        RECT 110.555 109.890 110.725 110.060 ;
        RECT 110.555 109.530 110.725 109.700 ;
        RECT 111.925 110.970 112.095 111.140 ;
        RECT 111.925 110.610 112.095 110.780 ;
        RECT 111.925 110.250 112.095 110.420 ;
        RECT 111.925 109.890 112.095 110.060 ;
        RECT 111.925 109.530 112.095 109.700 ;
        RECT 113.845 110.780 114.015 110.950 ;
        RECT 113.845 110.420 114.015 110.590 ;
        RECT 113.845 110.060 114.015 110.230 ;
        RECT 113.845 109.700 114.015 109.870 ;
        RECT 108.635 109.170 108.805 109.340 ;
        RECT 113.845 109.340 114.015 109.510 ;
        RECT 114.925 113.215 115.095 113.385 ;
        RECT 115.535 113.275 115.705 113.445 ;
        RECT 115.895 113.275 116.065 113.445 ;
        RECT 116.255 113.275 116.425 113.445 ;
        RECT 116.615 113.275 116.785 113.445 ;
        RECT 116.975 113.275 117.145 113.445 ;
        RECT 117.335 113.275 117.505 113.445 ;
        RECT 114.925 112.855 115.095 113.025 ;
        RECT 114.925 112.495 115.095 112.665 ;
        RECT 115.980 112.605 116.150 112.775 ;
        RECT 116.340 112.605 116.510 112.775 ;
        RECT 117.395 112.655 117.565 112.825 ;
        RECT 114.925 112.135 115.095 112.305 ;
        RECT 115.475 112.175 115.645 112.345 ;
        RECT 115.980 112.175 116.150 112.345 ;
        RECT 116.340 112.175 116.510 112.345 ;
        RECT 117.395 112.295 117.565 112.465 ;
        RECT 114.925 111.775 115.095 111.945 ;
        RECT 117.395 111.935 117.565 112.105 ;
        RECT 115.980 111.745 116.150 111.915 ;
        RECT 116.340 111.745 116.510 111.915 ;
        RECT 117.395 111.575 117.565 111.745 ;
        RECT 115.980 111.315 116.150 111.485 ;
        RECT 116.340 111.315 116.510 111.485 ;
        RECT 116.845 111.315 117.015 111.485 ;
        RECT 114.925 111.135 115.095 111.305 ;
        RECT 117.395 111.215 117.565 111.385 ;
        RECT 114.925 110.775 115.095 110.945 ;
        RECT 115.980 110.885 116.150 111.055 ;
        RECT 116.340 110.885 116.510 111.055 ;
        RECT 117.395 110.855 117.565 111.025 ;
        RECT 114.925 110.415 115.095 110.585 ;
        RECT 115.475 110.455 115.645 110.625 ;
        RECT 115.980 110.455 116.150 110.625 ;
        RECT 116.340 110.455 116.510 110.625 ;
        RECT 117.395 110.495 117.565 110.665 ;
        RECT 114.925 110.055 115.095 110.225 ;
        RECT 115.980 110.025 116.150 110.195 ;
        RECT 116.340 110.025 116.510 110.195 ;
        RECT 117.395 110.135 117.565 110.305 ;
        RECT 117.395 109.775 117.565 109.945 ;
        RECT 114.985 109.355 115.155 109.525 ;
        RECT 115.345 109.355 115.515 109.525 ;
        RECT 115.705 109.355 115.875 109.525 ;
        RECT 116.065 109.355 116.235 109.525 ;
        RECT 116.425 109.355 116.595 109.525 ;
        RECT 116.785 109.355 116.955 109.525 ;
        RECT 117.395 109.415 117.565 109.585 ;
        RECT 118.195 113.420 118.365 113.590 ;
        RECT 120.965 113.550 121.135 113.720 ;
        RECT 118.195 113.060 118.365 113.230 ;
        RECT 119.400 113.170 119.570 113.340 ;
        RECT 119.760 113.170 119.930 113.340 ;
        RECT 120.415 113.170 120.585 113.340 ;
        RECT 120.965 113.190 121.135 113.360 ;
        RECT 118.195 112.700 118.365 112.870 ;
        RECT 119.400 112.740 119.570 112.910 ;
        RECT 119.760 112.740 119.930 112.910 ;
        RECT 120.965 112.830 121.135 113.000 ;
        RECT 118.195 112.340 118.365 112.510 ;
        RECT 118.745 112.310 118.915 112.480 ;
        RECT 119.400 112.310 119.570 112.480 ;
        RECT 119.760 112.310 119.930 112.480 ;
        RECT 120.965 112.470 121.135 112.640 ;
        RECT 118.195 111.980 118.365 112.150 ;
        RECT 120.965 112.110 121.135 112.280 ;
        RECT 119.400 111.880 119.570 112.050 ;
        RECT 119.760 111.880 119.930 112.050 ;
        RECT 118.195 111.620 118.365 111.790 ;
        RECT 120.965 111.750 121.135 111.920 ;
        RECT 118.745 111.450 118.915 111.620 ;
        RECT 119.400 111.450 119.570 111.620 ;
        RECT 119.760 111.450 119.930 111.620 ;
        RECT 118.195 111.260 118.365 111.430 ;
        RECT 120.965 111.390 121.135 111.560 ;
        RECT 118.195 110.900 118.365 111.070 ;
        RECT 119.400 111.020 119.570 111.190 ;
        RECT 119.760 111.020 119.930 111.190 ;
        RECT 120.965 111.030 121.135 111.200 ;
        RECT 118.195 110.540 118.365 110.710 ;
        RECT 118.745 110.590 118.915 110.760 ;
        RECT 119.400 110.590 119.570 110.760 ;
        RECT 119.760 110.590 119.930 110.760 ;
        RECT 120.965 110.670 121.135 110.840 ;
        RECT 118.195 110.180 118.365 110.350 ;
        RECT 119.400 110.160 119.570 110.330 ;
        RECT 119.760 110.160 119.930 110.330 ;
        RECT 120.965 110.310 121.135 110.480 ;
        RECT 120.965 109.950 121.135 110.120 ;
        RECT 118.255 109.530 118.425 109.700 ;
        RECT 118.615 109.530 118.785 109.700 ;
        RECT 118.975 109.530 119.145 109.700 ;
        RECT 119.335 109.530 119.505 109.700 ;
        RECT 119.695 109.530 119.865 109.700 ;
        RECT 120.055 109.530 120.225 109.700 ;
        RECT 120.415 109.530 120.585 109.700 ;
        RECT 120.965 109.590 121.135 109.760 ;
        RECT 121.840 117.810 122.010 117.980 ;
        RECT 121.840 117.450 122.010 117.620 ;
        RECT 121.840 117.090 122.010 117.260 ;
        RECT 121.840 116.730 122.010 116.900 ;
        RECT 121.840 116.370 122.010 116.540 ;
        RECT 122.390 117.810 122.560 117.980 ;
        RECT 122.390 117.450 122.560 117.620 ;
        RECT 122.390 117.090 122.560 117.260 ;
        RECT 122.390 116.730 122.560 116.900 ;
        RECT 122.390 116.370 122.560 116.540 ;
        RECT 123.760 117.810 123.930 117.980 ;
        RECT 123.760 117.450 123.930 117.620 ;
        RECT 123.760 117.090 123.930 117.260 ;
        RECT 123.760 116.730 123.930 116.900 ;
        RECT 123.760 116.370 123.930 116.540 ;
        RECT 125.130 117.810 125.300 117.980 ;
        RECT 125.130 117.450 125.300 117.620 ;
        RECT 125.130 117.090 125.300 117.260 ;
        RECT 125.130 116.730 125.300 116.900 ;
        RECT 125.130 116.370 125.300 116.540 ;
        RECT 125.680 117.660 125.850 117.830 ;
        RECT 125.680 117.300 125.850 117.470 ;
        RECT 125.680 116.940 125.850 117.110 ;
        RECT 125.680 116.580 125.850 116.750 ;
        RECT 121.840 116.010 122.010 116.180 ;
        RECT 125.680 116.220 125.850 116.390 ;
        RECT 122.895 115.950 123.065 116.120 ;
        RECT 123.255 115.950 123.425 116.120 ;
        RECT 124.265 115.950 124.435 116.120 ;
        RECT 124.625 115.950 124.795 116.120 ;
        RECT 121.840 115.650 122.010 115.820 ;
        RECT 125.680 115.860 125.850 116.030 ;
        RECT 121.840 115.290 122.010 115.460 ;
        RECT 121.840 114.930 122.010 115.100 ;
        RECT 121.840 114.570 122.010 114.740 ;
        RECT 121.840 114.210 122.010 114.380 ;
        RECT 122.390 115.530 122.560 115.700 ;
        RECT 122.390 115.170 122.560 115.340 ;
        RECT 122.390 114.810 122.560 114.980 ;
        RECT 122.390 114.450 122.560 114.620 ;
        RECT 122.390 114.090 122.560 114.260 ;
        RECT 123.760 115.530 123.930 115.700 ;
        RECT 123.760 115.170 123.930 115.340 ;
        RECT 123.760 114.810 123.930 114.980 ;
        RECT 123.760 114.450 123.930 114.620 ;
        RECT 123.760 114.090 123.930 114.260 ;
        RECT 125.130 115.530 125.300 115.700 ;
        RECT 125.130 115.170 125.300 115.340 ;
        RECT 125.130 114.810 125.300 114.980 ;
        RECT 125.130 114.450 125.300 114.620 ;
        RECT 125.130 114.090 125.300 114.260 ;
        RECT 125.680 115.500 125.850 115.670 ;
        RECT 125.680 115.140 125.850 115.310 ;
        RECT 125.680 114.780 125.850 114.950 ;
        RECT 125.680 114.420 125.850 114.590 ;
        RECT 121.840 113.850 122.010 114.020 ;
        RECT 125.680 114.060 125.850 114.230 ;
        RECT 122.895 113.670 123.065 113.840 ;
        RECT 123.255 113.670 123.425 113.840 ;
        RECT 124.265 113.670 124.435 113.840 ;
        RECT 124.625 113.670 124.795 113.840 ;
        RECT 125.680 113.700 125.850 113.870 ;
        RECT 121.840 113.490 122.010 113.660 ;
        RECT 121.840 113.130 122.010 113.300 ;
        RECT 121.840 112.770 122.010 112.940 ;
        RECT 121.840 112.410 122.010 112.580 ;
        RECT 121.840 112.050 122.010 112.220 ;
        RECT 121.840 111.690 122.010 111.860 ;
        RECT 122.390 113.250 122.560 113.420 ;
        RECT 122.390 112.890 122.560 113.060 ;
        RECT 122.390 112.530 122.560 112.700 ;
        RECT 122.390 112.170 122.560 112.340 ;
        RECT 122.390 111.810 122.560 111.980 ;
        RECT 123.760 113.250 123.930 113.420 ;
        RECT 123.760 112.890 123.930 113.060 ;
        RECT 123.760 112.530 123.930 112.700 ;
        RECT 123.760 112.170 123.930 112.340 ;
        RECT 123.760 111.810 123.930 111.980 ;
        RECT 125.130 113.250 125.300 113.420 ;
        RECT 125.130 112.890 125.300 113.060 ;
        RECT 125.130 112.530 125.300 112.700 ;
        RECT 125.130 112.170 125.300 112.340 ;
        RECT 125.130 111.810 125.300 111.980 ;
        RECT 125.680 113.340 125.850 113.510 ;
        RECT 125.680 112.980 125.850 113.150 ;
        RECT 125.680 112.620 125.850 112.790 ;
        RECT 125.680 112.260 125.850 112.430 ;
        RECT 125.680 111.900 125.850 112.070 ;
        RECT 121.840 111.330 122.010 111.500 ;
        RECT 122.895 111.390 123.065 111.560 ;
        RECT 123.255 111.390 123.425 111.560 ;
        RECT 124.265 111.390 124.435 111.560 ;
        RECT 124.625 111.390 124.795 111.560 ;
        RECT 125.680 111.540 125.850 111.710 ;
        RECT 125.680 111.180 125.850 111.350 ;
        RECT 121.840 110.970 122.010 111.140 ;
        RECT 121.840 110.610 122.010 110.780 ;
        RECT 121.840 110.250 122.010 110.420 ;
        RECT 121.840 109.890 122.010 110.060 ;
        RECT 121.840 109.530 122.010 109.700 ;
        RECT 122.390 110.970 122.560 111.140 ;
        RECT 122.390 110.610 122.560 110.780 ;
        RECT 122.390 110.250 122.560 110.420 ;
        RECT 122.390 109.890 122.560 110.060 ;
        RECT 122.390 109.530 122.560 109.700 ;
        RECT 123.760 110.970 123.930 111.140 ;
        RECT 123.760 110.610 123.930 110.780 ;
        RECT 123.760 110.250 123.930 110.420 ;
        RECT 123.760 109.890 123.930 110.060 ;
        RECT 123.760 109.530 123.930 109.700 ;
        RECT 125.130 110.970 125.300 111.140 ;
        RECT 125.130 110.610 125.300 110.780 ;
        RECT 125.130 110.250 125.300 110.420 ;
        RECT 125.130 109.890 125.300 110.060 ;
        RECT 125.130 109.530 125.300 109.700 ;
        RECT 125.680 110.820 125.850 110.990 ;
        RECT 125.680 110.460 125.850 110.630 ;
        RECT 125.680 110.100 125.850 110.270 ;
        RECT 125.680 109.740 125.850 109.910 ;
        RECT 109.690 109.110 109.860 109.280 ;
        RECT 110.050 109.110 110.220 109.280 ;
        RECT 111.060 109.110 111.230 109.280 ;
        RECT 111.420 109.110 111.590 109.280 ;
        RECT 112.430 109.110 112.600 109.280 ;
        RECT 112.790 109.110 112.960 109.280 ;
        RECT 108.635 108.810 108.805 108.980 ;
        RECT 113.845 108.980 114.015 109.150 ;
        RECT 108.635 108.450 108.805 108.620 ;
        RECT 108.635 108.090 108.805 108.260 ;
        RECT 108.635 107.730 108.805 107.900 ;
        RECT 108.635 107.370 108.805 107.540 ;
        RECT 110.555 108.690 110.725 108.860 ;
        RECT 110.555 108.330 110.725 108.500 ;
        RECT 110.555 107.970 110.725 108.140 ;
        RECT 110.555 107.610 110.725 107.780 ;
        RECT 110.555 107.250 110.725 107.420 ;
        RECT 111.925 108.690 112.095 108.860 ;
        RECT 111.925 108.330 112.095 108.500 ;
        RECT 111.925 107.970 112.095 108.140 ;
        RECT 111.925 107.610 112.095 107.780 ;
        RECT 111.925 107.250 112.095 107.420 ;
        RECT 113.845 108.620 114.015 108.790 ;
        RECT 113.845 108.260 114.015 108.430 ;
        RECT 113.845 107.900 114.015 108.070 ;
        RECT 113.845 107.540 114.015 107.710 ;
        RECT 108.635 107.010 108.805 107.180 ;
        RECT 113.845 107.180 114.015 107.350 ;
        RECT 109.690 106.830 109.860 107.000 ;
        RECT 110.050 106.830 110.220 107.000 ;
        RECT 111.060 106.830 111.230 107.000 ;
        RECT 111.420 106.830 111.590 107.000 ;
        RECT 112.430 106.830 112.600 107.000 ;
        RECT 112.790 106.830 112.960 107.000 ;
        RECT 108.635 106.650 108.805 106.820 ;
        RECT 113.845 106.820 114.015 106.990 ;
        RECT 108.635 106.290 108.805 106.460 ;
        RECT 108.635 105.930 108.805 106.100 ;
        RECT 108.635 105.570 108.805 105.740 ;
        RECT 108.635 105.210 108.805 105.380 ;
        RECT 108.635 104.850 108.805 105.020 ;
        RECT 110.555 106.410 110.725 106.580 ;
        RECT 110.555 106.050 110.725 106.220 ;
        RECT 110.555 105.690 110.725 105.860 ;
        RECT 110.555 105.330 110.725 105.500 ;
        RECT 110.555 104.970 110.725 105.140 ;
        RECT 111.925 106.410 112.095 106.580 ;
        RECT 111.925 106.050 112.095 106.220 ;
        RECT 111.925 105.690 112.095 105.860 ;
        RECT 111.925 105.330 112.095 105.500 ;
        RECT 111.925 104.970 112.095 105.140 ;
        RECT 113.845 106.460 114.015 106.630 ;
        RECT 113.845 106.100 114.015 106.270 ;
        RECT 113.845 105.740 114.015 105.910 ;
        RECT 113.845 105.380 114.015 105.550 ;
        RECT 113.845 105.020 114.015 105.190 ;
        RECT 108.635 104.490 108.805 104.660 ;
        RECT 109.690 104.550 109.860 104.720 ;
        RECT 110.050 104.550 110.220 104.720 ;
        RECT 111.060 104.550 111.230 104.720 ;
        RECT 111.420 104.550 111.590 104.720 ;
        RECT 112.430 104.550 112.600 104.720 ;
        RECT 112.790 104.550 112.960 104.720 ;
        RECT 113.845 104.660 114.015 104.830 ;
        RECT 113.845 104.300 114.015 104.470 ;
        RECT 108.635 104.130 108.805 104.300 ;
        RECT 108.635 103.770 108.805 103.940 ;
        RECT 108.635 103.410 108.805 103.580 ;
        RECT 108.635 103.050 108.805 103.220 ;
        RECT 108.635 102.690 108.805 102.860 ;
        RECT 110.555 104.130 110.725 104.300 ;
        RECT 110.555 103.770 110.725 103.940 ;
        RECT 110.555 103.410 110.725 103.580 ;
        RECT 110.555 103.050 110.725 103.220 ;
        RECT 110.555 102.690 110.725 102.860 ;
        RECT 111.925 104.130 112.095 104.300 ;
        RECT 111.925 103.770 112.095 103.940 ;
        RECT 111.925 103.410 112.095 103.580 ;
        RECT 111.925 103.050 112.095 103.220 ;
        RECT 111.925 102.690 112.095 102.860 ;
        RECT 113.845 103.940 114.015 104.110 ;
        RECT 113.845 103.580 114.015 103.750 ;
        RECT 113.845 103.220 114.015 103.390 ;
        RECT 113.845 102.860 114.015 103.030 ;
        RECT 108.635 102.330 108.805 102.500 ;
        RECT 113.845 102.500 114.015 102.670 ;
        RECT 109.690 102.270 109.860 102.440 ;
        RECT 110.050 102.270 110.220 102.440 ;
        RECT 111.060 102.270 111.230 102.440 ;
        RECT 111.420 102.270 111.590 102.440 ;
        RECT 112.430 102.270 112.600 102.440 ;
        RECT 112.790 102.270 112.960 102.440 ;
        RECT 108.635 101.970 108.805 102.140 ;
        RECT 113.845 102.140 114.015 102.310 ;
        RECT 108.635 101.610 108.805 101.780 ;
        RECT 108.635 101.250 108.805 101.420 ;
        RECT 108.635 100.890 108.805 101.060 ;
        RECT 108.635 100.530 108.805 100.700 ;
        RECT 110.555 101.850 110.725 102.020 ;
        RECT 110.555 101.490 110.725 101.660 ;
        RECT 110.555 101.130 110.725 101.300 ;
        RECT 110.555 100.770 110.725 100.940 ;
        RECT 110.555 100.410 110.725 100.580 ;
        RECT 111.925 101.850 112.095 102.020 ;
        RECT 111.925 101.490 112.095 101.660 ;
        RECT 111.925 101.130 112.095 101.300 ;
        RECT 111.925 100.770 112.095 100.940 ;
        RECT 111.925 100.410 112.095 100.580 ;
        RECT 113.845 101.780 114.015 101.950 ;
        RECT 113.845 101.420 114.015 101.590 ;
        RECT 113.845 101.060 114.015 101.230 ;
        RECT 113.845 100.700 114.015 100.870 ;
        RECT 108.635 100.170 108.805 100.340 ;
        RECT 113.845 100.340 114.015 100.510 ;
        RECT 109.690 99.990 109.860 100.160 ;
        RECT 110.050 99.990 110.220 100.160 ;
        RECT 111.060 99.990 111.230 100.160 ;
        RECT 111.420 99.990 111.590 100.160 ;
        RECT 112.430 99.990 112.600 100.160 ;
        RECT 112.790 99.990 112.960 100.160 ;
        RECT 108.635 99.810 108.805 99.980 ;
        RECT 113.845 99.980 114.015 100.150 ;
        RECT 108.635 99.450 108.805 99.620 ;
        RECT 108.635 99.090 108.805 99.260 ;
        RECT 108.635 98.730 108.805 98.900 ;
        RECT 108.635 98.370 108.805 98.540 ;
        RECT 108.635 98.010 108.805 98.180 ;
        RECT 110.555 99.570 110.725 99.740 ;
        RECT 110.555 99.210 110.725 99.380 ;
        RECT 110.555 98.850 110.725 99.020 ;
        RECT 110.555 98.490 110.725 98.660 ;
        RECT 110.555 98.130 110.725 98.300 ;
        RECT 111.925 99.570 112.095 99.740 ;
        RECT 111.925 99.210 112.095 99.380 ;
        RECT 111.925 98.850 112.095 99.020 ;
        RECT 111.925 98.490 112.095 98.660 ;
        RECT 111.925 98.130 112.095 98.300 ;
        RECT 113.845 99.620 114.015 99.790 ;
        RECT 113.845 99.260 114.015 99.430 ;
        RECT 113.845 98.900 114.015 99.070 ;
        RECT 113.845 98.540 114.015 98.710 ;
        RECT 113.845 98.180 114.015 98.350 ;
        RECT 108.635 97.650 108.805 97.820 ;
        RECT 109.690 97.710 109.860 97.880 ;
        RECT 110.050 97.710 110.220 97.880 ;
        RECT 111.060 97.710 111.230 97.880 ;
        RECT 111.420 97.710 111.590 97.880 ;
        RECT 112.430 97.710 112.600 97.880 ;
        RECT 112.790 97.710 112.960 97.880 ;
        RECT 113.845 97.820 114.015 97.990 ;
        RECT 113.845 97.460 114.015 97.630 ;
        RECT 108.635 97.290 108.805 97.460 ;
        RECT 108.635 96.930 108.805 97.100 ;
        RECT 108.635 96.570 108.805 96.740 ;
        RECT 108.635 96.210 108.805 96.380 ;
        RECT 108.635 95.850 108.805 96.020 ;
        RECT 110.555 97.290 110.725 97.460 ;
        RECT 110.555 96.930 110.725 97.100 ;
        RECT 110.555 96.570 110.725 96.740 ;
        RECT 110.555 96.210 110.725 96.380 ;
        RECT 110.555 95.850 110.725 96.020 ;
        RECT 111.925 97.290 112.095 97.460 ;
        RECT 111.925 96.930 112.095 97.100 ;
        RECT 111.925 96.570 112.095 96.740 ;
        RECT 111.925 96.210 112.095 96.380 ;
        RECT 111.925 95.850 112.095 96.020 ;
        RECT 113.845 97.100 114.015 97.270 ;
        RECT 113.845 96.740 114.015 96.910 ;
        RECT 113.845 96.380 114.015 96.550 ;
        RECT 113.845 96.020 114.015 96.190 ;
        RECT 108.635 95.490 108.805 95.660 ;
        RECT 113.845 95.660 114.015 95.830 ;
        RECT 109.690 95.430 109.860 95.600 ;
        RECT 110.050 95.430 110.220 95.600 ;
        RECT 111.060 95.430 111.230 95.600 ;
        RECT 111.420 95.430 111.590 95.600 ;
        RECT 112.430 95.430 112.600 95.600 ;
        RECT 112.790 95.430 112.960 95.600 ;
        RECT 108.635 95.130 108.805 95.300 ;
        RECT 113.845 95.300 114.015 95.470 ;
        RECT 108.635 94.770 108.805 94.940 ;
        RECT 108.635 94.410 108.805 94.580 ;
        RECT 108.635 94.050 108.805 94.220 ;
        RECT 108.635 93.690 108.805 93.860 ;
        RECT 110.555 95.010 110.725 95.180 ;
        RECT 110.555 94.650 110.725 94.820 ;
        RECT 110.555 94.290 110.725 94.460 ;
        RECT 110.555 93.930 110.725 94.100 ;
        RECT 110.555 93.570 110.725 93.740 ;
        RECT 111.925 95.010 112.095 95.180 ;
        RECT 111.925 94.650 112.095 94.820 ;
        RECT 111.925 94.290 112.095 94.460 ;
        RECT 111.925 93.930 112.095 94.100 ;
        RECT 111.925 93.570 112.095 93.740 ;
        RECT 113.845 94.940 114.015 95.110 ;
        RECT 113.845 94.580 114.015 94.750 ;
        RECT 113.845 94.220 114.015 94.390 ;
        RECT 113.845 93.860 114.015 94.030 ;
        RECT 108.635 93.330 108.805 93.500 ;
        RECT 113.845 93.500 114.015 93.670 ;
        RECT 109.690 93.150 109.860 93.320 ;
        RECT 110.050 93.150 110.220 93.320 ;
        RECT 111.060 93.150 111.230 93.320 ;
        RECT 111.420 93.150 111.590 93.320 ;
        RECT 112.430 93.150 112.600 93.320 ;
        RECT 112.790 93.150 112.960 93.320 ;
        RECT 108.635 92.970 108.805 93.140 ;
        RECT 113.845 93.140 114.015 93.310 ;
        RECT 108.635 92.610 108.805 92.780 ;
        RECT 108.635 92.250 108.805 92.420 ;
        RECT 108.635 91.890 108.805 92.060 ;
        RECT 108.635 91.530 108.805 91.700 ;
        RECT 108.635 91.170 108.805 91.340 ;
        RECT 110.555 92.730 110.725 92.900 ;
        RECT 110.555 92.370 110.725 92.540 ;
        RECT 110.555 92.010 110.725 92.180 ;
        RECT 110.555 91.650 110.725 91.820 ;
        RECT 110.555 91.290 110.725 91.460 ;
        RECT 111.925 92.730 112.095 92.900 ;
        RECT 111.925 92.370 112.095 92.540 ;
        RECT 111.925 92.010 112.095 92.180 ;
        RECT 111.925 91.650 112.095 91.820 ;
        RECT 111.925 91.290 112.095 91.460 ;
        RECT 113.845 92.780 114.015 92.950 ;
        RECT 113.845 92.420 114.015 92.590 ;
        RECT 113.845 92.060 114.015 92.230 ;
        RECT 113.845 91.700 114.015 91.870 ;
        RECT 113.845 91.340 114.015 91.510 ;
        RECT 108.635 90.810 108.805 90.980 ;
        RECT 109.690 90.870 109.860 91.040 ;
        RECT 110.050 90.870 110.220 91.040 ;
        RECT 111.060 90.870 111.230 91.040 ;
        RECT 111.420 90.870 111.590 91.040 ;
        RECT 112.430 90.870 112.600 91.040 ;
        RECT 112.790 90.870 112.960 91.040 ;
        RECT 113.845 90.980 114.015 91.150 ;
        RECT 113.845 90.620 114.015 90.790 ;
        RECT 108.635 90.450 108.805 90.620 ;
        RECT 108.635 90.090 108.805 90.260 ;
        RECT 108.635 89.730 108.805 89.900 ;
        RECT 108.635 89.370 108.805 89.540 ;
        RECT 108.635 89.010 108.805 89.180 ;
        RECT 110.555 90.450 110.725 90.620 ;
        RECT 110.555 90.090 110.725 90.260 ;
        RECT 110.555 89.730 110.725 89.900 ;
        RECT 110.555 89.370 110.725 89.540 ;
        RECT 110.555 89.010 110.725 89.180 ;
        RECT 111.925 90.450 112.095 90.620 ;
        RECT 111.925 90.090 112.095 90.260 ;
        RECT 111.925 89.730 112.095 89.900 ;
        RECT 111.925 89.370 112.095 89.540 ;
        RECT 111.925 89.010 112.095 89.180 ;
        RECT 113.845 90.260 114.015 90.430 ;
        RECT 113.845 89.900 114.015 90.070 ;
        RECT 113.845 89.540 114.015 89.710 ;
        RECT 113.845 89.180 114.015 89.350 ;
        RECT 108.635 88.650 108.805 88.820 ;
        RECT 113.845 88.820 114.015 88.990 ;
        RECT 109.690 88.590 109.860 88.760 ;
        RECT 110.050 88.590 110.220 88.760 ;
        RECT 111.060 88.590 111.230 88.760 ;
        RECT 111.420 88.590 111.590 88.760 ;
        RECT 112.430 88.590 112.600 88.760 ;
        RECT 112.790 88.590 112.960 88.760 ;
        RECT 108.635 88.290 108.805 88.460 ;
        RECT 113.845 88.460 114.015 88.630 ;
        RECT 108.635 87.930 108.805 88.100 ;
        RECT 108.635 87.570 108.805 87.740 ;
        RECT 108.635 87.210 108.805 87.380 ;
        RECT 108.635 86.850 108.805 87.020 ;
        RECT 110.555 88.170 110.725 88.340 ;
        RECT 110.555 87.810 110.725 87.980 ;
        RECT 110.555 87.450 110.725 87.620 ;
        RECT 110.555 87.090 110.725 87.260 ;
        RECT 110.555 86.730 110.725 86.900 ;
        RECT 111.925 88.170 112.095 88.340 ;
        RECT 111.925 87.810 112.095 87.980 ;
        RECT 111.925 87.450 112.095 87.620 ;
        RECT 111.925 87.090 112.095 87.260 ;
        RECT 111.925 86.730 112.095 86.900 ;
        RECT 113.845 88.100 114.015 88.270 ;
        RECT 113.845 87.740 114.015 87.910 ;
        RECT 113.845 87.380 114.015 87.550 ;
        RECT 113.845 87.020 114.015 87.190 ;
        RECT 108.635 86.490 108.805 86.660 ;
        RECT 113.845 86.660 114.015 86.830 ;
        RECT 109.690 86.310 109.860 86.480 ;
        RECT 110.050 86.310 110.220 86.480 ;
        RECT 111.060 86.310 111.230 86.480 ;
        RECT 111.420 86.310 111.590 86.480 ;
        RECT 112.430 86.310 112.600 86.480 ;
        RECT 112.790 86.310 112.960 86.480 ;
        RECT 108.635 86.130 108.805 86.300 ;
        RECT 113.845 86.300 114.015 86.470 ;
        RECT 108.635 85.770 108.805 85.940 ;
        RECT 108.635 85.410 108.805 85.580 ;
        RECT 108.635 85.050 108.805 85.220 ;
        RECT 108.635 84.690 108.805 84.860 ;
        RECT 108.635 84.330 108.805 84.500 ;
        RECT 110.555 85.890 110.725 86.060 ;
        RECT 110.555 85.530 110.725 85.700 ;
        RECT 110.555 85.170 110.725 85.340 ;
        RECT 110.555 84.810 110.725 84.980 ;
        RECT 110.555 84.450 110.725 84.620 ;
        RECT 111.925 85.890 112.095 86.060 ;
        RECT 111.925 85.530 112.095 85.700 ;
        RECT 111.925 85.170 112.095 85.340 ;
        RECT 111.925 84.810 112.095 84.980 ;
        RECT 111.925 84.450 112.095 84.620 ;
        RECT 113.845 85.940 114.015 86.110 ;
        RECT 113.845 85.580 114.015 85.750 ;
        RECT 113.845 85.220 114.015 85.390 ;
        RECT 113.845 84.860 114.015 85.030 ;
        RECT 113.845 84.500 114.015 84.670 ;
        RECT 108.635 83.970 108.805 84.140 ;
        RECT 109.690 84.030 109.860 84.200 ;
        RECT 110.050 84.030 110.220 84.200 ;
        RECT 111.060 84.030 111.230 84.200 ;
        RECT 111.420 84.030 111.590 84.200 ;
        RECT 112.430 84.030 112.600 84.200 ;
        RECT 112.790 84.030 112.960 84.200 ;
        RECT 113.845 84.140 114.015 84.310 ;
        RECT 113.845 83.780 114.015 83.950 ;
        RECT 121.840 109.170 122.010 109.340 ;
        RECT 125.680 109.380 125.850 109.550 ;
        RECT 122.895 109.110 123.065 109.280 ;
        RECT 123.255 109.110 123.425 109.280 ;
        RECT 124.265 109.110 124.435 109.280 ;
        RECT 124.625 109.110 124.795 109.280 ;
        RECT 121.840 108.810 122.010 108.980 ;
        RECT 125.680 109.020 125.850 109.190 ;
        RECT 121.840 108.450 122.010 108.620 ;
        RECT 121.840 108.090 122.010 108.260 ;
        RECT 121.840 107.730 122.010 107.900 ;
        RECT 121.840 107.370 122.010 107.540 ;
        RECT 122.390 108.690 122.560 108.860 ;
        RECT 122.390 108.330 122.560 108.500 ;
        RECT 122.390 107.970 122.560 108.140 ;
        RECT 122.390 107.610 122.560 107.780 ;
        RECT 122.390 107.250 122.560 107.420 ;
        RECT 123.760 108.690 123.930 108.860 ;
        RECT 123.760 108.330 123.930 108.500 ;
        RECT 123.760 107.970 123.930 108.140 ;
        RECT 123.760 107.610 123.930 107.780 ;
        RECT 123.760 107.250 123.930 107.420 ;
        RECT 125.130 108.690 125.300 108.860 ;
        RECT 125.130 108.330 125.300 108.500 ;
        RECT 125.130 107.970 125.300 108.140 ;
        RECT 125.130 107.610 125.300 107.780 ;
        RECT 125.130 107.250 125.300 107.420 ;
        RECT 125.680 108.660 125.850 108.830 ;
        RECT 125.680 108.300 125.850 108.470 ;
        RECT 125.680 107.940 125.850 108.110 ;
        RECT 125.680 107.580 125.850 107.750 ;
        RECT 121.840 107.010 122.010 107.180 ;
        RECT 125.680 107.220 125.850 107.390 ;
        RECT 122.895 106.830 123.065 107.000 ;
        RECT 123.255 106.830 123.425 107.000 ;
        RECT 124.265 106.830 124.435 107.000 ;
        RECT 124.625 106.830 124.795 107.000 ;
        RECT 125.680 106.860 125.850 107.030 ;
        RECT 121.840 106.650 122.010 106.820 ;
        RECT 121.840 106.290 122.010 106.460 ;
        RECT 121.840 105.930 122.010 106.100 ;
        RECT 121.840 105.570 122.010 105.740 ;
        RECT 121.840 105.210 122.010 105.380 ;
        RECT 121.840 104.850 122.010 105.020 ;
        RECT 122.390 106.410 122.560 106.580 ;
        RECT 122.390 106.050 122.560 106.220 ;
        RECT 122.390 105.690 122.560 105.860 ;
        RECT 122.390 105.330 122.560 105.500 ;
        RECT 122.390 104.970 122.560 105.140 ;
        RECT 123.760 106.410 123.930 106.580 ;
        RECT 123.760 106.050 123.930 106.220 ;
        RECT 123.760 105.690 123.930 105.860 ;
        RECT 123.760 105.330 123.930 105.500 ;
        RECT 123.760 104.970 123.930 105.140 ;
        RECT 125.130 106.410 125.300 106.580 ;
        RECT 125.130 106.050 125.300 106.220 ;
        RECT 125.130 105.690 125.300 105.860 ;
        RECT 125.130 105.330 125.300 105.500 ;
        RECT 125.130 104.970 125.300 105.140 ;
        RECT 125.680 106.500 125.850 106.670 ;
        RECT 125.680 106.140 125.850 106.310 ;
        RECT 125.680 105.780 125.850 105.950 ;
        RECT 125.680 105.420 125.850 105.590 ;
        RECT 125.680 105.060 125.850 105.230 ;
        RECT 121.840 104.490 122.010 104.660 ;
        RECT 122.895 104.550 123.065 104.720 ;
        RECT 123.255 104.550 123.425 104.720 ;
        RECT 124.265 104.550 124.435 104.720 ;
        RECT 124.625 104.550 124.795 104.720 ;
        RECT 125.680 104.700 125.850 104.870 ;
        RECT 125.680 104.340 125.850 104.510 ;
        RECT 121.840 104.130 122.010 104.300 ;
        RECT 121.840 103.770 122.010 103.940 ;
        RECT 121.840 103.410 122.010 103.580 ;
        RECT 121.840 103.050 122.010 103.220 ;
        RECT 121.840 102.690 122.010 102.860 ;
        RECT 122.390 104.130 122.560 104.300 ;
        RECT 122.390 103.770 122.560 103.940 ;
        RECT 122.390 103.410 122.560 103.580 ;
        RECT 122.390 103.050 122.560 103.220 ;
        RECT 122.390 102.690 122.560 102.860 ;
        RECT 123.760 104.130 123.930 104.300 ;
        RECT 123.760 103.770 123.930 103.940 ;
        RECT 123.760 103.410 123.930 103.580 ;
        RECT 123.760 103.050 123.930 103.220 ;
        RECT 123.760 102.690 123.930 102.860 ;
        RECT 125.130 104.130 125.300 104.300 ;
        RECT 125.130 103.770 125.300 103.940 ;
        RECT 125.130 103.410 125.300 103.580 ;
        RECT 125.130 103.050 125.300 103.220 ;
        RECT 125.130 102.690 125.300 102.860 ;
        RECT 125.680 103.980 125.850 104.150 ;
        RECT 125.680 103.620 125.850 103.790 ;
        RECT 125.680 103.260 125.850 103.430 ;
        RECT 125.680 102.900 125.850 103.070 ;
        RECT 121.840 102.330 122.010 102.500 ;
        RECT 125.680 102.540 125.850 102.710 ;
        RECT 122.895 102.270 123.065 102.440 ;
        RECT 123.255 102.270 123.425 102.440 ;
        RECT 124.265 102.270 124.435 102.440 ;
        RECT 124.625 102.270 124.795 102.440 ;
        RECT 121.840 101.970 122.010 102.140 ;
        RECT 125.680 102.180 125.850 102.350 ;
        RECT 121.840 101.610 122.010 101.780 ;
        RECT 121.840 101.250 122.010 101.420 ;
        RECT 121.840 100.890 122.010 101.060 ;
        RECT 121.840 100.530 122.010 100.700 ;
        RECT 122.390 101.850 122.560 102.020 ;
        RECT 122.390 101.490 122.560 101.660 ;
        RECT 122.390 101.130 122.560 101.300 ;
        RECT 122.390 100.770 122.560 100.940 ;
        RECT 122.390 100.410 122.560 100.580 ;
        RECT 123.760 101.850 123.930 102.020 ;
        RECT 123.760 101.490 123.930 101.660 ;
        RECT 123.760 101.130 123.930 101.300 ;
        RECT 123.760 100.770 123.930 100.940 ;
        RECT 123.760 100.410 123.930 100.580 ;
        RECT 125.130 101.850 125.300 102.020 ;
        RECT 125.130 101.490 125.300 101.660 ;
        RECT 125.130 101.130 125.300 101.300 ;
        RECT 125.130 100.770 125.300 100.940 ;
        RECT 125.130 100.410 125.300 100.580 ;
        RECT 125.680 101.820 125.850 101.990 ;
        RECT 125.680 101.460 125.850 101.630 ;
        RECT 125.680 101.100 125.850 101.270 ;
        RECT 125.680 100.740 125.850 100.910 ;
        RECT 121.840 100.170 122.010 100.340 ;
        RECT 125.680 100.380 125.850 100.550 ;
        RECT 122.895 99.990 123.065 100.160 ;
        RECT 123.255 99.990 123.425 100.160 ;
        RECT 124.265 99.990 124.435 100.160 ;
        RECT 124.625 99.990 124.795 100.160 ;
        RECT 125.680 100.020 125.850 100.190 ;
        RECT 121.840 99.810 122.010 99.980 ;
        RECT 121.840 99.450 122.010 99.620 ;
        RECT 121.840 99.090 122.010 99.260 ;
        RECT 121.840 98.730 122.010 98.900 ;
        RECT 121.840 98.370 122.010 98.540 ;
        RECT 121.840 98.010 122.010 98.180 ;
        RECT 122.390 99.570 122.560 99.740 ;
        RECT 122.390 99.210 122.560 99.380 ;
        RECT 122.390 98.850 122.560 99.020 ;
        RECT 122.390 98.490 122.560 98.660 ;
        RECT 122.390 98.130 122.560 98.300 ;
        RECT 123.760 99.570 123.930 99.740 ;
        RECT 123.760 99.210 123.930 99.380 ;
        RECT 123.760 98.850 123.930 99.020 ;
        RECT 123.760 98.490 123.930 98.660 ;
        RECT 123.760 98.130 123.930 98.300 ;
        RECT 125.130 99.570 125.300 99.740 ;
        RECT 125.130 99.210 125.300 99.380 ;
        RECT 125.130 98.850 125.300 99.020 ;
        RECT 125.130 98.490 125.300 98.660 ;
        RECT 125.130 98.130 125.300 98.300 ;
        RECT 125.680 99.660 125.850 99.830 ;
        RECT 125.680 99.300 125.850 99.470 ;
        RECT 125.680 98.940 125.850 99.110 ;
        RECT 125.680 98.580 125.850 98.750 ;
        RECT 125.680 98.220 125.850 98.390 ;
        RECT 121.840 97.650 122.010 97.820 ;
        RECT 122.895 97.710 123.065 97.880 ;
        RECT 123.255 97.710 123.425 97.880 ;
        RECT 124.265 97.710 124.435 97.880 ;
        RECT 124.625 97.710 124.795 97.880 ;
        RECT 125.680 97.860 125.850 98.030 ;
        RECT 125.680 97.500 125.850 97.670 ;
        RECT 121.840 97.290 122.010 97.460 ;
        RECT 121.840 96.930 122.010 97.100 ;
        RECT 121.840 96.570 122.010 96.740 ;
        RECT 121.840 96.210 122.010 96.380 ;
        RECT 121.840 95.850 122.010 96.020 ;
        RECT 122.390 97.290 122.560 97.460 ;
        RECT 122.390 96.930 122.560 97.100 ;
        RECT 122.390 96.570 122.560 96.740 ;
        RECT 122.390 96.210 122.560 96.380 ;
        RECT 122.390 95.850 122.560 96.020 ;
        RECT 123.760 97.290 123.930 97.460 ;
        RECT 123.760 96.930 123.930 97.100 ;
        RECT 123.760 96.570 123.930 96.740 ;
        RECT 123.760 96.210 123.930 96.380 ;
        RECT 123.760 95.850 123.930 96.020 ;
        RECT 125.130 97.290 125.300 97.460 ;
        RECT 125.130 96.930 125.300 97.100 ;
        RECT 125.130 96.570 125.300 96.740 ;
        RECT 125.130 96.210 125.300 96.380 ;
        RECT 125.130 95.850 125.300 96.020 ;
        RECT 125.680 97.140 125.850 97.310 ;
        RECT 125.680 96.780 125.850 96.950 ;
        RECT 125.680 96.420 125.850 96.590 ;
        RECT 125.680 96.060 125.850 96.230 ;
        RECT 121.840 95.490 122.010 95.660 ;
        RECT 125.680 95.700 125.850 95.870 ;
        RECT 122.895 95.430 123.065 95.600 ;
        RECT 123.255 95.430 123.425 95.600 ;
        RECT 124.265 95.430 124.435 95.600 ;
        RECT 124.625 95.430 124.795 95.600 ;
        RECT 121.840 95.130 122.010 95.300 ;
        RECT 125.680 95.340 125.850 95.510 ;
        RECT 121.840 94.770 122.010 94.940 ;
        RECT 121.840 94.410 122.010 94.580 ;
        RECT 121.840 94.050 122.010 94.220 ;
        RECT 121.840 93.690 122.010 93.860 ;
        RECT 122.390 95.010 122.560 95.180 ;
        RECT 122.390 94.650 122.560 94.820 ;
        RECT 122.390 94.290 122.560 94.460 ;
        RECT 122.390 93.930 122.560 94.100 ;
        RECT 122.390 93.570 122.560 93.740 ;
        RECT 123.760 95.010 123.930 95.180 ;
        RECT 123.760 94.650 123.930 94.820 ;
        RECT 123.760 94.290 123.930 94.460 ;
        RECT 123.760 93.930 123.930 94.100 ;
        RECT 123.760 93.570 123.930 93.740 ;
        RECT 125.130 95.010 125.300 95.180 ;
        RECT 125.130 94.650 125.300 94.820 ;
        RECT 125.130 94.290 125.300 94.460 ;
        RECT 125.130 93.930 125.300 94.100 ;
        RECT 125.130 93.570 125.300 93.740 ;
        RECT 125.680 94.980 125.850 95.150 ;
        RECT 125.680 94.620 125.850 94.790 ;
        RECT 125.680 94.260 125.850 94.430 ;
        RECT 125.680 93.900 125.850 94.070 ;
        RECT 121.840 93.330 122.010 93.500 ;
        RECT 125.680 93.540 125.850 93.710 ;
        RECT 122.895 93.150 123.065 93.320 ;
        RECT 123.255 93.150 123.425 93.320 ;
        RECT 124.265 93.150 124.435 93.320 ;
        RECT 124.625 93.150 124.795 93.320 ;
        RECT 125.680 93.180 125.850 93.350 ;
        RECT 121.840 92.970 122.010 93.140 ;
        RECT 121.840 92.610 122.010 92.780 ;
        RECT 121.840 92.250 122.010 92.420 ;
        RECT 121.840 91.890 122.010 92.060 ;
        RECT 121.840 91.530 122.010 91.700 ;
        RECT 121.840 91.170 122.010 91.340 ;
        RECT 122.390 92.730 122.560 92.900 ;
        RECT 122.390 92.370 122.560 92.540 ;
        RECT 122.390 92.010 122.560 92.180 ;
        RECT 122.390 91.650 122.560 91.820 ;
        RECT 122.390 91.290 122.560 91.460 ;
        RECT 123.760 92.730 123.930 92.900 ;
        RECT 123.760 92.370 123.930 92.540 ;
        RECT 123.760 92.010 123.930 92.180 ;
        RECT 123.760 91.650 123.930 91.820 ;
        RECT 123.760 91.290 123.930 91.460 ;
        RECT 125.130 92.730 125.300 92.900 ;
        RECT 125.130 92.370 125.300 92.540 ;
        RECT 125.130 92.010 125.300 92.180 ;
        RECT 125.130 91.650 125.300 91.820 ;
        RECT 125.130 91.290 125.300 91.460 ;
        RECT 125.680 92.820 125.850 92.990 ;
        RECT 125.680 92.460 125.850 92.630 ;
        RECT 125.680 92.100 125.850 92.270 ;
        RECT 125.680 91.740 125.850 91.910 ;
        RECT 125.680 91.380 125.850 91.550 ;
        RECT 121.840 90.810 122.010 90.980 ;
        RECT 122.895 90.870 123.065 91.040 ;
        RECT 123.255 90.870 123.425 91.040 ;
        RECT 124.265 90.870 124.435 91.040 ;
        RECT 124.625 90.870 124.795 91.040 ;
        RECT 125.680 91.020 125.850 91.190 ;
        RECT 125.680 90.660 125.850 90.830 ;
        RECT 121.840 90.450 122.010 90.620 ;
        RECT 121.840 90.090 122.010 90.260 ;
        RECT 121.840 89.730 122.010 89.900 ;
        RECT 121.840 89.370 122.010 89.540 ;
        RECT 121.840 89.010 122.010 89.180 ;
        RECT 122.390 90.450 122.560 90.620 ;
        RECT 122.390 90.090 122.560 90.260 ;
        RECT 122.390 89.730 122.560 89.900 ;
        RECT 122.390 89.370 122.560 89.540 ;
        RECT 122.390 89.010 122.560 89.180 ;
        RECT 125.130 90.450 125.300 90.620 ;
        RECT 125.130 90.090 125.300 90.260 ;
        RECT 125.130 89.730 125.300 89.900 ;
        RECT 125.130 89.370 125.300 89.540 ;
        RECT 125.130 89.010 125.300 89.180 ;
        RECT 125.680 90.300 125.850 90.470 ;
        RECT 125.680 89.940 125.850 90.110 ;
        RECT 125.680 89.580 125.850 89.750 ;
        RECT 125.680 89.220 125.850 89.390 ;
        RECT 121.840 88.650 122.010 88.820 ;
        RECT 125.680 88.860 125.850 89.030 ;
        RECT 122.895 88.590 123.065 88.760 ;
        RECT 123.255 88.590 123.425 88.760 ;
        RECT 124.265 88.590 124.435 88.760 ;
        RECT 124.625 88.590 124.795 88.760 ;
        RECT 121.840 88.290 122.010 88.460 ;
        RECT 125.680 88.500 125.850 88.670 ;
        RECT 121.840 87.930 122.010 88.100 ;
        RECT 121.840 87.570 122.010 87.740 ;
        RECT 121.840 87.210 122.010 87.380 ;
        RECT 121.840 86.850 122.010 87.020 ;
        RECT 122.390 88.170 122.560 88.340 ;
        RECT 122.390 87.810 122.560 87.980 ;
        RECT 122.390 87.450 122.560 87.620 ;
        RECT 122.390 87.090 122.560 87.260 ;
        RECT 122.390 86.730 122.560 86.900 ;
        RECT 125.130 88.170 125.300 88.340 ;
        RECT 125.130 87.810 125.300 87.980 ;
        RECT 125.130 87.450 125.300 87.620 ;
        RECT 125.130 87.090 125.300 87.260 ;
        RECT 125.130 86.730 125.300 86.900 ;
        RECT 125.680 88.140 125.850 88.310 ;
        RECT 125.680 87.780 125.850 87.950 ;
        RECT 125.680 87.420 125.850 87.590 ;
        RECT 125.680 87.060 125.850 87.230 ;
        RECT 121.840 86.490 122.010 86.660 ;
        RECT 125.680 86.700 125.850 86.870 ;
        RECT 122.895 86.310 123.065 86.480 ;
        RECT 123.255 86.310 123.425 86.480 ;
        RECT 124.265 86.310 124.435 86.480 ;
        RECT 124.625 86.310 124.795 86.480 ;
        RECT 125.680 86.340 125.850 86.510 ;
        RECT 121.840 86.130 122.010 86.300 ;
        RECT 121.840 85.770 122.010 85.940 ;
        RECT 121.840 85.410 122.010 85.580 ;
        RECT 121.840 85.050 122.010 85.220 ;
        RECT 121.840 84.690 122.010 84.860 ;
        RECT 121.840 84.330 122.010 84.500 ;
        RECT 122.390 85.890 122.560 86.060 ;
        RECT 122.390 85.530 122.560 85.700 ;
        RECT 122.390 85.170 122.560 85.340 ;
        RECT 122.390 84.810 122.560 84.980 ;
        RECT 122.390 84.450 122.560 84.620 ;
        RECT 125.130 85.890 125.300 86.060 ;
        RECT 125.130 85.530 125.300 85.700 ;
        RECT 125.130 85.170 125.300 85.340 ;
        RECT 125.130 84.810 125.300 84.980 ;
        RECT 125.130 84.450 125.300 84.620 ;
        RECT 125.680 85.980 125.850 86.150 ;
        RECT 125.680 85.620 125.850 85.790 ;
        RECT 125.680 85.260 125.850 85.430 ;
        RECT 125.680 84.900 125.850 85.070 ;
        RECT 125.680 84.540 125.850 84.710 ;
        RECT 121.840 83.970 122.010 84.140 ;
        RECT 122.895 84.030 123.065 84.200 ;
        RECT 123.255 84.030 123.425 84.200 ;
        RECT 124.265 84.030 124.435 84.200 ;
        RECT 124.625 84.030 124.795 84.200 ;
        RECT 125.680 84.180 125.850 84.350 ;
        RECT 108.635 83.610 108.805 83.780 ;
        RECT 108.635 83.250 108.805 83.420 ;
        RECT 88.805 82.770 88.975 82.940 ;
        RECT 89.165 82.770 89.335 82.940 ;
        RECT 89.525 82.770 89.695 82.940 ;
        RECT 89.885 82.770 90.055 82.940 ;
        RECT 90.245 82.770 90.415 82.940 ;
        RECT 90.605 82.770 90.775 82.940 ;
        RECT 92.100 82.770 92.270 82.940 ;
        RECT 92.460 82.770 92.630 82.940 ;
        RECT 92.820 82.770 92.990 82.940 ;
        RECT 93.180 82.770 93.350 82.940 ;
        RECT 93.540 82.770 93.710 82.940 ;
        RECT 93.900 82.770 94.070 82.940 ;
        RECT 94.260 82.770 94.430 82.940 ;
        RECT 94.620 82.770 94.790 82.940 ;
        RECT 71.775 82.420 71.945 82.590 ;
        RECT 72.135 82.420 72.305 82.590 ;
        RECT 72.495 82.420 72.665 82.590 ;
        RECT 72.855 82.420 73.025 82.590 ;
        RECT 73.215 82.420 73.385 82.590 ;
        RECT 73.575 82.420 73.745 82.590 ;
        RECT 75.295 82.420 75.465 82.590 ;
        RECT 75.655 82.420 75.825 82.590 ;
        RECT 76.015 82.420 76.185 82.590 ;
        RECT 76.375 82.420 76.545 82.590 ;
        RECT 76.735 82.420 76.905 82.590 ;
        RECT 77.095 82.420 77.265 82.590 ;
        RECT 77.455 82.420 77.625 82.590 ;
        RECT 77.815 82.420 77.985 82.590 ;
        RECT 78.175 82.420 78.345 82.590 ;
        RECT 78.535 82.420 78.705 82.590 ;
        RECT 78.895 82.420 79.065 82.590 ;
        RECT 79.495 82.420 79.665 82.590 ;
        RECT 79.855 82.420 80.025 82.590 ;
        RECT 80.215 82.420 80.385 82.590 ;
        RECT 80.575 82.420 80.745 82.590 ;
        RECT 80.935 82.420 81.105 82.590 ;
        RECT 81.295 82.420 81.465 82.590 ;
        RECT 81.655 82.420 81.825 82.590 ;
        RECT 82.015 82.420 82.185 82.590 ;
        RECT 82.375 82.420 82.545 82.590 ;
        RECT 82.735 82.420 82.905 82.590 ;
        RECT 83.095 82.420 83.265 82.590 ;
        RECT 84.815 82.420 84.985 82.590 ;
        RECT 85.175 82.420 85.345 82.590 ;
        RECT 85.535 82.420 85.705 82.590 ;
        RECT 85.895 82.420 86.065 82.590 ;
        RECT 86.255 82.420 86.425 82.590 ;
        RECT 86.615 82.420 86.785 82.590 ;
        RECT 71.475 82.070 71.645 82.240 ;
        RECT 79.195 82.070 79.365 82.240 ;
        RECT 71.475 81.710 71.645 81.880 ;
        RECT 72.680 81.750 72.850 81.920 ;
        RECT 73.040 81.750 73.210 81.920 ;
        RECT 75.980 81.750 76.150 81.920 ;
        RECT 76.340 81.750 76.510 81.920 ;
        RECT 77.630 81.750 77.800 81.920 ;
        RECT 77.990 81.750 78.160 81.920 ;
        RECT 86.915 82.070 87.085 82.240 ;
        RECT 79.195 81.710 79.365 81.880 ;
        RECT 80.400 81.750 80.570 81.920 ;
        RECT 80.760 81.750 80.930 81.920 ;
        RECT 82.050 81.750 82.220 81.920 ;
        RECT 82.410 81.750 82.580 81.920 ;
        RECT 85.350 81.750 85.520 81.920 ;
        RECT 85.710 81.750 85.880 81.920 ;
        RECT 71.475 81.350 71.645 81.520 ;
        RECT 71.475 80.990 71.645 81.160 ;
        RECT 72.025 81.500 72.195 81.670 ;
        RECT 73.695 81.500 73.865 81.670 ;
        RECT 72.680 81.320 72.850 81.490 ;
        RECT 73.040 81.320 73.210 81.490 ;
        RECT 72.025 81.140 72.195 81.310 ;
        RECT 73.695 81.140 73.865 81.310 ;
        RECT 75.325 81.500 75.495 81.670 ;
        RECT 78.645 81.500 78.815 81.670 ;
        RECT 75.980 81.320 76.150 81.490 ;
        RECT 76.340 81.320 76.510 81.490 ;
        RECT 77.630 81.320 77.800 81.490 ;
        RECT 77.990 81.320 78.160 81.490 ;
        RECT 75.325 81.140 75.495 81.310 ;
        RECT 78.645 81.140 78.815 81.310 ;
        RECT 86.915 81.710 87.085 81.880 ;
        RECT 79.195 81.350 79.365 81.520 ;
        RECT 72.680 80.890 72.850 81.060 ;
        RECT 73.040 80.890 73.210 81.060 ;
        RECT 75.980 80.890 76.150 81.060 ;
        RECT 76.340 80.890 76.510 81.060 ;
        RECT 77.630 80.890 77.800 81.060 ;
        RECT 77.990 80.890 78.160 81.060 ;
        RECT 79.195 80.990 79.365 81.160 ;
        RECT 79.745 81.500 79.915 81.670 ;
        RECT 83.065 81.500 83.235 81.670 ;
        RECT 80.400 81.320 80.570 81.490 ;
        RECT 80.760 81.320 80.930 81.490 ;
        RECT 82.050 81.320 82.220 81.490 ;
        RECT 82.410 81.320 82.580 81.490 ;
        RECT 79.745 81.140 79.915 81.310 ;
        RECT 83.065 81.140 83.235 81.310 ;
        RECT 84.695 81.500 84.865 81.670 ;
        RECT 86.365 81.500 86.535 81.670 ;
        RECT 85.350 81.320 85.520 81.490 ;
        RECT 85.710 81.320 85.880 81.490 ;
        RECT 84.695 81.140 84.865 81.310 ;
        RECT 86.365 81.140 86.535 81.310 ;
        RECT 86.915 81.350 87.085 81.520 ;
        RECT 71.475 80.630 71.645 80.800 ;
        RECT 71.475 80.270 71.645 80.440 ;
        RECT 72.025 80.640 72.195 80.810 ;
        RECT 73.695 80.640 73.865 80.810 ;
        RECT 72.680 80.460 72.850 80.630 ;
        RECT 73.040 80.460 73.210 80.630 ;
        RECT 72.025 80.280 72.195 80.450 ;
        RECT 73.695 80.280 73.865 80.450 ;
        RECT 75.325 80.640 75.495 80.810 ;
        RECT 78.645 80.640 78.815 80.810 ;
        RECT 75.980 80.460 76.150 80.630 ;
        RECT 76.340 80.460 76.510 80.630 ;
        RECT 77.630 80.460 77.800 80.630 ;
        RECT 77.990 80.460 78.160 80.630 ;
        RECT 75.325 80.280 75.495 80.450 ;
        RECT 78.645 80.280 78.815 80.450 ;
        RECT 80.400 80.890 80.570 81.060 ;
        RECT 80.760 80.890 80.930 81.060 ;
        RECT 82.050 80.890 82.220 81.060 ;
        RECT 82.410 80.890 82.580 81.060 ;
        RECT 85.350 80.890 85.520 81.060 ;
        RECT 85.710 80.890 85.880 81.060 ;
        RECT 86.915 80.990 87.085 81.160 ;
        RECT 79.195 80.630 79.365 80.800 ;
        RECT 79.195 80.270 79.365 80.440 ;
        RECT 79.745 80.640 79.915 80.810 ;
        RECT 83.065 80.640 83.235 80.810 ;
        RECT 80.400 80.460 80.570 80.630 ;
        RECT 80.760 80.460 80.930 80.630 ;
        RECT 82.050 80.460 82.220 80.630 ;
        RECT 82.410 80.460 82.580 80.630 ;
        RECT 79.745 80.280 79.915 80.450 ;
        RECT 83.065 80.280 83.235 80.450 ;
        RECT 84.695 80.640 84.865 80.810 ;
        RECT 86.365 80.640 86.535 80.810 ;
        RECT 85.350 80.460 85.520 80.630 ;
        RECT 85.710 80.460 85.880 80.630 ;
        RECT 84.695 80.280 84.865 80.450 ;
        RECT 86.365 80.280 86.535 80.450 ;
        RECT 86.915 80.630 87.085 80.800 ;
        RECT 71.475 79.910 71.645 80.080 ;
        RECT 72.680 80.030 72.850 80.200 ;
        RECT 73.040 80.030 73.210 80.200 ;
        RECT 75.980 80.030 76.150 80.200 ;
        RECT 76.340 80.030 76.510 80.200 ;
        RECT 77.630 80.030 77.800 80.200 ;
        RECT 77.990 80.030 78.160 80.200 ;
        RECT 86.915 80.270 87.085 80.440 ;
        RECT 71.475 79.550 71.645 79.720 ;
        RECT 72.025 79.780 72.195 79.950 ;
        RECT 73.695 79.780 73.865 79.950 ;
        RECT 72.680 79.600 72.850 79.770 ;
        RECT 73.040 79.600 73.210 79.770 ;
        RECT 72.025 79.420 72.195 79.590 ;
        RECT 73.695 79.420 73.865 79.590 ;
        RECT 75.325 79.780 75.495 79.950 ;
        RECT 78.645 79.780 78.815 79.950 ;
        RECT 75.980 79.600 76.150 79.770 ;
        RECT 76.340 79.600 76.510 79.770 ;
        RECT 77.630 79.600 77.800 79.770 ;
        RECT 77.990 79.600 78.160 79.770 ;
        RECT 75.325 79.420 75.495 79.590 ;
        RECT 78.645 79.420 78.815 79.590 ;
        RECT 79.195 79.910 79.365 80.080 ;
        RECT 80.400 80.030 80.570 80.200 ;
        RECT 80.760 80.030 80.930 80.200 ;
        RECT 82.050 80.030 82.220 80.200 ;
        RECT 82.410 80.030 82.580 80.200 ;
        RECT 85.350 80.030 85.520 80.200 ;
        RECT 85.710 80.030 85.880 80.200 ;
        RECT 79.195 79.550 79.365 79.720 ;
        RECT 71.475 79.190 71.645 79.360 ;
        RECT 79.745 79.780 79.915 79.950 ;
        RECT 83.065 79.780 83.235 79.950 ;
        RECT 80.400 79.600 80.570 79.770 ;
        RECT 80.760 79.600 80.930 79.770 ;
        RECT 82.050 79.600 82.220 79.770 ;
        RECT 82.410 79.600 82.580 79.770 ;
        RECT 79.745 79.420 79.915 79.590 ;
        RECT 83.065 79.420 83.235 79.590 ;
        RECT 84.695 79.780 84.865 79.950 ;
        RECT 86.365 79.780 86.535 79.950 ;
        RECT 85.350 79.600 85.520 79.770 ;
        RECT 85.710 79.600 85.880 79.770 ;
        RECT 84.695 79.420 84.865 79.590 ;
        RECT 86.365 79.420 86.535 79.590 ;
        RECT 86.915 79.910 87.085 80.080 ;
        RECT 86.915 79.550 87.085 79.720 ;
        RECT 72.680 79.170 72.850 79.340 ;
        RECT 73.040 79.170 73.210 79.340 ;
        RECT 75.980 79.170 76.150 79.340 ;
        RECT 76.340 79.170 76.510 79.340 ;
        RECT 77.630 79.170 77.800 79.340 ;
        RECT 77.990 79.170 78.160 79.340 ;
        RECT 79.195 79.190 79.365 79.360 ;
        RECT 71.475 78.830 71.645 79.000 ;
        RECT 71.475 78.470 71.645 78.640 ;
        RECT 72.025 78.920 72.195 79.090 ;
        RECT 73.695 78.920 73.865 79.090 ;
        RECT 72.680 78.740 72.850 78.910 ;
        RECT 73.040 78.740 73.210 78.910 ;
        RECT 72.025 78.560 72.195 78.730 ;
        RECT 73.695 78.560 73.865 78.730 ;
        RECT 75.325 78.920 75.495 79.090 ;
        RECT 78.645 78.920 78.815 79.090 ;
        RECT 75.980 78.740 76.150 78.910 ;
        RECT 76.340 78.740 76.510 78.910 ;
        RECT 77.630 78.740 77.800 78.910 ;
        RECT 77.990 78.740 78.160 78.910 ;
        RECT 75.325 78.560 75.495 78.730 ;
        RECT 78.645 78.560 78.815 78.730 ;
        RECT 80.400 79.170 80.570 79.340 ;
        RECT 80.760 79.170 80.930 79.340 ;
        RECT 82.050 79.170 82.220 79.340 ;
        RECT 82.410 79.170 82.580 79.340 ;
        RECT 85.350 79.170 85.520 79.340 ;
        RECT 85.710 79.170 85.880 79.340 ;
        RECT 86.915 79.190 87.085 79.360 ;
        RECT 79.195 78.830 79.365 79.000 ;
        RECT 72.680 78.310 72.850 78.480 ;
        RECT 73.040 78.310 73.210 78.480 ;
        RECT 75.980 78.310 76.150 78.480 ;
        RECT 76.340 78.310 76.510 78.480 ;
        RECT 77.630 78.310 77.800 78.480 ;
        RECT 77.990 78.310 78.160 78.480 ;
        RECT 79.195 78.470 79.365 78.640 ;
        RECT 79.745 78.920 79.915 79.090 ;
        RECT 83.065 78.920 83.235 79.090 ;
        RECT 80.400 78.740 80.570 78.910 ;
        RECT 80.760 78.740 80.930 78.910 ;
        RECT 82.050 78.740 82.220 78.910 ;
        RECT 82.410 78.740 82.580 78.910 ;
        RECT 79.745 78.560 79.915 78.730 ;
        RECT 83.065 78.560 83.235 78.730 ;
        RECT 84.695 78.920 84.865 79.090 ;
        RECT 86.365 78.920 86.535 79.090 ;
        RECT 85.350 78.740 85.520 78.910 ;
        RECT 85.710 78.740 85.880 78.910 ;
        RECT 84.695 78.560 84.865 78.730 ;
        RECT 86.365 78.560 86.535 78.730 ;
        RECT 86.915 78.830 87.085 79.000 ;
        RECT 71.475 78.110 71.645 78.280 ;
        RECT 80.400 78.310 80.570 78.480 ;
        RECT 80.760 78.310 80.930 78.480 ;
        RECT 82.050 78.310 82.220 78.480 ;
        RECT 82.410 78.310 82.580 78.480 ;
        RECT 85.350 78.310 85.520 78.480 ;
        RECT 85.710 78.310 85.880 78.480 ;
        RECT 86.915 78.470 87.085 78.640 ;
        RECT 79.195 78.110 79.365 78.280 ;
        RECT 86.915 78.110 87.085 78.280 ;
        RECT 88.505 82.420 88.675 82.590 ;
        RECT 94.920 82.420 95.090 82.590 ;
        RECT 88.505 82.060 88.675 82.230 ;
        RECT 89.345 82.100 89.515 82.270 ;
        RECT 89.705 82.100 89.875 82.270 ;
        RECT 92.655 82.100 92.825 82.270 ;
        RECT 93.015 82.100 93.185 82.270 ;
        RECT 93.375 82.100 93.545 82.270 ;
        RECT 93.735 82.100 93.905 82.270 ;
        RECT 94.095 82.100 94.265 82.270 ;
        RECT 94.920 82.060 95.090 82.230 ;
        RECT 88.505 81.700 88.675 81.870 ;
        RECT 90.360 81.850 90.530 82.020 ;
        RECT 89.345 81.670 89.515 81.840 ;
        RECT 89.705 81.670 89.875 81.840 ;
        RECT 88.505 81.340 88.675 81.510 ;
        RECT 90.360 81.490 90.530 81.660 ;
        RECT 92.040 81.850 92.210 82.020 ;
        RECT 92.655 81.670 92.825 81.840 ;
        RECT 93.015 81.670 93.185 81.840 ;
        RECT 93.375 81.670 93.545 81.840 ;
        RECT 93.735 81.670 93.905 81.840 ;
        RECT 94.095 81.670 94.265 81.840 ;
        RECT 94.920 81.700 95.090 81.870 ;
        RECT 92.040 81.490 92.210 81.660 ;
        RECT 89.345 81.240 89.515 81.410 ;
        RECT 89.705 81.240 89.875 81.410 ;
        RECT 92.655 81.240 92.825 81.410 ;
        RECT 93.015 81.240 93.185 81.410 ;
        RECT 93.375 81.240 93.545 81.410 ;
        RECT 93.735 81.240 93.905 81.410 ;
        RECT 94.095 81.240 94.265 81.410 ;
        RECT 94.920 81.340 95.090 81.510 ;
        RECT 88.505 80.980 88.675 81.150 ;
        RECT 90.360 80.990 90.530 81.160 ;
        RECT 89.345 80.810 89.515 80.980 ;
        RECT 89.705 80.810 89.875 80.980 ;
        RECT 88.505 80.620 88.675 80.790 ;
        RECT 90.360 80.630 90.530 80.800 ;
        RECT 92.040 80.990 92.210 81.160 ;
        RECT 94.920 80.980 95.090 81.150 ;
        RECT 92.655 80.810 92.825 80.980 ;
        RECT 93.015 80.810 93.185 80.980 ;
        RECT 93.375 80.810 93.545 80.980 ;
        RECT 93.735 80.810 93.905 80.980 ;
        RECT 94.095 80.810 94.265 80.980 ;
        RECT 92.040 80.630 92.210 80.800 ;
        RECT 94.920 80.620 95.090 80.790 ;
        RECT 88.505 80.260 88.675 80.430 ;
        RECT 89.345 80.380 89.515 80.550 ;
        RECT 89.705 80.380 89.875 80.550 ;
        RECT 92.655 80.380 92.825 80.550 ;
        RECT 93.015 80.380 93.185 80.550 ;
        RECT 93.375 80.380 93.545 80.550 ;
        RECT 93.735 80.380 93.905 80.550 ;
        RECT 94.095 80.380 94.265 80.550 ;
        RECT 90.360 80.130 90.530 80.300 ;
        RECT 88.505 79.900 88.675 80.070 ;
        RECT 89.345 79.950 89.515 80.120 ;
        RECT 89.705 79.950 89.875 80.120 ;
        RECT 90.360 79.770 90.530 79.940 ;
        RECT 92.040 80.130 92.210 80.300 ;
        RECT 94.920 80.260 95.090 80.430 ;
        RECT 92.655 79.950 92.825 80.120 ;
        RECT 93.015 79.950 93.185 80.120 ;
        RECT 93.375 79.950 93.545 80.120 ;
        RECT 93.735 79.950 93.905 80.120 ;
        RECT 94.095 79.950 94.265 80.120 ;
        RECT 92.040 79.770 92.210 79.940 ;
        RECT 94.920 79.900 95.090 80.070 ;
        RECT 88.505 79.540 88.675 79.710 ;
        RECT 89.345 79.520 89.515 79.690 ;
        RECT 89.705 79.520 89.875 79.690 ;
        RECT 92.655 79.520 92.825 79.690 ;
        RECT 93.015 79.520 93.185 79.690 ;
        RECT 93.375 79.520 93.545 79.690 ;
        RECT 93.735 79.520 93.905 79.690 ;
        RECT 94.095 79.520 94.265 79.690 ;
        RECT 94.920 79.540 95.090 79.710 ;
        RECT 88.505 79.180 88.675 79.350 ;
        RECT 90.360 79.270 90.530 79.440 ;
        RECT 89.345 79.090 89.515 79.260 ;
        RECT 89.705 79.090 89.875 79.260 ;
        RECT 88.505 78.820 88.675 78.990 ;
        RECT 90.360 78.910 90.530 79.080 ;
        RECT 92.040 79.270 92.210 79.440 ;
        RECT 92.655 79.090 92.825 79.260 ;
        RECT 93.015 79.090 93.185 79.260 ;
        RECT 93.375 79.090 93.545 79.260 ;
        RECT 93.735 79.090 93.905 79.260 ;
        RECT 94.095 79.090 94.265 79.260 ;
        RECT 94.920 79.180 95.090 79.350 ;
        RECT 92.040 78.910 92.210 79.080 ;
        RECT 89.345 78.660 89.515 78.830 ;
        RECT 89.705 78.660 89.875 78.830 ;
        RECT 92.655 78.660 92.825 78.830 ;
        RECT 93.015 78.660 93.185 78.830 ;
        RECT 93.375 78.660 93.545 78.830 ;
        RECT 93.735 78.660 93.905 78.830 ;
        RECT 94.095 78.660 94.265 78.830 ;
        RECT 94.920 78.820 95.090 78.990 ;
        RECT 88.505 78.460 88.675 78.630 ;
        RECT 94.920 78.460 95.090 78.630 ;
        RECT 88.805 77.990 88.975 78.160 ;
        RECT 89.165 77.990 89.335 78.160 ;
        RECT 89.525 77.990 89.695 78.160 ;
        RECT 89.885 77.990 90.055 78.160 ;
        RECT 90.245 77.990 90.415 78.160 ;
        RECT 90.605 77.990 90.775 78.160 ;
        RECT 92.100 77.990 92.270 78.160 ;
        RECT 92.460 77.990 92.630 78.160 ;
        RECT 92.820 77.990 92.990 78.160 ;
        RECT 93.180 77.990 93.350 78.160 ;
        RECT 93.540 77.990 93.710 78.160 ;
        RECT 93.900 77.990 94.070 78.160 ;
        RECT 94.260 77.990 94.430 78.160 ;
        RECT 94.620 77.990 94.790 78.160 ;
        RECT 108.635 82.890 108.805 83.060 ;
        RECT 108.635 82.530 108.805 82.700 ;
        RECT 108.635 82.170 108.805 82.340 ;
        RECT 110.555 83.610 110.725 83.780 ;
        RECT 110.555 83.250 110.725 83.420 ;
        RECT 110.555 82.890 110.725 83.060 ;
        RECT 110.555 82.530 110.725 82.700 ;
        RECT 110.555 82.170 110.725 82.340 ;
        RECT 111.925 83.610 112.095 83.780 ;
        RECT 111.925 83.250 112.095 83.420 ;
        RECT 111.925 82.890 112.095 83.060 ;
        RECT 111.925 82.530 112.095 82.700 ;
        RECT 111.925 82.170 112.095 82.340 ;
        RECT 113.845 83.420 114.015 83.590 ;
        RECT 113.845 83.060 114.015 83.230 ;
        RECT 113.845 82.700 114.015 82.870 ;
        RECT 113.845 82.340 114.015 82.510 ;
        RECT 108.635 81.810 108.805 81.980 ;
        RECT 113.845 81.980 114.015 82.150 ;
        RECT 109.690 81.750 109.860 81.920 ;
        RECT 110.050 81.750 110.220 81.920 ;
        RECT 111.060 81.750 111.230 81.920 ;
        RECT 111.420 81.750 111.590 81.920 ;
        RECT 112.430 81.750 112.600 81.920 ;
        RECT 112.790 81.750 112.960 81.920 ;
        RECT 108.635 81.450 108.805 81.620 ;
        RECT 113.845 81.620 114.015 81.790 ;
        RECT 108.635 81.090 108.805 81.260 ;
        RECT 108.635 80.730 108.805 80.900 ;
        RECT 108.635 80.370 108.805 80.540 ;
        RECT 108.635 80.010 108.805 80.180 ;
        RECT 110.555 81.330 110.725 81.500 ;
        RECT 110.555 80.970 110.725 81.140 ;
        RECT 110.555 80.610 110.725 80.780 ;
        RECT 110.555 80.250 110.725 80.420 ;
        RECT 110.555 79.890 110.725 80.060 ;
        RECT 111.925 81.330 112.095 81.500 ;
        RECT 111.925 80.970 112.095 81.140 ;
        RECT 111.925 80.610 112.095 80.780 ;
        RECT 111.925 80.250 112.095 80.420 ;
        RECT 111.925 79.890 112.095 80.060 ;
        RECT 113.845 81.260 114.015 81.430 ;
        RECT 113.845 80.900 114.015 81.070 ;
        RECT 113.845 80.540 114.015 80.710 ;
        RECT 113.845 80.180 114.015 80.350 ;
        RECT 108.635 79.650 108.805 79.820 ;
        RECT 113.845 79.820 114.015 79.990 ;
        RECT 114.925 83.645 115.095 83.815 ;
        RECT 115.535 83.705 115.705 83.875 ;
        RECT 115.895 83.705 116.065 83.875 ;
        RECT 116.255 83.705 116.425 83.875 ;
        RECT 116.615 83.705 116.785 83.875 ;
        RECT 116.975 83.705 117.145 83.875 ;
        RECT 117.335 83.705 117.505 83.875 ;
        RECT 114.925 83.285 115.095 83.455 ;
        RECT 125.680 83.820 125.850 83.990 ;
        RECT 114.925 82.925 115.095 83.095 ;
        RECT 115.980 83.075 116.150 83.245 ;
        RECT 116.340 83.075 116.510 83.245 ;
        RECT 117.395 83.165 117.565 83.335 ;
        RECT 114.925 82.565 115.095 82.735 ;
        RECT 115.980 82.645 116.150 82.815 ;
        RECT 116.340 82.645 116.510 82.815 ;
        RECT 116.845 82.645 117.015 82.815 ;
        RECT 117.395 82.805 117.565 82.975 ;
        RECT 117.395 82.445 117.565 82.615 ;
        RECT 114.925 82.205 115.095 82.375 ;
        RECT 115.980 82.215 116.150 82.385 ;
        RECT 116.340 82.215 116.510 82.385 ;
        RECT 117.395 82.085 117.565 82.255 ;
        RECT 115.475 81.785 115.645 81.955 ;
        RECT 115.980 81.785 116.150 81.955 ;
        RECT 116.340 81.785 116.510 81.955 ;
        RECT 114.925 81.605 115.095 81.775 ;
        RECT 117.395 81.725 117.565 81.895 ;
        RECT 114.925 81.245 115.095 81.415 ;
        RECT 115.980 81.355 116.150 81.525 ;
        RECT 116.340 81.355 116.510 81.525 ;
        RECT 117.395 81.365 117.565 81.535 ;
        RECT 114.925 80.885 115.095 81.055 ;
        RECT 115.980 80.925 116.150 81.095 ;
        RECT 116.340 80.925 116.510 81.095 ;
        RECT 116.845 80.925 117.015 81.095 ;
        RECT 117.395 81.005 117.565 81.175 ;
        RECT 114.925 80.525 115.095 80.695 ;
        RECT 115.980 80.495 116.150 80.665 ;
        RECT 116.340 80.495 116.510 80.665 ;
        RECT 117.395 80.645 117.565 80.815 ;
        RECT 117.395 80.285 117.565 80.455 ;
        RECT 114.985 79.865 115.155 80.035 ;
        RECT 115.345 79.865 115.515 80.035 ;
        RECT 115.705 79.865 115.875 80.035 ;
        RECT 116.065 79.865 116.235 80.035 ;
        RECT 116.425 79.865 116.595 80.035 ;
        RECT 116.785 79.865 116.955 80.035 ;
        RECT 117.395 79.925 117.565 80.095 ;
        RECT 118.195 83.410 118.365 83.580 ;
        RECT 118.745 83.470 118.915 83.640 ;
        RECT 119.105 83.470 119.275 83.640 ;
        RECT 119.465 83.470 119.635 83.640 ;
        RECT 119.825 83.470 119.995 83.640 ;
        RECT 120.185 83.470 120.355 83.640 ;
        RECT 120.545 83.470 120.715 83.640 ;
        RECT 120.905 83.470 121.075 83.640 ;
        RECT 118.195 83.050 118.365 83.220 ;
        RECT 118.195 82.690 118.365 82.860 ;
        RECT 119.400 82.840 119.570 83.010 ;
        RECT 119.760 82.840 119.930 83.010 ;
        RECT 120.965 82.950 121.135 83.120 ;
        RECT 120.965 82.590 121.135 82.760 ;
        RECT 118.195 82.330 118.365 82.500 ;
        RECT 118.745 82.410 118.915 82.580 ;
        RECT 119.400 82.410 119.570 82.580 ;
        RECT 119.760 82.410 119.930 82.580 ;
        RECT 120.965 82.230 121.135 82.400 ;
        RECT 118.195 81.970 118.365 82.140 ;
        RECT 119.400 81.980 119.570 82.150 ;
        RECT 119.760 81.980 119.930 82.150 ;
        RECT 118.195 81.610 118.365 81.780 ;
        RECT 120.965 81.870 121.135 82.040 ;
        RECT 118.745 81.550 118.915 81.720 ;
        RECT 119.400 81.550 119.570 81.720 ;
        RECT 119.760 81.550 119.930 81.720 ;
        RECT 118.195 81.250 118.365 81.420 ;
        RECT 120.965 81.510 121.135 81.680 ;
        RECT 119.400 81.120 119.570 81.290 ;
        RECT 119.760 81.120 119.930 81.290 ;
        RECT 120.965 81.150 121.135 81.320 ;
        RECT 118.195 80.890 118.365 81.060 ;
        RECT 118.195 80.530 118.365 80.700 ;
        RECT 118.745 80.690 118.915 80.860 ;
        RECT 119.400 80.690 119.570 80.860 ;
        RECT 119.760 80.690 119.930 80.860 ;
        RECT 120.965 80.790 121.135 80.960 ;
        RECT 120.965 80.430 121.135 80.600 ;
        RECT 118.195 80.170 118.365 80.340 ;
        RECT 119.400 80.260 119.570 80.430 ;
        RECT 119.760 80.260 119.930 80.430 ;
        RECT 120.965 80.070 121.135 80.240 ;
        RECT 109.690 79.470 109.860 79.640 ;
        RECT 110.050 79.470 110.220 79.640 ;
        RECT 111.060 79.470 111.230 79.640 ;
        RECT 111.420 79.470 111.590 79.640 ;
        RECT 112.430 79.470 112.600 79.640 ;
        RECT 112.790 79.470 112.960 79.640 ;
        RECT 108.635 79.290 108.805 79.460 ;
        RECT 113.845 79.460 114.015 79.630 ;
        RECT 108.635 78.930 108.805 79.100 ;
        RECT 108.635 78.570 108.805 78.740 ;
        RECT 108.635 78.210 108.805 78.380 ;
        RECT 71.775 77.640 71.945 77.810 ;
        RECT 72.135 77.640 72.305 77.810 ;
        RECT 72.495 77.640 72.665 77.810 ;
        RECT 72.855 77.640 73.025 77.810 ;
        RECT 73.215 77.640 73.385 77.810 ;
        RECT 73.575 77.640 73.745 77.810 ;
        RECT 75.295 77.640 75.465 77.810 ;
        RECT 75.655 77.640 75.825 77.810 ;
        RECT 76.015 77.640 76.185 77.810 ;
        RECT 76.375 77.640 76.545 77.810 ;
        RECT 76.735 77.640 76.905 77.810 ;
        RECT 77.095 77.640 77.265 77.810 ;
        RECT 77.455 77.640 77.625 77.810 ;
        RECT 77.815 77.640 77.985 77.810 ;
        RECT 78.175 77.640 78.345 77.810 ;
        RECT 78.535 77.640 78.705 77.810 ;
        RECT 78.895 77.640 79.065 77.810 ;
        RECT 79.495 77.640 79.665 77.810 ;
        RECT 79.855 77.640 80.025 77.810 ;
        RECT 80.215 77.640 80.385 77.810 ;
        RECT 80.575 77.640 80.745 77.810 ;
        RECT 80.935 77.640 81.105 77.810 ;
        RECT 81.295 77.640 81.465 77.810 ;
        RECT 81.655 77.640 81.825 77.810 ;
        RECT 82.015 77.640 82.185 77.810 ;
        RECT 82.375 77.640 82.545 77.810 ;
        RECT 82.735 77.640 82.905 77.810 ;
        RECT 83.095 77.640 83.265 77.810 ;
        RECT 84.815 77.640 84.985 77.810 ;
        RECT 85.175 77.640 85.345 77.810 ;
        RECT 85.535 77.640 85.705 77.810 ;
        RECT 85.895 77.640 86.065 77.810 ;
        RECT 86.255 77.640 86.425 77.810 ;
        RECT 86.615 77.640 86.785 77.810 ;
        RECT 108.635 77.850 108.805 78.020 ;
        RECT 108.635 77.490 108.805 77.660 ;
        RECT 110.555 79.050 110.725 79.220 ;
        RECT 110.555 78.690 110.725 78.860 ;
        RECT 110.555 78.330 110.725 78.500 ;
        RECT 110.555 77.970 110.725 78.140 ;
        RECT 110.555 77.610 110.725 77.780 ;
        RECT 111.925 79.050 112.095 79.220 ;
        RECT 111.925 78.690 112.095 78.860 ;
        RECT 111.925 78.330 112.095 78.500 ;
        RECT 111.925 77.970 112.095 78.140 ;
        RECT 111.925 77.610 112.095 77.780 ;
        RECT 113.845 79.100 114.015 79.270 ;
        RECT 118.195 79.810 118.365 79.980 ;
        RECT 119.400 79.830 119.570 80.000 ;
        RECT 119.760 79.830 119.930 80.000 ;
        RECT 120.415 79.830 120.585 80.000 ;
        RECT 120.965 79.710 121.135 79.880 ;
        RECT 119.400 79.400 119.570 79.570 ;
        RECT 119.760 79.400 119.930 79.570 ;
        RECT 113.845 78.740 114.015 78.910 ;
        RECT 113.845 78.380 114.015 78.550 ;
        RECT 113.845 78.020 114.015 78.190 ;
        RECT 113.845 77.660 114.015 77.830 ;
        RECT 108.635 77.130 108.805 77.300 ;
        RECT 109.690 77.190 109.860 77.360 ;
        RECT 110.050 77.190 110.220 77.360 ;
        RECT 111.060 77.190 111.230 77.360 ;
        RECT 111.420 77.190 111.590 77.360 ;
        RECT 112.430 77.190 112.600 77.360 ;
        RECT 112.790 77.190 112.960 77.360 ;
        RECT 113.845 77.300 114.015 77.470 ;
        RECT 113.845 76.940 114.015 77.110 ;
        RECT 108.635 76.770 108.805 76.940 ;
        RECT 108.635 76.410 108.805 76.580 ;
        RECT 108.635 76.050 108.805 76.220 ;
        RECT 108.635 75.690 108.805 75.860 ;
        RECT 108.635 75.330 108.805 75.500 ;
        RECT 110.555 76.770 110.725 76.940 ;
        RECT 110.555 76.410 110.725 76.580 ;
        RECT 110.555 76.050 110.725 76.220 ;
        RECT 110.555 75.690 110.725 75.860 ;
        RECT 110.555 75.330 110.725 75.500 ;
        RECT 111.925 76.770 112.095 76.940 ;
        RECT 111.925 76.410 112.095 76.580 ;
        RECT 111.925 76.050 112.095 76.220 ;
        RECT 111.925 75.690 112.095 75.860 ;
        RECT 111.925 75.330 112.095 75.500 ;
        RECT 113.845 76.580 114.015 76.750 ;
        RECT 113.845 76.220 114.015 76.390 ;
        RECT 113.845 75.860 114.015 76.030 ;
        RECT 113.845 75.500 114.015 75.670 ;
        RECT 108.635 74.970 108.805 75.140 ;
        RECT 113.845 75.140 114.015 75.310 ;
        RECT 114.925 79.015 115.095 79.185 ;
        RECT 115.535 79.075 115.705 79.245 ;
        RECT 115.895 79.075 116.065 79.245 ;
        RECT 116.255 79.075 116.425 79.245 ;
        RECT 116.615 79.075 116.785 79.245 ;
        RECT 116.975 79.075 117.145 79.245 ;
        RECT 117.335 79.075 117.505 79.245 ;
        RECT 114.925 78.655 115.095 78.825 ;
        RECT 114.925 78.295 115.095 78.465 ;
        RECT 115.980 78.405 116.150 78.575 ;
        RECT 116.340 78.405 116.510 78.575 ;
        RECT 117.395 78.455 117.565 78.625 ;
        RECT 114.925 77.935 115.095 78.105 ;
        RECT 115.475 77.975 115.645 78.145 ;
        RECT 115.980 77.975 116.150 78.145 ;
        RECT 116.340 77.975 116.510 78.145 ;
        RECT 117.395 78.095 117.565 78.265 ;
        RECT 114.925 77.575 115.095 77.745 ;
        RECT 117.395 77.735 117.565 77.905 ;
        RECT 115.980 77.545 116.150 77.715 ;
        RECT 116.340 77.545 116.510 77.715 ;
        RECT 117.395 77.375 117.565 77.545 ;
        RECT 115.980 77.115 116.150 77.285 ;
        RECT 116.340 77.115 116.510 77.285 ;
        RECT 116.845 77.115 117.015 77.285 ;
        RECT 114.925 76.935 115.095 77.105 ;
        RECT 117.395 77.015 117.565 77.185 ;
        RECT 114.925 76.575 115.095 76.745 ;
        RECT 115.980 76.685 116.150 76.855 ;
        RECT 116.340 76.685 116.510 76.855 ;
        RECT 117.395 76.655 117.565 76.825 ;
        RECT 114.925 76.215 115.095 76.385 ;
        RECT 115.475 76.255 115.645 76.425 ;
        RECT 115.980 76.255 116.150 76.425 ;
        RECT 116.340 76.255 116.510 76.425 ;
        RECT 117.395 76.295 117.565 76.465 ;
        RECT 114.925 75.855 115.095 76.025 ;
        RECT 115.980 75.825 116.150 75.995 ;
        RECT 116.340 75.825 116.510 75.995 ;
        RECT 117.395 75.935 117.565 76.105 ;
        RECT 117.395 75.575 117.565 75.745 ;
        RECT 114.985 75.155 115.155 75.325 ;
        RECT 115.345 75.155 115.515 75.325 ;
        RECT 115.705 75.155 115.875 75.325 ;
        RECT 116.065 75.155 116.235 75.325 ;
        RECT 116.425 75.155 116.595 75.325 ;
        RECT 116.785 75.155 116.955 75.325 ;
        RECT 117.395 75.215 117.565 75.385 ;
        RECT 118.195 79.220 118.365 79.390 ;
        RECT 120.965 79.350 121.135 79.520 ;
        RECT 118.195 78.860 118.365 79.030 ;
        RECT 119.400 78.970 119.570 79.140 ;
        RECT 119.760 78.970 119.930 79.140 ;
        RECT 120.415 78.970 120.585 79.140 ;
        RECT 120.965 78.990 121.135 79.160 ;
        RECT 118.195 78.500 118.365 78.670 ;
        RECT 119.400 78.540 119.570 78.710 ;
        RECT 119.760 78.540 119.930 78.710 ;
        RECT 120.965 78.630 121.135 78.800 ;
        RECT 118.195 78.140 118.365 78.310 ;
        RECT 118.745 78.110 118.915 78.280 ;
        RECT 119.400 78.110 119.570 78.280 ;
        RECT 119.760 78.110 119.930 78.280 ;
        RECT 120.965 78.270 121.135 78.440 ;
        RECT 118.195 77.780 118.365 77.950 ;
        RECT 120.965 77.910 121.135 78.080 ;
        RECT 119.400 77.680 119.570 77.850 ;
        RECT 119.760 77.680 119.930 77.850 ;
        RECT 118.195 77.420 118.365 77.590 ;
        RECT 120.965 77.550 121.135 77.720 ;
        RECT 118.745 77.250 118.915 77.420 ;
        RECT 119.400 77.250 119.570 77.420 ;
        RECT 119.760 77.250 119.930 77.420 ;
        RECT 118.195 77.060 118.365 77.230 ;
        RECT 120.965 77.190 121.135 77.360 ;
        RECT 118.195 76.700 118.365 76.870 ;
        RECT 119.400 76.820 119.570 76.990 ;
        RECT 119.760 76.820 119.930 76.990 ;
        RECT 120.965 76.830 121.135 77.000 ;
        RECT 118.195 76.340 118.365 76.510 ;
        RECT 118.745 76.390 118.915 76.560 ;
        RECT 119.400 76.390 119.570 76.560 ;
        RECT 119.760 76.390 119.930 76.560 ;
        RECT 120.965 76.470 121.135 76.640 ;
        RECT 121.840 83.610 122.010 83.780 ;
        RECT 121.840 83.250 122.010 83.420 ;
        RECT 121.840 82.890 122.010 83.060 ;
        RECT 121.840 82.530 122.010 82.700 ;
        RECT 121.840 82.170 122.010 82.340 ;
        RECT 122.390 83.610 122.560 83.780 ;
        RECT 122.390 83.250 122.560 83.420 ;
        RECT 122.390 82.890 122.560 83.060 ;
        RECT 122.390 82.530 122.560 82.700 ;
        RECT 122.390 82.170 122.560 82.340 ;
        RECT 125.130 83.610 125.300 83.780 ;
        RECT 125.130 83.250 125.300 83.420 ;
        RECT 125.130 82.890 125.300 83.060 ;
        RECT 125.130 82.530 125.300 82.700 ;
        RECT 125.130 82.170 125.300 82.340 ;
        RECT 125.680 83.460 125.850 83.630 ;
        RECT 125.680 83.100 125.850 83.270 ;
        RECT 125.680 82.740 125.850 82.910 ;
        RECT 125.680 82.380 125.850 82.550 ;
        RECT 121.840 81.810 122.010 81.980 ;
        RECT 125.680 82.020 125.850 82.190 ;
        RECT 122.895 81.750 123.065 81.920 ;
        RECT 123.255 81.750 123.425 81.920 ;
        RECT 124.265 81.750 124.435 81.920 ;
        RECT 124.625 81.750 124.795 81.920 ;
        RECT 121.840 81.450 122.010 81.620 ;
        RECT 125.680 81.660 125.850 81.830 ;
        RECT 121.840 81.090 122.010 81.260 ;
        RECT 121.840 80.730 122.010 80.900 ;
        RECT 121.840 80.370 122.010 80.540 ;
        RECT 121.840 80.010 122.010 80.180 ;
        RECT 122.390 81.330 122.560 81.500 ;
        RECT 122.390 80.970 122.560 81.140 ;
        RECT 122.390 80.610 122.560 80.780 ;
        RECT 122.390 80.250 122.560 80.420 ;
        RECT 122.390 79.890 122.560 80.060 ;
        RECT 125.130 81.330 125.300 81.500 ;
        RECT 125.130 80.970 125.300 81.140 ;
        RECT 125.130 80.610 125.300 80.780 ;
        RECT 125.130 80.250 125.300 80.420 ;
        RECT 125.130 79.890 125.300 80.060 ;
        RECT 125.680 81.300 125.850 81.470 ;
        RECT 125.680 80.940 125.850 81.110 ;
        RECT 125.680 80.580 125.850 80.750 ;
        RECT 125.680 80.220 125.850 80.390 ;
        RECT 121.840 79.650 122.010 79.820 ;
        RECT 125.680 79.860 125.850 80.030 ;
        RECT 122.895 79.470 123.065 79.640 ;
        RECT 123.255 79.470 123.425 79.640 ;
        RECT 124.265 79.470 124.435 79.640 ;
        RECT 124.625 79.470 124.795 79.640 ;
        RECT 125.680 79.500 125.850 79.670 ;
        RECT 121.840 79.290 122.010 79.460 ;
        RECT 121.840 78.930 122.010 79.100 ;
        RECT 121.840 78.570 122.010 78.740 ;
        RECT 121.840 78.210 122.010 78.380 ;
        RECT 121.840 77.850 122.010 78.020 ;
        RECT 121.840 77.490 122.010 77.660 ;
        RECT 122.390 79.050 122.560 79.220 ;
        RECT 122.390 78.690 122.560 78.860 ;
        RECT 122.390 78.330 122.560 78.500 ;
        RECT 122.390 77.970 122.560 78.140 ;
        RECT 122.390 77.610 122.560 77.780 ;
        RECT 123.760 79.050 123.930 79.220 ;
        RECT 123.760 78.690 123.930 78.860 ;
        RECT 123.760 78.330 123.930 78.500 ;
        RECT 123.760 77.970 123.930 78.140 ;
        RECT 123.760 77.610 123.930 77.780 ;
        RECT 125.130 79.050 125.300 79.220 ;
        RECT 125.130 78.690 125.300 78.860 ;
        RECT 125.130 78.330 125.300 78.500 ;
        RECT 125.130 77.970 125.300 78.140 ;
        RECT 125.130 77.610 125.300 77.780 ;
        RECT 125.680 79.140 125.850 79.310 ;
        RECT 125.680 78.780 125.850 78.950 ;
        RECT 125.680 78.420 125.850 78.590 ;
        RECT 125.680 78.060 125.850 78.230 ;
        RECT 125.680 77.700 125.850 77.870 ;
        RECT 121.840 77.130 122.010 77.300 ;
        RECT 122.895 77.190 123.065 77.360 ;
        RECT 123.255 77.190 123.425 77.360 ;
        RECT 124.265 77.190 124.435 77.360 ;
        RECT 124.625 77.190 124.795 77.360 ;
        RECT 125.680 77.340 125.850 77.510 ;
        RECT 125.680 76.980 125.850 77.150 ;
        RECT 121.900 76.560 122.070 76.730 ;
        RECT 122.260 76.560 122.430 76.730 ;
        RECT 122.620 76.560 122.790 76.730 ;
        RECT 122.980 76.560 123.150 76.730 ;
        RECT 123.340 76.560 123.510 76.730 ;
        RECT 123.700 76.560 123.870 76.730 ;
        RECT 124.060 76.560 124.230 76.730 ;
        RECT 124.420 76.560 124.590 76.730 ;
        RECT 124.780 76.560 124.950 76.730 ;
        RECT 125.140 76.560 125.310 76.730 ;
        RECT 125.680 76.620 125.850 76.790 ;
        RECT 118.195 75.980 118.365 76.150 ;
        RECT 119.400 75.960 119.570 76.130 ;
        RECT 119.760 75.960 119.930 76.130 ;
        RECT 120.965 76.110 121.135 76.280 ;
        RECT 120.965 75.750 121.135 75.920 ;
        RECT 118.255 75.330 118.425 75.500 ;
        RECT 118.615 75.330 118.785 75.500 ;
        RECT 118.975 75.330 119.145 75.500 ;
        RECT 119.335 75.330 119.505 75.500 ;
        RECT 119.695 75.330 119.865 75.500 ;
        RECT 120.055 75.330 120.225 75.500 ;
        RECT 120.415 75.330 120.585 75.500 ;
        RECT 120.965 75.390 121.135 75.560 ;
        RECT 109.690 74.910 109.860 75.080 ;
        RECT 110.050 74.910 110.220 75.080 ;
        RECT 111.060 74.910 111.230 75.080 ;
        RECT 111.420 74.910 111.590 75.080 ;
        RECT 112.430 74.910 112.600 75.080 ;
        RECT 112.790 74.910 112.960 75.080 ;
        RECT 108.635 74.610 108.805 74.780 ;
        RECT 113.845 74.780 114.015 74.950 ;
        RECT 108.635 74.250 108.805 74.420 ;
        RECT 108.635 73.890 108.805 74.060 ;
        RECT 108.635 73.530 108.805 73.700 ;
        RECT 108.635 73.170 108.805 73.340 ;
        RECT 110.555 74.490 110.725 74.660 ;
        RECT 110.555 74.130 110.725 74.300 ;
        RECT 110.555 73.770 110.725 73.940 ;
        RECT 110.555 73.410 110.725 73.580 ;
        RECT 110.555 73.050 110.725 73.220 ;
        RECT 111.925 74.490 112.095 74.660 ;
        RECT 111.925 74.130 112.095 74.300 ;
        RECT 111.925 73.770 112.095 73.940 ;
        RECT 111.925 73.410 112.095 73.580 ;
        RECT 111.925 73.050 112.095 73.220 ;
        RECT 113.845 74.420 114.015 74.590 ;
        RECT 113.845 74.060 114.015 74.230 ;
        RECT 113.845 73.700 114.015 73.870 ;
        RECT 113.845 73.340 114.015 73.510 ;
        RECT 108.635 72.810 108.805 72.980 ;
        RECT 113.845 72.980 114.015 73.150 ;
        RECT 109.690 72.630 109.860 72.800 ;
        RECT 110.050 72.630 110.220 72.800 ;
        RECT 111.060 72.630 111.230 72.800 ;
        RECT 111.420 72.630 111.590 72.800 ;
        RECT 112.430 72.630 112.600 72.800 ;
        RECT 112.790 72.630 112.960 72.800 ;
        RECT 108.635 72.450 108.805 72.620 ;
        RECT 65.025 72.110 65.195 72.280 ;
        RECT 65.385 72.110 65.555 72.280 ;
        RECT 65.745 72.110 65.915 72.280 ;
        RECT 66.105 72.110 66.275 72.280 ;
        RECT 66.465 72.110 66.635 72.280 ;
        RECT 66.825 72.110 66.995 72.280 ;
        RECT 68.320 72.110 68.490 72.280 ;
        RECT 68.680 72.110 68.850 72.280 ;
        RECT 69.040 72.110 69.210 72.280 ;
        RECT 69.400 72.110 69.570 72.280 ;
        RECT 69.760 72.110 69.930 72.280 ;
        RECT 70.120 72.110 70.290 72.280 ;
        RECT 70.480 72.110 70.650 72.280 ;
        RECT 70.840 72.110 71.010 72.280 ;
        RECT 64.725 71.760 64.895 71.930 ;
        RECT 71.140 71.760 71.310 71.930 ;
        RECT 64.725 71.400 64.895 71.570 ;
        RECT 65.565 71.440 65.735 71.610 ;
        RECT 65.925 71.440 66.095 71.610 ;
        RECT 68.875 71.440 69.045 71.610 ;
        RECT 69.235 71.440 69.405 71.610 ;
        RECT 69.595 71.440 69.765 71.610 ;
        RECT 69.955 71.440 70.125 71.610 ;
        RECT 70.315 71.440 70.485 71.610 ;
        RECT 71.140 71.400 71.310 71.570 ;
        RECT 64.725 71.040 64.895 71.210 ;
        RECT 66.580 71.190 66.750 71.360 ;
        RECT 65.565 71.010 65.735 71.180 ;
        RECT 65.925 71.010 66.095 71.180 ;
        RECT 64.725 70.680 64.895 70.850 ;
        RECT 66.580 70.830 66.750 71.000 ;
        RECT 68.260 71.190 68.430 71.360 ;
        RECT 68.875 71.010 69.045 71.180 ;
        RECT 69.235 71.010 69.405 71.180 ;
        RECT 69.595 71.010 69.765 71.180 ;
        RECT 69.955 71.010 70.125 71.180 ;
        RECT 70.315 71.010 70.485 71.180 ;
        RECT 71.140 71.040 71.310 71.210 ;
        RECT 68.260 70.830 68.430 71.000 ;
        RECT 65.565 70.580 65.735 70.750 ;
        RECT 65.925 70.580 66.095 70.750 ;
        RECT 68.875 70.580 69.045 70.750 ;
        RECT 69.235 70.580 69.405 70.750 ;
        RECT 69.595 70.580 69.765 70.750 ;
        RECT 69.955 70.580 70.125 70.750 ;
        RECT 70.315 70.580 70.485 70.750 ;
        RECT 71.140 70.680 71.310 70.850 ;
        RECT 64.725 70.320 64.895 70.490 ;
        RECT 66.580 70.330 66.750 70.500 ;
        RECT 65.565 70.150 65.735 70.320 ;
        RECT 65.925 70.150 66.095 70.320 ;
        RECT 64.725 69.960 64.895 70.130 ;
        RECT 66.580 69.970 66.750 70.140 ;
        RECT 68.260 70.330 68.430 70.500 ;
        RECT 71.140 70.320 71.310 70.490 ;
        RECT 68.875 70.150 69.045 70.320 ;
        RECT 69.235 70.150 69.405 70.320 ;
        RECT 69.595 70.150 69.765 70.320 ;
        RECT 69.955 70.150 70.125 70.320 ;
        RECT 70.315 70.150 70.485 70.320 ;
        RECT 68.260 69.970 68.430 70.140 ;
        RECT 71.140 69.960 71.310 70.130 ;
        RECT 64.725 69.600 64.895 69.770 ;
        RECT 65.565 69.720 65.735 69.890 ;
        RECT 65.925 69.720 66.095 69.890 ;
        RECT 68.875 69.720 69.045 69.890 ;
        RECT 69.235 69.720 69.405 69.890 ;
        RECT 69.595 69.720 69.765 69.890 ;
        RECT 69.955 69.720 70.125 69.890 ;
        RECT 70.315 69.720 70.485 69.890 ;
        RECT 66.580 69.470 66.750 69.640 ;
        RECT 64.725 69.240 64.895 69.410 ;
        RECT 65.565 69.290 65.735 69.460 ;
        RECT 65.925 69.290 66.095 69.460 ;
        RECT 66.580 69.110 66.750 69.280 ;
        RECT 68.260 69.470 68.430 69.640 ;
        RECT 71.140 69.600 71.310 69.770 ;
        RECT 68.875 69.290 69.045 69.460 ;
        RECT 69.235 69.290 69.405 69.460 ;
        RECT 69.595 69.290 69.765 69.460 ;
        RECT 69.955 69.290 70.125 69.460 ;
        RECT 70.315 69.290 70.485 69.460 ;
        RECT 68.260 69.110 68.430 69.280 ;
        RECT 71.140 69.240 71.310 69.410 ;
        RECT 64.725 68.880 64.895 69.050 ;
        RECT 65.565 68.860 65.735 69.030 ;
        RECT 65.925 68.860 66.095 69.030 ;
        RECT 68.875 68.860 69.045 69.030 ;
        RECT 69.235 68.860 69.405 69.030 ;
        RECT 69.595 68.860 69.765 69.030 ;
        RECT 69.955 68.860 70.125 69.030 ;
        RECT 70.315 68.860 70.485 69.030 ;
        RECT 71.140 68.880 71.310 69.050 ;
        RECT 64.725 68.520 64.895 68.690 ;
        RECT 66.580 68.610 66.750 68.780 ;
        RECT 65.565 68.430 65.735 68.600 ;
        RECT 65.925 68.430 66.095 68.600 ;
        RECT 64.725 68.160 64.895 68.330 ;
        RECT 66.580 68.250 66.750 68.420 ;
        RECT 68.260 68.610 68.430 68.780 ;
        RECT 68.875 68.430 69.045 68.600 ;
        RECT 69.235 68.430 69.405 68.600 ;
        RECT 69.595 68.430 69.765 68.600 ;
        RECT 69.955 68.430 70.125 68.600 ;
        RECT 70.315 68.430 70.485 68.600 ;
        RECT 71.140 68.520 71.310 68.690 ;
        RECT 68.260 68.250 68.430 68.420 ;
        RECT 65.565 68.000 65.735 68.170 ;
        RECT 65.925 68.000 66.095 68.170 ;
        RECT 68.875 68.000 69.045 68.170 ;
        RECT 69.235 68.000 69.405 68.170 ;
        RECT 69.595 68.000 69.765 68.170 ;
        RECT 69.955 68.000 70.125 68.170 ;
        RECT 70.315 68.000 70.485 68.170 ;
        RECT 71.140 68.160 71.310 68.330 ;
        RECT 64.725 67.800 64.895 67.970 ;
        RECT 66.580 67.750 66.750 67.920 ;
        RECT 64.725 67.440 64.895 67.610 ;
        RECT 65.565 67.570 65.735 67.740 ;
        RECT 65.925 67.570 66.095 67.740 ;
        RECT 66.580 67.390 66.750 67.560 ;
        RECT 68.260 67.750 68.430 67.920 ;
        RECT 71.140 67.800 71.310 67.970 ;
        RECT 68.875 67.570 69.045 67.740 ;
        RECT 69.235 67.570 69.405 67.740 ;
        RECT 69.595 67.570 69.765 67.740 ;
        RECT 69.955 67.570 70.125 67.740 ;
        RECT 70.315 67.570 70.485 67.740 ;
        RECT 68.260 67.390 68.430 67.560 ;
        RECT 71.140 67.440 71.310 67.610 ;
        RECT 64.725 67.080 64.895 67.250 ;
        RECT 65.565 67.140 65.735 67.310 ;
        RECT 65.925 67.140 66.095 67.310 ;
        RECT 68.875 67.140 69.045 67.310 ;
        RECT 69.235 67.140 69.405 67.310 ;
        RECT 69.595 67.140 69.765 67.310 ;
        RECT 69.955 67.140 70.125 67.310 ;
        RECT 70.315 67.140 70.485 67.310 ;
        RECT 71.140 67.080 71.310 67.250 ;
        RECT 64.725 66.720 64.895 66.890 ;
        RECT 66.580 66.890 66.750 67.060 ;
        RECT 65.565 66.710 65.735 66.880 ;
        RECT 65.925 66.710 66.095 66.880 ;
        RECT 66.580 66.530 66.750 66.700 ;
        RECT 68.260 66.890 68.430 67.060 ;
        RECT 68.875 66.710 69.045 66.880 ;
        RECT 69.235 66.710 69.405 66.880 ;
        RECT 69.595 66.710 69.765 66.880 ;
        RECT 69.955 66.710 70.125 66.880 ;
        RECT 70.315 66.710 70.485 66.880 ;
        RECT 71.140 66.720 71.310 66.890 ;
        RECT 68.260 66.530 68.430 66.700 ;
        RECT 64.725 66.360 64.895 66.530 ;
        RECT 65.565 66.280 65.735 66.450 ;
        RECT 65.925 66.280 66.095 66.450 ;
        RECT 68.875 66.280 69.045 66.450 ;
        RECT 69.235 66.280 69.405 66.450 ;
        RECT 69.595 66.280 69.765 66.450 ;
        RECT 69.955 66.280 70.125 66.450 ;
        RECT 70.315 66.280 70.485 66.450 ;
        RECT 71.140 66.360 71.310 66.530 ;
        RECT 64.725 66.000 64.895 66.170 ;
        RECT 66.580 66.030 66.750 66.200 ;
        RECT 65.565 65.850 65.735 66.020 ;
        RECT 65.925 65.850 66.095 66.020 ;
        RECT 64.725 65.640 64.895 65.810 ;
        RECT 66.580 65.670 66.750 65.840 ;
        RECT 68.260 66.030 68.430 66.200 ;
        RECT 68.875 65.850 69.045 66.020 ;
        RECT 69.235 65.850 69.405 66.020 ;
        RECT 69.595 65.850 69.765 66.020 ;
        RECT 69.955 65.850 70.125 66.020 ;
        RECT 70.315 65.850 70.485 66.020 ;
        RECT 71.140 66.000 71.310 66.170 ;
        RECT 68.260 65.670 68.430 65.840 ;
        RECT 71.140 65.640 71.310 65.810 ;
        RECT 64.725 65.280 64.895 65.450 ;
        RECT 65.565 65.420 65.735 65.590 ;
        RECT 65.925 65.420 66.095 65.590 ;
        RECT 68.875 65.420 69.045 65.590 ;
        RECT 69.235 65.420 69.405 65.590 ;
        RECT 69.595 65.420 69.765 65.590 ;
        RECT 69.955 65.420 70.125 65.590 ;
        RECT 70.315 65.420 70.485 65.590 ;
        RECT 66.580 65.170 66.750 65.340 ;
        RECT 64.725 64.920 64.895 65.090 ;
        RECT 65.565 64.990 65.735 65.160 ;
        RECT 65.925 64.990 66.095 65.160 ;
        RECT 66.580 64.810 66.750 64.980 ;
        RECT 68.260 65.170 68.430 65.340 ;
        RECT 71.140 65.280 71.310 65.450 ;
        RECT 68.875 64.990 69.045 65.160 ;
        RECT 69.235 64.990 69.405 65.160 ;
        RECT 69.595 64.990 69.765 65.160 ;
        RECT 69.955 64.990 70.125 65.160 ;
        RECT 70.315 64.990 70.485 65.160 ;
        RECT 68.260 64.810 68.430 64.980 ;
        RECT 71.140 64.920 71.310 65.090 ;
        RECT 64.725 64.560 64.895 64.730 ;
        RECT 65.565 64.560 65.735 64.730 ;
        RECT 65.925 64.560 66.095 64.730 ;
        RECT 68.875 64.560 69.045 64.730 ;
        RECT 69.235 64.560 69.405 64.730 ;
        RECT 69.595 64.560 69.765 64.730 ;
        RECT 69.955 64.560 70.125 64.730 ;
        RECT 70.315 64.560 70.485 64.730 ;
        RECT 71.140 64.560 71.310 64.730 ;
        RECT 64.725 64.200 64.895 64.370 ;
        RECT 66.580 64.310 66.750 64.480 ;
        RECT 65.565 64.130 65.735 64.300 ;
        RECT 65.925 64.130 66.095 64.300 ;
        RECT 64.725 63.840 64.895 64.010 ;
        RECT 66.580 63.950 66.750 64.120 ;
        RECT 68.260 64.310 68.430 64.480 ;
        RECT 68.875 64.130 69.045 64.300 ;
        RECT 69.235 64.130 69.405 64.300 ;
        RECT 69.595 64.130 69.765 64.300 ;
        RECT 69.955 64.130 70.125 64.300 ;
        RECT 70.315 64.130 70.485 64.300 ;
        RECT 71.140 64.200 71.310 64.370 ;
        RECT 68.260 63.950 68.430 64.120 ;
        RECT 65.565 63.700 65.735 63.870 ;
        RECT 65.925 63.700 66.095 63.870 ;
        RECT 68.875 63.700 69.045 63.870 ;
        RECT 69.235 63.700 69.405 63.870 ;
        RECT 69.595 63.700 69.765 63.870 ;
        RECT 69.955 63.700 70.125 63.870 ;
        RECT 70.315 63.700 70.485 63.870 ;
        RECT 71.140 63.840 71.310 64.010 ;
        RECT 64.725 63.480 64.895 63.650 ;
        RECT 71.140 63.480 71.310 63.650 ;
        RECT 65.025 63.030 65.195 63.200 ;
        RECT 65.385 63.030 65.555 63.200 ;
        RECT 65.745 63.030 65.915 63.200 ;
        RECT 66.105 63.030 66.275 63.200 ;
        RECT 66.465 63.030 66.635 63.200 ;
        RECT 66.825 63.030 66.995 63.200 ;
        RECT 68.320 63.030 68.490 63.200 ;
        RECT 68.680 63.030 68.850 63.200 ;
        RECT 69.040 63.030 69.210 63.200 ;
        RECT 69.400 63.030 69.570 63.200 ;
        RECT 69.760 63.030 69.930 63.200 ;
        RECT 70.120 63.030 70.290 63.200 ;
        RECT 70.480 63.030 70.650 63.200 ;
        RECT 70.840 63.030 71.010 63.200 ;
        RECT 74.045 72.110 74.215 72.280 ;
        RECT 74.405 72.110 74.575 72.280 ;
        RECT 74.765 72.110 74.935 72.280 ;
        RECT 75.125 72.110 75.295 72.280 ;
        RECT 75.485 72.110 75.655 72.280 ;
        RECT 75.845 72.110 76.015 72.280 ;
        RECT 77.340 72.110 77.510 72.280 ;
        RECT 77.700 72.110 77.870 72.280 ;
        RECT 78.060 72.110 78.230 72.280 ;
        RECT 78.420 72.110 78.590 72.280 ;
        RECT 78.780 72.110 78.950 72.280 ;
        RECT 79.140 72.110 79.310 72.280 ;
        RECT 79.500 72.110 79.670 72.280 ;
        RECT 79.860 72.110 80.030 72.280 ;
        RECT 80.460 72.110 80.630 72.280 ;
        RECT 80.820 72.110 80.990 72.280 ;
        RECT 81.180 72.110 81.350 72.280 ;
        RECT 81.540 72.110 81.710 72.280 ;
        RECT 81.900 72.110 82.070 72.280 ;
        RECT 82.260 72.110 82.430 72.280 ;
        RECT 82.620 72.110 82.790 72.280 ;
        RECT 82.980 72.110 83.150 72.280 ;
        RECT 84.475 72.110 84.645 72.280 ;
        RECT 84.835 72.110 85.005 72.280 ;
        RECT 85.195 72.110 85.365 72.280 ;
        RECT 85.555 72.110 85.725 72.280 ;
        RECT 85.915 72.110 86.085 72.280 ;
        RECT 86.275 72.110 86.445 72.280 ;
        RECT 73.745 71.760 73.915 71.930 ;
        RECT 80.160 71.760 80.330 71.930 ;
        RECT 73.745 71.400 73.915 71.570 ;
        RECT 74.585 71.440 74.755 71.610 ;
        RECT 74.945 71.440 75.115 71.610 ;
        RECT 77.895 71.440 78.065 71.610 ;
        RECT 78.255 71.440 78.425 71.610 ;
        RECT 78.615 71.440 78.785 71.610 ;
        RECT 78.975 71.440 79.145 71.610 ;
        RECT 79.335 71.440 79.505 71.610 ;
        RECT 86.575 71.760 86.745 71.930 ;
        RECT 80.160 71.400 80.330 71.570 ;
        RECT 80.985 71.440 81.155 71.610 ;
        RECT 81.345 71.440 81.515 71.610 ;
        RECT 81.705 71.440 81.875 71.610 ;
        RECT 82.065 71.440 82.235 71.610 ;
        RECT 82.425 71.440 82.595 71.610 ;
        RECT 85.375 71.440 85.545 71.610 ;
        RECT 85.735 71.440 85.905 71.610 ;
        RECT 73.745 71.040 73.915 71.210 ;
        RECT 75.600 71.190 75.770 71.360 ;
        RECT 74.585 71.010 74.755 71.180 ;
        RECT 74.945 71.010 75.115 71.180 ;
        RECT 73.745 70.680 73.915 70.850 ;
        RECT 75.600 70.830 75.770 71.000 ;
        RECT 77.280 71.190 77.450 71.360 ;
        RECT 86.575 71.400 86.745 71.570 ;
        RECT 77.895 71.010 78.065 71.180 ;
        RECT 78.255 71.010 78.425 71.180 ;
        RECT 78.615 71.010 78.785 71.180 ;
        RECT 78.975 71.010 79.145 71.180 ;
        RECT 79.335 71.010 79.505 71.180 ;
        RECT 80.160 71.040 80.330 71.210 ;
        RECT 83.040 71.190 83.210 71.360 ;
        RECT 77.280 70.830 77.450 71.000 ;
        RECT 80.985 71.010 81.155 71.180 ;
        RECT 81.345 71.010 81.515 71.180 ;
        RECT 81.705 71.010 81.875 71.180 ;
        RECT 82.065 71.010 82.235 71.180 ;
        RECT 82.425 71.010 82.595 71.180 ;
        RECT 74.585 70.580 74.755 70.750 ;
        RECT 74.945 70.580 75.115 70.750 ;
        RECT 77.895 70.580 78.065 70.750 ;
        RECT 78.255 70.580 78.425 70.750 ;
        RECT 78.615 70.580 78.785 70.750 ;
        RECT 78.975 70.580 79.145 70.750 ;
        RECT 79.335 70.580 79.505 70.750 ;
        RECT 80.160 70.680 80.330 70.850 ;
        RECT 83.040 70.830 83.210 71.000 ;
        RECT 84.720 71.190 84.890 71.360 ;
        RECT 85.375 71.010 85.545 71.180 ;
        RECT 85.735 71.010 85.905 71.180 ;
        RECT 86.575 71.040 86.745 71.210 ;
        RECT 84.720 70.830 84.890 71.000 ;
        RECT 73.745 70.320 73.915 70.490 ;
        RECT 75.600 70.330 75.770 70.500 ;
        RECT 74.585 70.150 74.755 70.320 ;
        RECT 74.945 70.150 75.115 70.320 ;
        RECT 73.745 69.960 73.915 70.130 ;
        RECT 75.600 69.970 75.770 70.140 ;
        RECT 77.280 70.330 77.450 70.500 ;
        RECT 80.985 70.580 81.155 70.750 ;
        RECT 81.345 70.580 81.515 70.750 ;
        RECT 81.705 70.580 81.875 70.750 ;
        RECT 82.065 70.580 82.235 70.750 ;
        RECT 82.425 70.580 82.595 70.750 ;
        RECT 85.375 70.580 85.545 70.750 ;
        RECT 85.735 70.580 85.905 70.750 ;
        RECT 86.575 70.680 86.745 70.850 ;
        RECT 80.160 70.320 80.330 70.490 ;
        RECT 83.040 70.330 83.210 70.500 ;
        RECT 77.895 70.150 78.065 70.320 ;
        RECT 78.255 70.150 78.425 70.320 ;
        RECT 78.615 70.150 78.785 70.320 ;
        RECT 78.975 70.150 79.145 70.320 ;
        RECT 79.335 70.150 79.505 70.320 ;
        RECT 77.280 69.970 77.450 70.140 ;
        RECT 80.985 70.150 81.155 70.320 ;
        RECT 81.345 70.150 81.515 70.320 ;
        RECT 81.705 70.150 81.875 70.320 ;
        RECT 82.065 70.150 82.235 70.320 ;
        RECT 82.425 70.150 82.595 70.320 ;
        RECT 80.160 69.960 80.330 70.130 ;
        RECT 83.040 69.970 83.210 70.140 ;
        RECT 84.720 70.330 84.890 70.500 ;
        RECT 86.575 70.320 86.745 70.490 ;
        RECT 85.375 70.150 85.545 70.320 ;
        RECT 85.735 70.150 85.905 70.320 ;
        RECT 84.720 69.970 84.890 70.140 ;
        RECT 73.745 69.600 73.915 69.770 ;
        RECT 74.585 69.720 74.755 69.890 ;
        RECT 74.945 69.720 75.115 69.890 ;
        RECT 77.895 69.720 78.065 69.890 ;
        RECT 78.255 69.720 78.425 69.890 ;
        RECT 78.615 69.720 78.785 69.890 ;
        RECT 78.975 69.720 79.145 69.890 ;
        RECT 79.335 69.720 79.505 69.890 ;
        RECT 86.575 69.960 86.745 70.130 ;
        RECT 75.600 69.470 75.770 69.640 ;
        RECT 73.745 69.240 73.915 69.410 ;
        RECT 74.585 69.290 74.755 69.460 ;
        RECT 74.945 69.290 75.115 69.460 ;
        RECT 75.600 69.110 75.770 69.280 ;
        RECT 77.280 69.470 77.450 69.640 ;
        RECT 80.160 69.600 80.330 69.770 ;
        RECT 80.985 69.720 81.155 69.890 ;
        RECT 81.345 69.720 81.515 69.890 ;
        RECT 81.705 69.720 81.875 69.890 ;
        RECT 82.065 69.720 82.235 69.890 ;
        RECT 82.425 69.720 82.595 69.890 ;
        RECT 85.375 69.720 85.545 69.890 ;
        RECT 85.735 69.720 85.905 69.890 ;
        RECT 77.895 69.290 78.065 69.460 ;
        RECT 78.255 69.290 78.425 69.460 ;
        RECT 78.615 69.290 78.785 69.460 ;
        RECT 78.975 69.290 79.145 69.460 ;
        RECT 79.335 69.290 79.505 69.460 ;
        RECT 83.040 69.470 83.210 69.640 ;
        RECT 77.280 69.110 77.450 69.280 ;
        RECT 80.160 69.240 80.330 69.410 ;
        RECT 80.985 69.290 81.155 69.460 ;
        RECT 81.345 69.290 81.515 69.460 ;
        RECT 81.705 69.290 81.875 69.460 ;
        RECT 82.065 69.290 82.235 69.460 ;
        RECT 82.425 69.290 82.595 69.460 ;
        RECT 73.745 68.880 73.915 69.050 ;
        RECT 83.040 69.110 83.210 69.280 ;
        RECT 84.720 69.470 84.890 69.640 ;
        RECT 86.575 69.600 86.745 69.770 ;
        RECT 85.375 69.290 85.545 69.460 ;
        RECT 85.735 69.290 85.905 69.460 ;
        RECT 84.720 69.110 84.890 69.280 ;
        RECT 86.575 69.240 86.745 69.410 ;
        RECT 74.585 68.860 74.755 69.030 ;
        RECT 74.945 68.860 75.115 69.030 ;
        RECT 77.895 68.860 78.065 69.030 ;
        RECT 78.255 68.860 78.425 69.030 ;
        RECT 78.615 68.860 78.785 69.030 ;
        RECT 78.975 68.860 79.145 69.030 ;
        RECT 79.335 68.860 79.505 69.030 ;
        RECT 80.160 68.880 80.330 69.050 ;
        RECT 73.745 68.520 73.915 68.690 ;
        RECT 75.600 68.610 75.770 68.780 ;
        RECT 74.585 68.430 74.755 68.600 ;
        RECT 74.945 68.430 75.115 68.600 ;
        RECT 73.745 68.160 73.915 68.330 ;
        RECT 75.600 68.250 75.770 68.420 ;
        RECT 77.280 68.610 77.450 68.780 ;
        RECT 80.985 68.860 81.155 69.030 ;
        RECT 81.345 68.860 81.515 69.030 ;
        RECT 81.705 68.860 81.875 69.030 ;
        RECT 82.065 68.860 82.235 69.030 ;
        RECT 82.425 68.860 82.595 69.030 ;
        RECT 85.375 68.860 85.545 69.030 ;
        RECT 85.735 68.860 85.905 69.030 ;
        RECT 86.575 68.880 86.745 69.050 ;
        RECT 77.895 68.430 78.065 68.600 ;
        RECT 78.255 68.430 78.425 68.600 ;
        RECT 78.615 68.430 78.785 68.600 ;
        RECT 78.975 68.430 79.145 68.600 ;
        RECT 79.335 68.430 79.505 68.600 ;
        RECT 80.160 68.520 80.330 68.690 ;
        RECT 83.040 68.610 83.210 68.780 ;
        RECT 77.280 68.250 77.450 68.420 ;
        RECT 80.985 68.430 81.155 68.600 ;
        RECT 81.345 68.430 81.515 68.600 ;
        RECT 81.705 68.430 81.875 68.600 ;
        RECT 82.065 68.430 82.235 68.600 ;
        RECT 82.425 68.430 82.595 68.600 ;
        RECT 74.585 68.000 74.755 68.170 ;
        RECT 74.945 68.000 75.115 68.170 ;
        RECT 77.895 68.000 78.065 68.170 ;
        RECT 78.255 68.000 78.425 68.170 ;
        RECT 78.615 68.000 78.785 68.170 ;
        RECT 78.975 68.000 79.145 68.170 ;
        RECT 79.335 68.000 79.505 68.170 ;
        RECT 80.160 68.160 80.330 68.330 ;
        RECT 83.040 68.250 83.210 68.420 ;
        RECT 84.720 68.610 84.890 68.780 ;
        RECT 85.375 68.430 85.545 68.600 ;
        RECT 85.735 68.430 85.905 68.600 ;
        RECT 86.575 68.520 86.745 68.690 ;
        RECT 84.720 68.250 84.890 68.420 ;
        RECT 73.745 67.800 73.915 67.970 ;
        RECT 80.985 68.000 81.155 68.170 ;
        RECT 81.345 68.000 81.515 68.170 ;
        RECT 81.705 68.000 81.875 68.170 ;
        RECT 82.065 68.000 82.235 68.170 ;
        RECT 82.425 68.000 82.595 68.170 ;
        RECT 85.375 68.000 85.545 68.170 ;
        RECT 85.735 68.000 85.905 68.170 ;
        RECT 86.575 68.160 86.745 68.330 ;
        RECT 75.600 67.750 75.770 67.920 ;
        RECT 73.745 67.440 73.915 67.610 ;
        RECT 74.585 67.570 74.755 67.740 ;
        RECT 74.945 67.570 75.115 67.740 ;
        RECT 75.600 67.390 75.770 67.560 ;
        RECT 77.280 67.750 77.450 67.920 ;
        RECT 80.160 67.800 80.330 67.970 ;
        RECT 77.895 67.570 78.065 67.740 ;
        RECT 78.255 67.570 78.425 67.740 ;
        RECT 78.615 67.570 78.785 67.740 ;
        RECT 78.975 67.570 79.145 67.740 ;
        RECT 79.335 67.570 79.505 67.740 ;
        RECT 83.040 67.750 83.210 67.920 ;
        RECT 77.280 67.390 77.450 67.560 ;
        RECT 80.160 67.440 80.330 67.610 ;
        RECT 80.985 67.570 81.155 67.740 ;
        RECT 81.345 67.570 81.515 67.740 ;
        RECT 81.705 67.570 81.875 67.740 ;
        RECT 82.065 67.570 82.235 67.740 ;
        RECT 82.425 67.570 82.595 67.740 ;
        RECT 73.745 67.080 73.915 67.250 ;
        RECT 74.585 67.140 74.755 67.310 ;
        RECT 74.945 67.140 75.115 67.310 ;
        RECT 77.895 67.140 78.065 67.310 ;
        RECT 78.255 67.140 78.425 67.310 ;
        RECT 78.615 67.140 78.785 67.310 ;
        RECT 78.975 67.140 79.145 67.310 ;
        RECT 79.335 67.140 79.505 67.310 ;
        RECT 83.040 67.390 83.210 67.560 ;
        RECT 84.720 67.750 84.890 67.920 ;
        RECT 86.575 67.800 86.745 67.970 ;
        RECT 85.375 67.570 85.545 67.740 ;
        RECT 85.735 67.570 85.905 67.740 ;
        RECT 84.720 67.390 84.890 67.560 ;
        RECT 86.575 67.440 86.745 67.610 ;
        RECT 80.160 67.080 80.330 67.250 ;
        RECT 80.985 67.140 81.155 67.310 ;
        RECT 81.345 67.140 81.515 67.310 ;
        RECT 81.705 67.140 81.875 67.310 ;
        RECT 82.065 67.140 82.235 67.310 ;
        RECT 82.425 67.140 82.595 67.310 ;
        RECT 85.375 67.140 85.545 67.310 ;
        RECT 85.735 67.140 85.905 67.310 ;
        RECT 73.745 66.720 73.915 66.890 ;
        RECT 75.600 66.890 75.770 67.060 ;
        RECT 74.585 66.710 74.755 66.880 ;
        RECT 74.945 66.710 75.115 66.880 ;
        RECT 75.600 66.530 75.770 66.700 ;
        RECT 77.280 66.890 77.450 67.060 ;
        RECT 86.575 67.080 86.745 67.250 ;
        RECT 77.895 66.710 78.065 66.880 ;
        RECT 78.255 66.710 78.425 66.880 ;
        RECT 78.615 66.710 78.785 66.880 ;
        RECT 78.975 66.710 79.145 66.880 ;
        RECT 79.335 66.710 79.505 66.880 ;
        RECT 80.160 66.720 80.330 66.890 ;
        RECT 83.040 66.890 83.210 67.060 ;
        RECT 77.280 66.530 77.450 66.700 ;
        RECT 80.985 66.710 81.155 66.880 ;
        RECT 81.345 66.710 81.515 66.880 ;
        RECT 81.705 66.710 81.875 66.880 ;
        RECT 82.065 66.710 82.235 66.880 ;
        RECT 82.425 66.710 82.595 66.880 ;
        RECT 83.040 66.530 83.210 66.700 ;
        RECT 84.720 66.890 84.890 67.060 ;
        RECT 85.375 66.710 85.545 66.880 ;
        RECT 85.735 66.710 85.905 66.880 ;
        RECT 86.575 66.720 86.745 66.890 ;
        RECT 84.720 66.530 84.890 66.700 ;
        RECT 73.745 66.360 73.915 66.530 ;
        RECT 74.585 66.280 74.755 66.450 ;
        RECT 74.945 66.280 75.115 66.450 ;
        RECT 77.895 66.280 78.065 66.450 ;
        RECT 78.255 66.280 78.425 66.450 ;
        RECT 78.615 66.280 78.785 66.450 ;
        RECT 78.975 66.280 79.145 66.450 ;
        RECT 79.335 66.280 79.505 66.450 ;
        RECT 80.160 66.360 80.330 66.530 ;
        RECT 73.745 66.000 73.915 66.170 ;
        RECT 75.600 66.030 75.770 66.200 ;
        RECT 74.585 65.850 74.755 66.020 ;
        RECT 74.945 65.850 75.115 66.020 ;
        RECT 73.745 65.640 73.915 65.810 ;
        RECT 75.600 65.670 75.770 65.840 ;
        RECT 77.280 66.030 77.450 66.200 ;
        RECT 80.985 66.280 81.155 66.450 ;
        RECT 81.345 66.280 81.515 66.450 ;
        RECT 81.705 66.280 81.875 66.450 ;
        RECT 82.065 66.280 82.235 66.450 ;
        RECT 82.425 66.280 82.595 66.450 ;
        RECT 85.375 66.280 85.545 66.450 ;
        RECT 85.735 66.280 85.905 66.450 ;
        RECT 86.575 66.360 86.745 66.530 ;
        RECT 77.895 65.850 78.065 66.020 ;
        RECT 78.255 65.850 78.425 66.020 ;
        RECT 78.615 65.850 78.785 66.020 ;
        RECT 78.975 65.850 79.145 66.020 ;
        RECT 79.335 65.850 79.505 66.020 ;
        RECT 80.160 66.000 80.330 66.170 ;
        RECT 83.040 66.030 83.210 66.200 ;
        RECT 77.280 65.670 77.450 65.840 ;
        RECT 80.985 65.850 81.155 66.020 ;
        RECT 81.345 65.850 81.515 66.020 ;
        RECT 81.705 65.850 81.875 66.020 ;
        RECT 82.065 65.850 82.235 66.020 ;
        RECT 82.425 65.850 82.595 66.020 ;
        RECT 80.160 65.640 80.330 65.810 ;
        RECT 83.040 65.670 83.210 65.840 ;
        RECT 84.720 66.030 84.890 66.200 ;
        RECT 85.375 65.850 85.545 66.020 ;
        RECT 85.735 65.850 85.905 66.020 ;
        RECT 86.575 66.000 86.745 66.170 ;
        RECT 84.720 65.670 84.890 65.840 ;
        RECT 73.745 65.280 73.915 65.450 ;
        RECT 74.585 65.420 74.755 65.590 ;
        RECT 74.945 65.420 75.115 65.590 ;
        RECT 77.895 65.420 78.065 65.590 ;
        RECT 78.255 65.420 78.425 65.590 ;
        RECT 78.615 65.420 78.785 65.590 ;
        RECT 78.975 65.420 79.145 65.590 ;
        RECT 79.335 65.420 79.505 65.590 ;
        RECT 86.575 65.640 86.745 65.810 ;
        RECT 75.600 65.170 75.770 65.340 ;
        RECT 73.745 64.920 73.915 65.090 ;
        RECT 74.585 64.990 74.755 65.160 ;
        RECT 74.945 64.990 75.115 65.160 ;
        RECT 75.600 64.810 75.770 64.980 ;
        RECT 77.280 65.170 77.450 65.340 ;
        RECT 80.160 65.280 80.330 65.450 ;
        RECT 80.985 65.420 81.155 65.590 ;
        RECT 81.345 65.420 81.515 65.590 ;
        RECT 81.705 65.420 81.875 65.590 ;
        RECT 82.065 65.420 82.235 65.590 ;
        RECT 82.425 65.420 82.595 65.590 ;
        RECT 85.375 65.420 85.545 65.590 ;
        RECT 85.735 65.420 85.905 65.590 ;
        RECT 77.895 64.990 78.065 65.160 ;
        RECT 78.255 64.990 78.425 65.160 ;
        RECT 78.615 64.990 78.785 65.160 ;
        RECT 78.975 64.990 79.145 65.160 ;
        RECT 79.335 64.990 79.505 65.160 ;
        RECT 83.040 65.170 83.210 65.340 ;
        RECT 77.280 64.810 77.450 64.980 ;
        RECT 80.160 64.920 80.330 65.090 ;
        RECT 80.985 64.990 81.155 65.160 ;
        RECT 81.345 64.990 81.515 65.160 ;
        RECT 81.705 64.990 81.875 65.160 ;
        RECT 82.065 64.990 82.235 65.160 ;
        RECT 82.425 64.990 82.595 65.160 ;
        RECT 83.040 64.810 83.210 64.980 ;
        RECT 84.720 65.170 84.890 65.340 ;
        RECT 86.575 65.280 86.745 65.450 ;
        RECT 85.375 64.990 85.545 65.160 ;
        RECT 85.735 64.990 85.905 65.160 ;
        RECT 84.720 64.810 84.890 64.980 ;
        RECT 86.575 64.920 86.745 65.090 ;
        RECT 73.745 64.560 73.915 64.730 ;
        RECT 74.585 64.560 74.755 64.730 ;
        RECT 74.945 64.560 75.115 64.730 ;
        RECT 77.895 64.560 78.065 64.730 ;
        RECT 78.255 64.560 78.425 64.730 ;
        RECT 78.615 64.560 78.785 64.730 ;
        RECT 78.975 64.560 79.145 64.730 ;
        RECT 79.335 64.560 79.505 64.730 ;
        RECT 80.160 64.560 80.330 64.730 ;
        RECT 80.985 64.560 81.155 64.730 ;
        RECT 81.345 64.560 81.515 64.730 ;
        RECT 81.705 64.560 81.875 64.730 ;
        RECT 82.065 64.560 82.235 64.730 ;
        RECT 82.425 64.560 82.595 64.730 ;
        RECT 85.375 64.560 85.545 64.730 ;
        RECT 85.735 64.560 85.905 64.730 ;
        RECT 86.575 64.560 86.745 64.730 ;
        RECT 73.745 64.200 73.915 64.370 ;
        RECT 75.600 64.310 75.770 64.480 ;
        RECT 74.585 64.130 74.755 64.300 ;
        RECT 74.945 64.130 75.115 64.300 ;
        RECT 73.745 63.840 73.915 64.010 ;
        RECT 75.600 63.950 75.770 64.120 ;
        RECT 77.280 64.310 77.450 64.480 ;
        RECT 77.895 64.130 78.065 64.300 ;
        RECT 78.255 64.130 78.425 64.300 ;
        RECT 78.615 64.130 78.785 64.300 ;
        RECT 78.975 64.130 79.145 64.300 ;
        RECT 79.335 64.130 79.505 64.300 ;
        RECT 80.160 64.200 80.330 64.370 ;
        RECT 83.040 64.310 83.210 64.480 ;
        RECT 77.280 63.950 77.450 64.120 ;
        RECT 80.985 64.130 81.155 64.300 ;
        RECT 81.345 64.130 81.515 64.300 ;
        RECT 81.705 64.130 81.875 64.300 ;
        RECT 82.065 64.130 82.235 64.300 ;
        RECT 82.425 64.130 82.595 64.300 ;
        RECT 74.585 63.700 74.755 63.870 ;
        RECT 74.945 63.700 75.115 63.870 ;
        RECT 77.895 63.700 78.065 63.870 ;
        RECT 78.255 63.700 78.425 63.870 ;
        RECT 78.615 63.700 78.785 63.870 ;
        RECT 78.975 63.700 79.145 63.870 ;
        RECT 79.335 63.700 79.505 63.870 ;
        RECT 80.160 63.840 80.330 64.010 ;
        RECT 83.040 63.950 83.210 64.120 ;
        RECT 84.720 64.310 84.890 64.480 ;
        RECT 85.375 64.130 85.545 64.300 ;
        RECT 85.735 64.130 85.905 64.300 ;
        RECT 86.575 64.200 86.745 64.370 ;
        RECT 84.720 63.950 84.890 64.120 ;
        RECT 73.745 63.480 73.915 63.650 ;
        RECT 80.985 63.700 81.155 63.870 ;
        RECT 81.345 63.700 81.515 63.870 ;
        RECT 81.705 63.700 81.875 63.870 ;
        RECT 82.065 63.700 82.235 63.870 ;
        RECT 82.425 63.700 82.595 63.870 ;
        RECT 85.375 63.700 85.545 63.870 ;
        RECT 85.735 63.700 85.905 63.870 ;
        RECT 86.575 63.840 86.745 64.010 ;
        RECT 80.160 63.480 80.330 63.650 ;
        RECT 86.575 63.480 86.745 63.650 ;
        RECT 74.045 63.030 74.215 63.200 ;
        RECT 74.405 63.030 74.575 63.200 ;
        RECT 74.765 63.030 74.935 63.200 ;
        RECT 75.125 63.030 75.295 63.200 ;
        RECT 75.485 63.030 75.655 63.200 ;
        RECT 75.845 63.030 76.015 63.200 ;
        RECT 77.340 63.030 77.510 63.200 ;
        RECT 77.700 63.030 77.870 63.200 ;
        RECT 78.060 63.030 78.230 63.200 ;
        RECT 78.420 63.030 78.590 63.200 ;
        RECT 78.780 63.030 78.950 63.200 ;
        RECT 79.140 63.030 79.310 63.200 ;
        RECT 79.500 63.030 79.670 63.200 ;
        RECT 79.860 63.030 80.030 63.200 ;
        RECT 80.460 63.030 80.630 63.200 ;
        RECT 80.820 63.030 80.990 63.200 ;
        RECT 81.180 63.030 81.350 63.200 ;
        RECT 81.540 63.030 81.710 63.200 ;
        RECT 81.900 63.030 82.070 63.200 ;
        RECT 82.260 63.030 82.430 63.200 ;
        RECT 82.620 63.030 82.790 63.200 ;
        RECT 82.980 63.030 83.150 63.200 ;
        RECT 84.475 63.030 84.645 63.200 ;
        RECT 84.835 63.030 85.005 63.200 ;
        RECT 85.195 63.030 85.365 63.200 ;
        RECT 85.555 63.030 85.725 63.200 ;
        RECT 85.915 63.030 86.085 63.200 ;
        RECT 86.275 63.030 86.445 63.200 ;
        RECT 88.805 72.110 88.975 72.280 ;
        RECT 89.165 72.110 89.335 72.280 ;
        RECT 89.525 72.110 89.695 72.280 ;
        RECT 89.885 72.110 90.055 72.280 ;
        RECT 90.245 72.110 90.415 72.280 ;
        RECT 90.605 72.110 90.775 72.280 ;
        RECT 92.100 72.110 92.270 72.280 ;
        RECT 92.460 72.110 92.630 72.280 ;
        RECT 92.820 72.110 92.990 72.280 ;
        RECT 93.180 72.110 93.350 72.280 ;
        RECT 93.540 72.110 93.710 72.280 ;
        RECT 93.900 72.110 94.070 72.280 ;
        RECT 94.260 72.110 94.430 72.280 ;
        RECT 94.620 72.110 94.790 72.280 ;
        RECT 88.505 71.760 88.675 71.930 ;
        RECT 94.920 71.760 95.090 71.930 ;
        RECT 88.505 71.400 88.675 71.570 ;
        RECT 89.345 71.440 89.515 71.610 ;
        RECT 89.705 71.440 89.875 71.610 ;
        RECT 92.655 71.440 92.825 71.610 ;
        RECT 93.015 71.440 93.185 71.610 ;
        RECT 93.375 71.440 93.545 71.610 ;
        RECT 93.735 71.440 93.905 71.610 ;
        RECT 94.095 71.440 94.265 71.610 ;
        RECT 94.920 71.400 95.090 71.570 ;
        RECT 88.505 71.040 88.675 71.210 ;
        RECT 90.360 71.190 90.530 71.360 ;
        RECT 89.345 71.010 89.515 71.180 ;
        RECT 89.705 71.010 89.875 71.180 ;
        RECT 88.505 70.680 88.675 70.850 ;
        RECT 90.360 70.830 90.530 71.000 ;
        RECT 92.040 71.190 92.210 71.360 ;
        RECT 92.655 71.010 92.825 71.180 ;
        RECT 93.015 71.010 93.185 71.180 ;
        RECT 93.375 71.010 93.545 71.180 ;
        RECT 93.735 71.010 93.905 71.180 ;
        RECT 94.095 71.010 94.265 71.180 ;
        RECT 94.920 71.040 95.090 71.210 ;
        RECT 92.040 70.830 92.210 71.000 ;
        RECT 89.345 70.580 89.515 70.750 ;
        RECT 89.705 70.580 89.875 70.750 ;
        RECT 92.655 70.580 92.825 70.750 ;
        RECT 93.015 70.580 93.185 70.750 ;
        RECT 93.375 70.580 93.545 70.750 ;
        RECT 93.735 70.580 93.905 70.750 ;
        RECT 94.095 70.580 94.265 70.750 ;
        RECT 94.920 70.680 95.090 70.850 ;
        RECT 88.505 70.320 88.675 70.490 ;
        RECT 90.360 70.330 90.530 70.500 ;
        RECT 89.345 70.150 89.515 70.320 ;
        RECT 89.705 70.150 89.875 70.320 ;
        RECT 88.505 69.960 88.675 70.130 ;
        RECT 90.360 69.970 90.530 70.140 ;
        RECT 92.040 70.330 92.210 70.500 ;
        RECT 94.920 70.320 95.090 70.490 ;
        RECT 92.655 70.150 92.825 70.320 ;
        RECT 93.015 70.150 93.185 70.320 ;
        RECT 93.375 70.150 93.545 70.320 ;
        RECT 93.735 70.150 93.905 70.320 ;
        RECT 94.095 70.150 94.265 70.320 ;
        RECT 92.040 69.970 92.210 70.140 ;
        RECT 94.920 69.960 95.090 70.130 ;
        RECT 88.505 69.600 88.675 69.770 ;
        RECT 89.345 69.720 89.515 69.890 ;
        RECT 89.705 69.720 89.875 69.890 ;
        RECT 92.655 69.720 92.825 69.890 ;
        RECT 93.015 69.720 93.185 69.890 ;
        RECT 93.375 69.720 93.545 69.890 ;
        RECT 93.735 69.720 93.905 69.890 ;
        RECT 94.095 69.720 94.265 69.890 ;
        RECT 90.360 69.470 90.530 69.640 ;
        RECT 88.505 69.240 88.675 69.410 ;
        RECT 89.345 69.290 89.515 69.460 ;
        RECT 89.705 69.290 89.875 69.460 ;
        RECT 90.360 69.110 90.530 69.280 ;
        RECT 92.040 69.470 92.210 69.640 ;
        RECT 94.920 69.600 95.090 69.770 ;
        RECT 92.655 69.290 92.825 69.460 ;
        RECT 93.015 69.290 93.185 69.460 ;
        RECT 93.375 69.290 93.545 69.460 ;
        RECT 93.735 69.290 93.905 69.460 ;
        RECT 94.095 69.290 94.265 69.460 ;
        RECT 92.040 69.110 92.210 69.280 ;
        RECT 94.920 69.240 95.090 69.410 ;
        RECT 88.505 68.880 88.675 69.050 ;
        RECT 89.345 68.860 89.515 69.030 ;
        RECT 89.705 68.860 89.875 69.030 ;
        RECT 92.655 68.860 92.825 69.030 ;
        RECT 93.015 68.860 93.185 69.030 ;
        RECT 93.375 68.860 93.545 69.030 ;
        RECT 93.735 68.860 93.905 69.030 ;
        RECT 94.095 68.860 94.265 69.030 ;
        RECT 94.920 68.880 95.090 69.050 ;
        RECT 88.505 68.520 88.675 68.690 ;
        RECT 90.360 68.610 90.530 68.780 ;
        RECT 89.345 68.430 89.515 68.600 ;
        RECT 89.705 68.430 89.875 68.600 ;
        RECT 88.505 68.160 88.675 68.330 ;
        RECT 90.360 68.250 90.530 68.420 ;
        RECT 92.040 68.610 92.210 68.780 ;
        RECT 92.655 68.430 92.825 68.600 ;
        RECT 93.015 68.430 93.185 68.600 ;
        RECT 93.375 68.430 93.545 68.600 ;
        RECT 93.735 68.430 93.905 68.600 ;
        RECT 94.095 68.430 94.265 68.600 ;
        RECT 94.920 68.520 95.090 68.690 ;
        RECT 92.040 68.250 92.210 68.420 ;
        RECT 89.345 68.000 89.515 68.170 ;
        RECT 89.705 68.000 89.875 68.170 ;
        RECT 92.655 68.000 92.825 68.170 ;
        RECT 93.015 68.000 93.185 68.170 ;
        RECT 93.375 68.000 93.545 68.170 ;
        RECT 93.735 68.000 93.905 68.170 ;
        RECT 94.095 68.000 94.265 68.170 ;
        RECT 94.920 68.160 95.090 68.330 ;
        RECT 88.505 67.800 88.675 67.970 ;
        RECT 90.360 67.750 90.530 67.920 ;
        RECT 88.505 67.440 88.675 67.610 ;
        RECT 89.345 67.570 89.515 67.740 ;
        RECT 89.705 67.570 89.875 67.740 ;
        RECT 90.360 67.390 90.530 67.560 ;
        RECT 92.040 67.750 92.210 67.920 ;
        RECT 94.920 67.800 95.090 67.970 ;
        RECT 92.655 67.570 92.825 67.740 ;
        RECT 93.015 67.570 93.185 67.740 ;
        RECT 93.375 67.570 93.545 67.740 ;
        RECT 93.735 67.570 93.905 67.740 ;
        RECT 94.095 67.570 94.265 67.740 ;
        RECT 92.040 67.390 92.210 67.560 ;
        RECT 94.920 67.440 95.090 67.610 ;
        RECT 88.505 67.080 88.675 67.250 ;
        RECT 89.345 67.140 89.515 67.310 ;
        RECT 89.705 67.140 89.875 67.310 ;
        RECT 92.655 67.140 92.825 67.310 ;
        RECT 93.015 67.140 93.185 67.310 ;
        RECT 93.375 67.140 93.545 67.310 ;
        RECT 93.735 67.140 93.905 67.310 ;
        RECT 94.095 67.140 94.265 67.310 ;
        RECT 94.920 67.080 95.090 67.250 ;
        RECT 88.505 66.720 88.675 66.890 ;
        RECT 90.360 66.890 90.530 67.060 ;
        RECT 89.345 66.710 89.515 66.880 ;
        RECT 89.705 66.710 89.875 66.880 ;
        RECT 90.360 66.530 90.530 66.700 ;
        RECT 92.040 66.890 92.210 67.060 ;
        RECT 92.655 66.710 92.825 66.880 ;
        RECT 93.015 66.710 93.185 66.880 ;
        RECT 93.375 66.710 93.545 66.880 ;
        RECT 93.735 66.710 93.905 66.880 ;
        RECT 94.095 66.710 94.265 66.880 ;
        RECT 94.920 66.720 95.090 66.890 ;
        RECT 92.040 66.530 92.210 66.700 ;
        RECT 88.505 66.360 88.675 66.530 ;
        RECT 89.345 66.280 89.515 66.450 ;
        RECT 89.705 66.280 89.875 66.450 ;
        RECT 92.655 66.280 92.825 66.450 ;
        RECT 93.015 66.280 93.185 66.450 ;
        RECT 93.375 66.280 93.545 66.450 ;
        RECT 93.735 66.280 93.905 66.450 ;
        RECT 94.095 66.280 94.265 66.450 ;
        RECT 94.920 66.360 95.090 66.530 ;
        RECT 88.505 66.000 88.675 66.170 ;
        RECT 90.360 66.030 90.530 66.200 ;
        RECT 89.345 65.850 89.515 66.020 ;
        RECT 89.705 65.850 89.875 66.020 ;
        RECT 88.505 65.640 88.675 65.810 ;
        RECT 90.360 65.670 90.530 65.840 ;
        RECT 92.040 66.030 92.210 66.200 ;
        RECT 92.655 65.850 92.825 66.020 ;
        RECT 93.015 65.850 93.185 66.020 ;
        RECT 93.375 65.850 93.545 66.020 ;
        RECT 93.735 65.850 93.905 66.020 ;
        RECT 94.095 65.850 94.265 66.020 ;
        RECT 94.920 66.000 95.090 66.170 ;
        RECT 92.040 65.670 92.210 65.840 ;
        RECT 94.920 65.640 95.090 65.810 ;
        RECT 88.505 65.280 88.675 65.450 ;
        RECT 89.345 65.420 89.515 65.590 ;
        RECT 89.705 65.420 89.875 65.590 ;
        RECT 92.655 65.420 92.825 65.590 ;
        RECT 93.015 65.420 93.185 65.590 ;
        RECT 93.375 65.420 93.545 65.590 ;
        RECT 93.735 65.420 93.905 65.590 ;
        RECT 94.095 65.420 94.265 65.590 ;
        RECT 90.360 65.170 90.530 65.340 ;
        RECT 88.505 64.920 88.675 65.090 ;
        RECT 89.345 64.990 89.515 65.160 ;
        RECT 89.705 64.990 89.875 65.160 ;
        RECT 90.360 64.810 90.530 64.980 ;
        RECT 92.040 65.170 92.210 65.340 ;
        RECT 94.920 65.280 95.090 65.450 ;
        RECT 92.655 64.990 92.825 65.160 ;
        RECT 93.015 64.990 93.185 65.160 ;
        RECT 93.375 64.990 93.545 65.160 ;
        RECT 93.735 64.990 93.905 65.160 ;
        RECT 94.095 64.990 94.265 65.160 ;
        RECT 92.040 64.810 92.210 64.980 ;
        RECT 94.920 64.920 95.090 65.090 ;
        RECT 88.505 64.560 88.675 64.730 ;
        RECT 89.345 64.560 89.515 64.730 ;
        RECT 89.705 64.560 89.875 64.730 ;
        RECT 92.655 64.560 92.825 64.730 ;
        RECT 93.015 64.560 93.185 64.730 ;
        RECT 93.375 64.560 93.545 64.730 ;
        RECT 93.735 64.560 93.905 64.730 ;
        RECT 94.095 64.560 94.265 64.730 ;
        RECT 94.920 64.560 95.090 64.730 ;
        RECT 88.505 64.200 88.675 64.370 ;
        RECT 90.360 64.310 90.530 64.480 ;
        RECT 89.345 64.130 89.515 64.300 ;
        RECT 89.705 64.130 89.875 64.300 ;
        RECT 88.505 63.840 88.675 64.010 ;
        RECT 90.360 63.950 90.530 64.120 ;
        RECT 92.040 64.310 92.210 64.480 ;
        RECT 92.655 64.130 92.825 64.300 ;
        RECT 93.015 64.130 93.185 64.300 ;
        RECT 93.375 64.130 93.545 64.300 ;
        RECT 93.735 64.130 93.905 64.300 ;
        RECT 94.095 64.130 94.265 64.300 ;
        RECT 94.920 64.200 95.090 64.370 ;
        RECT 92.040 63.950 92.210 64.120 ;
        RECT 89.345 63.700 89.515 63.870 ;
        RECT 89.705 63.700 89.875 63.870 ;
        RECT 92.655 63.700 92.825 63.870 ;
        RECT 93.015 63.700 93.185 63.870 ;
        RECT 93.375 63.700 93.545 63.870 ;
        RECT 93.735 63.700 93.905 63.870 ;
        RECT 94.095 63.700 94.265 63.870 ;
        RECT 94.920 63.840 95.090 64.010 ;
        RECT 88.505 63.480 88.675 63.650 ;
        RECT 94.920 63.480 95.090 63.650 ;
        RECT 88.805 63.030 88.975 63.200 ;
        RECT 89.165 63.030 89.335 63.200 ;
        RECT 89.525 63.030 89.695 63.200 ;
        RECT 89.885 63.030 90.055 63.200 ;
        RECT 90.245 63.030 90.415 63.200 ;
        RECT 90.605 63.030 90.775 63.200 ;
        RECT 92.100 63.030 92.270 63.200 ;
        RECT 92.460 63.030 92.630 63.200 ;
        RECT 92.820 63.030 92.990 63.200 ;
        RECT 93.180 63.030 93.350 63.200 ;
        RECT 93.540 63.030 93.710 63.200 ;
        RECT 93.900 63.030 94.070 63.200 ;
        RECT 94.260 63.030 94.430 63.200 ;
        RECT 94.620 63.030 94.790 63.200 ;
        RECT 113.845 72.620 114.015 72.790 ;
        RECT 108.635 72.090 108.805 72.260 ;
        RECT 108.635 71.730 108.805 71.900 ;
        RECT 108.635 71.370 108.805 71.540 ;
        RECT 108.635 71.010 108.805 71.180 ;
        RECT 108.635 70.650 108.805 70.820 ;
        RECT 110.555 72.210 110.725 72.380 ;
        RECT 110.555 71.850 110.725 72.020 ;
        RECT 110.555 71.490 110.725 71.660 ;
        RECT 110.555 71.130 110.725 71.300 ;
        RECT 110.555 70.770 110.725 70.940 ;
        RECT 111.925 72.210 112.095 72.380 ;
        RECT 111.925 71.850 112.095 72.020 ;
        RECT 111.925 71.490 112.095 71.660 ;
        RECT 111.925 71.130 112.095 71.300 ;
        RECT 111.925 70.770 112.095 70.940 ;
        RECT 113.845 72.260 114.015 72.430 ;
        RECT 113.845 71.900 114.015 72.070 ;
        RECT 113.845 71.540 114.015 71.710 ;
        RECT 113.845 71.180 114.015 71.350 ;
        RECT 113.845 70.820 114.015 70.990 ;
        RECT 108.635 70.290 108.805 70.460 ;
        RECT 109.690 70.350 109.860 70.520 ;
        RECT 110.050 70.350 110.220 70.520 ;
        RECT 111.060 70.350 111.230 70.520 ;
        RECT 111.420 70.350 111.590 70.520 ;
        RECT 112.430 70.350 112.600 70.520 ;
        RECT 112.790 70.350 112.960 70.520 ;
        RECT 113.845 70.460 114.015 70.630 ;
        RECT 113.845 70.100 114.015 70.270 ;
        RECT 108.635 69.930 108.805 70.100 ;
        RECT 108.635 69.570 108.805 69.740 ;
        RECT 108.635 69.210 108.805 69.380 ;
        RECT 108.635 68.850 108.805 69.020 ;
        RECT 108.635 68.490 108.805 68.660 ;
        RECT 110.555 69.930 110.725 70.100 ;
        RECT 110.555 69.570 110.725 69.740 ;
        RECT 110.555 69.210 110.725 69.380 ;
        RECT 110.555 68.850 110.725 69.020 ;
        RECT 110.555 68.490 110.725 68.660 ;
        RECT 111.925 69.930 112.095 70.100 ;
        RECT 111.925 69.570 112.095 69.740 ;
        RECT 111.925 69.210 112.095 69.380 ;
        RECT 111.925 68.850 112.095 69.020 ;
        RECT 111.925 68.490 112.095 68.660 ;
        RECT 113.845 69.740 114.015 69.910 ;
        RECT 113.845 69.380 114.015 69.550 ;
        RECT 113.845 69.020 114.015 69.190 ;
        RECT 113.845 68.660 114.015 68.830 ;
        RECT 108.635 68.130 108.805 68.300 ;
        RECT 113.845 68.300 114.015 68.470 ;
        RECT 109.690 68.070 109.860 68.240 ;
        RECT 110.050 68.070 110.220 68.240 ;
        RECT 111.060 68.070 111.230 68.240 ;
        RECT 111.420 68.070 111.590 68.240 ;
        RECT 112.430 68.070 112.600 68.240 ;
        RECT 112.790 68.070 112.960 68.240 ;
        RECT 108.635 67.770 108.805 67.940 ;
        RECT 113.845 67.940 114.015 68.110 ;
        RECT 108.635 67.410 108.805 67.580 ;
        RECT 108.635 67.050 108.805 67.220 ;
        RECT 108.635 66.690 108.805 66.860 ;
        RECT 108.635 66.330 108.805 66.500 ;
        RECT 110.555 67.650 110.725 67.820 ;
        RECT 110.555 67.290 110.725 67.460 ;
        RECT 110.555 66.930 110.725 67.100 ;
        RECT 110.555 66.570 110.725 66.740 ;
        RECT 110.555 66.210 110.725 66.380 ;
        RECT 111.925 67.650 112.095 67.820 ;
        RECT 111.925 67.290 112.095 67.460 ;
        RECT 111.925 66.930 112.095 67.100 ;
        RECT 111.925 66.570 112.095 66.740 ;
        RECT 111.925 66.210 112.095 66.380 ;
        RECT 113.845 67.580 114.015 67.750 ;
        RECT 113.845 67.220 114.015 67.390 ;
        RECT 113.845 66.860 114.015 67.030 ;
        RECT 113.845 66.500 114.015 66.670 ;
        RECT 108.635 65.970 108.805 66.140 ;
        RECT 113.845 66.140 114.015 66.310 ;
        RECT 109.690 65.790 109.860 65.960 ;
        RECT 110.050 65.790 110.220 65.960 ;
        RECT 111.060 65.790 111.230 65.960 ;
        RECT 111.420 65.790 111.590 65.960 ;
        RECT 112.430 65.790 112.600 65.960 ;
        RECT 112.790 65.790 112.960 65.960 ;
        RECT 108.635 65.610 108.805 65.780 ;
        RECT 113.845 65.780 114.015 65.950 ;
        RECT 108.635 65.250 108.805 65.420 ;
        RECT 108.635 64.890 108.805 65.060 ;
        RECT 108.635 64.530 108.805 64.700 ;
        RECT 108.635 64.170 108.805 64.340 ;
        RECT 108.635 63.810 108.805 63.980 ;
        RECT 110.555 65.370 110.725 65.540 ;
        RECT 110.555 65.010 110.725 65.180 ;
        RECT 110.555 64.650 110.725 64.820 ;
        RECT 110.555 64.290 110.725 64.460 ;
        RECT 110.555 63.930 110.725 64.100 ;
        RECT 111.925 65.370 112.095 65.540 ;
        RECT 111.925 65.010 112.095 65.180 ;
        RECT 111.925 64.650 112.095 64.820 ;
        RECT 111.925 64.290 112.095 64.460 ;
        RECT 111.925 63.930 112.095 64.100 ;
        RECT 113.845 65.420 114.015 65.590 ;
        RECT 113.845 65.060 114.015 65.230 ;
        RECT 113.845 64.700 114.015 64.870 ;
        RECT 113.845 64.340 114.015 64.510 ;
        RECT 113.845 63.980 114.015 64.150 ;
        RECT 108.635 63.450 108.805 63.620 ;
        RECT 109.690 63.510 109.860 63.680 ;
        RECT 110.050 63.510 110.220 63.680 ;
        RECT 111.060 63.510 111.230 63.680 ;
        RECT 111.420 63.510 111.590 63.680 ;
        RECT 112.430 63.510 112.600 63.680 ;
        RECT 112.790 63.510 112.960 63.680 ;
        RECT 113.845 63.620 114.015 63.790 ;
        RECT 113.845 63.260 114.015 63.430 ;
        RECT 108.695 62.840 108.865 63.010 ;
        RECT 109.055 62.840 109.225 63.010 ;
        RECT 109.415 62.840 109.585 63.010 ;
        RECT 109.775 62.840 109.945 63.010 ;
        RECT 110.135 62.840 110.305 63.010 ;
        RECT 110.495 62.840 110.665 63.010 ;
        RECT 110.855 62.840 111.025 63.010 ;
        RECT 111.215 62.840 111.385 63.010 ;
        RECT 111.575 62.840 111.745 63.010 ;
        RECT 111.935 62.840 112.105 63.010 ;
        RECT 112.295 62.840 112.465 63.010 ;
        RECT 112.655 62.840 112.825 63.010 ;
        RECT 113.015 62.840 113.185 63.010 ;
        RECT 113.375 62.840 113.545 63.010 ;
        RECT 113.845 62.900 114.015 63.070 ;
        RECT 114.775 70.320 114.945 70.490 ;
        RECT 115.385 70.380 115.555 70.550 ;
        RECT 115.745 70.380 115.915 70.550 ;
        RECT 116.105 70.380 116.275 70.550 ;
        RECT 116.465 70.380 116.635 70.550 ;
        RECT 116.825 70.380 116.995 70.550 ;
        RECT 117.185 70.380 117.355 70.550 ;
        RECT 114.775 69.960 114.945 70.130 ;
        RECT 114.775 69.600 114.945 69.770 ;
        RECT 115.830 69.710 116.000 69.880 ;
        RECT 116.190 69.710 116.360 69.880 ;
        RECT 117.245 69.700 117.415 69.870 ;
        RECT 114.775 69.240 114.945 69.410 ;
        RECT 114.775 68.880 114.945 69.050 ;
        RECT 114.775 68.520 114.945 68.690 ;
        RECT 114.775 68.160 114.945 68.330 ;
        RECT 114.775 67.800 114.945 67.970 ;
        RECT 116.695 69.290 116.865 69.460 ;
        RECT 116.695 68.930 116.865 69.100 ;
        RECT 116.695 68.570 116.865 68.740 ;
        RECT 116.695 68.210 116.865 68.380 ;
        RECT 116.695 67.850 116.865 68.020 ;
        RECT 117.245 69.340 117.415 69.510 ;
        RECT 117.245 68.980 117.415 69.150 ;
        RECT 117.245 68.620 117.415 68.790 ;
        RECT 117.245 68.260 117.415 68.430 ;
        RECT 117.245 67.900 117.415 68.070 ;
        RECT 114.775 67.440 114.945 67.610 ;
        RECT 115.830 67.430 116.000 67.600 ;
        RECT 116.190 67.430 116.360 67.600 ;
        RECT 117.245 67.540 117.415 67.710 ;
        RECT 114.775 67.080 114.945 67.250 ;
        RECT 117.245 67.180 117.415 67.350 ;
        RECT 114.775 66.720 114.945 66.890 ;
        RECT 114.775 66.360 114.945 66.530 ;
        RECT 114.775 66.000 114.945 66.170 ;
        RECT 114.775 65.640 114.945 65.810 ;
        RECT 115.325 67.010 115.495 67.180 ;
        RECT 115.325 66.650 115.495 66.820 ;
        RECT 115.325 66.290 115.495 66.460 ;
        RECT 115.325 65.930 115.495 66.100 ;
        RECT 115.325 65.570 115.495 65.740 ;
        RECT 117.245 66.820 117.415 66.990 ;
        RECT 117.245 66.460 117.415 66.630 ;
        RECT 117.245 66.100 117.415 66.270 ;
        RECT 117.245 65.740 117.415 65.910 ;
        RECT 117.245 65.380 117.415 65.550 ;
        RECT 115.830 65.150 116.000 65.320 ;
        RECT 116.190 65.150 116.360 65.320 ;
        RECT 118.470 70.040 118.640 70.210 ;
        RECT 119.080 70.100 119.250 70.270 ;
        RECT 119.440 70.100 119.610 70.270 ;
        RECT 119.800 70.100 119.970 70.270 ;
        RECT 120.160 70.100 120.330 70.270 ;
        RECT 120.520 70.100 120.690 70.270 ;
        RECT 120.880 70.100 121.050 70.270 ;
        RECT 121.435 70.100 121.605 70.270 ;
        RECT 121.795 70.100 121.965 70.270 ;
        RECT 122.155 70.100 122.325 70.270 ;
        RECT 122.515 70.100 122.685 70.270 ;
        RECT 122.875 70.100 123.045 70.270 ;
        RECT 123.235 70.100 123.405 70.270 ;
        RECT 123.595 70.100 123.765 70.270 ;
        RECT 118.470 69.680 118.640 69.850 ;
        RECT 123.655 69.700 123.825 69.870 ;
        RECT 118.470 69.320 118.640 69.490 ;
        RECT 119.525 69.430 119.695 69.600 ;
        RECT 119.885 69.430 120.055 69.600 ;
        RECT 122.240 69.430 122.410 69.600 ;
        RECT 122.600 69.430 122.770 69.600 ;
        RECT 123.655 69.340 123.825 69.510 ;
        RECT 118.470 68.960 118.640 69.130 ;
        RECT 119.020 69.000 119.190 69.170 ;
        RECT 119.525 69.000 119.695 69.170 ;
        RECT 119.885 69.000 120.055 69.170 ;
        RECT 121.735 69.000 121.905 69.170 ;
        RECT 122.240 69.000 122.410 69.170 ;
        RECT 122.600 69.000 122.770 69.170 ;
        RECT 118.470 68.600 118.640 68.770 ;
        RECT 123.655 68.980 123.825 69.150 ;
        RECT 119.525 68.570 119.695 68.740 ;
        RECT 119.885 68.570 120.055 68.740 ;
        RECT 122.240 68.570 122.410 68.740 ;
        RECT 122.600 68.570 122.770 68.740 ;
        RECT 123.655 68.620 123.825 68.790 ;
        RECT 118.470 68.240 118.640 68.410 ;
        RECT 119.525 68.140 119.695 68.310 ;
        RECT 119.885 68.140 120.055 68.310 ;
        RECT 120.390 68.140 120.560 68.310 ;
        RECT 122.240 68.140 122.410 68.310 ;
        RECT 122.600 68.140 122.770 68.310 ;
        RECT 123.105 68.140 123.275 68.310 ;
        RECT 123.655 68.260 123.825 68.430 ;
        RECT 118.470 67.880 118.640 68.050 ;
        RECT 123.655 67.900 123.825 68.070 ;
        RECT 119.525 67.710 119.695 67.880 ;
        RECT 119.885 67.710 120.055 67.880 ;
        RECT 122.240 67.710 122.410 67.880 ;
        RECT 122.600 67.710 122.770 67.880 ;
        RECT 118.470 67.520 118.640 67.690 ;
        RECT 123.655 67.540 123.825 67.710 ;
        RECT 118.470 67.160 118.640 67.330 ;
        RECT 119.525 67.280 119.695 67.450 ;
        RECT 119.885 67.280 120.055 67.450 ;
        RECT 120.390 67.280 120.560 67.450 ;
        RECT 122.240 67.280 122.410 67.450 ;
        RECT 122.600 67.280 122.770 67.450 ;
        RECT 123.105 67.280 123.275 67.450 ;
        RECT 123.655 67.180 123.825 67.350 ;
        RECT 118.470 66.800 118.640 66.970 ;
        RECT 119.525 66.850 119.695 67.020 ;
        RECT 119.885 66.850 120.055 67.020 ;
        RECT 122.240 66.850 122.410 67.020 ;
        RECT 122.600 66.850 122.770 67.020 ;
        RECT 118.470 66.440 118.640 66.610 ;
        RECT 123.655 66.820 123.825 66.990 ;
        RECT 119.020 66.420 119.190 66.590 ;
        RECT 119.525 66.420 119.695 66.590 ;
        RECT 119.885 66.420 120.055 66.590 ;
        RECT 121.735 66.420 121.905 66.590 ;
        RECT 122.240 66.420 122.410 66.590 ;
        RECT 122.600 66.420 122.770 66.590 ;
        RECT 123.655 66.460 123.825 66.630 ;
        RECT 118.470 66.080 118.640 66.250 ;
        RECT 119.525 65.990 119.695 66.160 ;
        RECT 119.885 65.990 120.055 66.160 ;
        RECT 122.240 65.990 122.410 66.160 ;
        RECT 122.600 65.990 122.770 66.160 ;
        RECT 123.655 66.100 123.825 66.270 ;
        RECT 118.470 65.720 118.640 65.890 ;
        RECT 123.655 65.740 123.825 65.910 ;
        RECT 118.530 65.320 118.700 65.490 ;
        RECT 118.890 65.320 119.060 65.490 ;
        RECT 119.250 65.320 119.420 65.490 ;
        RECT 119.610 65.320 119.780 65.490 ;
        RECT 119.970 65.320 120.140 65.490 ;
        RECT 120.330 65.320 120.500 65.490 ;
        RECT 120.690 65.320 120.860 65.490 ;
        RECT 121.050 65.320 121.220 65.490 ;
        RECT 121.410 65.320 121.580 65.490 ;
        RECT 121.770 65.320 121.940 65.490 ;
        RECT 122.130 65.320 122.300 65.490 ;
        RECT 122.490 65.320 122.660 65.490 ;
        RECT 122.850 65.320 123.020 65.490 ;
        RECT 123.210 65.320 123.380 65.490 ;
        RECT 123.655 65.380 123.825 65.550 ;
        RECT 124.455 70.000 124.625 70.170 ;
        RECT 125.065 70.060 125.235 70.230 ;
        RECT 125.425 70.060 125.595 70.230 ;
        RECT 125.785 70.060 125.955 70.230 ;
        RECT 126.145 70.060 126.315 70.230 ;
        RECT 126.505 70.060 126.675 70.230 ;
        RECT 126.865 70.060 127.035 70.230 ;
        RECT 124.455 69.640 124.625 69.810 ;
        RECT 126.925 69.620 127.095 69.790 ;
        RECT 124.455 69.280 124.625 69.450 ;
        RECT 125.510 69.430 125.680 69.600 ;
        RECT 125.870 69.430 126.040 69.600 ;
        RECT 126.925 69.260 127.095 69.430 ;
        RECT 124.455 68.920 124.625 69.090 ;
        RECT 125.005 69.000 125.175 69.170 ;
        RECT 125.510 69.000 125.680 69.170 ;
        RECT 125.870 69.000 126.040 69.170 ;
        RECT 126.925 68.900 127.095 69.070 ;
        RECT 124.455 68.560 124.625 68.730 ;
        RECT 125.510 68.570 125.680 68.740 ;
        RECT 125.870 68.570 126.040 68.740 ;
        RECT 124.455 68.200 124.625 68.370 ;
        RECT 126.925 68.540 127.095 68.710 ;
        RECT 125.005 68.140 125.175 68.310 ;
        RECT 125.510 68.140 125.680 68.310 ;
        RECT 125.870 68.140 126.040 68.310 ;
        RECT 126.925 68.180 127.095 68.350 ;
        RECT 124.455 67.840 124.625 68.010 ;
        RECT 125.510 67.710 125.680 67.880 ;
        RECT 125.870 67.710 126.040 67.880 ;
        RECT 126.925 67.820 127.095 67.990 ;
        RECT 124.455 67.480 124.625 67.650 ;
        RECT 126.925 67.460 127.095 67.630 ;
        RECT 124.455 67.120 124.625 67.290 ;
        RECT 125.005 67.280 125.175 67.450 ;
        RECT 125.510 67.280 125.680 67.450 ;
        RECT 125.870 67.280 126.040 67.450 ;
        RECT 126.925 67.100 127.095 67.270 ;
        RECT 124.455 66.760 124.625 66.930 ;
        RECT 125.510 66.850 125.680 67.020 ;
        RECT 125.870 66.850 126.040 67.020 ;
        RECT 126.925 66.740 127.095 66.910 ;
        RECT 124.455 66.400 124.625 66.570 ;
        RECT 125.005 66.420 125.175 66.590 ;
        RECT 125.510 66.420 125.680 66.590 ;
        RECT 125.870 66.420 126.040 66.590 ;
        RECT 124.455 66.040 124.625 66.210 ;
        RECT 126.925 66.380 127.095 66.550 ;
        RECT 125.510 65.990 125.680 66.160 ;
        RECT 125.870 65.990 126.040 66.160 ;
        RECT 126.925 66.020 127.095 66.190 ;
        RECT 124.455 65.680 124.625 65.850 ;
        RECT 125.510 65.560 125.680 65.730 ;
        RECT 125.870 65.560 126.040 65.730 ;
        RECT 126.375 65.560 126.545 65.730 ;
        RECT 126.925 65.660 127.095 65.830 ;
        RECT 124.455 65.320 124.625 65.490 ;
        RECT 114.775 64.970 114.945 65.140 ;
        RECT 117.245 65.020 117.415 65.190 ;
        RECT 114.775 64.610 114.945 64.780 ;
        RECT 114.775 64.250 114.945 64.420 ;
        RECT 114.775 63.890 114.945 64.060 ;
        RECT 114.775 63.530 114.945 63.700 ;
        RECT 114.775 63.170 114.945 63.340 ;
        RECT 115.325 64.730 115.495 64.900 ;
        RECT 115.325 64.370 115.495 64.540 ;
        RECT 115.325 64.010 115.495 64.180 ;
        RECT 115.325 63.650 115.495 63.820 ;
        RECT 115.325 63.290 115.495 63.460 ;
        RECT 126.925 65.300 127.095 65.470 ;
        RECT 125.510 65.130 125.680 65.300 ;
        RECT 125.870 65.130 126.040 65.300 ;
        RECT 117.245 64.660 117.415 64.830 ;
        RECT 117.245 64.300 117.415 64.470 ;
        RECT 117.245 63.940 117.415 64.110 ;
        RECT 117.245 63.580 117.415 63.750 ;
        RECT 117.245 63.220 117.415 63.390 ;
        RECT 114.775 62.810 114.945 62.980 ;
        RECT 115.830 62.870 116.000 63.040 ;
        RECT 116.190 62.870 116.360 63.040 ;
        RECT 117.245 62.860 117.415 63.030 ;
        RECT 114.775 62.450 114.945 62.620 ;
        RECT 114.775 62.090 114.945 62.260 ;
        RECT 114.775 61.730 114.945 61.900 ;
        RECT 114.775 61.370 114.945 61.540 ;
        RECT 114.775 61.010 114.945 61.180 ;
        RECT 116.695 62.450 116.865 62.620 ;
        RECT 116.695 62.090 116.865 62.260 ;
        RECT 116.695 61.730 116.865 61.900 ;
        RECT 116.695 61.370 116.865 61.540 ;
        RECT 116.695 61.010 116.865 61.180 ;
        RECT 117.245 62.500 117.415 62.670 ;
        RECT 117.245 62.140 117.415 62.310 ;
        RECT 117.245 61.780 117.415 61.950 ;
        RECT 117.245 61.420 117.415 61.590 ;
        RECT 117.245 61.060 117.415 61.230 ;
        RECT 114.775 60.650 114.945 60.820 ;
        RECT 115.830 60.590 116.000 60.760 ;
        RECT 116.190 60.590 116.360 60.760 ;
        RECT 117.245 60.700 117.415 60.870 ;
        RECT 114.775 60.290 114.945 60.460 ;
        RECT 117.245 60.340 117.415 60.510 ;
        RECT 114.835 59.920 115.005 60.090 ;
        RECT 115.195 59.920 115.365 60.090 ;
        RECT 115.555 59.920 115.725 60.090 ;
        RECT 115.915 59.920 116.085 60.090 ;
        RECT 116.275 59.920 116.445 60.090 ;
        RECT 116.635 59.920 116.805 60.090 ;
        RECT 117.245 59.980 117.415 60.150 ;
        RECT 118.470 64.750 118.640 64.920 ;
        RECT 119.080 64.810 119.250 64.980 ;
        RECT 119.440 64.810 119.610 64.980 ;
        RECT 119.800 64.810 119.970 64.980 ;
        RECT 120.160 64.810 120.330 64.980 ;
        RECT 120.520 64.810 120.690 64.980 ;
        RECT 120.880 64.810 121.050 64.980 ;
        RECT 121.435 64.810 121.605 64.980 ;
        RECT 121.795 64.810 121.965 64.980 ;
        RECT 122.155 64.810 122.325 64.980 ;
        RECT 122.515 64.810 122.685 64.980 ;
        RECT 122.875 64.810 123.045 64.980 ;
        RECT 123.235 64.810 123.405 64.980 ;
        RECT 123.595 64.810 123.765 64.980 ;
        RECT 118.470 64.390 118.640 64.560 ;
        RECT 118.470 64.030 118.640 64.200 ;
        RECT 119.525 64.180 119.695 64.350 ;
        RECT 119.885 64.180 120.055 64.350 ;
        RECT 122.240 64.180 122.410 64.350 ;
        RECT 122.600 64.180 122.770 64.350 ;
        RECT 123.655 64.130 123.825 64.300 ;
        RECT 118.470 63.670 118.640 63.840 ;
        RECT 119.020 63.750 119.190 63.920 ;
        RECT 119.525 63.750 119.695 63.920 ;
        RECT 119.885 63.750 120.055 63.920 ;
        RECT 121.735 63.750 121.905 63.920 ;
        RECT 122.240 63.750 122.410 63.920 ;
        RECT 122.600 63.750 122.770 63.920 ;
        RECT 123.655 63.770 123.825 63.940 ;
        RECT 118.470 63.310 118.640 63.480 ;
        RECT 119.525 63.320 119.695 63.490 ;
        RECT 119.885 63.320 120.055 63.490 ;
        RECT 122.240 63.320 122.410 63.490 ;
        RECT 122.600 63.320 122.770 63.490 ;
        RECT 123.655 63.410 123.825 63.580 ;
        RECT 118.470 62.950 118.640 63.120 ;
        RECT 119.525 62.890 119.695 63.060 ;
        RECT 119.885 62.890 120.055 63.060 ;
        RECT 120.390 62.890 120.560 63.060 ;
        RECT 122.240 62.890 122.410 63.060 ;
        RECT 122.600 62.890 122.770 63.060 ;
        RECT 123.105 62.890 123.275 63.060 ;
        RECT 123.655 63.050 123.825 63.220 ;
        RECT 118.470 62.590 118.640 62.760 ;
        RECT 123.655 62.690 123.825 62.860 ;
        RECT 119.525 62.460 119.695 62.630 ;
        RECT 119.885 62.460 120.055 62.630 ;
        RECT 122.240 62.460 122.410 62.630 ;
        RECT 122.600 62.460 122.770 62.630 ;
        RECT 118.470 62.230 118.640 62.400 ;
        RECT 123.655 62.330 123.825 62.500 ;
        RECT 118.470 61.870 118.640 62.040 ;
        RECT 119.525 62.030 119.695 62.200 ;
        RECT 119.885 62.030 120.055 62.200 ;
        RECT 120.390 62.030 120.560 62.200 ;
        RECT 122.240 62.030 122.410 62.200 ;
        RECT 122.600 62.030 122.770 62.200 ;
        RECT 123.105 62.030 123.275 62.200 ;
        RECT 123.655 61.970 123.825 62.140 ;
        RECT 118.470 61.510 118.640 61.680 ;
        RECT 119.525 61.600 119.695 61.770 ;
        RECT 119.885 61.600 120.055 61.770 ;
        RECT 122.240 61.600 122.410 61.770 ;
        RECT 122.600 61.600 122.770 61.770 ;
        RECT 123.655 61.610 123.825 61.780 ;
        RECT 118.470 61.150 118.640 61.320 ;
        RECT 119.020 61.170 119.190 61.340 ;
        RECT 119.525 61.170 119.695 61.340 ;
        RECT 119.885 61.170 120.055 61.340 ;
        RECT 121.735 61.170 121.905 61.340 ;
        RECT 122.240 61.170 122.410 61.340 ;
        RECT 122.600 61.170 122.770 61.340 ;
        RECT 123.655 61.250 123.825 61.420 ;
        RECT 118.470 60.790 118.640 60.960 ;
        RECT 119.525 60.740 119.695 60.910 ;
        RECT 119.885 60.740 120.055 60.910 ;
        RECT 122.240 60.740 122.410 60.910 ;
        RECT 122.600 60.740 122.770 60.910 ;
        RECT 123.655 60.890 123.825 61.060 ;
        RECT 123.655 60.530 123.825 60.700 ;
        RECT 118.530 60.110 118.700 60.280 ;
        RECT 118.890 60.110 119.060 60.280 ;
        RECT 119.250 60.110 119.420 60.280 ;
        RECT 119.610 60.110 119.780 60.280 ;
        RECT 119.970 60.110 120.140 60.280 ;
        RECT 120.330 60.110 120.500 60.280 ;
        RECT 120.690 60.110 120.860 60.280 ;
        RECT 121.050 60.110 121.220 60.280 ;
        RECT 121.410 60.110 121.580 60.280 ;
        RECT 121.770 60.110 121.940 60.280 ;
        RECT 122.130 60.110 122.300 60.280 ;
        RECT 122.490 60.110 122.660 60.280 ;
        RECT 122.850 60.110 123.020 60.280 ;
        RECT 123.210 60.110 123.380 60.280 ;
        RECT 123.655 60.170 123.825 60.340 ;
        RECT 124.455 64.950 124.625 65.120 ;
        RECT 126.925 64.940 127.095 65.110 ;
        RECT 124.455 64.590 124.625 64.760 ;
        RECT 125.510 64.700 125.680 64.870 ;
        RECT 125.870 64.700 126.040 64.870 ;
        RECT 126.375 64.700 126.545 64.870 ;
        RECT 126.925 64.580 127.095 64.750 ;
        RECT 124.455 64.230 124.625 64.400 ;
        RECT 125.510 64.270 125.680 64.440 ;
        RECT 125.870 64.270 126.040 64.440 ;
        RECT 124.455 63.870 124.625 64.040 ;
        RECT 126.925 64.220 127.095 64.390 ;
        RECT 125.005 63.840 125.175 64.010 ;
        RECT 125.510 63.840 125.680 64.010 ;
        RECT 125.870 63.840 126.040 64.010 ;
        RECT 126.925 63.860 127.095 64.030 ;
        RECT 124.455 63.510 124.625 63.680 ;
        RECT 125.510 63.410 125.680 63.580 ;
        RECT 125.870 63.410 126.040 63.580 ;
        RECT 126.925 63.500 127.095 63.670 ;
        RECT 124.455 63.150 124.625 63.320 ;
        RECT 125.005 62.980 125.175 63.150 ;
        RECT 125.510 62.980 125.680 63.150 ;
        RECT 125.870 62.980 126.040 63.150 ;
        RECT 126.925 63.140 127.095 63.310 ;
        RECT 124.455 62.790 124.625 62.960 ;
        RECT 126.925 62.780 127.095 62.950 ;
        RECT 124.455 62.430 124.625 62.600 ;
        RECT 125.510 62.550 125.680 62.720 ;
        RECT 125.870 62.550 126.040 62.720 ;
        RECT 126.925 62.420 127.095 62.590 ;
        RECT 124.455 62.070 124.625 62.240 ;
        RECT 125.005 62.120 125.175 62.290 ;
        RECT 125.510 62.120 125.680 62.290 ;
        RECT 125.870 62.120 126.040 62.290 ;
        RECT 124.455 61.710 124.625 61.880 ;
        RECT 126.925 62.060 127.095 62.230 ;
        RECT 125.510 61.690 125.680 61.860 ;
        RECT 125.870 61.690 126.040 61.860 ;
        RECT 126.925 61.700 127.095 61.870 ;
        RECT 124.455 61.350 124.625 61.520 ;
        RECT 125.005 61.260 125.175 61.430 ;
        RECT 125.510 61.260 125.680 61.430 ;
        RECT 125.870 61.260 126.040 61.430 ;
        RECT 126.925 61.340 127.095 61.510 ;
        RECT 124.455 60.990 124.625 61.160 ;
        RECT 125.510 60.830 125.680 61.000 ;
        RECT 125.870 60.830 126.040 61.000 ;
        RECT 126.925 60.980 127.095 61.150 ;
        RECT 124.455 60.630 124.625 60.800 ;
        RECT 126.925 60.620 127.095 60.790 ;
        RECT 124.515 60.200 124.685 60.370 ;
        RECT 124.875 60.200 125.045 60.370 ;
        RECT 125.235 60.200 125.405 60.370 ;
        RECT 125.595 60.200 125.765 60.370 ;
        RECT 125.955 60.200 126.125 60.370 ;
        RECT 126.315 60.200 126.485 60.370 ;
        RECT 126.925 60.260 127.095 60.430 ;
      LAYER met1 ;
        RECT 107.530 173.590 110.225 173.880 ;
        RECT 110.515 173.590 114.235 173.880 ;
        RECT 107.530 169.100 107.820 173.590 ;
        RECT 108.195 172.935 109.195 173.195 ;
        RECT 108.195 172.505 109.195 172.765 ;
        RECT 109.385 172.340 109.675 173.590 ;
        RECT 108.195 172.075 109.195 172.335 ;
        RECT 108.195 171.645 109.195 171.905 ;
        RECT 109.385 171.510 109.675 172.070 ;
        RECT 110.205 171.510 110.535 173.185 ;
        RECT 111.065 172.340 111.355 173.590 ;
        RECT 112.045 173.180 113.045 173.195 ;
        RECT 111.545 172.950 113.545 173.180 ;
        RECT 112.045 172.935 113.045 172.950 ;
        RECT 112.045 172.750 113.045 172.765 ;
        RECT 111.545 172.520 113.545 172.750 ;
        RECT 112.045 172.505 113.045 172.520 ;
        RECT 112.045 172.320 113.045 172.335 ;
        RECT 111.545 172.090 113.545 172.320 ;
        RECT 112.045 172.075 113.045 172.090 ;
        RECT 111.065 171.510 111.355 172.070 ;
        RECT 111.545 171.645 113.545 171.905 ;
        RECT 108.195 171.215 109.195 171.475 ;
        RECT 109.385 171.180 111.355 171.510 ;
        RECT 112.045 171.460 113.045 171.475 ;
        RECT 111.545 171.230 113.545 171.460 ;
        RECT 112.045 171.215 113.045 171.230 ;
        RECT 108.195 170.785 109.195 171.045 ;
        RECT 109.385 170.620 109.675 171.180 ;
        RECT 111.065 170.620 111.355 171.180 ;
        RECT 111.545 170.785 113.545 171.045 ;
        RECT 108.195 170.355 109.195 170.615 ;
        RECT 112.045 170.600 113.045 170.615 ;
        RECT 111.545 170.370 113.545 170.600 ;
        RECT 112.045 170.355 113.045 170.370 ;
        RECT 108.195 169.925 109.195 170.185 ;
        RECT 108.195 169.495 109.195 169.755 ;
        RECT 109.385 169.100 109.675 170.350 ;
        RECT 111.065 169.100 111.355 170.350 ;
        RECT 112.045 170.170 113.045 170.185 ;
        RECT 111.545 169.940 113.545 170.170 ;
        RECT 112.045 169.925 113.045 169.940 ;
        RECT 112.045 169.740 113.045 169.755 ;
        RECT 111.545 169.510 113.545 169.740 ;
        RECT 112.045 169.495 113.045 169.510 ;
        RECT 113.945 169.100 114.235 173.590 ;
        RECT 107.530 168.810 110.225 169.100 ;
        RECT 110.515 168.810 114.235 169.100 ;
        RECT 108.575 164.440 114.075 164.730 ;
        RECT 56.120 151.190 62.770 151.480 ;
        RECT 56.120 111.980 56.410 151.190 ;
        RECT 57.150 141.295 58.150 141.555 ;
        RECT 57.150 139.015 58.150 139.275 ;
        RECT 57.150 136.735 58.150 136.995 ;
        RECT 57.150 134.455 58.150 134.715 ;
        RECT 57.150 132.175 58.150 132.435 ;
        RECT 58.340 130.330 58.630 151.190 ;
        RECT 60.260 149.410 60.550 151.190 ;
        RECT 60.740 150.535 61.740 150.795 ;
        RECT 60.740 149.755 61.740 150.015 ;
        RECT 60.740 148.975 61.740 149.235 ;
        RECT 60.740 146.695 61.740 146.955 ;
        RECT 61.930 144.850 62.260 148.800 ;
        RECT 60.740 144.415 61.740 144.675 ;
        RECT 60.260 143.910 60.550 144.240 ;
        RECT 60.260 143.620 61.740 143.910 ;
        RECT 60.260 143.130 60.550 143.620 ;
        RECT 60.260 142.840 61.740 143.130 ;
        RECT 60.260 142.350 60.550 142.840 ;
        RECT 60.260 142.060 61.740 142.350 ;
        RECT 60.260 141.730 60.550 142.060 ;
        RECT 60.740 141.295 61.740 141.555 ;
        RECT 60.260 139.450 60.550 141.120 ;
        RECT 60.740 139.015 61.740 139.275 ;
        RECT 60.260 137.170 60.550 138.840 ;
        RECT 60.740 136.735 61.740 136.995 ;
        RECT 60.260 134.890 60.550 136.560 ;
        RECT 60.740 134.455 61.740 134.715 ;
        RECT 60.260 132.610 60.550 134.280 ;
        RECT 60.740 132.175 61.740 132.435 ;
        RECT 60.260 130.330 60.550 132.000 ;
        RECT 57.150 129.895 58.150 130.155 ;
        RECT 60.740 129.895 61.740 130.155 ;
        RECT 56.630 125.770 56.960 129.720 ;
        RECT 60.260 128.050 60.550 129.720 ;
        RECT 61.930 128.050 62.260 141.120 ;
        RECT 57.150 127.615 58.150 127.875 ;
        RECT 60.740 127.615 61.740 127.875 ;
        RECT 60.260 125.770 60.550 127.440 ;
        RECT 57.150 125.335 58.150 125.595 ;
        RECT 60.740 125.335 61.740 125.595 ;
        RECT 57.150 123.055 58.150 123.315 ;
        RECT 57.150 120.775 58.150 121.035 ;
        RECT 57.150 118.495 58.150 118.755 ;
        RECT 57.150 116.215 58.150 116.475 ;
        RECT 57.150 113.935 58.150 114.195 ;
        RECT 58.340 111.980 58.630 125.160 ;
        RECT 60.260 123.490 60.550 125.160 ;
        RECT 60.740 123.055 61.740 123.315 ;
        RECT 60.260 121.210 60.550 122.880 ;
        RECT 60.740 120.775 61.740 121.035 ;
        RECT 60.260 118.930 60.550 120.600 ;
        RECT 60.740 118.495 61.740 118.755 ;
        RECT 60.260 116.650 60.550 118.320 ;
        RECT 60.740 116.215 61.740 116.475 ;
        RECT 60.260 114.370 60.550 116.040 ;
        RECT 61.930 114.370 62.260 127.440 ;
        RECT 60.740 113.935 61.740 114.195 ;
        RECT 60.260 111.980 60.550 113.760 ;
        RECT 60.740 113.155 61.740 113.415 ;
        RECT 60.740 112.375 61.740 112.635 ;
        RECT 62.480 111.980 62.770 151.190 ;
        RECT 64.375 151.190 66.935 151.480 ;
        RECT 64.375 142.460 64.665 151.190 ;
        RECT 65.405 150.535 65.905 150.795 ;
        RECT 65.405 149.755 65.905 150.015 ;
        RECT 66.095 149.410 66.385 151.190 ;
        RECT 65.405 148.975 65.905 149.235 ;
        RECT 64.885 144.850 65.215 148.800 ;
        RECT 65.405 146.695 65.905 146.955 ;
        RECT 65.405 144.415 65.905 144.675 ;
        RECT 65.405 143.635 65.905 143.895 ;
        RECT 65.405 142.855 65.905 143.115 ;
        RECT 66.095 142.460 66.385 144.240 ;
        RECT 66.645 142.460 66.935 151.190 ;
        RECT 91.855 151.190 94.415 151.480 ;
        RECT 64.375 142.170 66.935 142.460 ;
        RECT 72.530 142.470 77.830 142.760 ;
        RECT 64.375 137.980 66.935 138.270 ;
        RECT 64.375 117.570 64.665 137.980 ;
        RECT 64.925 135.155 65.215 137.980 ;
        RECT 65.405 137.325 65.905 137.585 ;
        RECT 66.075 137.185 66.365 137.980 ;
        RECT 65.405 136.045 65.905 136.305 ;
        RECT 66.075 135.155 66.385 137.185 ;
        RECT 65.405 134.765 65.905 135.025 ;
        RECT 64.885 132.765 65.215 134.725 ;
        RECT 66.095 132.765 66.425 134.590 ;
        RECT 64.885 132.475 66.425 132.765 ;
        RECT 64.885 130.640 65.215 132.475 ;
        RECT 66.095 130.640 66.425 132.475 ;
        RECT 65.405 130.205 65.905 130.465 ;
        RECT 64.925 129.195 65.215 130.065 ;
        RECT 66.075 129.195 66.385 130.065 ;
        RECT 64.925 128.915 66.385 129.195 ;
        RECT 64.925 127.915 65.215 128.915 ;
        RECT 66.075 128.035 66.385 128.915 ;
        RECT 66.075 127.915 66.365 128.035 ;
        RECT 64.925 127.635 66.365 127.915 ;
        RECT 64.925 126.635 65.215 127.635 ;
        RECT 66.075 127.505 66.365 127.635 ;
        RECT 66.075 126.635 66.385 127.505 ;
        RECT 64.925 126.355 66.385 126.635 ;
        RECT 64.925 125.475 65.215 126.355 ;
        RECT 66.075 125.475 66.385 126.355 ;
        RECT 65.405 125.085 65.905 125.345 ;
        RECT 64.880 123.240 65.215 124.910 ;
        RECT 64.880 122.630 65.210 123.240 ;
        RECT 65.405 122.805 65.905 123.065 ;
        RECT 64.880 120.960 65.215 122.630 ;
        RECT 65.405 120.525 65.905 120.785 ;
        RECT 64.925 117.570 65.215 120.385 ;
        RECT 65.405 119.245 65.905 119.505 ;
        RECT 66.075 118.355 66.385 120.385 ;
        RECT 65.405 117.965 65.905 118.225 ;
        RECT 66.075 117.570 66.365 118.355 ;
        RECT 66.645 117.570 66.935 137.980 ;
        RECT 64.375 117.280 66.935 117.570 ;
        RECT 68.130 137.980 71.190 138.270 ;
        RECT 68.130 117.570 68.420 137.980 ;
        RECT 68.700 137.185 68.990 137.980 ;
        RECT 69.160 137.325 70.160 137.585 ;
        RECT 68.680 135.155 68.990 137.185 ;
        RECT 70.330 137.185 70.620 137.980 ;
        RECT 69.160 136.045 70.160 136.305 ;
        RECT 70.330 135.155 70.640 137.185 ;
        RECT 69.160 134.765 70.160 135.025 ;
        RECT 68.640 130.640 68.970 134.590 ;
        RECT 70.330 132.730 70.660 134.590 ;
        RECT 69.160 132.465 70.660 132.730 ;
        RECT 70.330 130.640 70.660 132.465 ;
        RECT 69.160 130.205 70.160 130.465 ;
        RECT 68.680 129.195 68.990 130.065 ;
        RECT 70.330 129.195 70.640 130.065 ;
        RECT 68.680 128.915 70.640 129.195 ;
        RECT 68.680 128.035 68.990 128.915 ;
        RECT 68.700 127.915 68.990 128.035 ;
        RECT 70.330 128.035 70.640 128.915 ;
        RECT 70.330 127.915 70.620 128.035 ;
        RECT 68.700 127.635 70.620 127.915 ;
        RECT 68.700 127.505 68.990 127.635 ;
        RECT 68.680 126.635 68.990 127.505 ;
        RECT 70.330 127.505 70.620 127.635 ;
        RECT 70.330 126.635 70.640 127.505 ;
        RECT 68.680 126.355 70.640 126.635 ;
        RECT 68.680 125.475 68.990 126.355 ;
        RECT 70.330 125.475 70.640 126.355 ;
        RECT 69.160 125.085 70.160 125.345 ;
        RECT 70.330 123.050 70.660 124.910 ;
        RECT 69.160 122.775 70.660 123.050 ;
        RECT 70.330 120.960 70.660 122.775 ;
        RECT 69.160 120.525 70.160 120.785 ;
        RECT 68.680 118.355 68.990 120.385 ;
        RECT 69.160 119.245 70.160 119.505 ;
        RECT 68.700 117.570 68.990 118.355 ;
        RECT 70.330 118.355 70.640 120.385 ;
        RECT 69.160 117.965 70.160 118.225 ;
        RECT 70.330 117.570 70.620 118.355 ;
        RECT 70.900 117.570 71.190 137.980 ;
        RECT 68.130 117.280 71.190 117.570 ;
        RECT 56.120 111.690 62.770 111.980 ;
        RECT 63.625 113.030 67.345 113.320 ;
        RECT 67.610 113.030 70.305 113.320 ;
        RECT 63.625 89.180 63.915 113.030 ;
        RECT 64.315 112.375 65.315 112.635 ;
        RECT 64.315 110.095 65.315 110.355 ;
        RECT 65.505 108.250 65.795 113.030 ;
        RECT 68.635 108.250 68.925 113.030 ;
        RECT 69.115 112.375 69.615 112.635 ;
        RECT 69.115 110.095 69.615 110.355 ;
        RECT 64.315 107.815 65.315 108.075 ;
        RECT 69.115 107.815 69.615 108.075 ;
        RECT 64.315 105.535 65.315 105.795 ;
        RECT 65.505 103.690 65.835 107.640 ;
        RECT 67.025 105.525 67.985 105.805 ;
        RECT 64.315 103.255 65.315 103.515 ;
        RECT 67.340 103.080 67.670 105.525 ;
        RECT 68.595 103.690 68.925 107.640 ;
        RECT 69.115 105.535 69.615 105.795 ;
        RECT 69.115 103.255 69.615 103.515 ;
        RECT 65.505 102.750 68.925 103.080 ;
        RECT 64.315 100.975 65.315 101.235 ;
        RECT 65.505 99.130 65.835 102.750 ;
        RECT 67.025 100.965 67.985 101.245 ;
        RECT 64.315 98.695 65.315 98.955 ;
        RECT 67.340 98.520 67.670 100.965 ;
        RECT 68.595 99.130 68.925 102.750 ;
        RECT 69.115 100.975 69.615 101.235 ;
        RECT 69.115 98.695 69.615 98.955 ;
        RECT 65.505 98.190 68.925 98.520 ;
        RECT 64.315 96.415 65.315 96.675 ;
        RECT 65.505 94.570 65.835 98.190 ;
        RECT 68.595 94.570 68.925 98.190 ;
        RECT 69.115 96.415 69.615 96.675 ;
        RECT 64.315 94.135 65.315 94.395 ;
        RECT 69.115 94.135 69.615 94.395 ;
        RECT 64.315 91.855 65.315 92.115 ;
        RECT 64.315 89.575 65.315 89.835 ;
        RECT 65.505 89.180 65.795 93.960 ;
        RECT 68.635 89.180 68.925 93.960 ;
        RECT 69.115 91.855 69.615 92.115 ;
        RECT 69.115 89.575 69.615 89.835 ;
        RECT 70.015 89.180 70.305 113.030 ;
        RECT 72.530 113.020 72.820 142.470 ;
        RECT 73.560 141.855 74.060 142.115 ;
        RECT 73.040 130.610 73.370 141.120 ;
        RECT 74.250 140.820 74.540 142.470 ;
        RECT 73.560 140.590 74.540 140.820 ;
        RECT 74.250 139.685 74.540 140.590 ;
        RECT 73.560 139.295 74.060 139.555 ;
        RECT 74.250 137.450 74.540 139.120 ;
        RECT 73.560 137.015 74.060 137.275 ;
        RECT 74.250 135.170 74.540 136.840 ;
        RECT 75.820 135.285 76.110 142.470 ;
        RECT 76.300 141.455 76.800 141.715 ;
        RECT 76.300 138.175 76.800 138.435 ;
        RECT 76.990 135.285 77.280 142.470 ;
        RECT 73.560 134.735 74.060 134.995 ;
        RECT 76.300 134.895 76.800 135.155 ;
        RECT 74.250 132.890 74.540 134.560 ;
        RECT 73.560 132.455 74.060 132.715 ;
        RECT 74.250 130.610 74.540 132.280 ;
        RECT 73.560 130.175 74.060 130.435 ;
        RECT 73.080 129.165 73.370 130.035 ;
        RECT 74.250 129.165 74.540 130.035 ;
        RECT 73.080 128.885 74.540 129.165 ;
        RECT 73.080 127.885 73.370 128.885 ;
        RECT 74.250 127.885 74.540 128.885 ;
        RECT 73.080 127.605 74.540 127.885 ;
        RECT 76.300 127.615 76.800 127.875 ;
        RECT 73.080 126.605 73.370 127.605 ;
        RECT 74.250 126.605 74.540 127.605 ;
        RECT 73.080 126.325 74.540 126.605 ;
        RECT 73.080 125.445 73.370 126.325 ;
        RECT 74.250 125.445 74.540 126.325 ;
        RECT 73.560 125.055 74.060 125.315 ;
        RECT 73.040 114.370 73.370 124.880 ;
        RECT 74.250 123.210 74.540 124.880 ;
        RECT 73.560 122.775 74.060 123.035 ;
        RECT 74.250 120.930 74.540 122.600 ;
        RECT 73.560 120.495 74.060 120.755 ;
        RECT 76.990 120.750 77.320 134.740 ;
        RECT 76.300 120.335 76.800 120.595 ;
        RECT 74.250 118.650 74.540 120.320 ;
        RECT 73.560 118.215 74.060 118.475 ;
        RECT 74.250 116.370 74.540 118.040 ;
        RECT 73.560 115.935 74.060 116.195 ;
        RECT 74.250 114.900 74.540 115.795 ;
        RECT 73.560 114.670 74.540 114.900 ;
        RECT 73.560 113.375 74.060 113.635 ;
        RECT 74.250 113.020 74.540 114.670 ;
        RECT 75.820 113.020 76.110 120.195 ;
        RECT 76.300 117.055 76.800 117.315 ;
        RECT 76.300 113.775 76.800 114.035 ;
        RECT 76.990 113.020 77.280 120.195 ;
        RECT 77.540 113.020 77.830 142.470 ;
        RECT 72.530 112.730 77.830 113.020 ;
        RECT 80.960 142.470 86.260 142.760 ;
        RECT 80.960 113.020 81.250 142.470 ;
        RECT 81.510 135.285 81.800 142.470 ;
        RECT 81.990 141.455 82.490 141.715 ;
        RECT 81.990 138.175 82.490 138.435 ;
        RECT 82.680 135.285 82.970 142.470 ;
        RECT 84.250 140.820 84.540 142.470 ;
        RECT 84.730 141.855 85.230 142.115 ;
        RECT 84.250 140.590 85.230 140.820 ;
        RECT 84.250 139.685 84.540 140.590 ;
        RECT 84.730 139.295 85.230 139.555 ;
        RECT 84.250 137.450 84.540 139.120 ;
        RECT 84.730 137.015 85.230 137.275 ;
        RECT 84.250 135.170 84.540 136.840 ;
        RECT 81.990 134.895 82.490 135.155 ;
        RECT 81.470 120.750 81.800 134.740 ;
        RECT 84.730 134.735 85.230 134.995 ;
        RECT 84.250 132.890 84.540 134.560 ;
        RECT 84.730 132.455 85.230 132.715 ;
        RECT 84.250 130.610 84.540 132.280 ;
        RECT 85.420 130.610 85.750 141.120 ;
        RECT 84.730 130.175 85.230 130.435 ;
        RECT 84.250 129.165 84.540 130.035 ;
        RECT 85.420 129.165 85.710 130.035 ;
        RECT 84.250 128.885 85.710 129.165 ;
        RECT 84.250 127.885 84.540 128.885 ;
        RECT 85.420 127.885 85.710 128.885 ;
        RECT 81.990 127.615 82.490 127.875 ;
        RECT 84.250 127.605 85.710 127.885 ;
        RECT 84.250 126.605 84.540 127.605 ;
        RECT 85.420 126.605 85.710 127.605 ;
        RECT 84.250 126.325 85.710 126.605 ;
        RECT 84.250 125.445 84.540 126.325 ;
        RECT 85.420 125.445 85.710 126.325 ;
        RECT 84.730 125.055 85.230 125.315 ;
        RECT 84.250 123.210 84.540 124.880 ;
        RECT 84.730 122.775 85.230 123.035 ;
        RECT 84.250 120.930 84.540 122.600 ;
        RECT 81.990 120.335 82.490 120.595 ;
        RECT 84.730 120.495 85.230 120.755 ;
        RECT 81.510 113.020 81.800 120.195 ;
        RECT 81.990 117.055 82.490 117.315 ;
        RECT 81.990 113.775 82.490 114.035 ;
        RECT 82.680 113.020 82.970 120.195 ;
        RECT 84.250 118.650 84.540 120.320 ;
        RECT 84.730 118.215 85.230 118.475 ;
        RECT 84.250 116.370 84.540 118.040 ;
        RECT 84.730 115.935 85.230 116.195 ;
        RECT 84.250 114.900 84.540 115.795 ;
        RECT 84.250 114.670 85.230 114.900 ;
        RECT 84.250 113.020 84.540 114.670 ;
        RECT 85.420 114.370 85.750 124.880 ;
        RECT 84.730 113.375 85.230 113.635 ;
        RECT 85.970 113.020 86.260 142.470 ;
        RECT 91.855 142.460 92.145 151.190 ;
        RECT 92.405 149.410 92.695 151.190 ;
        RECT 92.885 150.535 93.385 150.795 ;
        RECT 92.885 149.755 93.385 150.015 ;
        RECT 92.885 148.975 93.385 149.235 ;
        RECT 92.885 146.695 93.385 146.955 ;
        RECT 93.575 144.850 93.905 148.800 ;
        RECT 92.885 144.415 93.385 144.675 ;
        RECT 92.405 142.460 92.695 144.240 ;
        RECT 92.885 143.635 93.385 143.895 ;
        RECT 92.885 142.855 93.385 143.115 ;
        RECT 94.125 142.460 94.415 151.190 ;
        RECT 91.855 142.170 94.415 142.460 ;
        RECT 96.020 151.190 102.670 151.480 ;
        RECT 87.600 137.980 90.660 138.270 ;
        RECT 87.600 117.570 87.890 137.980 ;
        RECT 88.170 137.185 88.460 137.980 ;
        RECT 88.630 137.325 89.630 137.585 ;
        RECT 88.150 135.155 88.460 137.185 ;
        RECT 89.800 137.185 90.090 137.980 ;
        RECT 88.630 136.045 89.630 136.305 ;
        RECT 89.800 135.155 90.110 137.185 ;
        RECT 88.630 134.765 89.630 135.025 ;
        RECT 88.130 132.730 88.460 134.590 ;
        RECT 88.130 132.465 89.630 132.730 ;
        RECT 88.130 130.640 88.460 132.465 ;
        RECT 89.820 130.640 90.150 134.590 ;
        RECT 88.630 130.205 89.630 130.465 ;
        RECT 88.150 129.195 88.460 130.065 ;
        RECT 89.800 129.195 90.110 130.065 ;
        RECT 88.150 128.915 90.110 129.195 ;
        RECT 88.150 128.035 88.460 128.915 ;
        RECT 88.170 127.915 88.460 128.035 ;
        RECT 89.800 128.035 90.110 128.915 ;
        RECT 89.800 127.915 90.090 128.035 ;
        RECT 88.170 127.635 90.090 127.915 ;
        RECT 88.170 127.505 88.460 127.635 ;
        RECT 88.150 126.635 88.460 127.505 ;
        RECT 89.800 127.505 90.090 127.635 ;
        RECT 89.800 126.635 90.110 127.505 ;
        RECT 88.150 126.355 90.110 126.635 ;
        RECT 88.150 125.475 88.460 126.355 ;
        RECT 89.800 125.475 90.110 126.355 ;
        RECT 88.630 125.085 89.630 125.345 ;
        RECT 88.130 123.050 88.460 124.910 ;
        RECT 88.130 122.775 89.630 123.050 ;
        RECT 88.130 120.960 88.460 122.775 ;
        RECT 88.630 120.525 89.630 120.785 ;
        RECT 88.150 118.355 88.460 120.385 ;
        RECT 88.630 119.245 89.630 119.505 ;
        RECT 88.170 117.570 88.460 118.355 ;
        RECT 89.800 118.355 90.110 120.385 ;
        RECT 88.630 117.965 89.630 118.225 ;
        RECT 89.800 117.570 90.090 118.355 ;
        RECT 90.370 117.570 90.660 137.980 ;
        RECT 87.600 117.280 90.660 117.570 ;
        RECT 91.855 137.980 94.415 138.270 ;
        RECT 91.855 117.570 92.145 137.980 ;
        RECT 92.425 137.185 92.715 137.980 ;
        RECT 92.885 137.325 93.385 137.585 ;
        RECT 92.405 135.155 92.715 137.185 ;
        RECT 92.885 136.045 93.385 136.305 ;
        RECT 93.575 135.155 93.865 137.980 ;
        RECT 92.885 134.765 93.385 135.025 ;
        RECT 92.365 132.765 92.695 134.590 ;
        RECT 93.575 132.765 93.905 134.725 ;
        RECT 92.365 132.475 93.905 132.765 ;
        RECT 92.365 130.640 92.695 132.475 ;
        RECT 93.575 130.640 93.905 132.475 ;
        RECT 92.885 130.205 93.385 130.465 ;
        RECT 92.405 129.195 92.715 130.065 ;
        RECT 93.575 129.195 93.865 130.065 ;
        RECT 92.405 128.915 93.865 129.195 ;
        RECT 92.405 128.035 92.715 128.915 ;
        RECT 92.425 127.915 92.715 128.035 ;
        RECT 93.575 127.915 93.865 128.915 ;
        RECT 92.425 127.635 93.865 127.915 ;
        RECT 92.425 127.505 92.715 127.635 ;
        RECT 92.405 126.635 92.715 127.505 ;
        RECT 93.575 126.635 93.865 127.635 ;
        RECT 92.405 126.355 93.865 126.635 ;
        RECT 92.405 125.475 92.715 126.355 ;
        RECT 93.575 125.475 93.865 126.355 ;
        RECT 92.885 125.085 93.385 125.345 ;
        RECT 93.575 123.240 93.910 124.910 ;
        RECT 92.885 122.805 93.385 123.065 ;
        RECT 93.580 122.630 93.910 123.240 ;
        RECT 93.575 120.960 93.910 122.630 ;
        RECT 92.885 120.525 93.385 120.785 ;
        RECT 92.405 118.355 92.715 120.385 ;
        RECT 92.885 119.245 93.385 119.505 ;
        RECT 92.425 117.570 92.715 118.355 ;
        RECT 92.885 117.965 93.385 118.225 ;
        RECT 93.575 117.570 93.865 120.385 ;
        RECT 94.125 117.570 94.415 137.980 ;
        RECT 91.855 117.280 94.415 117.570 ;
        RECT 80.960 112.730 86.260 113.020 ;
        RECT 88.485 113.030 91.180 113.320 ;
        RECT 91.445 113.030 95.165 113.320 ;
        RECT 63.625 88.890 67.345 89.180 ;
        RECT 67.610 88.890 70.305 89.180 ;
        RECT 88.485 89.180 88.775 113.030 ;
        RECT 89.175 112.375 89.675 112.635 ;
        RECT 89.175 110.095 89.675 110.355 ;
        RECT 89.865 108.250 90.155 113.030 ;
        RECT 92.995 108.250 93.285 113.030 ;
        RECT 93.475 112.375 94.475 112.635 ;
        RECT 93.475 110.095 94.475 110.355 ;
        RECT 89.175 107.815 89.675 108.075 ;
        RECT 93.475 107.815 94.475 108.075 ;
        RECT 89.175 105.535 89.675 105.795 ;
        RECT 89.865 103.690 90.195 107.640 ;
        RECT 90.805 105.525 91.765 105.805 ;
        RECT 89.175 103.255 89.675 103.515 ;
        RECT 91.120 103.080 91.450 105.525 ;
        RECT 92.955 103.690 93.285 107.640 ;
        RECT 93.475 105.535 94.475 105.795 ;
        RECT 93.475 103.255 94.475 103.515 ;
        RECT 89.865 102.750 93.285 103.080 ;
        RECT 89.175 100.975 89.675 101.235 ;
        RECT 89.865 99.130 90.195 102.750 ;
        RECT 90.805 100.965 91.765 101.245 ;
        RECT 89.175 98.695 89.675 98.955 ;
        RECT 91.120 98.520 91.450 100.965 ;
        RECT 92.955 99.130 93.285 102.750 ;
        RECT 93.475 100.975 94.475 101.235 ;
        RECT 93.475 98.695 94.475 98.955 ;
        RECT 89.865 98.190 93.285 98.520 ;
        RECT 89.175 96.415 89.675 96.675 ;
        RECT 89.865 94.570 90.195 98.190 ;
        RECT 92.955 94.570 93.285 98.190 ;
        RECT 93.475 96.415 94.475 96.675 ;
        RECT 89.175 94.135 89.675 94.395 ;
        RECT 93.475 94.135 94.475 94.395 ;
        RECT 89.175 91.855 89.675 92.115 ;
        RECT 89.175 89.575 89.675 89.835 ;
        RECT 89.865 89.180 90.155 93.960 ;
        RECT 92.995 89.180 93.285 93.960 ;
        RECT 93.475 91.855 94.475 92.115 ;
        RECT 93.475 89.575 94.475 89.835 ;
        RECT 94.875 89.180 95.165 113.030 ;
        RECT 96.020 111.980 96.310 151.190 ;
        RECT 97.050 150.535 98.050 150.795 ;
        RECT 97.050 149.755 98.050 150.015 ;
        RECT 98.240 149.410 98.530 151.190 ;
        RECT 97.050 148.975 98.050 149.235 ;
        RECT 96.530 144.850 96.860 148.800 ;
        RECT 97.050 146.695 98.050 146.955 ;
        RECT 97.050 144.415 98.050 144.675 ;
        RECT 98.240 143.910 98.530 144.240 ;
        RECT 97.050 143.620 98.530 143.910 ;
        RECT 98.240 143.130 98.530 143.620 ;
        RECT 97.050 142.840 98.530 143.130 ;
        RECT 98.240 142.350 98.530 142.840 ;
        RECT 97.050 142.060 98.530 142.350 ;
        RECT 98.240 141.730 98.530 142.060 ;
        RECT 97.050 141.295 98.050 141.555 ;
        RECT 96.530 128.050 96.860 141.120 ;
        RECT 98.240 139.450 98.530 141.120 ;
        RECT 97.050 139.015 98.050 139.275 ;
        RECT 98.240 137.170 98.530 138.840 ;
        RECT 97.050 136.735 98.050 136.995 ;
        RECT 98.240 134.890 98.530 136.560 ;
        RECT 97.050 134.455 98.050 134.715 ;
        RECT 98.240 132.610 98.530 134.280 ;
        RECT 97.050 132.175 98.050 132.435 ;
        RECT 98.240 130.330 98.530 132.000 ;
        RECT 100.160 130.330 100.450 151.190 ;
        RECT 100.640 141.295 101.640 141.555 ;
        RECT 100.640 139.015 101.640 139.275 ;
        RECT 100.640 136.735 101.640 136.995 ;
        RECT 100.640 134.455 101.640 134.715 ;
        RECT 100.640 132.175 101.640 132.435 ;
        RECT 97.050 129.895 98.050 130.155 ;
        RECT 100.640 129.895 101.640 130.155 ;
        RECT 98.240 128.050 98.530 129.720 ;
        RECT 97.050 127.615 98.050 127.875 ;
        RECT 100.640 127.615 101.640 127.875 ;
        RECT 96.530 114.370 96.860 127.440 ;
        RECT 98.240 125.770 98.530 127.440 ;
        RECT 101.830 125.770 102.160 129.720 ;
        RECT 97.050 125.335 98.050 125.595 ;
        RECT 100.640 125.335 101.640 125.595 ;
        RECT 98.240 123.490 98.530 125.160 ;
        RECT 97.050 123.055 98.050 123.315 ;
        RECT 98.240 121.210 98.530 122.880 ;
        RECT 97.050 120.775 98.050 121.035 ;
        RECT 98.240 118.930 98.530 120.600 ;
        RECT 97.050 118.495 98.050 118.755 ;
        RECT 98.240 116.650 98.530 118.320 ;
        RECT 97.050 116.215 98.050 116.475 ;
        RECT 98.240 114.370 98.530 116.040 ;
        RECT 97.050 113.935 98.050 114.195 ;
        RECT 97.050 113.155 98.050 113.415 ;
        RECT 97.050 112.375 98.050 112.635 ;
        RECT 98.240 111.980 98.530 113.760 ;
        RECT 100.160 111.980 100.450 125.160 ;
        RECT 100.640 123.055 101.640 123.315 ;
        RECT 100.640 120.775 101.640 121.035 ;
        RECT 100.640 118.495 101.640 118.755 ;
        RECT 100.640 116.215 101.640 116.475 ;
        RECT 100.640 113.935 101.640 114.195 ;
        RECT 102.380 111.980 102.670 151.190 ;
        RECT 96.020 111.690 102.670 111.980 ;
        RECT 88.485 88.890 91.180 89.180 ;
        RECT 91.445 88.890 95.165 89.180 ;
        RECT 88.445 82.710 91.140 83.000 ;
        RECT 91.430 82.710 95.150 83.000 ;
        RECT 71.415 82.360 74.390 82.650 ;
        RECT 74.800 82.360 83.760 82.650 ;
        RECT 84.170 82.360 87.145 82.650 ;
        RECT 71.415 77.870 71.705 82.360 ;
        RECT 72.595 81.950 73.445 81.965 ;
        RECT 72.445 81.720 73.445 81.950 ;
        RECT 72.595 81.705 73.445 81.720 ;
        RECT 71.965 81.110 72.255 81.700 ;
        RECT 72.595 81.520 73.445 81.535 ;
        RECT 72.445 81.290 73.445 81.520 ;
        RECT 72.595 81.275 73.445 81.290 ;
        RECT 73.635 81.110 73.925 82.360 ;
        RECT 72.595 81.090 73.445 81.105 ;
        RECT 72.445 80.860 73.445 81.090 ;
        RECT 72.595 80.845 73.445 80.860 ;
        RECT 71.925 80.250 72.255 80.840 ;
        RECT 72.445 80.415 73.445 80.675 ;
        RECT 73.635 80.250 73.925 80.840 ;
        RECT 72.595 80.230 73.445 80.245 ;
        RECT 72.445 80.000 73.445 80.230 ;
        RECT 72.595 79.985 73.445 80.000 ;
        RECT 71.965 79.390 72.255 79.980 ;
        RECT 73.635 79.850 73.925 79.980 ;
        RECT 74.430 79.850 74.760 81.895 ;
        RECT 75.265 81.110 75.555 82.360 ;
        RECT 75.820 81.950 76.670 81.965 ;
        RECT 77.395 81.950 78.245 81.965 ;
        RECT 75.745 81.720 76.745 81.950 ;
        RECT 77.395 81.720 78.395 81.950 ;
        RECT 75.820 81.705 76.670 81.720 ;
        RECT 77.395 81.705 78.245 81.720 ;
        RECT 78.625 81.700 78.915 82.360 ;
        RECT 75.820 81.520 76.670 81.535 ;
        RECT 77.395 81.520 78.245 81.535 ;
        RECT 75.745 81.290 76.745 81.520 ;
        RECT 77.395 81.290 78.395 81.520 ;
        RECT 75.820 81.275 76.670 81.290 ;
        RECT 77.395 81.275 78.245 81.290 ;
        RECT 78.585 81.110 78.915 81.700 ;
        RECT 75.745 80.845 76.745 81.105 ;
        RECT 77.395 81.090 78.245 81.105 ;
        RECT 77.395 80.860 78.395 81.090 ;
        RECT 77.395 80.845 78.245 80.860 ;
        RECT 75.225 79.850 75.555 80.840 ;
        RECT 75.745 80.415 76.745 80.675 ;
        RECT 77.395 80.415 78.395 80.675 ;
        RECT 75.745 79.985 76.745 80.245 ;
        RECT 77.395 80.230 78.245 80.245 ;
        RECT 77.395 80.000 78.395 80.230 ;
        RECT 77.395 79.985 78.245 80.000 ;
        RECT 72.445 79.555 73.445 79.815 ;
        RECT 73.635 79.520 75.555 79.850 ;
        RECT 75.745 79.555 76.745 79.815 ;
        RECT 77.395 79.555 78.395 79.815 ;
        RECT 73.635 79.390 73.925 79.520 ;
        RECT 75.225 79.390 75.555 79.520 ;
        RECT 78.585 79.390 78.915 80.840 ;
        RECT 72.595 79.370 73.445 79.385 ;
        RECT 72.445 79.140 73.445 79.370 ;
        RECT 72.595 79.125 73.445 79.140 ;
        RECT 75.745 79.125 76.745 79.385 ;
        RECT 77.395 79.370 78.245 79.385 ;
        RECT 77.395 79.140 78.395 79.370 ;
        RECT 77.395 79.125 78.245 79.140 ;
        RECT 71.965 78.530 72.255 79.120 ;
        RECT 72.595 78.940 73.445 78.955 ;
        RECT 72.445 78.710 73.445 78.940 ;
        RECT 72.595 78.695 73.445 78.710 ;
        RECT 72.595 78.510 73.445 78.525 ;
        RECT 72.445 78.280 73.445 78.510 ;
        RECT 72.595 78.265 73.445 78.280 ;
        RECT 72.595 77.870 73.445 77.875 ;
        RECT 73.635 77.870 73.925 79.120 ;
        RECT 75.265 77.870 75.555 79.120 ;
        RECT 75.820 78.940 76.670 78.955 ;
        RECT 77.395 78.940 78.245 78.955 ;
        RECT 75.745 78.710 76.745 78.940 ;
        RECT 77.395 78.710 78.395 78.940 ;
        RECT 75.820 78.695 76.670 78.710 ;
        RECT 77.395 78.695 78.245 78.710 ;
        RECT 78.585 78.530 78.915 79.120 ;
        RECT 75.820 78.510 76.670 78.525 ;
        RECT 77.395 78.510 78.245 78.525 ;
        RECT 75.745 78.280 76.745 78.510 ;
        RECT 77.395 78.280 78.395 78.510 ;
        RECT 75.820 78.265 76.670 78.280 ;
        RECT 77.395 78.265 78.245 78.280 ;
        RECT 75.820 77.870 76.670 77.875 ;
        RECT 77.395 77.870 78.245 77.875 ;
        RECT 78.625 77.870 78.915 78.530 ;
        RECT 79.135 77.870 79.425 82.360 ;
        RECT 79.645 81.700 79.935 82.360 ;
        RECT 80.315 81.950 81.165 81.965 ;
        RECT 81.890 81.950 82.740 81.965 ;
        RECT 80.165 81.720 81.165 81.950 ;
        RECT 81.815 81.720 82.815 81.950 ;
        RECT 80.315 81.705 81.165 81.720 ;
        RECT 81.890 81.705 82.740 81.720 ;
        RECT 79.645 81.110 79.975 81.700 ;
        RECT 80.315 81.520 81.165 81.535 ;
        RECT 81.890 81.520 82.740 81.535 ;
        RECT 80.165 81.290 81.165 81.520 ;
        RECT 81.815 81.290 82.815 81.520 ;
        RECT 80.315 81.275 81.165 81.290 ;
        RECT 81.890 81.275 82.740 81.290 ;
        RECT 83.005 81.110 83.295 82.360 ;
        RECT 80.315 81.090 81.165 81.105 ;
        RECT 80.165 80.860 81.165 81.090 ;
        RECT 80.315 80.845 81.165 80.860 ;
        RECT 81.815 80.845 82.815 81.105 ;
        RECT 79.645 79.390 79.975 80.840 ;
        RECT 80.165 80.415 81.165 80.675 ;
        RECT 81.815 80.415 82.815 80.675 ;
        RECT 80.315 80.230 81.165 80.245 ;
        RECT 80.165 80.000 81.165 80.230 ;
        RECT 80.315 79.985 81.165 80.000 ;
        RECT 81.815 79.985 82.815 80.245 ;
        RECT 83.005 79.850 83.335 80.840 ;
        RECT 83.800 79.850 84.130 81.895 ;
        RECT 84.635 81.110 84.925 82.360 ;
        RECT 85.115 81.950 85.965 81.965 ;
        RECT 85.115 81.720 86.115 81.950 ;
        RECT 85.115 81.705 85.965 81.720 ;
        RECT 85.115 81.520 85.965 81.535 ;
        RECT 85.115 81.290 86.115 81.520 ;
        RECT 85.115 81.275 85.965 81.290 ;
        RECT 86.305 81.110 86.595 81.700 ;
        RECT 85.115 81.090 85.965 81.105 ;
        RECT 85.115 80.860 86.115 81.090 ;
        RECT 85.115 80.845 85.965 80.860 ;
        RECT 84.635 80.250 84.925 80.840 ;
        RECT 85.115 80.415 86.115 80.675 ;
        RECT 86.305 80.250 86.635 80.840 ;
        RECT 85.115 80.230 85.965 80.245 ;
        RECT 85.115 80.000 86.115 80.230 ;
        RECT 85.115 79.985 85.965 80.000 ;
        RECT 84.635 79.850 84.925 79.980 ;
        RECT 80.165 79.555 81.165 79.815 ;
        RECT 81.815 79.555 82.815 79.815 ;
        RECT 83.005 79.520 84.925 79.850 ;
        RECT 85.115 79.555 86.115 79.815 ;
        RECT 83.005 79.390 83.335 79.520 ;
        RECT 84.635 79.390 84.925 79.520 ;
        RECT 86.305 79.390 86.595 79.980 ;
        RECT 80.315 79.370 81.165 79.385 ;
        RECT 80.165 79.140 81.165 79.370 ;
        RECT 80.315 79.125 81.165 79.140 ;
        RECT 81.815 79.125 82.815 79.385 ;
        RECT 85.115 79.370 85.965 79.385 ;
        RECT 85.115 79.140 86.115 79.370 ;
        RECT 85.115 79.125 85.965 79.140 ;
        RECT 79.645 78.530 79.975 79.120 ;
        RECT 80.315 78.940 81.165 78.955 ;
        RECT 81.890 78.940 82.740 78.955 ;
        RECT 80.165 78.710 81.165 78.940 ;
        RECT 81.815 78.710 82.815 78.940 ;
        RECT 80.315 78.695 81.165 78.710 ;
        RECT 81.890 78.695 82.740 78.710 ;
        RECT 79.645 77.870 79.935 78.530 ;
        RECT 80.315 78.510 81.165 78.525 ;
        RECT 81.890 78.510 82.740 78.525 ;
        RECT 80.165 78.280 81.165 78.510 ;
        RECT 81.815 78.280 82.815 78.510 ;
        RECT 80.315 78.265 81.165 78.280 ;
        RECT 81.890 78.265 82.740 78.280 ;
        RECT 80.315 77.870 81.165 77.875 ;
        RECT 81.890 77.870 82.740 77.875 ;
        RECT 83.005 77.870 83.295 79.120 ;
        RECT 84.635 77.870 84.925 79.120 ;
        RECT 85.115 78.940 85.965 78.955 ;
        RECT 85.115 78.710 86.115 78.940 ;
        RECT 85.115 78.695 85.965 78.710 ;
        RECT 86.305 78.530 86.595 79.120 ;
        RECT 85.115 78.510 85.965 78.525 ;
        RECT 85.115 78.280 86.115 78.510 ;
        RECT 85.115 78.265 85.965 78.280 ;
        RECT 85.115 77.870 85.965 77.875 ;
        RECT 86.855 77.870 87.145 82.360 ;
        RECT 88.445 78.220 88.735 82.710 ;
        RECT 89.110 82.055 90.110 82.315 ;
        RECT 89.110 81.625 90.110 81.885 ;
        RECT 90.300 81.460 90.590 82.710 ;
        RECT 89.110 81.195 90.110 81.455 ;
        RECT 89.110 80.765 90.110 81.025 ;
        RECT 90.300 80.630 90.590 81.190 ;
        RECT 91.120 80.630 91.450 82.305 ;
        RECT 91.980 81.460 92.270 82.710 ;
        RECT 92.960 82.300 93.960 82.315 ;
        RECT 92.460 82.070 94.460 82.300 ;
        RECT 92.960 82.055 93.960 82.070 ;
        RECT 92.960 81.870 93.960 81.885 ;
        RECT 92.460 81.640 94.460 81.870 ;
        RECT 92.960 81.625 93.960 81.640 ;
        RECT 92.960 81.440 93.960 81.455 ;
        RECT 92.460 81.210 94.460 81.440 ;
        RECT 92.960 81.195 93.960 81.210 ;
        RECT 91.980 80.630 92.270 81.190 ;
        RECT 92.460 80.765 94.460 81.025 ;
        RECT 89.110 80.335 90.110 80.595 ;
        RECT 90.300 80.300 92.270 80.630 ;
        RECT 92.960 80.580 93.960 80.595 ;
        RECT 92.460 80.350 94.460 80.580 ;
        RECT 92.960 80.335 93.960 80.350 ;
        RECT 89.110 79.905 90.110 80.165 ;
        RECT 90.300 79.740 90.590 80.300 ;
        RECT 91.980 79.740 92.270 80.300 ;
        RECT 92.460 79.905 94.460 80.165 ;
        RECT 89.110 79.475 90.110 79.735 ;
        RECT 92.960 79.720 93.960 79.735 ;
        RECT 92.460 79.490 94.460 79.720 ;
        RECT 92.960 79.475 93.960 79.490 ;
        RECT 89.110 79.045 90.110 79.305 ;
        RECT 89.110 78.615 90.110 78.875 ;
        RECT 90.300 78.220 90.590 79.470 ;
        RECT 91.980 78.220 92.270 79.470 ;
        RECT 92.960 79.290 93.960 79.305 ;
        RECT 92.460 79.060 94.460 79.290 ;
        RECT 92.960 79.045 93.960 79.060 ;
        RECT 92.960 78.860 93.960 78.875 ;
        RECT 92.460 78.630 94.460 78.860 ;
        RECT 92.960 78.615 93.960 78.630 ;
        RECT 94.860 78.220 95.150 82.710 ;
        RECT 88.445 77.930 91.140 78.220 ;
        RECT 91.430 77.930 95.150 78.220 ;
        RECT 71.415 77.580 74.390 77.870 ;
        RECT 74.800 77.580 83.760 77.870 ;
        RECT 84.170 77.580 87.145 77.870 ;
        RECT 64.665 72.050 67.360 72.340 ;
        RECT 67.650 72.050 71.370 72.340 ;
        RECT 64.665 63.260 64.955 72.050 ;
        RECT 65.330 71.395 66.330 71.655 ;
        RECT 65.330 70.965 66.330 71.225 ;
        RECT 66.520 70.800 66.810 72.050 ;
        RECT 65.330 70.535 66.330 70.795 ;
        RECT 65.330 70.105 66.330 70.365 ;
        RECT 66.520 69.985 66.810 70.530 ;
        RECT 67.340 69.985 67.670 71.645 ;
        RECT 68.200 70.800 68.490 72.050 ;
        RECT 69.180 71.640 70.180 71.655 ;
        RECT 68.680 71.410 70.680 71.640 ;
        RECT 69.180 71.395 70.180 71.410 ;
        RECT 69.180 71.210 70.180 71.225 ;
        RECT 68.680 70.980 70.680 71.210 ;
        RECT 69.180 70.965 70.180 70.980 ;
        RECT 69.180 70.780 70.180 70.795 ;
        RECT 68.680 70.550 70.680 70.780 ;
        RECT 69.180 70.535 70.180 70.550 ;
        RECT 68.200 69.985 68.490 70.530 ;
        RECT 68.680 70.105 70.680 70.365 ;
        RECT 65.330 69.675 66.330 69.935 ;
        RECT 66.520 69.655 68.490 69.985 ;
        RECT 69.180 69.920 70.180 69.935 ;
        RECT 68.680 69.690 70.680 69.920 ;
        RECT 69.180 69.675 70.180 69.690 ;
        RECT 65.330 69.245 66.330 69.505 ;
        RECT 66.520 69.080 66.810 69.655 ;
        RECT 67.025 69.235 67.985 69.515 ;
        RECT 65.330 68.815 66.330 69.075 ;
        RECT 65.330 68.385 66.330 68.645 ;
        RECT 65.330 67.955 66.330 68.215 ;
        RECT 65.330 67.525 66.330 67.785 ;
        RECT 65.330 67.095 66.330 67.355 ;
        RECT 66.520 66.960 66.810 68.810 ;
        RECT 67.340 66.960 67.670 69.235 ;
        RECT 68.200 69.080 68.490 69.655 ;
        RECT 68.680 69.245 70.680 69.505 ;
        RECT 69.180 69.060 70.180 69.075 ;
        RECT 68.680 68.830 70.680 69.060 ;
        RECT 69.180 68.815 70.180 68.830 ;
        RECT 68.200 66.960 68.490 68.810 ;
        RECT 68.680 68.385 70.680 68.645 ;
        RECT 69.180 68.200 70.180 68.215 ;
        RECT 68.680 67.970 70.680 68.200 ;
        RECT 69.180 67.955 70.180 67.970 ;
        RECT 68.680 67.525 70.680 67.785 ;
        RECT 69.180 67.340 70.180 67.355 ;
        RECT 68.680 67.110 70.680 67.340 ;
        RECT 69.180 67.095 70.180 67.110 ;
        RECT 65.330 66.665 66.330 66.925 ;
        RECT 66.520 66.630 68.490 66.960 ;
        RECT 68.680 66.665 70.680 66.925 ;
        RECT 65.330 66.235 66.330 66.495 ;
        RECT 65.330 65.805 66.330 66.065 ;
        RECT 65.330 65.375 66.330 65.635 ;
        RECT 65.330 64.945 66.330 65.205 ;
        RECT 66.520 64.780 66.810 66.630 ;
        RECT 68.200 64.780 68.490 66.630 ;
        RECT 69.180 66.480 70.180 66.495 ;
        RECT 68.680 66.250 70.680 66.480 ;
        RECT 69.180 66.235 70.180 66.250 ;
        RECT 68.680 65.805 70.680 66.065 ;
        RECT 69.180 65.620 70.180 65.635 ;
        RECT 68.680 65.390 70.680 65.620 ;
        RECT 69.180 65.375 70.180 65.390 ;
        RECT 68.680 64.945 70.680 65.205 ;
        RECT 65.330 64.515 66.330 64.775 ;
        RECT 69.180 64.760 70.180 64.775 ;
        RECT 68.680 64.530 70.680 64.760 ;
        RECT 69.180 64.515 70.180 64.530 ;
        RECT 65.330 64.085 66.330 64.345 ;
        RECT 65.330 63.655 66.330 63.915 ;
        RECT 66.520 63.260 66.810 64.510 ;
        RECT 68.200 63.260 68.490 64.510 ;
        RECT 69.180 64.330 70.180 64.345 ;
        RECT 68.680 64.100 70.680 64.330 ;
        RECT 69.180 64.085 70.180 64.100 ;
        RECT 69.180 63.900 70.180 63.915 ;
        RECT 68.680 63.670 70.680 63.900 ;
        RECT 69.180 63.655 70.180 63.670 ;
        RECT 71.080 63.260 71.370 72.050 ;
        RECT 64.665 62.970 67.360 63.260 ;
        RECT 67.650 62.970 71.370 63.260 ;
        RECT 73.685 72.050 76.380 72.340 ;
        RECT 76.670 72.050 83.820 72.340 ;
        RECT 84.110 72.050 86.805 72.340 ;
        RECT 73.685 63.260 73.975 72.050 ;
        RECT 74.350 71.395 75.350 71.655 ;
        RECT 74.350 70.965 75.350 71.225 ;
        RECT 75.540 70.800 75.830 72.050 ;
        RECT 74.350 70.535 75.350 70.795 ;
        RECT 74.350 70.105 75.350 70.365 ;
        RECT 75.540 69.985 75.830 70.530 ;
        RECT 76.360 69.985 76.690 71.645 ;
        RECT 77.220 70.800 77.510 72.050 ;
        RECT 78.200 71.640 79.200 71.655 ;
        RECT 77.700 71.410 79.700 71.640 ;
        RECT 78.200 71.395 79.200 71.410 ;
        RECT 78.200 71.210 79.200 71.225 ;
        RECT 77.700 70.980 79.700 71.210 ;
        RECT 78.200 70.965 79.200 70.980 ;
        RECT 78.200 70.780 79.200 70.795 ;
        RECT 77.700 70.550 79.700 70.780 ;
        RECT 78.200 70.535 79.200 70.550 ;
        RECT 77.220 69.985 77.510 70.530 ;
        RECT 77.700 70.105 79.700 70.365 ;
        RECT 74.350 69.675 75.350 69.935 ;
        RECT 75.540 69.655 77.510 69.985 ;
        RECT 78.200 69.920 79.200 69.935 ;
        RECT 77.700 69.690 79.700 69.920 ;
        RECT 78.200 69.675 79.200 69.690 ;
        RECT 74.350 69.245 75.350 69.505 ;
        RECT 75.540 69.080 75.830 69.655 ;
        RECT 76.045 69.235 77.005 69.515 ;
        RECT 74.350 68.815 75.350 69.075 ;
        RECT 74.350 68.385 75.350 68.645 ;
        RECT 74.350 67.955 75.350 68.215 ;
        RECT 74.350 67.525 75.350 67.785 ;
        RECT 74.350 67.095 75.350 67.355 ;
        RECT 75.540 66.960 75.830 68.810 ;
        RECT 76.360 66.960 76.690 69.235 ;
        RECT 77.220 69.080 77.510 69.655 ;
        RECT 77.700 69.245 79.700 69.505 ;
        RECT 78.200 69.060 79.200 69.075 ;
        RECT 77.700 68.830 79.700 69.060 ;
        RECT 78.200 68.815 79.200 68.830 ;
        RECT 77.220 66.960 77.510 68.810 ;
        RECT 77.700 68.385 79.700 68.645 ;
        RECT 78.200 68.200 79.200 68.215 ;
        RECT 77.700 67.970 79.700 68.200 ;
        RECT 78.200 67.955 79.200 67.970 ;
        RECT 77.700 67.525 79.700 67.785 ;
        RECT 78.200 67.340 79.200 67.355 ;
        RECT 77.700 67.110 79.700 67.340 ;
        RECT 78.200 67.095 79.200 67.110 ;
        RECT 74.350 66.665 75.350 66.925 ;
        RECT 75.540 66.630 77.510 66.960 ;
        RECT 77.700 66.665 79.700 66.925 ;
        RECT 74.350 66.235 75.350 66.495 ;
        RECT 74.350 65.805 75.350 66.065 ;
        RECT 74.350 65.375 75.350 65.635 ;
        RECT 74.350 64.945 75.350 65.205 ;
        RECT 75.540 64.780 75.830 66.630 ;
        RECT 77.220 64.780 77.510 66.630 ;
        RECT 78.200 66.480 79.200 66.495 ;
        RECT 77.700 66.250 79.700 66.480 ;
        RECT 78.200 66.235 79.200 66.250 ;
        RECT 77.700 65.805 79.700 66.065 ;
        RECT 78.200 65.620 79.200 65.635 ;
        RECT 77.700 65.390 79.700 65.620 ;
        RECT 78.200 65.375 79.200 65.390 ;
        RECT 77.700 64.945 79.700 65.205 ;
        RECT 74.350 64.515 75.350 64.775 ;
        RECT 78.200 64.760 79.200 64.775 ;
        RECT 77.700 64.530 79.700 64.760 ;
        RECT 78.200 64.515 79.200 64.530 ;
        RECT 74.350 64.085 75.350 64.345 ;
        RECT 74.350 63.655 75.350 63.915 ;
        RECT 75.540 63.260 75.830 64.510 ;
        RECT 77.220 63.260 77.510 64.510 ;
        RECT 78.200 64.330 79.200 64.345 ;
        RECT 77.700 64.100 79.700 64.330 ;
        RECT 78.200 64.085 79.200 64.100 ;
        RECT 78.200 63.900 79.200 63.915 ;
        RECT 77.700 63.670 79.700 63.900 ;
        RECT 78.200 63.655 79.200 63.670 ;
        RECT 80.100 63.260 80.390 72.050 ;
        RECT 81.290 71.640 82.290 71.655 ;
        RECT 80.790 71.410 82.790 71.640 ;
        RECT 81.290 71.395 82.290 71.410 ;
        RECT 81.290 71.210 82.290 71.225 ;
        RECT 80.790 70.980 82.790 71.210 ;
        RECT 81.290 70.965 82.290 70.980 ;
        RECT 82.980 70.800 83.270 72.050 ;
        RECT 81.290 70.780 82.290 70.795 ;
        RECT 80.790 70.550 82.790 70.780 ;
        RECT 81.290 70.535 82.290 70.550 ;
        RECT 80.790 70.105 82.790 70.365 ;
        RECT 82.980 69.985 83.270 70.530 ;
        RECT 83.800 69.985 84.130 71.645 ;
        RECT 84.660 70.800 84.950 72.050 ;
        RECT 85.140 71.395 86.140 71.655 ;
        RECT 85.140 70.965 86.140 71.225 ;
        RECT 85.140 70.535 86.140 70.795 ;
        RECT 84.660 69.985 84.950 70.530 ;
        RECT 85.140 70.105 86.140 70.365 ;
        RECT 81.290 69.920 82.290 69.935 ;
        RECT 80.790 69.690 82.790 69.920 ;
        RECT 81.290 69.675 82.290 69.690 ;
        RECT 82.980 69.655 84.950 69.985 ;
        RECT 85.140 69.675 86.140 69.935 ;
        RECT 80.790 69.245 82.790 69.505 ;
        RECT 82.980 69.080 83.270 69.655 ;
        RECT 83.485 69.235 84.445 69.515 ;
        RECT 81.290 69.060 82.290 69.075 ;
        RECT 80.790 68.830 82.790 69.060 ;
        RECT 81.290 68.815 82.290 68.830 ;
        RECT 80.790 68.385 82.790 68.645 ;
        RECT 81.290 68.200 82.290 68.215 ;
        RECT 80.790 67.970 82.790 68.200 ;
        RECT 81.290 67.955 82.290 67.970 ;
        RECT 80.790 67.525 82.790 67.785 ;
        RECT 81.290 67.340 82.290 67.355 ;
        RECT 80.790 67.110 82.790 67.340 ;
        RECT 81.290 67.095 82.290 67.110 ;
        RECT 82.980 66.960 83.270 68.810 ;
        RECT 83.800 66.960 84.130 69.235 ;
        RECT 84.660 69.080 84.950 69.655 ;
        RECT 85.140 69.245 86.140 69.505 ;
        RECT 85.140 68.815 86.140 69.075 ;
        RECT 84.660 66.960 84.950 68.810 ;
        RECT 85.140 68.385 86.140 68.645 ;
        RECT 85.140 67.955 86.140 68.215 ;
        RECT 85.140 67.525 86.140 67.785 ;
        RECT 85.140 67.095 86.140 67.355 ;
        RECT 80.790 66.665 82.790 66.925 ;
        RECT 82.980 66.630 84.950 66.960 ;
        RECT 85.140 66.665 86.140 66.925 ;
        RECT 81.290 66.480 82.290 66.495 ;
        RECT 80.790 66.250 82.790 66.480 ;
        RECT 81.290 66.235 82.290 66.250 ;
        RECT 80.790 65.805 82.790 66.065 ;
        RECT 81.290 65.620 82.290 65.635 ;
        RECT 80.790 65.390 82.790 65.620 ;
        RECT 81.290 65.375 82.290 65.390 ;
        RECT 80.790 64.945 82.790 65.205 ;
        RECT 82.980 64.780 83.270 66.630 ;
        RECT 84.660 64.780 84.950 66.630 ;
        RECT 85.140 66.235 86.140 66.495 ;
        RECT 85.140 65.805 86.140 66.065 ;
        RECT 85.140 65.375 86.140 65.635 ;
        RECT 85.140 64.945 86.140 65.205 ;
        RECT 81.290 64.760 82.290 64.775 ;
        RECT 80.790 64.530 82.790 64.760 ;
        RECT 81.290 64.515 82.290 64.530 ;
        RECT 85.140 64.515 86.140 64.775 ;
        RECT 81.290 64.330 82.290 64.345 ;
        RECT 80.790 64.100 82.790 64.330 ;
        RECT 81.290 64.085 82.290 64.100 ;
        RECT 81.290 63.900 82.290 63.915 ;
        RECT 80.790 63.670 82.790 63.900 ;
        RECT 81.290 63.655 82.290 63.670 ;
        RECT 82.980 63.260 83.270 64.510 ;
        RECT 84.660 63.260 84.950 64.510 ;
        RECT 85.140 64.085 86.140 64.345 ;
        RECT 85.140 63.655 86.140 63.915 ;
        RECT 86.515 63.260 86.805 72.050 ;
        RECT 73.685 62.970 76.380 63.260 ;
        RECT 76.670 62.970 83.820 63.260 ;
        RECT 84.110 62.970 86.805 63.260 ;
        RECT 88.445 72.050 91.140 72.340 ;
        RECT 91.430 72.050 95.150 72.340 ;
        RECT 88.445 63.260 88.735 72.050 ;
        RECT 89.110 71.395 90.110 71.655 ;
        RECT 89.110 70.965 90.110 71.225 ;
        RECT 90.300 70.800 90.590 72.050 ;
        RECT 89.110 70.535 90.110 70.795 ;
        RECT 89.110 70.105 90.110 70.365 ;
        RECT 90.300 69.985 90.590 70.530 ;
        RECT 91.120 69.985 91.450 71.645 ;
        RECT 91.980 70.800 92.270 72.050 ;
        RECT 92.960 71.640 93.960 71.655 ;
        RECT 92.460 71.410 94.460 71.640 ;
        RECT 92.960 71.395 93.960 71.410 ;
        RECT 92.960 71.210 93.960 71.225 ;
        RECT 92.460 70.980 94.460 71.210 ;
        RECT 92.960 70.965 93.960 70.980 ;
        RECT 92.960 70.780 93.960 70.795 ;
        RECT 92.460 70.550 94.460 70.780 ;
        RECT 92.960 70.535 93.960 70.550 ;
        RECT 91.980 69.985 92.270 70.530 ;
        RECT 92.460 70.105 94.460 70.365 ;
        RECT 89.110 69.675 90.110 69.935 ;
        RECT 90.300 69.655 92.270 69.985 ;
        RECT 92.960 69.920 93.960 69.935 ;
        RECT 92.460 69.690 94.460 69.920 ;
        RECT 92.960 69.675 93.960 69.690 ;
        RECT 89.110 69.245 90.110 69.505 ;
        RECT 90.300 69.080 90.590 69.655 ;
        RECT 90.805 69.235 91.765 69.515 ;
        RECT 89.110 68.815 90.110 69.075 ;
        RECT 89.110 68.385 90.110 68.645 ;
        RECT 89.110 67.955 90.110 68.215 ;
        RECT 89.110 67.525 90.110 67.785 ;
        RECT 89.110 67.095 90.110 67.355 ;
        RECT 90.300 66.960 90.590 68.810 ;
        RECT 91.120 66.960 91.450 69.235 ;
        RECT 91.980 69.080 92.270 69.655 ;
        RECT 92.460 69.245 94.460 69.505 ;
        RECT 92.960 69.060 93.960 69.075 ;
        RECT 92.460 68.830 94.460 69.060 ;
        RECT 92.960 68.815 93.960 68.830 ;
        RECT 91.980 66.960 92.270 68.810 ;
        RECT 92.460 68.385 94.460 68.645 ;
        RECT 92.960 68.200 93.960 68.215 ;
        RECT 92.460 67.970 94.460 68.200 ;
        RECT 92.960 67.955 93.960 67.970 ;
        RECT 92.460 67.525 94.460 67.785 ;
        RECT 92.960 67.340 93.960 67.355 ;
        RECT 92.460 67.110 94.460 67.340 ;
        RECT 92.960 67.095 93.960 67.110 ;
        RECT 89.110 66.665 90.110 66.925 ;
        RECT 90.300 66.630 92.270 66.960 ;
        RECT 92.460 66.665 94.460 66.925 ;
        RECT 89.110 66.235 90.110 66.495 ;
        RECT 89.110 65.805 90.110 66.065 ;
        RECT 89.110 65.375 90.110 65.635 ;
        RECT 89.110 64.945 90.110 65.205 ;
        RECT 90.300 64.780 90.590 66.630 ;
        RECT 91.980 64.780 92.270 66.630 ;
        RECT 92.960 66.480 93.960 66.495 ;
        RECT 92.460 66.250 94.460 66.480 ;
        RECT 92.960 66.235 93.960 66.250 ;
        RECT 92.460 65.805 94.460 66.065 ;
        RECT 92.960 65.620 93.960 65.635 ;
        RECT 92.460 65.390 94.460 65.620 ;
        RECT 92.960 65.375 93.960 65.390 ;
        RECT 92.460 64.945 94.460 65.205 ;
        RECT 89.110 64.515 90.110 64.775 ;
        RECT 92.960 64.760 93.960 64.775 ;
        RECT 92.460 64.530 94.460 64.760 ;
        RECT 92.960 64.515 93.960 64.530 ;
        RECT 89.110 64.085 90.110 64.345 ;
        RECT 89.110 63.655 90.110 63.915 ;
        RECT 90.300 63.260 90.590 64.510 ;
        RECT 91.980 63.260 92.270 64.510 ;
        RECT 92.960 64.330 93.960 64.345 ;
        RECT 92.460 64.100 94.460 64.330 ;
        RECT 92.960 64.085 93.960 64.100 ;
        RECT 92.960 63.900 93.960 63.915 ;
        RECT 92.460 63.670 94.460 63.900 ;
        RECT 92.960 63.655 93.960 63.670 ;
        RECT 94.860 63.260 95.150 72.050 ;
        RECT 88.445 62.970 91.140 63.260 ;
        RECT 91.430 62.970 95.150 63.260 ;
        RECT 108.575 63.070 108.865 164.440 ;
        RECT 109.605 163.785 110.305 164.045 ;
        RECT 109.605 161.505 110.305 161.765 ;
        RECT 110.495 159.660 110.785 164.440 ;
        RECT 110.975 163.785 111.675 164.045 ;
        RECT 110.975 161.505 111.675 161.765 ;
        RECT 111.865 159.660 112.155 164.440 ;
        RECT 112.345 163.785 113.045 164.045 ;
        RECT 112.345 161.505 113.045 161.765 ;
        RECT 109.605 159.225 110.305 159.485 ;
        RECT 110.975 159.225 111.675 159.485 ;
        RECT 112.345 159.225 113.045 159.485 ;
        RECT 110.475 157.215 110.805 159.050 ;
        RECT 111.845 157.215 112.175 159.050 ;
        RECT 109.605 156.935 113.045 157.215 ;
        RECT 109.605 154.665 110.305 154.925 ;
        RECT 110.475 152.655 110.805 156.935 ;
        RECT 110.975 154.665 111.675 154.925 ;
        RECT 111.845 152.655 112.175 156.935 ;
        RECT 112.345 154.665 113.045 154.925 ;
        RECT 109.605 152.375 113.045 152.655 ;
        RECT 109.605 150.105 110.305 150.365 ;
        RECT 110.475 148.095 110.805 152.375 ;
        RECT 110.975 150.105 111.675 150.365 ;
        RECT 111.845 148.095 112.175 152.375 ;
        RECT 112.345 150.105 113.045 150.365 ;
        RECT 109.605 147.815 113.045 148.095 ;
        RECT 109.605 145.545 110.305 145.805 ;
        RECT 110.475 143.535 110.805 147.815 ;
        RECT 110.975 145.545 111.675 145.805 ;
        RECT 111.845 143.535 112.175 147.815 ;
        RECT 112.345 145.545 113.045 145.805 ;
        RECT 109.605 143.255 113.045 143.535 ;
        RECT 109.605 140.985 110.305 141.245 ;
        RECT 110.475 138.975 110.805 143.255 ;
        RECT 110.975 140.985 111.675 141.245 ;
        RECT 111.845 138.975 112.175 143.255 ;
        RECT 112.345 140.985 113.045 141.245 ;
        RECT 109.605 138.695 113.045 138.975 ;
        RECT 109.605 136.425 110.305 136.685 ;
        RECT 109.605 134.145 110.305 134.405 ;
        RECT 109.605 131.865 110.305 132.125 ;
        RECT 109.605 129.585 110.305 129.845 ;
        RECT 109.605 127.305 110.305 127.565 ;
        RECT 109.605 125.025 110.305 125.285 ;
        RECT 109.605 122.745 110.305 123.005 ;
        RECT 109.605 120.465 110.305 120.725 ;
        RECT 109.605 118.185 110.305 118.445 ;
        RECT 109.605 115.905 110.305 116.165 ;
        RECT 109.605 113.625 110.305 113.885 ;
        RECT 109.605 111.345 110.305 111.605 ;
        RECT 109.605 109.065 110.305 109.325 ;
        RECT 109.605 106.785 110.305 107.045 ;
        RECT 109.605 104.505 110.305 104.765 ;
        RECT 109.605 102.225 110.305 102.485 ;
        RECT 109.605 99.945 110.305 100.205 ;
        RECT 109.605 97.665 110.305 97.925 ;
        RECT 109.605 95.385 110.305 95.645 ;
        RECT 109.605 93.105 110.305 93.365 ;
        RECT 109.605 90.825 110.305 91.085 ;
        RECT 109.605 88.545 110.305 88.805 ;
        RECT 109.605 86.265 110.305 86.525 ;
        RECT 109.605 83.985 110.305 84.245 ;
        RECT 109.605 81.705 110.305 81.965 ;
        RECT 109.605 79.425 110.305 79.685 ;
        RECT 109.605 77.145 110.305 77.405 ;
        RECT 109.605 74.865 110.305 75.125 ;
        RECT 109.605 72.585 110.305 72.845 ;
        RECT 109.605 70.305 110.305 70.565 ;
        RECT 110.475 68.460 110.805 138.695 ;
        RECT 110.975 136.425 111.675 136.685 ;
        RECT 110.975 134.145 111.675 134.405 ;
        RECT 110.975 131.865 111.675 132.125 ;
        RECT 110.975 129.585 111.675 129.845 ;
        RECT 110.975 127.305 111.675 127.565 ;
        RECT 110.975 125.025 111.675 125.285 ;
        RECT 110.975 122.745 111.675 123.005 ;
        RECT 110.975 120.465 111.675 120.725 ;
        RECT 110.975 118.185 111.675 118.445 ;
        RECT 110.975 115.905 111.675 116.165 ;
        RECT 110.975 113.625 111.675 113.885 ;
        RECT 110.975 111.345 111.675 111.605 ;
        RECT 110.975 109.065 111.675 109.325 ;
        RECT 110.975 106.785 111.675 107.045 ;
        RECT 110.975 104.505 111.675 104.765 ;
        RECT 110.975 102.225 111.675 102.485 ;
        RECT 110.975 99.945 111.675 100.205 ;
        RECT 110.975 97.665 111.675 97.925 ;
        RECT 110.975 95.385 111.675 95.645 ;
        RECT 110.975 93.105 111.675 93.365 ;
        RECT 110.975 90.825 111.675 91.085 ;
        RECT 110.975 88.545 111.675 88.805 ;
        RECT 110.975 86.265 111.675 86.525 ;
        RECT 110.975 83.985 111.675 84.245 ;
        RECT 110.975 81.705 111.675 81.965 ;
        RECT 110.975 79.425 111.675 79.685 ;
        RECT 110.975 77.145 111.675 77.405 ;
        RECT 110.975 74.865 111.675 75.125 ;
        RECT 110.975 72.585 111.675 72.845 ;
        RECT 110.975 70.305 111.675 70.565 ;
        RECT 111.845 68.460 112.175 138.695 ;
        RECT 112.345 136.425 113.045 136.685 ;
        RECT 112.345 134.145 113.045 134.405 ;
        RECT 112.345 131.865 113.045 132.125 ;
        RECT 112.345 129.585 113.045 129.845 ;
        RECT 112.345 127.305 113.045 127.565 ;
        RECT 112.345 125.025 113.045 125.285 ;
        RECT 112.345 122.745 113.045 123.005 ;
        RECT 112.345 120.465 113.045 120.725 ;
        RECT 112.345 118.185 113.045 118.445 ;
        RECT 112.345 115.905 113.045 116.165 ;
        RECT 112.345 113.625 113.045 113.885 ;
        RECT 113.785 113.505 114.075 164.440 ;
        RECT 121.780 164.400 125.910 164.690 ;
        RECT 114.865 117.845 117.625 118.135 ;
        RECT 114.865 114.295 115.155 117.845 ;
        RECT 116.100 117.475 116.390 117.845 ;
        RECT 115.895 117.245 116.595 117.475 ;
        RECT 115.375 115.930 115.705 117.170 ;
        RECT 116.100 117.045 116.390 117.245 ;
        RECT 115.895 116.815 116.595 117.045 ;
        RECT 116.785 116.815 117.075 117.845 ;
        RECT 115.895 116.370 116.595 116.630 ;
        RECT 115.895 115.940 116.595 116.200 ;
        RECT 115.895 115.510 116.595 115.770 ;
        RECT 115.895 115.095 116.595 115.325 ;
        RECT 116.100 114.895 116.390 115.095 ;
        RECT 115.895 114.665 116.595 114.895 ;
        RECT 116.100 114.295 116.390 114.665 ;
        RECT 116.785 114.295 117.075 115.325 ;
        RECT 117.335 114.840 117.625 117.845 ;
        RECT 118.135 117.610 121.195 117.900 ;
        RECT 118.135 114.840 118.425 117.610 ;
        RECT 118.685 114.860 118.975 117.610 ;
        RECT 119.485 117.240 119.775 117.610 ;
        RECT 119.165 117.010 120.165 117.240 ;
        RECT 119.485 116.810 119.775 117.010 ;
        RECT 119.165 116.580 120.165 116.810 ;
        RECT 119.485 116.380 119.775 116.580 ;
        RECT 119.165 116.150 120.165 116.380 ;
        RECT 119.485 115.950 119.775 116.150 ;
        RECT 119.165 115.720 120.165 115.950 ;
        RECT 119.485 115.520 119.775 115.720 ;
        RECT 119.165 115.290 120.165 115.520 ;
        RECT 119.485 115.090 119.775 115.290 ;
        RECT 120.905 115.185 121.195 117.610 ;
        RECT 121.780 115.185 122.070 164.400 ;
        RECT 122.330 159.660 122.620 164.400 ;
        RECT 122.810 163.785 123.510 164.045 ;
        RECT 122.810 161.505 123.510 161.765 ;
        RECT 122.810 159.225 123.510 159.485 ;
        RECT 122.330 157.380 122.620 159.050 ;
        RECT 122.810 156.945 123.510 157.205 ;
        RECT 122.330 155.100 122.620 156.770 ;
        RECT 122.810 154.665 123.510 154.925 ;
        RECT 122.330 152.820 122.620 154.490 ;
        RECT 122.810 152.385 123.510 152.645 ;
        RECT 122.330 150.540 122.620 152.210 ;
        RECT 122.810 150.105 123.510 150.365 ;
        RECT 122.330 148.260 122.620 149.930 ;
        RECT 122.810 147.825 123.510 148.085 ;
        RECT 122.330 145.980 122.620 147.650 ;
        RECT 122.810 145.545 123.510 145.805 ;
        RECT 122.330 143.700 122.620 145.370 ;
        RECT 122.810 143.265 123.510 143.525 ;
        RECT 122.330 141.420 122.620 143.090 ;
        RECT 122.810 140.985 123.510 141.245 ;
        RECT 122.330 139.140 122.620 140.810 ;
        RECT 122.810 138.705 123.510 138.965 ;
        RECT 122.330 136.860 122.620 138.530 ;
        RECT 122.810 136.425 123.510 136.685 ;
        RECT 122.330 134.580 122.620 136.250 ;
        RECT 122.810 134.145 123.510 134.405 ;
        RECT 122.330 132.300 122.620 133.970 ;
        RECT 122.810 131.865 123.510 132.125 ;
        RECT 122.330 130.020 122.620 131.690 ;
        RECT 122.810 129.585 123.510 129.845 ;
        RECT 122.330 127.740 122.620 129.410 ;
        RECT 122.810 127.305 123.510 127.565 ;
        RECT 122.330 125.460 122.620 127.130 ;
        RECT 122.810 125.025 123.510 125.285 ;
        RECT 122.330 123.180 122.620 124.850 ;
        RECT 122.810 122.745 123.510 123.005 ;
        RECT 122.330 120.900 122.620 122.570 ;
        RECT 122.810 120.465 123.510 120.725 ;
        RECT 122.330 118.620 122.620 120.290 ;
        RECT 122.810 118.185 123.510 118.445 ;
        RECT 122.330 116.340 122.620 118.010 ;
        RECT 122.810 115.905 123.510 116.165 ;
        RECT 119.165 114.860 120.165 115.090 ;
        RECT 117.335 114.295 118.425 114.840 ;
        RECT 119.485 114.660 119.775 114.860 ;
        RECT 119.165 114.430 120.165 114.660 ;
        RECT 114.865 114.005 118.425 114.295 ;
        RECT 118.135 113.800 118.425 114.005 ;
        RECT 119.165 113.985 120.165 114.245 ;
        RECT 118.135 113.570 120.165 113.800 ;
        RECT 113.785 113.215 117.625 113.505 ;
        RECT 112.345 111.345 113.045 111.605 ;
        RECT 113.785 111.385 115.155 113.215 ;
        RECT 115.415 112.145 115.705 113.215 ;
        RECT 116.100 112.805 116.390 113.215 ;
        RECT 115.895 112.575 116.595 112.805 ;
        RECT 116.100 112.375 116.390 112.575 ;
        RECT 115.895 112.145 116.595 112.375 ;
        RECT 115.895 111.700 116.595 111.960 ;
        RECT 112.345 109.065 113.045 109.325 ;
        RECT 112.345 106.785 113.045 107.045 ;
        RECT 112.345 104.505 113.045 104.765 ;
        RECT 112.345 102.225 113.045 102.485 ;
        RECT 112.345 99.945 113.045 100.205 ;
        RECT 112.345 97.665 113.045 97.925 ;
        RECT 112.345 95.385 113.045 95.645 ;
        RECT 112.345 93.105 113.045 93.365 ;
        RECT 112.345 90.825 113.045 91.085 ;
        RECT 112.345 88.545 113.045 88.805 ;
        RECT 112.345 86.265 113.045 86.525 ;
        RECT 112.345 83.985 113.045 84.245 ;
        RECT 112.345 81.705 113.045 81.965 ;
        RECT 112.345 79.425 113.045 79.685 ;
        RECT 113.785 79.305 114.075 111.385 ;
        RECT 114.865 109.585 115.155 111.385 ;
        RECT 115.895 111.270 116.595 111.530 ;
        RECT 115.895 110.840 116.595 111.100 ;
        RECT 115.415 109.585 115.705 110.655 ;
        RECT 115.895 110.425 116.595 110.655 ;
        RECT 116.100 110.225 116.390 110.425 ;
        RECT 115.895 109.995 116.595 110.225 ;
        RECT 116.100 109.585 116.390 109.995 ;
        RECT 116.785 109.870 117.115 111.515 ;
        RECT 117.335 109.585 117.625 113.215 ;
        RECT 114.865 109.295 117.625 109.585 ;
        RECT 118.135 109.760 118.425 113.570 ;
        RECT 119.165 113.125 120.165 113.385 ;
        RECT 120.355 113.140 120.685 114.235 ;
        RECT 120.905 113.185 122.070 115.185 ;
        RECT 122.330 114.060 122.620 115.730 ;
        RECT 122.810 113.625 123.510 113.885 ;
        RECT 119.165 112.710 120.165 112.940 ;
        RECT 119.485 112.510 119.775 112.710 ;
        RECT 118.685 109.760 118.975 112.510 ;
        RECT 119.165 112.280 120.165 112.510 ;
        RECT 119.485 112.080 119.775 112.280 ;
        RECT 119.165 111.850 120.165 112.080 ;
        RECT 119.485 111.650 119.775 111.850 ;
        RECT 119.165 111.420 120.165 111.650 ;
        RECT 119.485 111.220 119.775 111.420 ;
        RECT 119.165 110.990 120.165 111.220 ;
        RECT 119.485 110.790 119.775 110.990 ;
        RECT 119.165 110.560 120.165 110.790 ;
        RECT 119.485 110.360 119.775 110.560 ;
        RECT 119.165 110.130 120.165 110.360 ;
        RECT 119.485 109.760 119.775 110.130 ;
        RECT 120.905 109.760 121.195 113.185 ;
        RECT 118.135 109.470 121.195 109.760 ;
        RECT 114.865 83.645 117.625 83.935 ;
        RECT 114.865 80.095 115.155 83.645 ;
        RECT 116.100 83.275 116.390 83.645 ;
        RECT 115.895 83.045 116.595 83.275 ;
        RECT 115.375 81.730 115.705 82.970 ;
        RECT 116.100 82.845 116.390 83.045 ;
        RECT 115.895 82.615 116.595 82.845 ;
        RECT 116.785 82.615 117.075 83.645 ;
        RECT 115.895 82.170 116.595 82.430 ;
        RECT 115.895 81.740 116.595 82.000 ;
        RECT 115.895 81.310 116.595 81.570 ;
        RECT 115.895 80.895 116.595 81.125 ;
        RECT 116.100 80.695 116.390 80.895 ;
        RECT 115.895 80.465 116.595 80.695 ;
        RECT 116.100 80.095 116.390 80.465 ;
        RECT 116.785 80.095 117.075 81.125 ;
        RECT 117.335 80.640 117.625 83.645 ;
        RECT 118.135 83.410 121.195 83.700 ;
        RECT 118.135 80.640 118.425 83.410 ;
        RECT 118.685 80.660 118.975 83.410 ;
        RECT 119.485 83.040 119.775 83.410 ;
        RECT 119.165 82.810 120.165 83.040 ;
        RECT 119.485 82.610 119.775 82.810 ;
        RECT 119.165 82.380 120.165 82.610 ;
        RECT 119.485 82.180 119.775 82.380 ;
        RECT 119.165 81.950 120.165 82.180 ;
        RECT 119.485 81.750 119.775 81.950 ;
        RECT 119.165 81.520 120.165 81.750 ;
        RECT 119.485 81.320 119.775 81.520 ;
        RECT 119.165 81.090 120.165 81.320 ;
        RECT 119.485 80.890 119.775 81.090 ;
        RECT 119.165 80.660 120.165 80.890 ;
        RECT 117.335 80.095 118.425 80.640 ;
        RECT 119.485 80.460 119.775 80.660 ;
        RECT 119.165 80.230 120.165 80.460 ;
        RECT 114.865 79.805 118.425 80.095 ;
        RECT 118.135 79.600 118.425 79.805 ;
        RECT 119.165 79.785 120.165 80.045 ;
        RECT 118.135 79.370 120.165 79.600 ;
        RECT 113.785 79.015 117.625 79.305 ;
        RECT 112.345 77.145 113.045 77.405 ;
        RECT 113.785 77.185 115.155 79.015 ;
        RECT 115.415 77.945 115.705 79.015 ;
        RECT 116.100 78.605 116.390 79.015 ;
        RECT 115.895 78.375 116.595 78.605 ;
        RECT 116.100 78.175 116.390 78.375 ;
        RECT 115.895 77.945 116.595 78.175 ;
        RECT 115.895 77.500 116.595 77.760 ;
        RECT 112.345 74.865 113.045 75.125 ;
        RECT 112.345 72.585 113.045 72.845 ;
        RECT 112.345 70.305 113.045 70.565 ;
        RECT 109.605 68.025 110.305 68.285 ;
        RECT 110.975 68.025 111.675 68.285 ;
        RECT 112.345 68.025 113.045 68.285 ;
        RECT 109.605 65.745 110.305 66.005 ;
        RECT 109.605 63.465 110.305 63.725 ;
        RECT 110.495 63.070 110.785 67.850 ;
        RECT 110.975 65.745 111.675 66.005 ;
        RECT 110.975 63.465 111.675 63.725 ;
        RECT 111.865 63.070 112.155 67.850 ;
        RECT 112.345 65.745 113.045 66.005 ;
        RECT 112.345 63.465 113.045 63.725 ;
        RECT 113.785 63.070 114.075 77.185 ;
        RECT 114.865 75.385 115.155 77.185 ;
        RECT 115.895 77.070 116.595 77.330 ;
        RECT 115.895 76.640 116.595 76.900 ;
        RECT 115.415 75.385 115.705 76.455 ;
        RECT 115.895 76.225 116.595 76.455 ;
        RECT 116.100 76.025 116.390 76.225 ;
        RECT 115.895 75.795 116.595 76.025 ;
        RECT 116.100 75.385 116.390 75.795 ;
        RECT 116.785 75.670 117.115 77.315 ;
        RECT 117.335 75.385 117.625 79.015 ;
        RECT 114.865 75.095 117.625 75.385 ;
        RECT 118.135 75.560 118.425 79.370 ;
        RECT 119.165 78.925 120.165 79.185 ;
        RECT 120.355 78.940 120.685 80.035 ;
        RECT 120.905 79.185 121.195 83.410 ;
        RECT 121.780 79.185 122.070 113.185 ;
        RECT 122.330 111.780 122.620 113.450 ;
        RECT 122.810 111.345 123.510 111.605 ;
        RECT 122.330 109.500 122.620 111.170 ;
        RECT 122.810 109.065 123.510 109.325 ;
        RECT 122.330 107.220 122.620 108.890 ;
        RECT 122.810 106.785 123.510 107.045 ;
        RECT 122.330 104.940 122.620 106.610 ;
        RECT 122.810 104.505 123.510 104.765 ;
        RECT 122.330 102.660 122.620 104.330 ;
        RECT 122.810 102.225 123.510 102.485 ;
        RECT 122.330 100.380 122.620 102.050 ;
        RECT 122.810 99.945 123.510 100.205 ;
        RECT 122.330 98.100 122.620 99.770 ;
        RECT 122.810 97.665 123.510 97.925 ;
        RECT 122.330 95.820 122.620 97.490 ;
        RECT 122.810 95.385 123.510 95.645 ;
        RECT 122.330 93.540 122.620 95.210 ;
        RECT 122.810 93.105 123.510 93.365 ;
        RECT 122.330 91.260 122.620 92.930 ;
        RECT 122.810 90.825 123.510 91.085 ;
        RECT 122.330 88.790 122.620 90.650 ;
        RECT 122.810 88.790 123.510 88.805 ;
        RECT 122.330 88.560 123.510 88.790 ;
        RECT 122.330 86.510 122.620 88.560 ;
        RECT 122.810 88.545 123.510 88.560 ;
        RECT 122.810 86.510 123.510 86.525 ;
        RECT 122.330 86.280 123.510 86.510 ;
        RECT 122.330 84.420 122.620 86.280 ;
        RECT 122.810 86.265 123.510 86.280 ;
        RECT 122.810 83.985 123.510 84.245 ;
        RECT 122.330 79.860 122.620 83.810 ;
        RECT 123.680 82.520 124.010 163.910 ;
        RECT 124.180 163.785 124.880 164.045 ;
        RECT 124.180 161.505 124.880 161.765 ;
        RECT 125.070 159.660 125.360 164.400 ;
        RECT 124.180 159.225 124.880 159.485 ;
        RECT 125.070 157.380 125.360 159.050 ;
        RECT 124.180 156.945 124.880 157.205 ;
        RECT 125.070 155.100 125.360 156.770 ;
        RECT 124.180 154.665 124.880 154.925 ;
        RECT 125.070 152.820 125.360 154.490 ;
        RECT 124.180 152.385 124.880 152.645 ;
        RECT 125.070 150.540 125.360 152.210 ;
        RECT 124.180 150.105 124.880 150.365 ;
        RECT 125.070 148.260 125.360 149.930 ;
        RECT 124.180 147.825 124.880 148.085 ;
        RECT 125.070 145.980 125.360 147.650 ;
        RECT 124.180 145.545 124.880 145.805 ;
        RECT 125.070 143.700 125.360 145.370 ;
        RECT 124.180 143.265 124.880 143.525 ;
        RECT 125.070 141.420 125.360 143.090 ;
        RECT 124.180 140.985 124.880 141.245 ;
        RECT 125.070 139.140 125.360 140.810 ;
        RECT 124.180 138.705 124.880 138.965 ;
        RECT 125.070 136.860 125.360 138.530 ;
        RECT 124.180 136.425 124.880 136.685 ;
        RECT 125.070 134.580 125.360 136.250 ;
        RECT 124.180 134.145 124.880 134.405 ;
        RECT 125.070 132.300 125.360 133.970 ;
        RECT 124.180 131.865 124.880 132.125 ;
        RECT 125.070 130.020 125.360 131.690 ;
        RECT 124.180 129.585 124.880 129.845 ;
        RECT 125.070 127.740 125.360 129.410 ;
        RECT 124.180 127.305 124.880 127.565 ;
        RECT 125.070 125.460 125.360 127.130 ;
        RECT 124.180 125.025 124.880 125.285 ;
        RECT 125.070 123.180 125.360 124.850 ;
        RECT 124.180 122.745 124.880 123.005 ;
        RECT 125.070 120.900 125.360 122.570 ;
        RECT 124.180 120.465 124.880 120.725 ;
        RECT 125.070 118.620 125.360 120.290 ;
        RECT 124.180 118.185 124.880 118.445 ;
        RECT 125.070 116.340 125.360 118.010 ;
        RECT 124.180 115.905 124.880 116.165 ;
        RECT 125.070 114.060 125.360 115.730 ;
        RECT 124.180 113.625 124.880 113.885 ;
        RECT 125.070 111.780 125.360 113.450 ;
        RECT 124.180 111.345 124.880 111.605 ;
        RECT 125.070 109.500 125.360 111.170 ;
        RECT 124.180 109.065 124.880 109.325 ;
        RECT 125.070 107.220 125.360 108.890 ;
        RECT 124.180 106.785 124.880 107.045 ;
        RECT 125.070 104.940 125.360 106.610 ;
        RECT 124.180 104.505 124.880 104.765 ;
        RECT 125.070 102.660 125.360 104.330 ;
        RECT 124.180 102.225 124.880 102.485 ;
        RECT 125.070 100.380 125.360 102.050 ;
        RECT 124.180 99.945 124.880 100.205 ;
        RECT 125.070 98.100 125.360 99.770 ;
        RECT 124.180 97.665 124.880 97.925 ;
        RECT 125.070 95.820 125.360 97.490 ;
        RECT 124.180 95.385 124.880 95.645 ;
        RECT 125.070 93.540 125.360 95.210 ;
        RECT 124.180 93.105 124.880 93.365 ;
        RECT 125.070 91.260 125.360 92.930 ;
        RECT 124.180 90.825 124.880 91.085 ;
        RECT 124.180 88.790 124.880 88.805 ;
        RECT 125.070 88.790 125.360 90.650 ;
        RECT 124.180 88.560 125.360 88.790 ;
        RECT 124.180 88.545 124.880 88.560 ;
        RECT 124.180 86.510 124.880 86.525 ;
        RECT 125.070 86.510 125.360 88.560 ;
        RECT 124.180 86.280 125.360 86.510 ;
        RECT 124.180 86.265 124.880 86.280 ;
        RECT 124.180 84.230 124.880 84.245 ;
        RECT 125.070 84.230 125.360 86.280 ;
        RECT 124.180 84.000 125.360 84.230 ;
        RECT 124.180 83.985 124.880 84.000 ;
        RECT 122.810 81.705 123.510 81.965 ;
        RECT 124.180 81.950 124.880 81.965 ;
        RECT 125.070 81.950 125.360 84.000 ;
        RECT 124.180 81.720 125.360 81.950 ;
        RECT 124.180 81.705 124.880 81.720 ;
        RECT 122.810 79.425 123.510 79.685 ;
        RECT 124.180 79.425 124.880 79.685 ;
        RECT 119.165 78.510 120.165 78.740 ;
        RECT 119.485 78.310 119.775 78.510 ;
        RECT 118.685 75.560 118.975 78.310 ;
        RECT 119.165 78.080 120.165 78.310 ;
        RECT 119.485 77.880 119.775 78.080 ;
        RECT 119.165 77.650 120.165 77.880 ;
        RECT 119.485 77.450 119.775 77.650 ;
        RECT 119.165 77.220 120.165 77.450 ;
        RECT 119.485 77.020 119.775 77.220 ;
        RECT 120.905 77.185 122.070 79.185 ;
        RECT 119.165 76.790 120.165 77.020 ;
        RECT 119.485 76.590 119.775 76.790 ;
        RECT 119.165 76.360 120.165 76.590 ;
        RECT 119.485 76.160 119.775 76.360 ;
        RECT 119.165 75.930 120.165 76.160 ;
        RECT 119.485 75.560 119.775 75.930 ;
        RECT 120.905 75.560 121.195 77.185 ;
        RECT 121.780 76.790 122.070 77.185 ;
        RECT 122.330 76.790 122.620 79.250 ;
        RECT 122.810 77.145 123.510 77.405 ;
        RECT 123.700 76.790 123.990 79.250 ;
        RECT 124.180 77.145 124.880 77.405 ;
        RECT 125.070 76.790 125.360 81.720 ;
        RECT 125.620 76.790 125.910 164.400 ;
        RECT 121.780 76.500 125.910 76.790 ;
        RECT 118.135 75.270 121.195 75.560 ;
        RECT 108.575 62.780 114.075 63.070 ;
        RECT 114.715 70.330 117.475 70.610 ;
        RECT 114.715 70.320 123.885 70.330 ;
        RECT 114.715 60.150 115.005 70.320 ;
        RECT 115.745 69.665 116.445 69.925 ;
        RECT 115.225 63.260 115.555 69.440 ;
        RECT 116.635 67.820 116.925 70.320 ;
        RECT 117.185 70.040 123.885 70.320 ;
        RECT 117.185 67.810 118.700 70.040 ;
        RECT 118.960 68.970 119.250 70.040 ;
        RECT 119.440 69.385 120.140 69.645 ;
        RECT 119.440 68.955 120.140 69.215 ;
        RECT 119.440 68.525 120.140 68.785 ;
        RECT 119.440 68.110 120.140 68.370 ;
        RECT 115.745 67.385 116.445 67.645 ;
        RECT 115.745 65.105 116.445 65.365 ;
        RECT 115.745 62.825 116.445 63.085 ;
        RECT 115.745 60.545 116.445 60.805 ;
        RECT 116.635 60.150 116.925 62.650 ;
        RECT 117.185 60.150 117.475 67.810 ;
        RECT 118.410 65.550 118.700 67.810 ;
        RECT 119.440 67.665 120.140 67.925 ;
        RECT 119.440 67.250 120.140 67.510 ;
        RECT 120.330 67.250 120.660 69.730 ;
        RECT 121.675 68.970 121.965 70.040 ;
        RECT 122.360 69.630 122.650 70.040 ;
        RECT 122.155 69.400 122.855 69.630 ;
        RECT 122.360 69.200 122.650 69.400 ;
        RECT 122.155 68.970 122.855 69.200 ;
        RECT 122.155 68.525 122.855 68.785 ;
        RECT 122.155 68.095 122.855 68.355 ;
        RECT 122.155 67.665 122.855 67.925 ;
        RECT 122.155 67.235 122.855 67.495 ;
        RECT 123.045 67.250 123.375 69.805 ;
        RECT 119.440 66.805 120.140 67.065 ;
        RECT 122.155 66.805 122.855 67.065 ;
        RECT 118.960 65.550 119.250 66.620 ;
        RECT 119.440 66.375 120.140 66.635 ;
        RECT 119.440 65.945 120.140 66.205 ;
        RECT 121.675 65.550 121.965 66.620 ;
        RECT 122.155 66.390 122.855 66.620 ;
        RECT 122.360 66.190 122.650 66.390 ;
        RECT 122.155 65.960 122.855 66.190 ;
        RECT 122.360 65.550 122.650 65.960 ;
        RECT 123.595 65.550 123.885 70.040 ;
        RECT 118.410 65.260 123.885 65.550 ;
        RECT 124.395 70.000 127.155 70.290 ;
        RECT 114.715 59.860 117.475 60.150 ;
        RECT 118.410 64.750 123.885 65.040 ;
        RECT 118.410 60.340 118.700 64.750 ;
        RECT 118.960 63.720 119.250 64.750 ;
        RECT 119.440 64.135 120.140 64.395 ;
        RECT 119.440 63.705 120.140 63.965 ;
        RECT 119.440 63.275 120.140 63.535 ;
        RECT 120.330 63.375 120.770 64.465 ;
        RECT 121.675 63.720 121.965 64.750 ;
        RECT 122.360 64.380 122.650 64.750 ;
        RECT 122.155 64.150 122.855 64.380 ;
        RECT 122.360 63.950 122.650 64.150 ;
        RECT 122.155 63.720 122.855 63.950 ;
        RECT 119.440 62.860 120.140 63.120 ;
        RECT 119.440 62.415 120.140 62.675 ;
        RECT 119.440 62.000 120.140 62.260 ;
        RECT 120.330 62.000 120.660 63.375 ;
        RECT 122.155 63.275 122.855 63.535 ;
        RECT 123.595 63.115 123.885 64.750 ;
        RECT 124.395 63.115 124.685 70.000 ;
        RECT 124.945 66.390 125.235 70.000 ;
        RECT 125.425 69.385 126.125 69.645 ;
        RECT 125.425 68.955 126.125 69.215 ;
        RECT 125.425 68.525 126.125 68.785 ;
        RECT 125.425 68.095 126.125 68.355 ;
        RECT 125.425 67.665 126.125 67.925 ;
        RECT 125.425 67.235 126.125 67.495 ;
        RECT 125.425 66.805 126.125 67.065 ;
        RECT 125.425 66.375 126.125 66.635 ;
        RECT 125.425 65.945 126.125 66.205 ;
        RECT 125.425 65.515 126.125 65.775 ;
        RECT 125.425 65.085 126.125 65.345 ;
        RECT 125.425 64.655 126.125 64.915 ;
        RECT 126.315 64.670 126.610 65.760 ;
        RECT 125.425 64.225 126.125 64.485 ;
        RECT 122.155 62.845 122.855 63.105 ;
        RECT 122.155 62.415 122.855 62.675 ;
        RECT 122.155 61.985 122.855 62.245 ;
        RECT 119.440 61.555 120.140 61.815 ;
        RECT 122.155 61.555 122.855 61.815 ;
        RECT 118.960 60.340 119.250 61.370 ;
        RECT 119.440 61.125 120.140 61.385 ;
        RECT 119.440 60.695 120.140 60.955 ;
        RECT 121.675 60.340 121.965 61.370 ;
        RECT 122.155 61.140 122.855 61.370 ;
        RECT 122.360 60.940 122.650 61.140 ;
        RECT 122.155 60.710 122.855 60.940 ;
        RECT 122.360 60.340 122.650 60.710 ;
        RECT 123.045 60.685 123.375 63.090 ;
        RECT 123.595 61.975 124.685 63.115 ;
        RECT 123.595 60.340 123.885 61.975 ;
        RECT 118.410 60.050 123.885 60.340 ;
        RECT 124.395 60.430 124.685 61.975 ;
        RECT 124.945 60.430 125.235 64.040 ;
        RECT 125.425 63.795 126.125 64.055 ;
        RECT 125.425 63.365 126.125 63.625 ;
        RECT 125.425 62.935 126.125 63.195 ;
        RECT 125.425 62.505 126.125 62.765 ;
        RECT 125.425 62.075 126.125 62.335 ;
        RECT 125.425 61.645 126.125 61.905 ;
        RECT 125.425 61.215 126.125 61.475 ;
        RECT 125.425 60.785 126.125 61.045 ;
        RECT 126.865 60.430 127.155 70.000 ;
        RECT 124.395 60.140 127.155 60.430 ;
      LAYER via ;
        RECT 108.245 173.605 108.505 173.865 ;
        RECT 108.565 173.605 108.825 173.865 ;
        RECT 108.885 173.605 109.145 173.865 ;
        RECT 112.095 173.605 112.355 173.865 ;
        RECT 112.415 173.605 112.675 173.865 ;
        RECT 112.735 173.605 112.995 173.865 ;
        RECT 108.245 172.935 108.505 173.195 ;
        RECT 108.565 172.935 108.825 173.195 ;
        RECT 108.885 172.935 109.145 173.195 ;
        RECT 108.245 172.505 108.505 172.765 ;
        RECT 108.565 172.505 108.825 172.765 ;
        RECT 108.885 172.505 109.145 172.765 ;
        RECT 110.240 172.840 110.500 173.100 ;
        RECT 110.240 172.520 110.500 172.780 ;
        RECT 108.245 172.075 108.505 172.335 ;
        RECT 108.565 172.075 108.825 172.335 ;
        RECT 108.885 172.075 109.145 172.335 ;
        RECT 108.245 171.645 108.505 171.905 ;
        RECT 108.565 171.645 108.825 171.905 ;
        RECT 108.885 171.645 109.145 171.905 ;
        RECT 112.095 172.935 112.355 173.195 ;
        RECT 112.415 172.935 112.675 173.195 ;
        RECT 112.735 172.935 112.995 173.195 ;
        RECT 112.095 172.505 112.355 172.765 ;
        RECT 112.415 172.505 112.675 172.765 ;
        RECT 112.735 172.505 112.995 172.765 ;
        RECT 112.095 172.075 112.355 172.335 ;
        RECT 112.415 172.075 112.675 172.335 ;
        RECT 112.735 172.075 112.995 172.335 ;
        RECT 111.615 171.645 111.875 171.905 ;
        RECT 111.935 171.645 112.195 171.905 ;
        RECT 112.255 171.645 112.515 171.905 ;
        RECT 112.575 171.645 112.835 171.905 ;
        RECT 112.895 171.645 113.155 171.905 ;
        RECT 113.215 171.645 113.475 171.905 ;
        RECT 108.245 171.215 108.505 171.475 ;
        RECT 108.565 171.215 108.825 171.475 ;
        RECT 108.885 171.215 109.145 171.475 ;
        RECT 112.095 171.215 112.355 171.475 ;
        RECT 112.415 171.215 112.675 171.475 ;
        RECT 112.735 171.215 112.995 171.475 ;
        RECT 108.245 170.785 108.505 171.045 ;
        RECT 108.565 170.785 108.825 171.045 ;
        RECT 108.885 170.785 109.145 171.045 ;
        RECT 111.615 170.785 111.875 171.045 ;
        RECT 111.935 170.785 112.195 171.045 ;
        RECT 112.255 170.785 112.515 171.045 ;
        RECT 112.575 170.785 112.835 171.045 ;
        RECT 112.895 170.785 113.155 171.045 ;
        RECT 113.215 170.785 113.475 171.045 ;
        RECT 108.245 170.355 108.505 170.615 ;
        RECT 108.565 170.355 108.825 170.615 ;
        RECT 108.885 170.355 109.145 170.615 ;
        RECT 112.095 170.355 112.355 170.615 ;
        RECT 112.415 170.355 112.675 170.615 ;
        RECT 112.735 170.355 112.995 170.615 ;
        RECT 108.245 169.925 108.505 170.185 ;
        RECT 108.565 169.925 108.825 170.185 ;
        RECT 108.885 169.925 109.145 170.185 ;
        RECT 108.245 169.495 108.505 169.755 ;
        RECT 108.565 169.495 108.825 169.755 ;
        RECT 108.885 169.495 109.145 169.755 ;
        RECT 112.095 169.925 112.355 170.185 ;
        RECT 112.415 169.925 112.675 170.185 ;
        RECT 112.735 169.925 112.995 170.185 ;
        RECT 112.095 169.495 112.355 169.755 ;
        RECT 112.415 169.495 112.675 169.755 ;
        RECT 112.735 169.495 112.995 169.755 ;
        RECT 108.245 168.825 108.505 169.085 ;
        RECT 108.565 168.825 108.825 169.085 ;
        RECT 108.885 168.825 109.145 169.085 ;
        RECT 112.095 168.825 112.355 169.085 ;
        RECT 112.415 168.825 112.675 169.085 ;
        RECT 112.735 168.825 112.995 169.085 ;
        RECT 109.665 164.455 109.925 164.715 ;
        RECT 109.985 164.455 110.245 164.715 ;
        RECT 111.035 164.455 111.295 164.715 ;
        RECT 111.355 164.455 111.615 164.715 ;
        RECT 112.405 164.455 112.665 164.715 ;
        RECT 112.725 164.455 112.985 164.715 ;
        RECT 57.200 151.205 57.460 151.465 ;
        RECT 57.520 151.205 57.780 151.465 ;
        RECT 57.840 151.205 58.100 151.465 ;
        RECT 60.790 151.205 61.050 151.465 ;
        RECT 61.110 151.205 61.370 151.465 ;
        RECT 61.430 151.205 61.690 151.465 ;
        RECT 57.200 141.295 57.460 141.555 ;
        RECT 57.520 141.295 57.780 141.555 ;
        RECT 57.840 141.295 58.100 141.555 ;
        RECT 57.200 139.015 57.460 139.275 ;
        RECT 57.520 139.015 57.780 139.275 ;
        RECT 57.840 139.015 58.100 139.275 ;
        RECT 57.200 136.735 57.460 136.995 ;
        RECT 57.520 136.735 57.780 136.995 ;
        RECT 57.840 136.735 58.100 136.995 ;
        RECT 57.200 134.455 57.460 134.715 ;
        RECT 57.520 134.455 57.780 134.715 ;
        RECT 57.840 134.455 58.100 134.715 ;
        RECT 57.200 132.175 57.460 132.435 ;
        RECT 57.520 132.175 57.780 132.435 ;
        RECT 57.840 132.175 58.100 132.435 ;
        RECT 60.790 150.535 61.050 150.795 ;
        RECT 61.110 150.535 61.370 150.795 ;
        RECT 61.430 150.535 61.690 150.795 ;
        RECT 60.790 149.755 61.050 150.015 ;
        RECT 61.110 149.755 61.370 150.015 ;
        RECT 61.430 149.755 61.690 150.015 ;
        RECT 60.790 148.975 61.050 149.235 ;
        RECT 61.110 148.975 61.370 149.235 ;
        RECT 61.430 148.975 61.690 149.235 ;
        RECT 61.965 148.540 62.225 148.800 ;
        RECT 61.965 148.220 62.225 148.480 ;
        RECT 61.965 147.900 62.225 148.160 ;
        RECT 60.790 146.695 61.050 146.955 ;
        RECT 61.110 146.695 61.370 146.955 ;
        RECT 61.430 146.695 61.690 146.955 ;
        RECT 60.790 144.415 61.050 144.675 ;
        RECT 61.110 144.415 61.370 144.675 ;
        RECT 61.430 144.415 61.690 144.675 ;
        RECT 60.790 143.635 61.050 143.895 ;
        RECT 61.110 143.635 61.370 143.895 ;
        RECT 61.430 143.635 61.690 143.895 ;
        RECT 60.790 142.855 61.050 143.115 ;
        RECT 61.110 142.855 61.370 143.115 ;
        RECT 61.430 142.855 61.690 143.115 ;
        RECT 60.790 142.075 61.050 142.335 ;
        RECT 61.110 142.075 61.370 142.335 ;
        RECT 61.430 142.075 61.690 142.335 ;
        RECT 60.790 141.295 61.050 141.555 ;
        RECT 61.110 141.295 61.370 141.555 ;
        RECT 61.430 141.295 61.690 141.555 ;
        RECT 61.965 140.860 62.225 141.120 ;
        RECT 61.965 140.540 62.225 140.800 ;
        RECT 61.965 140.220 62.225 140.480 ;
        RECT 60.790 139.015 61.050 139.275 ;
        RECT 61.110 139.015 61.370 139.275 ;
        RECT 61.430 139.015 61.690 139.275 ;
        RECT 60.790 136.735 61.050 136.995 ;
        RECT 61.110 136.735 61.370 136.995 ;
        RECT 61.430 136.735 61.690 136.995 ;
        RECT 60.790 134.455 61.050 134.715 ;
        RECT 61.110 134.455 61.370 134.715 ;
        RECT 61.430 134.455 61.690 134.715 ;
        RECT 60.790 132.175 61.050 132.435 ;
        RECT 61.110 132.175 61.370 132.435 ;
        RECT 61.430 132.175 61.690 132.435 ;
        RECT 57.200 129.895 57.460 130.155 ;
        RECT 57.520 129.895 57.780 130.155 ;
        RECT 57.840 129.895 58.100 130.155 ;
        RECT 60.790 129.895 61.050 130.155 ;
        RECT 61.110 129.895 61.370 130.155 ;
        RECT 61.430 129.895 61.690 130.155 ;
        RECT 56.665 127.935 56.925 128.195 ;
        RECT 56.665 127.615 56.925 127.875 ;
        RECT 57.200 127.615 57.460 127.875 ;
        RECT 57.520 127.615 57.780 127.875 ;
        RECT 57.840 127.615 58.100 127.875 ;
        RECT 60.790 127.615 61.050 127.875 ;
        RECT 61.110 127.615 61.370 127.875 ;
        RECT 61.430 127.615 61.690 127.875 ;
        RECT 56.665 127.295 56.925 127.555 ;
        RECT 57.200 125.335 57.460 125.595 ;
        RECT 57.520 125.335 57.780 125.595 ;
        RECT 57.840 125.335 58.100 125.595 ;
        RECT 60.790 125.335 61.050 125.595 ;
        RECT 61.110 125.335 61.370 125.595 ;
        RECT 61.430 125.335 61.690 125.595 ;
        RECT 57.200 123.055 57.460 123.315 ;
        RECT 57.520 123.055 57.780 123.315 ;
        RECT 57.840 123.055 58.100 123.315 ;
        RECT 57.200 120.775 57.460 121.035 ;
        RECT 57.520 120.775 57.780 121.035 ;
        RECT 57.840 120.775 58.100 121.035 ;
        RECT 57.200 118.495 57.460 118.755 ;
        RECT 57.520 118.495 57.780 118.755 ;
        RECT 57.840 118.495 58.100 118.755 ;
        RECT 57.200 116.215 57.460 116.475 ;
        RECT 57.520 116.215 57.780 116.475 ;
        RECT 57.840 116.215 58.100 116.475 ;
        RECT 57.200 113.935 57.460 114.195 ;
        RECT 57.520 113.935 57.780 114.195 ;
        RECT 57.840 113.935 58.100 114.195 ;
        RECT 60.790 123.055 61.050 123.315 ;
        RECT 61.110 123.055 61.370 123.315 ;
        RECT 61.430 123.055 61.690 123.315 ;
        RECT 60.790 120.775 61.050 121.035 ;
        RECT 61.110 120.775 61.370 121.035 ;
        RECT 61.430 120.775 61.690 121.035 ;
        RECT 60.790 118.495 61.050 118.755 ;
        RECT 61.110 118.495 61.370 118.755 ;
        RECT 61.430 118.495 61.690 118.755 ;
        RECT 60.790 116.215 61.050 116.475 ;
        RECT 61.110 116.215 61.370 116.475 ;
        RECT 61.430 116.215 61.690 116.475 ;
        RECT 61.965 115.010 62.225 115.270 ;
        RECT 61.965 114.690 62.225 114.950 ;
        RECT 61.965 114.370 62.225 114.630 ;
        RECT 60.790 113.935 61.050 114.195 ;
        RECT 61.110 113.935 61.370 114.195 ;
        RECT 61.430 113.935 61.690 114.195 ;
        RECT 60.790 113.155 61.050 113.415 ;
        RECT 61.110 113.155 61.370 113.415 ;
        RECT 61.430 113.155 61.690 113.415 ;
        RECT 60.790 112.375 61.050 112.635 ;
        RECT 61.110 112.375 61.370 112.635 ;
        RECT 61.430 112.375 61.690 112.635 ;
        RECT 65.525 151.205 65.785 151.465 ;
        RECT 65.525 150.535 65.785 150.795 ;
        RECT 65.525 149.755 65.785 150.015 ;
        RECT 65.525 148.975 65.785 149.235 ;
        RECT 64.920 147.015 65.180 147.275 ;
        RECT 64.920 146.695 65.180 146.955 ;
        RECT 65.525 146.695 65.785 146.955 ;
        RECT 64.920 146.375 65.180 146.635 ;
        RECT 65.525 144.415 65.785 144.675 ;
        RECT 65.525 143.635 65.785 143.895 ;
        RECT 65.525 142.855 65.785 143.115 ;
        RECT 93.005 151.205 93.265 151.465 ;
        RECT 65.525 142.185 65.785 142.445 ;
        RECT 73.680 142.485 73.940 142.745 ;
        RECT 76.420 142.485 76.680 142.745 ;
        RECT 65.525 137.995 65.785 138.255 ;
        RECT 65.525 137.325 65.785 137.585 ;
        RECT 65.525 136.045 65.785 136.305 ;
        RECT 65.525 134.765 65.785 135.025 ;
        RECT 64.920 134.465 65.180 134.725 ;
        RECT 64.920 134.145 65.180 134.405 ;
        RECT 64.920 133.825 65.180 134.085 ;
        RECT 66.130 134.330 66.390 134.590 ;
        RECT 66.130 134.010 66.390 134.270 ;
        RECT 66.130 133.690 66.390 133.950 ;
        RECT 65.525 130.205 65.785 130.465 ;
        RECT 65.525 128.925 65.785 129.185 ;
        RECT 65.525 127.645 65.785 127.905 ;
        RECT 65.525 126.365 65.785 126.625 ;
        RECT 65.525 125.085 65.785 125.345 ;
        RECT 64.915 123.125 65.175 123.385 ;
        RECT 64.915 122.805 65.175 123.065 ;
        RECT 65.525 122.805 65.785 123.065 ;
        RECT 64.915 122.485 65.175 122.745 ;
        RECT 65.525 120.525 65.785 120.785 ;
        RECT 65.525 119.245 65.785 119.505 ;
        RECT 65.525 117.965 65.785 118.225 ;
        RECT 65.525 117.295 65.785 117.555 ;
        RECT 69.210 137.995 69.470 138.255 ;
        RECT 69.530 137.995 69.790 138.255 ;
        RECT 69.850 137.995 70.110 138.255 ;
        RECT 69.210 137.325 69.470 137.585 ;
        RECT 69.530 137.325 69.790 137.585 ;
        RECT 69.850 137.325 70.110 137.585 ;
        RECT 69.210 136.045 69.470 136.305 ;
        RECT 69.530 136.045 69.790 136.305 ;
        RECT 69.850 136.045 70.110 136.305 ;
        RECT 69.210 134.765 69.470 135.025 ;
        RECT 69.530 134.765 69.790 135.025 ;
        RECT 69.850 134.765 70.110 135.025 ;
        RECT 69.210 132.465 69.470 132.725 ;
        RECT 69.530 132.465 69.790 132.725 ;
        RECT 69.850 132.465 70.110 132.725 ;
        RECT 68.675 131.280 68.935 131.540 ;
        RECT 68.675 130.960 68.935 131.220 ;
        RECT 68.675 130.640 68.935 130.900 ;
        RECT 69.210 130.205 69.470 130.465 ;
        RECT 69.530 130.205 69.790 130.465 ;
        RECT 69.850 130.205 70.110 130.465 ;
        RECT 69.210 128.925 69.470 129.185 ;
        RECT 69.530 128.925 69.790 129.185 ;
        RECT 69.850 128.925 70.110 129.185 ;
        RECT 69.210 127.645 69.470 127.905 ;
        RECT 69.530 127.645 69.790 127.905 ;
        RECT 69.850 127.645 70.110 127.905 ;
        RECT 69.210 126.365 69.470 126.625 ;
        RECT 69.530 126.365 69.790 126.625 ;
        RECT 69.850 126.365 70.110 126.625 ;
        RECT 69.210 125.085 69.470 125.345 ;
        RECT 69.530 125.085 69.790 125.345 ;
        RECT 69.850 125.085 70.110 125.345 ;
        RECT 69.210 122.775 69.470 123.035 ;
        RECT 69.530 122.775 69.790 123.035 ;
        RECT 69.850 122.775 70.110 123.035 ;
        RECT 69.210 120.525 69.470 120.785 ;
        RECT 69.530 120.525 69.790 120.785 ;
        RECT 69.850 120.525 70.110 120.785 ;
        RECT 69.210 119.245 69.470 119.505 ;
        RECT 69.530 119.245 69.790 119.505 ;
        RECT 69.850 119.245 70.110 119.505 ;
        RECT 69.210 117.965 69.470 118.225 ;
        RECT 69.530 117.965 69.790 118.225 ;
        RECT 69.850 117.965 70.110 118.225 ;
        RECT 69.210 117.295 69.470 117.555 ;
        RECT 69.530 117.295 69.790 117.555 ;
        RECT 69.850 117.295 70.110 117.555 ;
        RECT 57.200 111.705 57.460 111.965 ;
        RECT 57.520 111.705 57.780 111.965 ;
        RECT 57.840 111.705 58.100 111.965 ;
        RECT 60.790 111.705 61.050 111.965 ;
        RECT 61.110 111.705 61.370 111.965 ;
        RECT 61.430 111.705 61.690 111.965 ;
        RECT 64.365 113.045 64.625 113.305 ;
        RECT 64.685 113.045 64.945 113.305 ;
        RECT 65.005 113.045 65.265 113.305 ;
        RECT 69.235 113.045 69.495 113.305 ;
        RECT 64.365 112.375 64.625 112.635 ;
        RECT 64.685 112.375 64.945 112.635 ;
        RECT 65.005 112.375 65.265 112.635 ;
        RECT 64.365 110.095 64.625 110.355 ;
        RECT 64.685 110.095 64.945 110.355 ;
        RECT 65.005 110.095 65.265 110.355 ;
        RECT 69.235 112.375 69.495 112.635 ;
        RECT 69.235 110.095 69.495 110.355 ;
        RECT 64.365 107.815 64.625 108.075 ;
        RECT 64.685 107.815 64.945 108.075 ;
        RECT 65.005 107.815 65.265 108.075 ;
        RECT 69.235 107.815 69.495 108.075 ;
        RECT 65.540 107.380 65.800 107.640 ;
        RECT 65.540 107.060 65.800 107.320 ;
        RECT 65.540 106.740 65.800 107.000 ;
        RECT 64.365 105.535 64.625 105.795 ;
        RECT 64.685 105.535 64.945 105.795 ;
        RECT 65.005 105.535 65.265 105.795 ;
        RECT 68.630 107.380 68.890 107.640 ;
        RECT 68.630 107.060 68.890 107.320 ;
        RECT 68.630 106.740 68.890 107.000 ;
        RECT 67.055 105.535 67.315 105.795 ;
        RECT 67.375 105.535 67.635 105.795 ;
        RECT 67.695 105.535 67.955 105.795 ;
        RECT 64.365 103.255 64.625 103.515 ;
        RECT 64.685 103.255 64.945 103.515 ;
        RECT 65.005 103.255 65.265 103.515 ;
        RECT 69.235 105.535 69.495 105.795 ;
        RECT 69.235 103.255 69.495 103.515 ;
        RECT 64.365 100.975 64.625 101.235 ;
        RECT 64.685 100.975 64.945 101.235 ;
        RECT 65.005 100.975 65.265 101.235 ;
        RECT 67.055 100.975 67.315 101.235 ;
        RECT 67.375 100.975 67.635 101.235 ;
        RECT 67.695 100.975 67.955 101.235 ;
        RECT 64.365 98.695 64.625 98.955 ;
        RECT 64.685 98.695 64.945 98.955 ;
        RECT 65.005 98.695 65.265 98.955 ;
        RECT 69.235 100.975 69.495 101.235 ;
        RECT 69.235 98.695 69.495 98.955 ;
        RECT 64.365 96.415 64.625 96.675 ;
        RECT 64.685 96.415 64.945 96.675 ;
        RECT 65.005 96.415 65.265 96.675 ;
        RECT 69.235 96.415 69.495 96.675 ;
        RECT 64.365 94.135 64.625 94.395 ;
        RECT 64.685 94.135 64.945 94.395 ;
        RECT 65.005 94.135 65.265 94.395 ;
        RECT 69.235 94.135 69.495 94.395 ;
        RECT 64.365 91.855 64.625 92.115 ;
        RECT 64.685 91.855 64.945 92.115 ;
        RECT 65.005 91.855 65.265 92.115 ;
        RECT 64.365 89.575 64.625 89.835 ;
        RECT 64.685 89.575 64.945 89.835 ;
        RECT 65.005 89.575 65.265 89.835 ;
        RECT 69.235 91.855 69.495 92.115 ;
        RECT 69.235 89.575 69.495 89.835 ;
        RECT 73.680 141.855 73.940 142.115 ;
        RECT 73.075 140.860 73.335 141.120 ;
        RECT 73.075 140.540 73.335 140.800 ;
        RECT 73.680 139.295 73.940 139.555 ;
        RECT 73.680 137.015 73.940 137.275 ;
        RECT 76.420 141.455 76.680 141.715 ;
        RECT 76.420 138.175 76.680 138.435 ;
        RECT 73.680 134.735 73.940 134.995 ;
        RECT 76.420 134.895 76.680 135.155 ;
        RECT 73.680 132.455 73.940 132.715 ;
        RECT 73.680 130.175 73.940 130.435 ;
        RECT 73.680 128.895 73.940 129.155 ;
        RECT 73.680 127.615 73.940 127.875 ;
        RECT 76.420 127.615 76.680 127.875 ;
        RECT 73.680 126.335 73.940 126.595 ;
        RECT 77.025 126.535 77.285 126.795 ;
        RECT 77.025 126.215 77.285 126.475 ;
        RECT 77.025 125.895 77.285 126.155 ;
        RECT 77.025 125.575 77.285 125.835 ;
        RECT 73.680 125.055 73.940 125.315 ;
        RECT 73.680 122.775 73.940 123.035 ;
        RECT 73.680 120.495 73.940 120.755 ;
        RECT 76.420 120.335 76.680 120.595 ;
        RECT 73.680 118.215 73.940 118.475 ;
        RECT 73.680 115.935 73.940 116.195 ;
        RECT 73.075 114.690 73.335 114.950 ;
        RECT 73.075 114.370 73.335 114.630 ;
        RECT 73.680 113.375 73.940 113.635 ;
        RECT 76.420 117.055 76.680 117.315 ;
        RECT 76.420 113.775 76.680 114.035 ;
        RECT 73.680 112.745 73.940 113.005 ;
        RECT 76.420 112.745 76.680 113.005 ;
        RECT 82.110 142.485 82.370 142.745 ;
        RECT 84.850 142.485 85.110 142.745 ;
        RECT 82.110 141.455 82.370 141.715 ;
        RECT 82.110 138.175 82.370 138.435 ;
        RECT 84.850 141.855 85.110 142.115 ;
        RECT 85.455 140.860 85.715 141.120 ;
        RECT 85.455 140.540 85.715 140.800 ;
        RECT 84.850 139.295 85.110 139.555 ;
        RECT 84.850 137.015 85.110 137.275 ;
        RECT 82.110 134.895 82.370 135.155 ;
        RECT 84.850 134.735 85.110 134.995 ;
        RECT 84.850 132.455 85.110 132.715 ;
        RECT 84.850 130.175 85.110 130.435 ;
        RECT 84.850 128.895 85.110 129.155 ;
        RECT 82.110 127.615 82.370 127.875 ;
        RECT 84.850 127.615 85.110 127.875 ;
        RECT 81.505 126.535 81.765 126.795 ;
        RECT 81.505 126.215 81.765 126.475 ;
        RECT 81.505 125.895 81.765 126.155 ;
        RECT 81.505 125.575 81.765 125.835 ;
        RECT 84.850 126.335 85.110 126.595 ;
        RECT 84.850 125.055 85.110 125.315 ;
        RECT 84.850 122.775 85.110 123.035 ;
        RECT 82.110 120.335 82.370 120.595 ;
        RECT 84.850 120.495 85.110 120.755 ;
        RECT 82.110 117.055 82.370 117.315 ;
        RECT 82.110 113.775 82.370 114.035 ;
        RECT 84.850 118.215 85.110 118.475 ;
        RECT 84.850 115.935 85.110 116.195 ;
        RECT 85.455 114.690 85.715 114.950 ;
        RECT 85.455 114.370 85.715 114.630 ;
        RECT 84.850 113.375 85.110 113.635 ;
        RECT 93.005 150.535 93.265 150.795 ;
        RECT 93.005 149.755 93.265 150.015 ;
        RECT 93.005 148.975 93.265 149.235 ;
        RECT 93.610 147.015 93.870 147.275 ;
        RECT 93.005 146.695 93.265 146.955 ;
        RECT 93.610 146.695 93.870 146.955 ;
        RECT 93.610 146.375 93.870 146.635 ;
        RECT 93.005 144.415 93.265 144.675 ;
        RECT 93.005 143.635 93.265 143.895 ;
        RECT 93.005 142.855 93.265 143.115 ;
        RECT 93.005 142.185 93.265 142.445 ;
        RECT 97.100 151.205 97.360 151.465 ;
        RECT 97.420 151.205 97.680 151.465 ;
        RECT 97.740 151.205 98.000 151.465 ;
        RECT 100.690 151.205 100.950 151.465 ;
        RECT 101.010 151.205 101.270 151.465 ;
        RECT 101.330 151.205 101.590 151.465 ;
        RECT 88.680 137.995 88.940 138.255 ;
        RECT 89.000 137.995 89.260 138.255 ;
        RECT 89.320 137.995 89.580 138.255 ;
        RECT 88.680 137.325 88.940 137.585 ;
        RECT 89.000 137.325 89.260 137.585 ;
        RECT 89.320 137.325 89.580 137.585 ;
        RECT 88.680 136.045 88.940 136.305 ;
        RECT 89.000 136.045 89.260 136.305 ;
        RECT 89.320 136.045 89.580 136.305 ;
        RECT 88.680 134.765 88.940 135.025 ;
        RECT 89.000 134.765 89.260 135.025 ;
        RECT 89.320 134.765 89.580 135.025 ;
        RECT 88.680 132.465 88.940 132.725 ;
        RECT 89.000 132.465 89.260 132.725 ;
        RECT 89.320 132.465 89.580 132.725 ;
        RECT 89.855 131.280 90.115 131.540 ;
        RECT 89.855 130.960 90.115 131.220 ;
        RECT 89.855 130.640 90.115 130.900 ;
        RECT 88.680 130.205 88.940 130.465 ;
        RECT 89.000 130.205 89.260 130.465 ;
        RECT 89.320 130.205 89.580 130.465 ;
        RECT 88.680 128.925 88.940 129.185 ;
        RECT 89.000 128.925 89.260 129.185 ;
        RECT 89.320 128.925 89.580 129.185 ;
        RECT 88.680 127.645 88.940 127.905 ;
        RECT 89.000 127.645 89.260 127.905 ;
        RECT 89.320 127.645 89.580 127.905 ;
        RECT 88.680 126.365 88.940 126.625 ;
        RECT 89.000 126.365 89.260 126.625 ;
        RECT 89.320 126.365 89.580 126.625 ;
        RECT 88.680 125.085 88.940 125.345 ;
        RECT 89.000 125.085 89.260 125.345 ;
        RECT 89.320 125.085 89.580 125.345 ;
        RECT 88.680 122.775 88.940 123.035 ;
        RECT 89.000 122.775 89.260 123.035 ;
        RECT 89.320 122.775 89.580 123.035 ;
        RECT 88.680 120.525 88.940 120.785 ;
        RECT 89.000 120.525 89.260 120.785 ;
        RECT 89.320 120.525 89.580 120.785 ;
        RECT 88.680 119.245 88.940 119.505 ;
        RECT 89.000 119.245 89.260 119.505 ;
        RECT 89.320 119.245 89.580 119.505 ;
        RECT 88.680 117.965 88.940 118.225 ;
        RECT 89.000 117.965 89.260 118.225 ;
        RECT 89.320 117.965 89.580 118.225 ;
        RECT 88.680 117.295 88.940 117.555 ;
        RECT 89.000 117.295 89.260 117.555 ;
        RECT 89.320 117.295 89.580 117.555 ;
        RECT 93.005 137.995 93.265 138.255 ;
        RECT 93.005 137.325 93.265 137.585 ;
        RECT 93.005 136.045 93.265 136.305 ;
        RECT 93.005 134.765 93.265 135.025 ;
        RECT 92.400 134.330 92.660 134.590 ;
        RECT 92.400 134.010 92.660 134.270 ;
        RECT 92.400 133.690 92.660 133.950 ;
        RECT 93.610 134.465 93.870 134.725 ;
        RECT 93.610 134.145 93.870 134.405 ;
        RECT 93.610 133.825 93.870 134.085 ;
        RECT 93.005 130.205 93.265 130.465 ;
        RECT 93.005 128.925 93.265 129.185 ;
        RECT 93.005 127.645 93.265 127.905 ;
        RECT 93.005 126.365 93.265 126.625 ;
        RECT 93.005 125.085 93.265 125.345 ;
        RECT 93.615 123.125 93.875 123.385 ;
        RECT 93.005 122.805 93.265 123.065 ;
        RECT 93.615 122.805 93.875 123.065 ;
        RECT 93.615 122.485 93.875 122.745 ;
        RECT 93.005 120.525 93.265 120.785 ;
        RECT 93.005 119.245 93.265 119.505 ;
        RECT 93.005 117.965 93.265 118.225 ;
        RECT 93.005 117.295 93.265 117.555 ;
        RECT 82.110 112.745 82.370 113.005 ;
        RECT 84.850 112.745 85.110 113.005 ;
        RECT 89.295 113.045 89.555 113.305 ;
        RECT 93.525 113.045 93.785 113.305 ;
        RECT 93.845 113.045 94.105 113.305 ;
        RECT 94.165 113.045 94.425 113.305 ;
        RECT 64.365 88.905 64.625 89.165 ;
        RECT 64.685 88.905 64.945 89.165 ;
        RECT 65.005 88.905 65.265 89.165 ;
        RECT 69.235 88.905 69.495 89.165 ;
        RECT 89.295 112.375 89.555 112.635 ;
        RECT 89.295 110.095 89.555 110.355 ;
        RECT 93.525 112.375 93.785 112.635 ;
        RECT 93.845 112.375 94.105 112.635 ;
        RECT 94.165 112.375 94.425 112.635 ;
        RECT 93.525 110.095 93.785 110.355 ;
        RECT 93.845 110.095 94.105 110.355 ;
        RECT 94.165 110.095 94.425 110.355 ;
        RECT 89.295 107.815 89.555 108.075 ;
        RECT 93.525 107.815 93.785 108.075 ;
        RECT 93.845 107.815 94.105 108.075 ;
        RECT 94.165 107.815 94.425 108.075 ;
        RECT 89.900 107.380 90.160 107.640 ;
        RECT 89.900 107.060 90.160 107.320 ;
        RECT 89.900 106.740 90.160 107.000 ;
        RECT 89.295 105.535 89.555 105.795 ;
        RECT 92.990 107.380 93.250 107.640 ;
        RECT 92.990 107.060 93.250 107.320 ;
        RECT 92.990 106.740 93.250 107.000 ;
        RECT 90.835 105.535 91.095 105.795 ;
        RECT 91.155 105.535 91.415 105.795 ;
        RECT 91.475 105.535 91.735 105.795 ;
        RECT 89.295 103.255 89.555 103.515 ;
        RECT 93.525 105.535 93.785 105.795 ;
        RECT 93.845 105.535 94.105 105.795 ;
        RECT 94.165 105.535 94.425 105.795 ;
        RECT 93.525 103.255 93.785 103.515 ;
        RECT 93.845 103.255 94.105 103.515 ;
        RECT 94.165 103.255 94.425 103.515 ;
        RECT 89.295 100.975 89.555 101.235 ;
        RECT 90.835 100.975 91.095 101.235 ;
        RECT 91.155 100.975 91.415 101.235 ;
        RECT 91.475 100.975 91.735 101.235 ;
        RECT 89.295 98.695 89.555 98.955 ;
        RECT 93.525 100.975 93.785 101.235 ;
        RECT 93.845 100.975 94.105 101.235 ;
        RECT 94.165 100.975 94.425 101.235 ;
        RECT 93.525 98.695 93.785 98.955 ;
        RECT 93.845 98.695 94.105 98.955 ;
        RECT 94.165 98.695 94.425 98.955 ;
        RECT 89.295 96.415 89.555 96.675 ;
        RECT 93.525 96.415 93.785 96.675 ;
        RECT 93.845 96.415 94.105 96.675 ;
        RECT 94.165 96.415 94.425 96.675 ;
        RECT 89.295 94.135 89.555 94.395 ;
        RECT 93.525 94.135 93.785 94.395 ;
        RECT 93.845 94.135 94.105 94.395 ;
        RECT 94.165 94.135 94.425 94.395 ;
        RECT 89.295 91.855 89.555 92.115 ;
        RECT 89.295 89.575 89.555 89.835 ;
        RECT 93.525 91.855 93.785 92.115 ;
        RECT 93.845 91.855 94.105 92.115 ;
        RECT 94.165 91.855 94.425 92.115 ;
        RECT 93.525 89.575 93.785 89.835 ;
        RECT 93.845 89.575 94.105 89.835 ;
        RECT 94.165 89.575 94.425 89.835 ;
        RECT 97.100 150.535 97.360 150.795 ;
        RECT 97.420 150.535 97.680 150.795 ;
        RECT 97.740 150.535 98.000 150.795 ;
        RECT 97.100 149.755 97.360 150.015 ;
        RECT 97.420 149.755 97.680 150.015 ;
        RECT 97.740 149.755 98.000 150.015 ;
        RECT 97.100 148.975 97.360 149.235 ;
        RECT 97.420 148.975 97.680 149.235 ;
        RECT 97.740 148.975 98.000 149.235 ;
        RECT 96.565 148.540 96.825 148.800 ;
        RECT 96.565 148.220 96.825 148.480 ;
        RECT 96.565 147.900 96.825 148.160 ;
        RECT 97.100 146.695 97.360 146.955 ;
        RECT 97.420 146.695 97.680 146.955 ;
        RECT 97.740 146.695 98.000 146.955 ;
        RECT 97.100 144.415 97.360 144.675 ;
        RECT 97.420 144.415 97.680 144.675 ;
        RECT 97.740 144.415 98.000 144.675 ;
        RECT 97.100 143.635 97.360 143.895 ;
        RECT 97.420 143.635 97.680 143.895 ;
        RECT 97.740 143.635 98.000 143.895 ;
        RECT 97.100 142.855 97.360 143.115 ;
        RECT 97.420 142.855 97.680 143.115 ;
        RECT 97.740 142.855 98.000 143.115 ;
        RECT 97.100 142.075 97.360 142.335 ;
        RECT 97.420 142.075 97.680 142.335 ;
        RECT 97.740 142.075 98.000 142.335 ;
        RECT 97.100 141.295 97.360 141.555 ;
        RECT 97.420 141.295 97.680 141.555 ;
        RECT 97.740 141.295 98.000 141.555 ;
        RECT 96.565 140.860 96.825 141.120 ;
        RECT 96.565 140.540 96.825 140.800 ;
        RECT 96.565 140.220 96.825 140.480 ;
        RECT 97.100 139.015 97.360 139.275 ;
        RECT 97.420 139.015 97.680 139.275 ;
        RECT 97.740 139.015 98.000 139.275 ;
        RECT 97.100 136.735 97.360 136.995 ;
        RECT 97.420 136.735 97.680 136.995 ;
        RECT 97.740 136.735 98.000 136.995 ;
        RECT 97.100 134.455 97.360 134.715 ;
        RECT 97.420 134.455 97.680 134.715 ;
        RECT 97.740 134.455 98.000 134.715 ;
        RECT 97.100 132.175 97.360 132.435 ;
        RECT 97.420 132.175 97.680 132.435 ;
        RECT 97.740 132.175 98.000 132.435 ;
        RECT 100.690 141.295 100.950 141.555 ;
        RECT 101.010 141.295 101.270 141.555 ;
        RECT 101.330 141.295 101.590 141.555 ;
        RECT 100.690 139.015 100.950 139.275 ;
        RECT 101.010 139.015 101.270 139.275 ;
        RECT 101.330 139.015 101.590 139.275 ;
        RECT 100.690 136.735 100.950 136.995 ;
        RECT 101.010 136.735 101.270 136.995 ;
        RECT 101.330 136.735 101.590 136.995 ;
        RECT 100.690 134.455 100.950 134.715 ;
        RECT 101.010 134.455 101.270 134.715 ;
        RECT 101.330 134.455 101.590 134.715 ;
        RECT 100.690 132.175 100.950 132.435 ;
        RECT 101.010 132.175 101.270 132.435 ;
        RECT 101.330 132.175 101.590 132.435 ;
        RECT 97.100 129.895 97.360 130.155 ;
        RECT 97.420 129.895 97.680 130.155 ;
        RECT 97.740 129.895 98.000 130.155 ;
        RECT 100.690 129.895 100.950 130.155 ;
        RECT 101.010 129.895 101.270 130.155 ;
        RECT 101.330 129.895 101.590 130.155 ;
        RECT 101.865 127.935 102.125 128.195 ;
        RECT 97.100 127.615 97.360 127.875 ;
        RECT 97.420 127.615 97.680 127.875 ;
        RECT 97.740 127.615 98.000 127.875 ;
        RECT 100.690 127.615 100.950 127.875 ;
        RECT 101.010 127.615 101.270 127.875 ;
        RECT 101.330 127.615 101.590 127.875 ;
        RECT 101.865 127.615 102.125 127.875 ;
        RECT 101.865 127.295 102.125 127.555 ;
        RECT 97.100 125.335 97.360 125.595 ;
        RECT 97.420 125.335 97.680 125.595 ;
        RECT 97.740 125.335 98.000 125.595 ;
        RECT 100.690 125.335 100.950 125.595 ;
        RECT 101.010 125.335 101.270 125.595 ;
        RECT 101.330 125.335 101.590 125.595 ;
        RECT 97.100 123.055 97.360 123.315 ;
        RECT 97.420 123.055 97.680 123.315 ;
        RECT 97.740 123.055 98.000 123.315 ;
        RECT 97.100 120.775 97.360 121.035 ;
        RECT 97.420 120.775 97.680 121.035 ;
        RECT 97.740 120.775 98.000 121.035 ;
        RECT 97.100 118.495 97.360 118.755 ;
        RECT 97.420 118.495 97.680 118.755 ;
        RECT 97.740 118.495 98.000 118.755 ;
        RECT 97.100 116.215 97.360 116.475 ;
        RECT 97.420 116.215 97.680 116.475 ;
        RECT 97.740 116.215 98.000 116.475 ;
        RECT 96.565 115.010 96.825 115.270 ;
        RECT 96.565 114.690 96.825 114.950 ;
        RECT 96.565 114.370 96.825 114.630 ;
        RECT 97.100 113.935 97.360 114.195 ;
        RECT 97.420 113.935 97.680 114.195 ;
        RECT 97.740 113.935 98.000 114.195 ;
        RECT 97.100 113.155 97.360 113.415 ;
        RECT 97.420 113.155 97.680 113.415 ;
        RECT 97.740 113.155 98.000 113.415 ;
        RECT 97.100 112.375 97.360 112.635 ;
        RECT 97.420 112.375 97.680 112.635 ;
        RECT 97.740 112.375 98.000 112.635 ;
        RECT 100.690 123.055 100.950 123.315 ;
        RECT 101.010 123.055 101.270 123.315 ;
        RECT 101.330 123.055 101.590 123.315 ;
        RECT 100.690 120.775 100.950 121.035 ;
        RECT 101.010 120.775 101.270 121.035 ;
        RECT 101.330 120.775 101.590 121.035 ;
        RECT 100.690 118.495 100.950 118.755 ;
        RECT 101.010 118.495 101.270 118.755 ;
        RECT 101.330 118.495 101.590 118.755 ;
        RECT 100.690 116.215 100.950 116.475 ;
        RECT 101.010 116.215 101.270 116.475 ;
        RECT 101.330 116.215 101.590 116.475 ;
        RECT 100.690 113.935 100.950 114.195 ;
        RECT 101.010 113.935 101.270 114.195 ;
        RECT 101.330 113.935 101.590 114.195 ;
        RECT 97.100 111.705 97.360 111.965 ;
        RECT 97.420 111.705 97.680 111.965 ;
        RECT 97.740 111.705 98.000 111.965 ;
        RECT 100.690 111.705 100.950 111.965 ;
        RECT 101.010 111.705 101.270 111.965 ;
        RECT 101.330 111.705 101.590 111.965 ;
        RECT 89.295 88.905 89.555 89.165 ;
        RECT 93.525 88.905 93.785 89.165 ;
        RECT 93.845 88.905 94.105 89.165 ;
        RECT 94.165 88.905 94.425 89.165 ;
        RECT 89.160 82.725 89.420 82.985 ;
        RECT 89.480 82.725 89.740 82.985 ;
        RECT 89.800 82.725 90.060 82.985 ;
        RECT 93.010 82.725 93.270 82.985 ;
        RECT 93.330 82.725 93.590 82.985 ;
        RECT 93.650 82.725 93.910 82.985 ;
        RECT 72.730 82.375 72.990 82.635 ;
        RECT 73.050 82.375 73.310 82.635 ;
        RECT 75.955 82.375 76.215 82.635 ;
        RECT 76.275 82.375 76.535 82.635 ;
        RECT 77.530 82.375 77.790 82.635 ;
        RECT 77.850 82.375 78.110 82.635 ;
        RECT 80.450 82.375 80.710 82.635 ;
        RECT 80.770 82.375 81.030 82.635 ;
        RECT 82.025 82.375 82.285 82.635 ;
        RECT 82.345 82.375 82.605 82.635 ;
        RECT 85.250 82.375 85.510 82.635 ;
        RECT 85.570 82.375 85.830 82.635 ;
        RECT 72.730 81.705 72.990 81.965 ;
        RECT 73.050 81.705 73.310 81.965 ;
        RECT 72.730 81.275 72.990 81.535 ;
        RECT 73.050 81.275 73.310 81.535 ;
        RECT 74.465 81.495 74.725 81.755 ;
        RECT 74.465 81.175 74.725 81.435 ;
        RECT 72.730 80.845 72.990 81.105 ;
        RECT 73.050 80.845 73.310 81.105 ;
        RECT 71.960 80.575 72.220 80.835 ;
        RECT 71.960 80.255 72.220 80.515 ;
        RECT 72.495 80.415 72.755 80.675 ;
        RECT 72.815 80.415 73.075 80.675 ;
        RECT 73.135 80.415 73.395 80.675 ;
        RECT 72.730 79.985 72.990 80.245 ;
        RECT 73.050 79.985 73.310 80.245 ;
        RECT 75.955 81.705 76.215 81.965 ;
        RECT 76.275 81.705 76.535 81.965 ;
        RECT 77.530 81.705 77.790 81.965 ;
        RECT 77.850 81.705 78.110 81.965 ;
        RECT 75.955 81.275 76.215 81.535 ;
        RECT 76.275 81.275 76.535 81.535 ;
        RECT 77.530 81.275 77.790 81.535 ;
        RECT 77.850 81.275 78.110 81.535 ;
        RECT 75.795 80.845 76.055 81.105 ;
        RECT 76.115 80.845 76.375 81.105 ;
        RECT 76.435 80.845 76.695 81.105 ;
        RECT 77.530 80.845 77.790 81.105 ;
        RECT 77.850 80.845 78.110 81.105 ;
        RECT 75.795 80.415 76.055 80.675 ;
        RECT 76.115 80.415 76.375 80.675 ;
        RECT 76.435 80.415 76.695 80.675 ;
        RECT 77.445 80.415 77.705 80.675 ;
        RECT 77.765 80.415 78.025 80.675 ;
        RECT 78.085 80.415 78.345 80.675 ;
        RECT 78.620 80.465 78.880 80.725 ;
        RECT 75.795 79.985 76.055 80.245 ;
        RECT 76.115 79.985 76.375 80.245 ;
        RECT 76.435 79.985 76.695 80.245 ;
        RECT 77.530 79.985 77.790 80.245 ;
        RECT 77.850 79.985 78.110 80.245 ;
        RECT 78.620 80.145 78.880 80.405 ;
        RECT 72.495 79.555 72.755 79.815 ;
        RECT 72.815 79.555 73.075 79.815 ;
        RECT 73.135 79.555 73.395 79.815 ;
        RECT 78.620 79.825 78.880 80.085 ;
        RECT 75.795 79.555 76.055 79.815 ;
        RECT 76.115 79.555 76.375 79.815 ;
        RECT 76.435 79.555 76.695 79.815 ;
        RECT 77.445 79.555 77.705 79.815 ;
        RECT 77.765 79.555 78.025 79.815 ;
        RECT 78.085 79.555 78.345 79.815 ;
        RECT 78.620 79.505 78.880 79.765 ;
        RECT 72.730 79.125 72.990 79.385 ;
        RECT 73.050 79.125 73.310 79.385 ;
        RECT 75.795 79.125 76.055 79.385 ;
        RECT 76.115 79.125 76.375 79.385 ;
        RECT 76.435 79.125 76.695 79.385 ;
        RECT 77.530 79.125 77.790 79.385 ;
        RECT 77.850 79.125 78.110 79.385 ;
        RECT 72.730 78.695 72.990 78.955 ;
        RECT 73.050 78.695 73.310 78.955 ;
        RECT 72.730 78.265 72.990 78.525 ;
        RECT 73.050 78.265 73.310 78.525 ;
        RECT 72.730 77.615 72.990 77.875 ;
        RECT 73.050 77.615 73.310 77.875 ;
        RECT 75.955 78.695 76.215 78.955 ;
        RECT 76.275 78.695 76.535 78.955 ;
        RECT 77.530 78.695 77.790 78.955 ;
        RECT 77.850 78.695 78.110 78.955 ;
        RECT 75.955 78.265 76.215 78.525 ;
        RECT 76.275 78.265 76.535 78.525 ;
        RECT 77.530 78.265 77.790 78.525 ;
        RECT 77.850 78.265 78.110 78.525 ;
        RECT 75.955 77.615 76.215 77.875 ;
        RECT 76.275 77.615 76.535 77.875 ;
        RECT 77.530 77.615 77.790 77.875 ;
        RECT 77.850 77.615 78.110 77.875 ;
        RECT 80.450 81.705 80.710 81.965 ;
        RECT 80.770 81.705 81.030 81.965 ;
        RECT 82.025 81.705 82.285 81.965 ;
        RECT 82.345 81.705 82.605 81.965 ;
        RECT 80.450 81.275 80.710 81.535 ;
        RECT 80.770 81.275 81.030 81.535 ;
        RECT 82.025 81.275 82.285 81.535 ;
        RECT 82.345 81.275 82.605 81.535 ;
        RECT 83.835 81.495 84.095 81.755 ;
        RECT 83.835 81.175 84.095 81.435 ;
        RECT 80.450 80.845 80.710 81.105 ;
        RECT 80.770 80.845 81.030 81.105 ;
        RECT 81.865 80.845 82.125 81.105 ;
        RECT 82.185 80.845 82.445 81.105 ;
        RECT 82.505 80.845 82.765 81.105 ;
        RECT 79.680 80.465 79.940 80.725 ;
        RECT 80.215 80.415 80.475 80.675 ;
        RECT 80.535 80.415 80.795 80.675 ;
        RECT 80.855 80.415 81.115 80.675 ;
        RECT 81.865 80.415 82.125 80.675 ;
        RECT 82.185 80.415 82.445 80.675 ;
        RECT 82.505 80.415 82.765 80.675 ;
        RECT 79.680 80.145 79.940 80.405 ;
        RECT 79.680 79.825 79.940 80.085 ;
        RECT 80.450 79.985 80.710 80.245 ;
        RECT 80.770 79.985 81.030 80.245 ;
        RECT 81.865 79.985 82.125 80.245 ;
        RECT 82.185 79.985 82.445 80.245 ;
        RECT 82.505 79.985 82.765 80.245 ;
        RECT 85.250 81.705 85.510 81.965 ;
        RECT 85.570 81.705 85.830 81.965 ;
        RECT 85.250 81.275 85.510 81.535 ;
        RECT 85.570 81.275 85.830 81.535 ;
        RECT 85.250 80.845 85.510 81.105 ;
        RECT 85.570 80.845 85.830 81.105 ;
        RECT 85.165 80.415 85.425 80.675 ;
        RECT 85.485 80.415 85.745 80.675 ;
        RECT 85.805 80.415 86.065 80.675 ;
        RECT 86.340 80.575 86.600 80.835 ;
        RECT 86.340 80.255 86.600 80.515 ;
        RECT 85.250 79.985 85.510 80.245 ;
        RECT 85.570 79.985 85.830 80.245 ;
        RECT 79.680 79.505 79.940 79.765 ;
        RECT 80.215 79.555 80.475 79.815 ;
        RECT 80.535 79.555 80.795 79.815 ;
        RECT 80.855 79.555 81.115 79.815 ;
        RECT 81.865 79.555 82.125 79.815 ;
        RECT 82.185 79.555 82.445 79.815 ;
        RECT 82.505 79.555 82.765 79.815 ;
        RECT 85.165 79.555 85.425 79.815 ;
        RECT 85.485 79.555 85.745 79.815 ;
        RECT 85.805 79.555 86.065 79.815 ;
        RECT 80.450 79.125 80.710 79.385 ;
        RECT 80.770 79.125 81.030 79.385 ;
        RECT 81.865 79.125 82.125 79.385 ;
        RECT 82.185 79.125 82.445 79.385 ;
        RECT 82.505 79.125 82.765 79.385 ;
        RECT 85.250 79.125 85.510 79.385 ;
        RECT 85.570 79.125 85.830 79.385 ;
        RECT 80.450 78.695 80.710 78.955 ;
        RECT 80.770 78.695 81.030 78.955 ;
        RECT 82.025 78.695 82.285 78.955 ;
        RECT 82.345 78.695 82.605 78.955 ;
        RECT 80.450 78.265 80.710 78.525 ;
        RECT 80.770 78.265 81.030 78.525 ;
        RECT 82.025 78.265 82.285 78.525 ;
        RECT 82.345 78.265 82.605 78.525 ;
        RECT 80.450 77.615 80.710 77.875 ;
        RECT 80.770 77.615 81.030 77.875 ;
        RECT 82.025 77.615 82.285 77.875 ;
        RECT 82.345 77.615 82.605 77.875 ;
        RECT 85.250 78.695 85.510 78.955 ;
        RECT 85.570 78.695 85.830 78.955 ;
        RECT 85.250 78.265 85.510 78.525 ;
        RECT 85.570 78.265 85.830 78.525 ;
        RECT 85.250 77.615 85.510 77.875 ;
        RECT 85.570 77.615 85.830 77.875 ;
        RECT 89.160 82.055 89.420 82.315 ;
        RECT 89.480 82.055 89.740 82.315 ;
        RECT 89.800 82.055 90.060 82.315 ;
        RECT 89.160 81.625 89.420 81.885 ;
        RECT 89.480 81.625 89.740 81.885 ;
        RECT 89.800 81.625 90.060 81.885 ;
        RECT 91.155 81.960 91.415 82.220 ;
        RECT 91.155 81.640 91.415 81.900 ;
        RECT 89.160 81.195 89.420 81.455 ;
        RECT 89.480 81.195 89.740 81.455 ;
        RECT 89.800 81.195 90.060 81.455 ;
        RECT 89.160 80.765 89.420 81.025 ;
        RECT 89.480 80.765 89.740 81.025 ;
        RECT 89.800 80.765 90.060 81.025 ;
        RECT 93.010 82.055 93.270 82.315 ;
        RECT 93.330 82.055 93.590 82.315 ;
        RECT 93.650 82.055 93.910 82.315 ;
        RECT 93.010 81.625 93.270 81.885 ;
        RECT 93.330 81.625 93.590 81.885 ;
        RECT 93.650 81.625 93.910 81.885 ;
        RECT 93.010 81.195 93.270 81.455 ;
        RECT 93.330 81.195 93.590 81.455 ;
        RECT 93.650 81.195 93.910 81.455 ;
        RECT 92.530 80.765 92.790 81.025 ;
        RECT 92.850 80.765 93.110 81.025 ;
        RECT 93.170 80.765 93.430 81.025 ;
        RECT 93.490 80.765 93.750 81.025 ;
        RECT 93.810 80.765 94.070 81.025 ;
        RECT 94.130 80.765 94.390 81.025 ;
        RECT 89.160 80.335 89.420 80.595 ;
        RECT 89.480 80.335 89.740 80.595 ;
        RECT 89.800 80.335 90.060 80.595 ;
        RECT 93.010 80.335 93.270 80.595 ;
        RECT 93.330 80.335 93.590 80.595 ;
        RECT 93.650 80.335 93.910 80.595 ;
        RECT 89.160 79.905 89.420 80.165 ;
        RECT 89.480 79.905 89.740 80.165 ;
        RECT 89.800 79.905 90.060 80.165 ;
        RECT 92.530 79.905 92.790 80.165 ;
        RECT 92.850 79.905 93.110 80.165 ;
        RECT 93.170 79.905 93.430 80.165 ;
        RECT 93.490 79.905 93.750 80.165 ;
        RECT 93.810 79.905 94.070 80.165 ;
        RECT 94.130 79.905 94.390 80.165 ;
        RECT 89.160 79.475 89.420 79.735 ;
        RECT 89.480 79.475 89.740 79.735 ;
        RECT 89.800 79.475 90.060 79.735 ;
        RECT 93.010 79.475 93.270 79.735 ;
        RECT 93.330 79.475 93.590 79.735 ;
        RECT 93.650 79.475 93.910 79.735 ;
        RECT 89.160 79.045 89.420 79.305 ;
        RECT 89.480 79.045 89.740 79.305 ;
        RECT 89.800 79.045 90.060 79.305 ;
        RECT 89.160 78.615 89.420 78.875 ;
        RECT 89.480 78.615 89.740 78.875 ;
        RECT 89.800 78.615 90.060 78.875 ;
        RECT 93.010 79.045 93.270 79.305 ;
        RECT 93.330 79.045 93.590 79.305 ;
        RECT 93.650 79.045 93.910 79.305 ;
        RECT 93.010 78.615 93.270 78.875 ;
        RECT 93.330 78.615 93.590 78.875 ;
        RECT 93.650 78.615 93.910 78.875 ;
        RECT 89.160 77.945 89.420 78.205 ;
        RECT 89.480 77.945 89.740 78.205 ;
        RECT 89.800 77.945 90.060 78.205 ;
        RECT 93.010 77.945 93.270 78.205 ;
        RECT 93.330 77.945 93.590 78.205 ;
        RECT 93.650 77.945 93.910 78.205 ;
        RECT 65.380 72.065 65.640 72.325 ;
        RECT 65.700 72.065 65.960 72.325 ;
        RECT 66.020 72.065 66.280 72.325 ;
        RECT 69.230 72.065 69.490 72.325 ;
        RECT 69.550 72.065 69.810 72.325 ;
        RECT 69.870 72.065 70.130 72.325 ;
        RECT 65.380 71.395 65.640 71.655 ;
        RECT 65.700 71.395 65.960 71.655 ;
        RECT 66.020 71.395 66.280 71.655 ;
        RECT 65.380 70.965 65.640 71.225 ;
        RECT 65.700 70.965 65.960 71.225 ;
        RECT 66.020 70.965 66.280 71.225 ;
        RECT 67.375 71.300 67.635 71.560 ;
        RECT 67.375 70.980 67.635 71.240 ;
        RECT 65.380 70.535 65.640 70.795 ;
        RECT 65.700 70.535 65.960 70.795 ;
        RECT 66.020 70.535 66.280 70.795 ;
        RECT 65.380 70.105 65.640 70.365 ;
        RECT 65.700 70.105 65.960 70.365 ;
        RECT 66.020 70.105 66.280 70.365 ;
        RECT 69.230 71.395 69.490 71.655 ;
        RECT 69.550 71.395 69.810 71.655 ;
        RECT 69.870 71.395 70.130 71.655 ;
        RECT 69.230 70.965 69.490 71.225 ;
        RECT 69.550 70.965 69.810 71.225 ;
        RECT 69.870 70.965 70.130 71.225 ;
        RECT 69.230 70.535 69.490 70.795 ;
        RECT 69.550 70.535 69.810 70.795 ;
        RECT 69.870 70.535 70.130 70.795 ;
        RECT 68.750 70.105 69.010 70.365 ;
        RECT 69.070 70.105 69.330 70.365 ;
        RECT 69.390 70.105 69.650 70.365 ;
        RECT 69.710 70.105 69.970 70.365 ;
        RECT 70.030 70.105 70.290 70.365 ;
        RECT 70.350 70.105 70.610 70.365 ;
        RECT 65.380 69.675 65.640 69.935 ;
        RECT 65.700 69.675 65.960 69.935 ;
        RECT 66.020 69.675 66.280 69.935 ;
        RECT 69.230 69.675 69.490 69.935 ;
        RECT 69.550 69.675 69.810 69.935 ;
        RECT 69.870 69.675 70.130 69.935 ;
        RECT 65.380 69.245 65.640 69.505 ;
        RECT 65.700 69.245 65.960 69.505 ;
        RECT 66.020 69.245 66.280 69.505 ;
        RECT 67.055 69.245 67.315 69.505 ;
        RECT 67.375 69.245 67.635 69.505 ;
        RECT 67.695 69.245 67.955 69.505 ;
        RECT 65.380 68.815 65.640 69.075 ;
        RECT 65.700 68.815 65.960 69.075 ;
        RECT 66.020 68.815 66.280 69.075 ;
        RECT 65.380 68.385 65.640 68.645 ;
        RECT 65.700 68.385 65.960 68.645 ;
        RECT 66.020 68.385 66.280 68.645 ;
        RECT 65.380 67.955 65.640 68.215 ;
        RECT 65.700 67.955 65.960 68.215 ;
        RECT 66.020 67.955 66.280 68.215 ;
        RECT 65.380 67.525 65.640 67.785 ;
        RECT 65.700 67.525 65.960 67.785 ;
        RECT 66.020 67.525 66.280 67.785 ;
        RECT 65.380 67.095 65.640 67.355 ;
        RECT 65.700 67.095 65.960 67.355 ;
        RECT 66.020 67.095 66.280 67.355 ;
        RECT 68.750 69.245 69.010 69.505 ;
        RECT 69.070 69.245 69.330 69.505 ;
        RECT 69.390 69.245 69.650 69.505 ;
        RECT 69.710 69.245 69.970 69.505 ;
        RECT 70.030 69.245 70.290 69.505 ;
        RECT 70.350 69.245 70.610 69.505 ;
        RECT 69.230 68.815 69.490 69.075 ;
        RECT 69.550 68.815 69.810 69.075 ;
        RECT 69.870 68.815 70.130 69.075 ;
        RECT 68.750 68.385 69.010 68.645 ;
        RECT 69.070 68.385 69.330 68.645 ;
        RECT 69.390 68.385 69.650 68.645 ;
        RECT 69.710 68.385 69.970 68.645 ;
        RECT 70.030 68.385 70.290 68.645 ;
        RECT 70.350 68.385 70.610 68.645 ;
        RECT 69.230 67.955 69.490 68.215 ;
        RECT 69.550 67.955 69.810 68.215 ;
        RECT 69.870 67.955 70.130 68.215 ;
        RECT 68.750 67.525 69.010 67.785 ;
        RECT 69.070 67.525 69.330 67.785 ;
        RECT 69.390 67.525 69.650 67.785 ;
        RECT 69.710 67.525 69.970 67.785 ;
        RECT 70.030 67.525 70.290 67.785 ;
        RECT 70.350 67.525 70.610 67.785 ;
        RECT 69.230 67.095 69.490 67.355 ;
        RECT 69.550 67.095 69.810 67.355 ;
        RECT 69.870 67.095 70.130 67.355 ;
        RECT 65.380 66.665 65.640 66.925 ;
        RECT 65.700 66.665 65.960 66.925 ;
        RECT 66.020 66.665 66.280 66.925 ;
        RECT 68.750 66.665 69.010 66.925 ;
        RECT 69.070 66.665 69.330 66.925 ;
        RECT 69.390 66.665 69.650 66.925 ;
        RECT 69.710 66.665 69.970 66.925 ;
        RECT 70.030 66.665 70.290 66.925 ;
        RECT 70.350 66.665 70.610 66.925 ;
        RECT 65.380 66.235 65.640 66.495 ;
        RECT 65.700 66.235 65.960 66.495 ;
        RECT 66.020 66.235 66.280 66.495 ;
        RECT 65.380 65.805 65.640 66.065 ;
        RECT 65.700 65.805 65.960 66.065 ;
        RECT 66.020 65.805 66.280 66.065 ;
        RECT 65.380 65.375 65.640 65.635 ;
        RECT 65.700 65.375 65.960 65.635 ;
        RECT 66.020 65.375 66.280 65.635 ;
        RECT 65.380 64.945 65.640 65.205 ;
        RECT 65.700 64.945 65.960 65.205 ;
        RECT 66.020 64.945 66.280 65.205 ;
        RECT 69.230 66.235 69.490 66.495 ;
        RECT 69.550 66.235 69.810 66.495 ;
        RECT 69.870 66.235 70.130 66.495 ;
        RECT 68.750 65.805 69.010 66.065 ;
        RECT 69.070 65.805 69.330 66.065 ;
        RECT 69.390 65.805 69.650 66.065 ;
        RECT 69.710 65.805 69.970 66.065 ;
        RECT 70.030 65.805 70.290 66.065 ;
        RECT 70.350 65.805 70.610 66.065 ;
        RECT 69.230 65.375 69.490 65.635 ;
        RECT 69.550 65.375 69.810 65.635 ;
        RECT 69.870 65.375 70.130 65.635 ;
        RECT 68.750 64.945 69.010 65.205 ;
        RECT 69.070 64.945 69.330 65.205 ;
        RECT 69.390 64.945 69.650 65.205 ;
        RECT 69.710 64.945 69.970 65.205 ;
        RECT 70.030 64.945 70.290 65.205 ;
        RECT 70.350 64.945 70.610 65.205 ;
        RECT 65.380 64.515 65.640 64.775 ;
        RECT 65.700 64.515 65.960 64.775 ;
        RECT 66.020 64.515 66.280 64.775 ;
        RECT 69.230 64.515 69.490 64.775 ;
        RECT 69.550 64.515 69.810 64.775 ;
        RECT 69.870 64.515 70.130 64.775 ;
        RECT 65.380 64.085 65.640 64.345 ;
        RECT 65.700 64.085 65.960 64.345 ;
        RECT 66.020 64.085 66.280 64.345 ;
        RECT 65.380 63.655 65.640 63.915 ;
        RECT 65.700 63.655 65.960 63.915 ;
        RECT 66.020 63.655 66.280 63.915 ;
        RECT 69.230 64.085 69.490 64.345 ;
        RECT 69.550 64.085 69.810 64.345 ;
        RECT 69.870 64.085 70.130 64.345 ;
        RECT 69.230 63.655 69.490 63.915 ;
        RECT 69.550 63.655 69.810 63.915 ;
        RECT 69.870 63.655 70.130 63.915 ;
        RECT 65.380 62.985 65.640 63.245 ;
        RECT 65.700 62.985 65.960 63.245 ;
        RECT 66.020 62.985 66.280 63.245 ;
        RECT 69.230 62.985 69.490 63.245 ;
        RECT 69.550 62.985 69.810 63.245 ;
        RECT 69.870 62.985 70.130 63.245 ;
        RECT 74.400 72.065 74.660 72.325 ;
        RECT 74.720 72.065 74.980 72.325 ;
        RECT 75.040 72.065 75.300 72.325 ;
        RECT 78.250 72.065 78.510 72.325 ;
        RECT 78.570 72.065 78.830 72.325 ;
        RECT 78.890 72.065 79.150 72.325 ;
        RECT 81.340 72.065 81.600 72.325 ;
        RECT 81.660 72.065 81.920 72.325 ;
        RECT 81.980 72.065 82.240 72.325 ;
        RECT 85.190 72.065 85.450 72.325 ;
        RECT 85.510 72.065 85.770 72.325 ;
        RECT 85.830 72.065 86.090 72.325 ;
        RECT 74.400 71.395 74.660 71.655 ;
        RECT 74.720 71.395 74.980 71.655 ;
        RECT 75.040 71.395 75.300 71.655 ;
        RECT 74.400 70.965 74.660 71.225 ;
        RECT 74.720 70.965 74.980 71.225 ;
        RECT 75.040 70.965 75.300 71.225 ;
        RECT 76.395 71.300 76.655 71.560 ;
        RECT 76.395 70.980 76.655 71.240 ;
        RECT 74.400 70.535 74.660 70.795 ;
        RECT 74.720 70.535 74.980 70.795 ;
        RECT 75.040 70.535 75.300 70.795 ;
        RECT 74.400 70.105 74.660 70.365 ;
        RECT 74.720 70.105 74.980 70.365 ;
        RECT 75.040 70.105 75.300 70.365 ;
        RECT 78.250 71.395 78.510 71.655 ;
        RECT 78.570 71.395 78.830 71.655 ;
        RECT 78.890 71.395 79.150 71.655 ;
        RECT 78.250 70.965 78.510 71.225 ;
        RECT 78.570 70.965 78.830 71.225 ;
        RECT 78.890 70.965 79.150 71.225 ;
        RECT 78.250 70.535 78.510 70.795 ;
        RECT 78.570 70.535 78.830 70.795 ;
        RECT 78.890 70.535 79.150 70.795 ;
        RECT 77.770 70.105 78.030 70.365 ;
        RECT 78.090 70.105 78.350 70.365 ;
        RECT 78.410 70.105 78.670 70.365 ;
        RECT 78.730 70.105 78.990 70.365 ;
        RECT 79.050 70.105 79.310 70.365 ;
        RECT 79.370 70.105 79.630 70.365 ;
        RECT 74.400 69.675 74.660 69.935 ;
        RECT 74.720 69.675 74.980 69.935 ;
        RECT 75.040 69.675 75.300 69.935 ;
        RECT 78.250 69.675 78.510 69.935 ;
        RECT 78.570 69.675 78.830 69.935 ;
        RECT 78.890 69.675 79.150 69.935 ;
        RECT 74.400 69.245 74.660 69.505 ;
        RECT 74.720 69.245 74.980 69.505 ;
        RECT 75.040 69.245 75.300 69.505 ;
        RECT 76.075 69.245 76.335 69.505 ;
        RECT 76.395 69.245 76.655 69.505 ;
        RECT 76.715 69.245 76.975 69.505 ;
        RECT 74.400 68.815 74.660 69.075 ;
        RECT 74.720 68.815 74.980 69.075 ;
        RECT 75.040 68.815 75.300 69.075 ;
        RECT 74.400 68.385 74.660 68.645 ;
        RECT 74.720 68.385 74.980 68.645 ;
        RECT 75.040 68.385 75.300 68.645 ;
        RECT 74.400 67.955 74.660 68.215 ;
        RECT 74.720 67.955 74.980 68.215 ;
        RECT 75.040 67.955 75.300 68.215 ;
        RECT 74.400 67.525 74.660 67.785 ;
        RECT 74.720 67.525 74.980 67.785 ;
        RECT 75.040 67.525 75.300 67.785 ;
        RECT 74.400 67.095 74.660 67.355 ;
        RECT 74.720 67.095 74.980 67.355 ;
        RECT 75.040 67.095 75.300 67.355 ;
        RECT 77.770 69.245 78.030 69.505 ;
        RECT 78.090 69.245 78.350 69.505 ;
        RECT 78.410 69.245 78.670 69.505 ;
        RECT 78.730 69.245 78.990 69.505 ;
        RECT 79.050 69.245 79.310 69.505 ;
        RECT 79.370 69.245 79.630 69.505 ;
        RECT 78.250 68.815 78.510 69.075 ;
        RECT 78.570 68.815 78.830 69.075 ;
        RECT 78.890 68.815 79.150 69.075 ;
        RECT 77.770 68.385 78.030 68.645 ;
        RECT 78.090 68.385 78.350 68.645 ;
        RECT 78.410 68.385 78.670 68.645 ;
        RECT 78.730 68.385 78.990 68.645 ;
        RECT 79.050 68.385 79.310 68.645 ;
        RECT 79.370 68.385 79.630 68.645 ;
        RECT 78.250 67.955 78.510 68.215 ;
        RECT 78.570 67.955 78.830 68.215 ;
        RECT 78.890 67.955 79.150 68.215 ;
        RECT 77.770 67.525 78.030 67.785 ;
        RECT 78.090 67.525 78.350 67.785 ;
        RECT 78.410 67.525 78.670 67.785 ;
        RECT 78.730 67.525 78.990 67.785 ;
        RECT 79.050 67.525 79.310 67.785 ;
        RECT 79.370 67.525 79.630 67.785 ;
        RECT 78.250 67.095 78.510 67.355 ;
        RECT 78.570 67.095 78.830 67.355 ;
        RECT 78.890 67.095 79.150 67.355 ;
        RECT 74.400 66.665 74.660 66.925 ;
        RECT 74.720 66.665 74.980 66.925 ;
        RECT 75.040 66.665 75.300 66.925 ;
        RECT 77.770 66.665 78.030 66.925 ;
        RECT 78.090 66.665 78.350 66.925 ;
        RECT 78.410 66.665 78.670 66.925 ;
        RECT 78.730 66.665 78.990 66.925 ;
        RECT 79.050 66.665 79.310 66.925 ;
        RECT 79.370 66.665 79.630 66.925 ;
        RECT 74.400 66.235 74.660 66.495 ;
        RECT 74.720 66.235 74.980 66.495 ;
        RECT 75.040 66.235 75.300 66.495 ;
        RECT 74.400 65.805 74.660 66.065 ;
        RECT 74.720 65.805 74.980 66.065 ;
        RECT 75.040 65.805 75.300 66.065 ;
        RECT 74.400 65.375 74.660 65.635 ;
        RECT 74.720 65.375 74.980 65.635 ;
        RECT 75.040 65.375 75.300 65.635 ;
        RECT 74.400 64.945 74.660 65.205 ;
        RECT 74.720 64.945 74.980 65.205 ;
        RECT 75.040 64.945 75.300 65.205 ;
        RECT 78.250 66.235 78.510 66.495 ;
        RECT 78.570 66.235 78.830 66.495 ;
        RECT 78.890 66.235 79.150 66.495 ;
        RECT 77.770 65.805 78.030 66.065 ;
        RECT 78.090 65.805 78.350 66.065 ;
        RECT 78.410 65.805 78.670 66.065 ;
        RECT 78.730 65.805 78.990 66.065 ;
        RECT 79.050 65.805 79.310 66.065 ;
        RECT 79.370 65.805 79.630 66.065 ;
        RECT 78.250 65.375 78.510 65.635 ;
        RECT 78.570 65.375 78.830 65.635 ;
        RECT 78.890 65.375 79.150 65.635 ;
        RECT 77.770 64.945 78.030 65.205 ;
        RECT 78.090 64.945 78.350 65.205 ;
        RECT 78.410 64.945 78.670 65.205 ;
        RECT 78.730 64.945 78.990 65.205 ;
        RECT 79.050 64.945 79.310 65.205 ;
        RECT 79.370 64.945 79.630 65.205 ;
        RECT 74.400 64.515 74.660 64.775 ;
        RECT 74.720 64.515 74.980 64.775 ;
        RECT 75.040 64.515 75.300 64.775 ;
        RECT 78.250 64.515 78.510 64.775 ;
        RECT 78.570 64.515 78.830 64.775 ;
        RECT 78.890 64.515 79.150 64.775 ;
        RECT 74.400 64.085 74.660 64.345 ;
        RECT 74.720 64.085 74.980 64.345 ;
        RECT 75.040 64.085 75.300 64.345 ;
        RECT 74.400 63.655 74.660 63.915 ;
        RECT 74.720 63.655 74.980 63.915 ;
        RECT 75.040 63.655 75.300 63.915 ;
        RECT 78.250 64.085 78.510 64.345 ;
        RECT 78.570 64.085 78.830 64.345 ;
        RECT 78.890 64.085 79.150 64.345 ;
        RECT 78.250 63.655 78.510 63.915 ;
        RECT 78.570 63.655 78.830 63.915 ;
        RECT 78.890 63.655 79.150 63.915 ;
        RECT 81.340 71.395 81.600 71.655 ;
        RECT 81.660 71.395 81.920 71.655 ;
        RECT 81.980 71.395 82.240 71.655 ;
        RECT 81.340 70.965 81.600 71.225 ;
        RECT 81.660 70.965 81.920 71.225 ;
        RECT 81.980 70.965 82.240 71.225 ;
        RECT 83.835 71.300 84.095 71.560 ;
        RECT 83.835 70.980 84.095 71.240 ;
        RECT 81.340 70.535 81.600 70.795 ;
        RECT 81.660 70.535 81.920 70.795 ;
        RECT 81.980 70.535 82.240 70.795 ;
        RECT 80.860 70.105 81.120 70.365 ;
        RECT 81.180 70.105 81.440 70.365 ;
        RECT 81.500 70.105 81.760 70.365 ;
        RECT 81.820 70.105 82.080 70.365 ;
        RECT 82.140 70.105 82.400 70.365 ;
        RECT 82.460 70.105 82.720 70.365 ;
        RECT 85.190 71.395 85.450 71.655 ;
        RECT 85.510 71.395 85.770 71.655 ;
        RECT 85.830 71.395 86.090 71.655 ;
        RECT 85.190 70.965 85.450 71.225 ;
        RECT 85.510 70.965 85.770 71.225 ;
        RECT 85.830 70.965 86.090 71.225 ;
        RECT 85.190 70.535 85.450 70.795 ;
        RECT 85.510 70.535 85.770 70.795 ;
        RECT 85.830 70.535 86.090 70.795 ;
        RECT 85.190 70.105 85.450 70.365 ;
        RECT 85.510 70.105 85.770 70.365 ;
        RECT 85.830 70.105 86.090 70.365 ;
        RECT 81.340 69.675 81.600 69.935 ;
        RECT 81.660 69.675 81.920 69.935 ;
        RECT 81.980 69.675 82.240 69.935 ;
        RECT 85.190 69.675 85.450 69.935 ;
        RECT 85.510 69.675 85.770 69.935 ;
        RECT 85.830 69.675 86.090 69.935 ;
        RECT 80.860 69.245 81.120 69.505 ;
        RECT 81.180 69.245 81.440 69.505 ;
        RECT 81.500 69.245 81.760 69.505 ;
        RECT 81.820 69.245 82.080 69.505 ;
        RECT 82.140 69.245 82.400 69.505 ;
        RECT 82.460 69.245 82.720 69.505 ;
        RECT 83.515 69.245 83.775 69.505 ;
        RECT 83.835 69.245 84.095 69.505 ;
        RECT 84.155 69.245 84.415 69.505 ;
        RECT 81.340 68.815 81.600 69.075 ;
        RECT 81.660 68.815 81.920 69.075 ;
        RECT 81.980 68.815 82.240 69.075 ;
        RECT 80.860 68.385 81.120 68.645 ;
        RECT 81.180 68.385 81.440 68.645 ;
        RECT 81.500 68.385 81.760 68.645 ;
        RECT 81.820 68.385 82.080 68.645 ;
        RECT 82.140 68.385 82.400 68.645 ;
        RECT 82.460 68.385 82.720 68.645 ;
        RECT 81.340 67.955 81.600 68.215 ;
        RECT 81.660 67.955 81.920 68.215 ;
        RECT 81.980 67.955 82.240 68.215 ;
        RECT 80.860 67.525 81.120 67.785 ;
        RECT 81.180 67.525 81.440 67.785 ;
        RECT 81.500 67.525 81.760 67.785 ;
        RECT 81.820 67.525 82.080 67.785 ;
        RECT 82.140 67.525 82.400 67.785 ;
        RECT 82.460 67.525 82.720 67.785 ;
        RECT 81.340 67.095 81.600 67.355 ;
        RECT 81.660 67.095 81.920 67.355 ;
        RECT 81.980 67.095 82.240 67.355 ;
        RECT 85.190 69.245 85.450 69.505 ;
        RECT 85.510 69.245 85.770 69.505 ;
        RECT 85.830 69.245 86.090 69.505 ;
        RECT 85.190 68.815 85.450 69.075 ;
        RECT 85.510 68.815 85.770 69.075 ;
        RECT 85.830 68.815 86.090 69.075 ;
        RECT 85.190 68.385 85.450 68.645 ;
        RECT 85.510 68.385 85.770 68.645 ;
        RECT 85.830 68.385 86.090 68.645 ;
        RECT 85.190 67.955 85.450 68.215 ;
        RECT 85.510 67.955 85.770 68.215 ;
        RECT 85.830 67.955 86.090 68.215 ;
        RECT 85.190 67.525 85.450 67.785 ;
        RECT 85.510 67.525 85.770 67.785 ;
        RECT 85.830 67.525 86.090 67.785 ;
        RECT 85.190 67.095 85.450 67.355 ;
        RECT 85.510 67.095 85.770 67.355 ;
        RECT 85.830 67.095 86.090 67.355 ;
        RECT 80.860 66.665 81.120 66.925 ;
        RECT 81.180 66.665 81.440 66.925 ;
        RECT 81.500 66.665 81.760 66.925 ;
        RECT 81.820 66.665 82.080 66.925 ;
        RECT 82.140 66.665 82.400 66.925 ;
        RECT 82.460 66.665 82.720 66.925 ;
        RECT 85.190 66.665 85.450 66.925 ;
        RECT 85.510 66.665 85.770 66.925 ;
        RECT 85.830 66.665 86.090 66.925 ;
        RECT 81.340 66.235 81.600 66.495 ;
        RECT 81.660 66.235 81.920 66.495 ;
        RECT 81.980 66.235 82.240 66.495 ;
        RECT 80.860 65.805 81.120 66.065 ;
        RECT 81.180 65.805 81.440 66.065 ;
        RECT 81.500 65.805 81.760 66.065 ;
        RECT 81.820 65.805 82.080 66.065 ;
        RECT 82.140 65.805 82.400 66.065 ;
        RECT 82.460 65.805 82.720 66.065 ;
        RECT 81.340 65.375 81.600 65.635 ;
        RECT 81.660 65.375 81.920 65.635 ;
        RECT 81.980 65.375 82.240 65.635 ;
        RECT 80.860 64.945 81.120 65.205 ;
        RECT 81.180 64.945 81.440 65.205 ;
        RECT 81.500 64.945 81.760 65.205 ;
        RECT 81.820 64.945 82.080 65.205 ;
        RECT 82.140 64.945 82.400 65.205 ;
        RECT 82.460 64.945 82.720 65.205 ;
        RECT 85.190 66.235 85.450 66.495 ;
        RECT 85.510 66.235 85.770 66.495 ;
        RECT 85.830 66.235 86.090 66.495 ;
        RECT 85.190 65.805 85.450 66.065 ;
        RECT 85.510 65.805 85.770 66.065 ;
        RECT 85.830 65.805 86.090 66.065 ;
        RECT 85.190 65.375 85.450 65.635 ;
        RECT 85.510 65.375 85.770 65.635 ;
        RECT 85.830 65.375 86.090 65.635 ;
        RECT 85.190 64.945 85.450 65.205 ;
        RECT 85.510 64.945 85.770 65.205 ;
        RECT 85.830 64.945 86.090 65.205 ;
        RECT 81.340 64.515 81.600 64.775 ;
        RECT 81.660 64.515 81.920 64.775 ;
        RECT 81.980 64.515 82.240 64.775 ;
        RECT 85.190 64.515 85.450 64.775 ;
        RECT 85.510 64.515 85.770 64.775 ;
        RECT 85.830 64.515 86.090 64.775 ;
        RECT 81.340 64.085 81.600 64.345 ;
        RECT 81.660 64.085 81.920 64.345 ;
        RECT 81.980 64.085 82.240 64.345 ;
        RECT 81.340 63.655 81.600 63.915 ;
        RECT 81.660 63.655 81.920 63.915 ;
        RECT 81.980 63.655 82.240 63.915 ;
        RECT 85.190 64.085 85.450 64.345 ;
        RECT 85.510 64.085 85.770 64.345 ;
        RECT 85.830 64.085 86.090 64.345 ;
        RECT 85.190 63.655 85.450 63.915 ;
        RECT 85.510 63.655 85.770 63.915 ;
        RECT 85.830 63.655 86.090 63.915 ;
        RECT 74.400 62.985 74.660 63.245 ;
        RECT 74.720 62.985 74.980 63.245 ;
        RECT 75.040 62.985 75.300 63.245 ;
        RECT 78.250 62.985 78.510 63.245 ;
        RECT 78.570 62.985 78.830 63.245 ;
        RECT 78.890 62.985 79.150 63.245 ;
        RECT 81.340 62.985 81.600 63.245 ;
        RECT 81.660 62.985 81.920 63.245 ;
        RECT 81.980 62.985 82.240 63.245 ;
        RECT 85.190 62.985 85.450 63.245 ;
        RECT 85.510 62.985 85.770 63.245 ;
        RECT 85.830 62.985 86.090 63.245 ;
        RECT 89.160 72.065 89.420 72.325 ;
        RECT 89.480 72.065 89.740 72.325 ;
        RECT 89.800 72.065 90.060 72.325 ;
        RECT 93.010 72.065 93.270 72.325 ;
        RECT 93.330 72.065 93.590 72.325 ;
        RECT 93.650 72.065 93.910 72.325 ;
        RECT 89.160 71.395 89.420 71.655 ;
        RECT 89.480 71.395 89.740 71.655 ;
        RECT 89.800 71.395 90.060 71.655 ;
        RECT 89.160 70.965 89.420 71.225 ;
        RECT 89.480 70.965 89.740 71.225 ;
        RECT 89.800 70.965 90.060 71.225 ;
        RECT 91.155 71.300 91.415 71.560 ;
        RECT 91.155 70.980 91.415 71.240 ;
        RECT 89.160 70.535 89.420 70.795 ;
        RECT 89.480 70.535 89.740 70.795 ;
        RECT 89.800 70.535 90.060 70.795 ;
        RECT 89.160 70.105 89.420 70.365 ;
        RECT 89.480 70.105 89.740 70.365 ;
        RECT 89.800 70.105 90.060 70.365 ;
        RECT 93.010 71.395 93.270 71.655 ;
        RECT 93.330 71.395 93.590 71.655 ;
        RECT 93.650 71.395 93.910 71.655 ;
        RECT 93.010 70.965 93.270 71.225 ;
        RECT 93.330 70.965 93.590 71.225 ;
        RECT 93.650 70.965 93.910 71.225 ;
        RECT 93.010 70.535 93.270 70.795 ;
        RECT 93.330 70.535 93.590 70.795 ;
        RECT 93.650 70.535 93.910 70.795 ;
        RECT 92.530 70.105 92.790 70.365 ;
        RECT 92.850 70.105 93.110 70.365 ;
        RECT 93.170 70.105 93.430 70.365 ;
        RECT 93.490 70.105 93.750 70.365 ;
        RECT 93.810 70.105 94.070 70.365 ;
        RECT 94.130 70.105 94.390 70.365 ;
        RECT 89.160 69.675 89.420 69.935 ;
        RECT 89.480 69.675 89.740 69.935 ;
        RECT 89.800 69.675 90.060 69.935 ;
        RECT 93.010 69.675 93.270 69.935 ;
        RECT 93.330 69.675 93.590 69.935 ;
        RECT 93.650 69.675 93.910 69.935 ;
        RECT 89.160 69.245 89.420 69.505 ;
        RECT 89.480 69.245 89.740 69.505 ;
        RECT 89.800 69.245 90.060 69.505 ;
        RECT 90.835 69.245 91.095 69.505 ;
        RECT 91.155 69.245 91.415 69.505 ;
        RECT 91.475 69.245 91.735 69.505 ;
        RECT 89.160 68.815 89.420 69.075 ;
        RECT 89.480 68.815 89.740 69.075 ;
        RECT 89.800 68.815 90.060 69.075 ;
        RECT 89.160 68.385 89.420 68.645 ;
        RECT 89.480 68.385 89.740 68.645 ;
        RECT 89.800 68.385 90.060 68.645 ;
        RECT 89.160 67.955 89.420 68.215 ;
        RECT 89.480 67.955 89.740 68.215 ;
        RECT 89.800 67.955 90.060 68.215 ;
        RECT 89.160 67.525 89.420 67.785 ;
        RECT 89.480 67.525 89.740 67.785 ;
        RECT 89.800 67.525 90.060 67.785 ;
        RECT 89.160 67.095 89.420 67.355 ;
        RECT 89.480 67.095 89.740 67.355 ;
        RECT 89.800 67.095 90.060 67.355 ;
        RECT 92.530 69.245 92.790 69.505 ;
        RECT 92.850 69.245 93.110 69.505 ;
        RECT 93.170 69.245 93.430 69.505 ;
        RECT 93.490 69.245 93.750 69.505 ;
        RECT 93.810 69.245 94.070 69.505 ;
        RECT 94.130 69.245 94.390 69.505 ;
        RECT 93.010 68.815 93.270 69.075 ;
        RECT 93.330 68.815 93.590 69.075 ;
        RECT 93.650 68.815 93.910 69.075 ;
        RECT 92.530 68.385 92.790 68.645 ;
        RECT 92.850 68.385 93.110 68.645 ;
        RECT 93.170 68.385 93.430 68.645 ;
        RECT 93.490 68.385 93.750 68.645 ;
        RECT 93.810 68.385 94.070 68.645 ;
        RECT 94.130 68.385 94.390 68.645 ;
        RECT 93.010 67.955 93.270 68.215 ;
        RECT 93.330 67.955 93.590 68.215 ;
        RECT 93.650 67.955 93.910 68.215 ;
        RECT 92.530 67.525 92.790 67.785 ;
        RECT 92.850 67.525 93.110 67.785 ;
        RECT 93.170 67.525 93.430 67.785 ;
        RECT 93.490 67.525 93.750 67.785 ;
        RECT 93.810 67.525 94.070 67.785 ;
        RECT 94.130 67.525 94.390 67.785 ;
        RECT 93.010 67.095 93.270 67.355 ;
        RECT 93.330 67.095 93.590 67.355 ;
        RECT 93.650 67.095 93.910 67.355 ;
        RECT 89.160 66.665 89.420 66.925 ;
        RECT 89.480 66.665 89.740 66.925 ;
        RECT 89.800 66.665 90.060 66.925 ;
        RECT 92.530 66.665 92.790 66.925 ;
        RECT 92.850 66.665 93.110 66.925 ;
        RECT 93.170 66.665 93.430 66.925 ;
        RECT 93.490 66.665 93.750 66.925 ;
        RECT 93.810 66.665 94.070 66.925 ;
        RECT 94.130 66.665 94.390 66.925 ;
        RECT 89.160 66.235 89.420 66.495 ;
        RECT 89.480 66.235 89.740 66.495 ;
        RECT 89.800 66.235 90.060 66.495 ;
        RECT 89.160 65.805 89.420 66.065 ;
        RECT 89.480 65.805 89.740 66.065 ;
        RECT 89.800 65.805 90.060 66.065 ;
        RECT 89.160 65.375 89.420 65.635 ;
        RECT 89.480 65.375 89.740 65.635 ;
        RECT 89.800 65.375 90.060 65.635 ;
        RECT 89.160 64.945 89.420 65.205 ;
        RECT 89.480 64.945 89.740 65.205 ;
        RECT 89.800 64.945 90.060 65.205 ;
        RECT 93.010 66.235 93.270 66.495 ;
        RECT 93.330 66.235 93.590 66.495 ;
        RECT 93.650 66.235 93.910 66.495 ;
        RECT 92.530 65.805 92.790 66.065 ;
        RECT 92.850 65.805 93.110 66.065 ;
        RECT 93.170 65.805 93.430 66.065 ;
        RECT 93.490 65.805 93.750 66.065 ;
        RECT 93.810 65.805 94.070 66.065 ;
        RECT 94.130 65.805 94.390 66.065 ;
        RECT 93.010 65.375 93.270 65.635 ;
        RECT 93.330 65.375 93.590 65.635 ;
        RECT 93.650 65.375 93.910 65.635 ;
        RECT 92.530 64.945 92.790 65.205 ;
        RECT 92.850 64.945 93.110 65.205 ;
        RECT 93.170 64.945 93.430 65.205 ;
        RECT 93.490 64.945 93.750 65.205 ;
        RECT 93.810 64.945 94.070 65.205 ;
        RECT 94.130 64.945 94.390 65.205 ;
        RECT 89.160 64.515 89.420 64.775 ;
        RECT 89.480 64.515 89.740 64.775 ;
        RECT 89.800 64.515 90.060 64.775 ;
        RECT 93.010 64.515 93.270 64.775 ;
        RECT 93.330 64.515 93.590 64.775 ;
        RECT 93.650 64.515 93.910 64.775 ;
        RECT 89.160 64.085 89.420 64.345 ;
        RECT 89.480 64.085 89.740 64.345 ;
        RECT 89.800 64.085 90.060 64.345 ;
        RECT 89.160 63.655 89.420 63.915 ;
        RECT 89.480 63.655 89.740 63.915 ;
        RECT 89.800 63.655 90.060 63.915 ;
        RECT 93.010 64.085 93.270 64.345 ;
        RECT 93.330 64.085 93.590 64.345 ;
        RECT 93.650 64.085 93.910 64.345 ;
        RECT 93.010 63.655 93.270 63.915 ;
        RECT 93.330 63.655 93.590 63.915 ;
        RECT 93.650 63.655 93.910 63.915 ;
        RECT 89.160 62.985 89.420 63.245 ;
        RECT 89.480 62.985 89.740 63.245 ;
        RECT 89.800 62.985 90.060 63.245 ;
        RECT 93.010 62.985 93.270 63.245 ;
        RECT 93.330 62.985 93.590 63.245 ;
        RECT 93.650 62.985 93.910 63.245 ;
        RECT 109.665 163.785 109.925 164.045 ;
        RECT 109.985 163.785 110.245 164.045 ;
        RECT 109.665 161.505 109.925 161.765 ;
        RECT 109.985 161.505 110.245 161.765 ;
        RECT 111.035 163.785 111.295 164.045 ;
        RECT 111.355 163.785 111.615 164.045 ;
        RECT 111.035 161.505 111.295 161.765 ;
        RECT 111.355 161.505 111.615 161.765 ;
        RECT 112.405 163.785 112.665 164.045 ;
        RECT 112.725 163.785 112.985 164.045 ;
        RECT 112.405 161.505 112.665 161.765 ;
        RECT 112.725 161.505 112.985 161.765 ;
        RECT 109.665 159.225 109.925 159.485 ;
        RECT 109.985 159.225 110.245 159.485 ;
        RECT 111.035 159.225 111.295 159.485 ;
        RECT 111.355 159.225 111.615 159.485 ;
        RECT 112.405 159.225 112.665 159.485 ;
        RECT 112.725 159.225 112.985 159.485 ;
        RECT 109.665 156.945 109.925 157.205 ;
        RECT 109.985 156.945 110.245 157.205 ;
        RECT 111.035 156.945 111.295 157.205 ;
        RECT 111.355 156.945 111.615 157.205 ;
        RECT 112.405 156.945 112.665 157.205 ;
        RECT 112.725 156.945 112.985 157.205 ;
        RECT 109.665 154.665 109.925 154.925 ;
        RECT 109.985 154.665 110.245 154.925 ;
        RECT 111.035 154.665 111.295 154.925 ;
        RECT 111.355 154.665 111.615 154.925 ;
        RECT 112.405 154.665 112.665 154.925 ;
        RECT 112.725 154.665 112.985 154.925 ;
        RECT 109.665 152.385 109.925 152.645 ;
        RECT 109.985 152.385 110.245 152.645 ;
        RECT 111.035 152.385 111.295 152.645 ;
        RECT 111.355 152.385 111.615 152.645 ;
        RECT 112.405 152.385 112.665 152.645 ;
        RECT 112.725 152.385 112.985 152.645 ;
        RECT 109.665 150.105 109.925 150.365 ;
        RECT 109.985 150.105 110.245 150.365 ;
        RECT 111.035 150.105 111.295 150.365 ;
        RECT 111.355 150.105 111.615 150.365 ;
        RECT 112.405 150.105 112.665 150.365 ;
        RECT 112.725 150.105 112.985 150.365 ;
        RECT 109.665 147.825 109.925 148.085 ;
        RECT 109.985 147.825 110.245 148.085 ;
        RECT 111.035 147.825 111.295 148.085 ;
        RECT 111.355 147.825 111.615 148.085 ;
        RECT 112.405 147.825 112.665 148.085 ;
        RECT 112.725 147.825 112.985 148.085 ;
        RECT 109.665 145.545 109.925 145.805 ;
        RECT 109.985 145.545 110.245 145.805 ;
        RECT 111.035 145.545 111.295 145.805 ;
        RECT 111.355 145.545 111.615 145.805 ;
        RECT 112.405 145.545 112.665 145.805 ;
        RECT 112.725 145.545 112.985 145.805 ;
        RECT 109.665 143.265 109.925 143.525 ;
        RECT 109.985 143.265 110.245 143.525 ;
        RECT 111.035 143.265 111.295 143.525 ;
        RECT 111.355 143.265 111.615 143.525 ;
        RECT 112.405 143.265 112.665 143.525 ;
        RECT 112.725 143.265 112.985 143.525 ;
        RECT 109.665 140.985 109.925 141.245 ;
        RECT 109.985 140.985 110.245 141.245 ;
        RECT 111.035 140.985 111.295 141.245 ;
        RECT 111.355 140.985 111.615 141.245 ;
        RECT 112.405 140.985 112.665 141.245 ;
        RECT 112.725 140.985 112.985 141.245 ;
        RECT 109.665 138.705 109.925 138.965 ;
        RECT 109.985 138.705 110.245 138.965 ;
        RECT 111.035 138.705 111.295 138.965 ;
        RECT 111.355 138.705 111.615 138.965 ;
        RECT 112.405 138.705 112.665 138.965 ;
        RECT 112.725 138.705 112.985 138.965 ;
        RECT 109.665 136.425 109.925 136.685 ;
        RECT 109.985 136.425 110.245 136.685 ;
        RECT 109.665 134.145 109.925 134.405 ;
        RECT 109.985 134.145 110.245 134.405 ;
        RECT 109.665 131.865 109.925 132.125 ;
        RECT 109.985 131.865 110.245 132.125 ;
        RECT 109.665 129.585 109.925 129.845 ;
        RECT 109.985 129.585 110.245 129.845 ;
        RECT 109.665 127.305 109.925 127.565 ;
        RECT 109.985 127.305 110.245 127.565 ;
        RECT 109.665 125.025 109.925 125.285 ;
        RECT 109.985 125.025 110.245 125.285 ;
        RECT 109.665 122.745 109.925 123.005 ;
        RECT 109.985 122.745 110.245 123.005 ;
        RECT 109.665 120.465 109.925 120.725 ;
        RECT 109.985 120.465 110.245 120.725 ;
        RECT 109.665 118.185 109.925 118.445 ;
        RECT 109.985 118.185 110.245 118.445 ;
        RECT 109.665 115.905 109.925 116.165 ;
        RECT 109.985 115.905 110.245 116.165 ;
        RECT 109.665 113.625 109.925 113.885 ;
        RECT 109.985 113.625 110.245 113.885 ;
        RECT 109.665 111.345 109.925 111.605 ;
        RECT 109.985 111.345 110.245 111.605 ;
        RECT 109.665 109.065 109.925 109.325 ;
        RECT 109.985 109.065 110.245 109.325 ;
        RECT 109.665 106.785 109.925 107.045 ;
        RECT 109.985 106.785 110.245 107.045 ;
        RECT 109.665 104.505 109.925 104.765 ;
        RECT 109.985 104.505 110.245 104.765 ;
        RECT 109.665 102.225 109.925 102.485 ;
        RECT 109.985 102.225 110.245 102.485 ;
        RECT 109.665 99.945 109.925 100.205 ;
        RECT 109.985 99.945 110.245 100.205 ;
        RECT 109.665 97.665 109.925 97.925 ;
        RECT 109.985 97.665 110.245 97.925 ;
        RECT 109.665 95.385 109.925 95.645 ;
        RECT 109.985 95.385 110.245 95.645 ;
        RECT 109.665 93.105 109.925 93.365 ;
        RECT 109.985 93.105 110.245 93.365 ;
        RECT 109.665 90.825 109.925 91.085 ;
        RECT 109.985 90.825 110.245 91.085 ;
        RECT 109.665 88.545 109.925 88.805 ;
        RECT 109.985 88.545 110.245 88.805 ;
        RECT 109.665 86.265 109.925 86.525 ;
        RECT 109.985 86.265 110.245 86.525 ;
        RECT 109.665 83.985 109.925 84.245 ;
        RECT 109.985 83.985 110.245 84.245 ;
        RECT 109.665 81.705 109.925 81.965 ;
        RECT 109.985 81.705 110.245 81.965 ;
        RECT 109.665 79.425 109.925 79.685 ;
        RECT 109.985 79.425 110.245 79.685 ;
        RECT 109.665 77.145 109.925 77.405 ;
        RECT 109.985 77.145 110.245 77.405 ;
        RECT 109.665 74.865 109.925 75.125 ;
        RECT 109.985 74.865 110.245 75.125 ;
        RECT 109.665 72.585 109.925 72.845 ;
        RECT 109.985 72.585 110.245 72.845 ;
        RECT 109.665 70.305 109.925 70.565 ;
        RECT 109.985 70.305 110.245 70.565 ;
        RECT 111.035 136.425 111.295 136.685 ;
        RECT 111.355 136.425 111.615 136.685 ;
        RECT 111.035 134.145 111.295 134.405 ;
        RECT 111.355 134.145 111.615 134.405 ;
        RECT 111.035 131.865 111.295 132.125 ;
        RECT 111.355 131.865 111.615 132.125 ;
        RECT 111.035 129.585 111.295 129.845 ;
        RECT 111.355 129.585 111.615 129.845 ;
        RECT 111.035 127.305 111.295 127.565 ;
        RECT 111.355 127.305 111.615 127.565 ;
        RECT 111.035 125.025 111.295 125.285 ;
        RECT 111.355 125.025 111.615 125.285 ;
        RECT 111.035 122.745 111.295 123.005 ;
        RECT 111.355 122.745 111.615 123.005 ;
        RECT 111.035 120.465 111.295 120.725 ;
        RECT 111.355 120.465 111.615 120.725 ;
        RECT 111.035 118.185 111.295 118.445 ;
        RECT 111.355 118.185 111.615 118.445 ;
        RECT 111.035 115.905 111.295 116.165 ;
        RECT 111.355 115.905 111.615 116.165 ;
        RECT 111.035 113.625 111.295 113.885 ;
        RECT 111.355 113.625 111.615 113.885 ;
        RECT 111.035 111.345 111.295 111.605 ;
        RECT 111.355 111.345 111.615 111.605 ;
        RECT 111.035 109.065 111.295 109.325 ;
        RECT 111.355 109.065 111.615 109.325 ;
        RECT 111.035 106.785 111.295 107.045 ;
        RECT 111.355 106.785 111.615 107.045 ;
        RECT 111.035 104.505 111.295 104.765 ;
        RECT 111.355 104.505 111.615 104.765 ;
        RECT 111.035 102.225 111.295 102.485 ;
        RECT 111.355 102.225 111.615 102.485 ;
        RECT 111.035 99.945 111.295 100.205 ;
        RECT 111.355 99.945 111.615 100.205 ;
        RECT 112.405 136.425 112.665 136.685 ;
        RECT 112.725 136.425 112.985 136.685 ;
        RECT 112.405 134.145 112.665 134.405 ;
        RECT 112.725 134.145 112.985 134.405 ;
        RECT 112.405 131.865 112.665 132.125 ;
        RECT 112.725 131.865 112.985 132.125 ;
        RECT 112.405 129.585 112.665 129.845 ;
        RECT 112.725 129.585 112.985 129.845 ;
        RECT 112.405 127.305 112.665 127.565 ;
        RECT 112.725 127.305 112.985 127.565 ;
        RECT 112.405 125.025 112.665 125.285 ;
        RECT 112.725 125.025 112.985 125.285 ;
        RECT 112.405 122.745 112.665 123.005 ;
        RECT 112.725 122.745 112.985 123.005 ;
        RECT 112.405 120.465 112.665 120.725 ;
        RECT 112.725 120.465 112.985 120.725 ;
        RECT 112.405 118.185 112.665 118.445 ;
        RECT 112.725 118.185 112.985 118.445 ;
        RECT 112.405 115.905 112.665 116.165 ;
        RECT 112.725 115.905 112.985 116.165 ;
        RECT 112.405 113.625 112.665 113.885 ;
        RECT 112.725 113.625 112.985 113.885 ;
        RECT 122.870 164.415 123.130 164.675 ;
        RECT 123.190 164.415 123.450 164.675 ;
        RECT 124.240 164.415 124.500 164.675 ;
        RECT 124.560 164.415 124.820 164.675 ;
        RECT 115.410 116.825 115.670 117.085 ;
        RECT 115.410 116.505 115.670 116.765 ;
        RECT 115.955 116.370 116.215 116.630 ;
        RECT 116.275 116.370 116.535 116.630 ;
        RECT 115.955 115.940 116.215 116.200 ;
        RECT 116.275 115.940 116.535 116.200 ;
        RECT 115.955 115.510 116.215 115.770 ;
        RECT 116.275 115.510 116.535 115.770 ;
        RECT 122.870 163.785 123.130 164.045 ;
        RECT 123.190 163.785 123.450 164.045 ;
        RECT 123.715 163.635 123.975 163.895 ;
        RECT 124.240 163.785 124.500 164.045 ;
        RECT 124.560 163.785 124.820 164.045 ;
        RECT 123.715 163.315 123.975 163.575 ;
        RECT 123.715 162.995 123.975 163.255 ;
        RECT 123.715 162.675 123.975 162.935 ;
        RECT 123.715 162.355 123.975 162.615 ;
        RECT 123.715 162.035 123.975 162.295 ;
        RECT 122.870 161.505 123.130 161.765 ;
        RECT 123.190 161.505 123.450 161.765 ;
        RECT 123.715 161.715 123.975 161.975 ;
        RECT 123.715 161.395 123.975 161.655 ;
        RECT 124.240 161.505 124.500 161.765 ;
        RECT 124.560 161.505 124.820 161.765 ;
        RECT 123.715 161.075 123.975 161.335 ;
        RECT 123.715 160.755 123.975 161.015 ;
        RECT 123.715 160.435 123.975 160.695 ;
        RECT 123.715 160.115 123.975 160.375 ;
        RECT 123.715 159.795 123.975 160.055 ;
        RECT 122.870 159.225 123.130 159.485 ;
        RECT 123.190 159.225 123.450 159.485 ;
        RECT 123.715 159.475 123.975 159.735 ;
        RECT 123.715 159.155 123.975 159.415 ;
        RECT 124.240 159.225 124.500 159.485 ;
        RECT 124.560 159.225 124.820 159.485 ;
        RECT 123.715 158.835 123.975 159.095 ;
        RECT 123.715 158.515 123.975 158.775 ;
        RECT 123.715 158.195 123.975 158.455 ;
        RECT 123.715 157.875 123.975 158.135 ;
        RECT 123.715 157.555 123.975 157.815 ;
        RECT 123.715 157.235 123.975 157.495 ;
        RECT 122.870 156.945 123.130 157.205 ;
        RECT 123.190 156.945 123.450 157.205 ;
        RECT 123.715 156.915 123.975 157.175 ;
        RECT 124.240 156.945 124.500 157.205 ;
        RECT 124.560 156.945 124.820 157.205 ;
        RECT 123.715 156.595 123.975 156.855 ;
        RECT 123.715 156.275 123.975 156.535 ;
        RECT 123.715 155.955 123.975 156.215 ;
        RECT 123.715 155.635 123.975 155.895 ;
        RECT 123.715 155.315 123.975 155.575 ;
        RECT 123.715 154.995 123.975 155.255 ;
        RECT 122.870 154.665 123.130 154.925 ;
        RECT 123.190 154.665 123.450 154.925 ;
        RECT 123.715 154.675 123.975 154.935 ;
        RECT 124.240 154.665 124.500 154.925 ;
        RECT 124.560 154.665 124.820 154.925 ;
        RECT 123.715 154.355 123.975 154.615 ;
        RECT 123.715 154.035 123.975 154.295 ;
        RECT 123.715 153.715 123.975 153.975 ;
        RECT 123.715 153.395 123.975 153.655 ;
        RECT 123.715 153.075 123.975 153.335 ;
        RECT 123.715 152.755 123.975 153.015 ;
        RECT 122.870 152.385 123.130 152.645 ;
        RECT 123.190 152.385 123.450 152.645 ;
        RECT 123.715 152.435 123.975 152.695 ;
        RECT 124.240 152.385 124.500 152.645 ;
        RECT 124.560 152.385 124.820 152.645 ;
        RECT 123.715 152.115 123.975 152.375 ;
        RECT 123.715 151.795 123.975 152.055 ;
        RECT 123.715 151.475 123.975 151.735 ;
        RECT 123.715 151.155 123.975 151.415 ;
        RECT 123.715 150.835 123.975 151.095 ;
        RECT 123.715 150.515 123.975 150.775 ;
        RECT 122.870 150.105 123.130 150.365 ;
        RECT 123.190 150.105 123.450 150.365 ;
        RECT 123.715 150.195 123.975 150.455 ;
        RECT 123.715 149.875 123.975 150.135 ;
        RECT 124.240 150.105 124.500 150.365 ;
        RECT 124.560 150.105 124.820 150.365 ;
        RECT 123.715 149.555 123.975 149.815 ;
        RECT 123.715 149.235 123.975 149.495 ;
        RECT 123.715 148.915 123.975 149.175 ;
        RECT 123.715 148.595 123.975 148.855 ;
        RECT 123.715 148.275 123.975 148.535 ;
        RECT 122.870 147.825 123.130 148.085 ;
        RECT 123.190 147.825 123.450 148.085 ;
        RECT 123.715 147.955 123.975 148.215 ;
        RECT 123.715 147.635 123.975 147.895 ;
        RECT 124.240 147.825 124.500 148.085 ;
        RECT 124.560 147.825 124.820 148.085 ;
        RECT 123.715 147.315 123.975 147.575 ;
        RECT 123.715 146.995 123.975 147.255 ;
        RECT 123.715 146.675 123.975 146.935 ;
        RECT 123.715 146.355 123.975 146.615 ;
        RECT 123.715 146.035 123.975 146.295 ;
        RECT 122.870 145.545 123.130 145.805 ;
        RECT 123.190 145.545 123.450 145.805 ;
        RECT 123.715 145.715 123.975 145.975 ;
        RECT 123.715 145.395 123.975 145.655 ;
        RECT 124.240 145.545 124.500 145.805 ;
        RECT 124.560 145.545 124.820 145.805 ;
        RECT 123.715 145.075 123.975 145.335 ;
        RECT 123.715 144.755 123.975 145.015 ;
        RECT 123.715 144.435 123.975 144.695 ;
        RECT 123.715 144.115 123.975 144.375 ;
        RECT 123.715 143.795 123.975 144.055 ;
        RECT 122.870 143.265 123.130 143.525 ;
        RECT 123.190 143.265 123.450 143.525 ;
        RECT 123.715 143.475 123.975 143.735 ;
        RECT 123.715 143.155 123.975 143.415 ;
        RECT 124.240 143.265 124.500 143.525 ;
        RECT 124.560 143.265 124.820 143.525 ;
        RECT 123.715 142.835 123.975 143.095 ;
        RECT 123.715 142.515 123.975 142.775 ;
        RECT 123.715 142.195 123.975 142.455 ;
        RECT 123.715 141.875 123.975 142.135 ;
        RECT 123.715 141.555 123.975 141.815 ;
        RECT 122.870 140.985 123.130 141.245 ;
        RECT 123.190 140.985 123.450 141.245 ;
        RECT 123.715 141.235 123.975 141.495 ;
        RECT 123.715 140.915 123.975 141.175 ;
        RECT 124.240 140.985 124.500 141.245 ;
        RECT 124.560 140.985 124.820 141.245 ;
        RECT 123.715 140.595 123.975 140.855 ;
        RECT 123.715 140.275 123.975 140.535 ;
        RECT 123.715 139.955 123.975 140.215 ;
        RECT 123.715 139.635 123.975 139.895 ;
        RECT 123.715 139.315 123.975 139.575 ;
        RECT 123.715 138.995 123.975 139.255 ;
        RECT 122.870 138.705 123.130 138.965 ;
        RECT 123.190 138.705 123.450 138.965 ;
        RECT 123.715 138.675 123.975 138.935 ;
        RECT 124.240 138.705 124.500 138.965 ;
        RECT 124.560 138.705 124.820 138.965 ;
        RECT 123.715 138.355 123.975 138.615 ;
        RECT 123.715 138.035 123.975 138.295 ;
        RECT 123.715 137.715 123.975 137.975 ;
        RECT 123.715 137.395 123.975 137.655 ;
        RECT 123.715 137.075 123.975 137.335 ;
        RECT 123.715 136.755 123.975 137.015 ;
        RECT 122.870 136.425 123.130 136.685 ;
        RECT 123.190 136.425 123.450 136.685 ;
        RECT 123.715 136.435 123.975 136.695 ;
        RECT 122.870 134.145 123.130 134.405 ;
        RECT 123.190 134.145 123.450 134.405 ;
        RECT 122.870 131.865 123.130 132.125 ;
        RECT 123.190 131.865 123.450 132.125 ;
        RECT 122.870 129.585 123.130 129.845 ;
        RECT 123.190 129.585 123.450 129.845 ;
        RECT 122.870 127.305 123.130 127.565 ;
        RECT 123.190 127.305 123.450 127.565 ;
        RECT 122.870 125.025 123.130 125.285 ;
        RECT 123.190 125.025 123.450 125.285 ;
        RECT 122.870 122.745 123.130 123.005 ;
        RECT 123.190 122.745 123.450 123.005 ;
        RECT 122.870 120.465 123.130 120.725 ;
        RECT 123.190 120.465 123.450 120.725 ;
        RECT 122.870 118.185 123.130 118.445 ;
        RECT 123.190 118.185 123.450 118.445 ;
        RECT 122.870 115.905 123.130 116.165 ;
        RECT 123.190 115.905 123.450 116.165 ;
        RECT 119.215 113.985 119.475 114.245 ;
        RECT 119.535 113.985 119.795 114.245 ;
        RECT 119.855 113.985 120.115 114.245 ;
        RECT 120.390 113.880 120.650 114.140 ;
        RECT 112.405 111.345 112.665 111.605 ;
        RECT 112.725 111.345 112.985 111.605 ;
        RECT 115.955 111.700 116.215 111.960 ;
        RECT 116.275 111.700 116.535 111.960 ;
        RECT 112.405 109.065 112.665 109.325 ;
        RECT 112.725 109.065 112.985 109.325 ;
        RECT 112.405 106.785 112.665 107.045 ;
        RECT 112.725 106.785 112.985 107.045 ;
        RECT 112.405 104.505 112.665 104.765 ;
        RECT 112.725 104.505 112.985 104.765 ;
        RECT 112.405 102.225 112.665 102.485 ;
        RECT 112.725 102.225 112.985 102.485 ;
        RECT 112.405 99.945 112.665 100.205 ;
        RECT 112.725 99.945 112.985 100.205 ;
        RECT 111.880 99.245 112.140 99.505 ;
        RECT 111.880 98.925 112.140 99.185 ;
        RECT 111.880 98.605 112.140 98.865 ;
        RECT 111.880 98.285 112.140 98.545 ;
        RECT 111.035 97.665 111.295 97.925 ;
        RECT 111.355 97.665 111.615 97.925 ;
        RECT 111.035 95.385 111.295 95.645 ;
        RECT 111.355 95.385 111.615 95.645 ;
        RECT 111.035 93.105 111.295 93.365 ;
        RECT 111.355 93.105 111.615 93.365 ;
        RECT 111.035 90.825 111.295 91.085 ;
        RECT 111.355 90.825 111.615 91.085 ;
        RECT 111.035 88.545 111.295 88.805 ;
        RECT 111.355 88.545 111.615 88.805 ;
        RECT 111.035 86.265 111.295 86.525 ;
        RECT 111.355 86.265 111.615 86.525 ;
        RECT 111.035 83.985 111.295 84.245 ;
        RECT 111.355 83.985 111.615 84.245 ;
        RECT 111.035 81.705 111.295 81.965 ;
        RECT 111.355 81.705 111.615 81.965 ;
        RECT 111.035 79.425 111.295 79.685 ;
        RECT 111.355 79.425 111.615 79.685 ;
        RECT 111.035 77.145 111.295 77.405 ;
        RECT 111.355 77.145 111.615 77.405 ;
        RECT 111.035 74.865 111.295 75.125 ;
        RECT 111.355 74.865 111.615 75.125 ;
        RECT 111.035 72.585 111.295 72.845 ;
        RECT 111.355 72.585 111.615 72.845 ;
        RECT 111.035 70.305 111.295 70.565 ;
        RECT 111.355 70.305 111.615 70.565 ;
        RECT 112.405 97.665 112.665 97.925 ;
        RECT 112.725 97.665 112.985 97.925 ;
        RECT 112.405 95.385 112.665 95.645 ;
        RECT 112.725 95.385 112.985 95.645 ;
        RECT 112.405 93.105 112.665 93.365 ;
        RECT 112.725 93.105 112.985 93.365 ;
        RECT 112.405 90.825 112.665 91.085 ;
        RECT 112.725 90.825 112.985 91.085 ;
        RECT 112.405 88.545 112.665 88.805 ;
        RECT 112.725 88.545 112.985 88.805 ;
        RECT 112.405 86.265 112.665 86.525 ;
        RECT 112.725 86.265 112.985 86.525 ;
        RECT 112.405 83.985 112.665 84.245 ;
        RECT 112.725 83.985 112.985 84.245 ;
        RECT 112.405 81.705 112.665 81.965 ;
        RECT 112.725 81.705 112.985 81.965 ;
        RECT 112.405 79.425 112.665 79.685 ;
        RECT 112.725 79.425 112.985 79.685 ;
        RECT 115.955 111.270 116.215 111.530 ;
        RECT 116.275 111.270 116.535 111.530 ;
        RECT 115.955 110.840 116.215 111.100 ;
        RECT 116.275 110.840 116.535 111.100 ;
        RECT 116.820 110.275 117.080 110.535 ;
        RECT 116.820 109.955 117.080 110.215 ;
        RECT 120.390 113.560 120.650 113.820 ;
        RECT 119.215 113.125 119.475 113.385 ;
        RECT 119.535 113.125 119.795 113.385 ;
        RECT 119.855 113.125 120.115 113.385 ;
        RECT 120.390 113.240 120.650 113.500 ;
        RECT 122.870 113.625 123.130 113.885 ;
        RECT 123.190 113.625 123.450 113.885 ;
        RECT 115.410 82.625 115.670 82.885 ;
        RECT 115.410 82.305 115.670 82.565 ;
        RECT 115.955 82.170 116.215 82.430 ;
        RECT 116.275 82.170 116.535 82.430 ;
        RECT 115.955 81.740 116.215 82.000 ;
        RECT 116.275 81.740 116.535 82.000 ;
        RECT 115.955 81.310 116.215 81.570 ;
        RECT 116.275 81.310 116.535 81.570 ;
        RECT 119.215 79.785 119.475 80.045 ;
        RECT 119.535 79.785 119.795 80.045 ;
        RECT 119.855 79.785 120.115 80.045 ;
        RECT 120.390 79.680 120.650 79.940 ;
        RECT 112.405 77.145 112.665 77.405 ;
        RECT 112.725 77.145 112.985 77.405 ;
        RECT 115.955 77.500 116.215 77.760 ;
        RECT 116.275 77.500 116.535 77.760 ;
        RECT 112.405 74.865 112.665 75.125 ;
        RECT 112.725 74.865 112.985 75.125 ;
        RECT 112.405 72.585 112.665 72.845 ;
        RECT 112.725 72.585 112.985 72.845 ;
        RECT 112.405 70.305 112.665 70.565 ;
        RECT 112.725 70.305 112.985 70.565 ;
        RECT 111.880 69.490 112.140 69.750 ;
        RECT 111.880 69.170 112.140 69.430 ;
        RECT 111.880 68.850 112.140 69.110 ;
        RECT 109.665 68.025 109.925 68.285 ;
        RECT 109.985 68.025 110.245 68.285 ;
        RECT 111.035 68.025 111.295 68.285 ;
        RECT 111.355 68.025 111.615 68.285 ;
        RECT 112.405 68.025 112.665 68.285 ;
        RECT 112.725 68.025 112.985 68.285 ;
        RECT 109.665 65.745 109.925 66.005 ;
        RECT 109.985 65.745 110.245 66.005 ;
        RECT 109.665 63.465 109.925 63.725 ;
        RECT 109.985 63.465 110.245 63.725 ;
        RECT 111.035 65.745 111.295 66.005 ;
        RECT 111.355 65.745 111.615 66.005 ;
        RECT 111.035 63.465 111.295 63.725 ;
        RECT 111.355 63.465 111.615 63.725 ;
        RECT 112.405 65.745 112.665 66.005 ;
        RECT 112.725 65.745 112.985 66.005 ;
        RECT 112.405 63.465 112.665 63.725 ;
        RECT 112.725 63.465 112.985 63.725 ;
        RECT 115.955 77.070 116.215 77.330 ;
        RECT 116.275 77.070 116.535 77.330 ;
        RECT 115.955 76.640 116.215 76.900 ;
        RECT 116.275 76.640 116.535 76.900 ;
        RECT 116.820 76.075 117.080 76.335 ;
        RECT 116.820 75.755 117.080 76.015 ;
        RECT 115.805 75.110 116.065 75.370 ;
        RECT 116.125 75.110 116.385 75.370 ;
        RECT 120.390 79.360 120.650 79.620 ;
        RECT 119.215 78.925 119.475 79.185 ;
        RECT 119.535 78.925 119.795 79.185 ;
        RECT 119.855 78.925 120.115 79.185 ;
        RECT 120.390 79.040 120.650 79.300 ;
        RECT 122.870 111.345 123.130 111.605 ;
        RECT 123.190 111.345 123.450 111.605 ;
        RECT 122.870 109.065 123.130 109.325 ;
        RECT 123.190 109.065 123.450 109.325 ;
        RECT 122.870 106.785 123.130 107.045 ;
        RECT 123.190 106.785 123.450 107.045 ;
        RECT 122.870 104.505 123.130 104.765 ;
        RECT 123.190 104.505 123.450 104.765 ;
        RECT 122.870 102.225 123.130 102.485 ;
        RECT 123.190 102.225 123.450 102.485 ;
        RECT 122.870 99.945 123.130 100.205 ;
        RECT 123.190 99.945 123.450 100.205 ;
        RECT 122.870 97.665 123.130 97.925 ;
        RECT 123.190 97.665 123.450 97.925 ;
        RECT 122.870 95.385 123.130 95.645 ;
        RECT 123.190 95.385 123.450 95.645 ;
        RECT 122.870 93.105 123.130 93.365 ;
        RECT 123.190 93.105 123.450 93.365 ;
        RECT 122.870 90.825 123.130 91.085 ;
        RECT 123.190 90.825 123.450 91.085 ;
        RECT 122.870 88.545 123.130 88.805 ;
        RECT 123.190 88.545 123.450 88.805 ;
        RECT 122.870 86.265 123.130 86.525 ;
        RECT 123.190 86.265 123.450 86.525 ;
        RECT 122.870 83.985 123.130 84.245 ;
        RECT 123.190 83.985 123.450 84.245 ;
        RECT 122.345 83.160 122.605 83.420 ;
        RECT 122.345 82.840 122.605 83.100 ;
        RECT 122.345 82.520 122.605 82.780 ;
        RECT 124.240 136.425 124.500 136.685 ;
        RECT 124.560 136.425 124.820 136.685 ;
        RECT 124.240 134.145 124.500 134.405 ;
        RECT 124.560 134.145 124.820 134.405 ;
        RECT 124.240 131.865 124.500 132.125 ;
        RECT 124.560 131.865 124.820 132.125 ;
        RECT 124.240 129.585 124.500 129.845 ;
        RECT 124.560 129.585 124.820 129.845 ;
        RECT 124.240 127.305 124.500 127.565 ;
        RECT 124.560 127.305 124.820 127.565 ;
        RECT 124.240 125.025 124.500 125.285 ;
        RECT 124.560 125.025 124.820 125.285 ;
        RECT 124.240 122.745 124.500 123.005 ;
        RECT 124.560 122.745 124.820 123.005 ;
        RECT 124.240 120.465 124.500 120.725 ;
        RECT 124.560 120.465 124.820 120.725 ;
        RECT 124.240 118.185 124.500 118.445 ;
        RECT 124.560 118.185 124.820 118.445 ;
        RECT 124.240 115.905 124.500 116.165 ;
        RECT 124.560 115.905 124.820 116.165 ;
        RECT 124.240 113.625 124.500 113.885 ;
        RECT 124.560 113.625 124.820 113.885 ;
        RECT 124.240 111.345 124.500 111.605 ;
        RECT 124.560 111.345 124.820 111.605 ;
        RECT 124.240 109.065 124.500 109.325 ;
        RECT 124.560 109.065 124.820 109.325 ;
        RECT 124.240 106.785 124.500 107.045 ;
        RECT 124.560 106.785 124.820 107.045 ;
        RECT 124.240 104.505 124.500 104.765 ;
        RECT 124.560 104.505 124.820 104.765 ;
        RECT 124.240 102.225 124.500 102.485 ;
        RECT 124.560 102.225 124.820 102.485 ;
        RECT 124.240 99.945 124.500 100.205 ;
        RECT 124.560 99.945 124.820 100.205 ;
        RECT 124.240 97.665 124.500 97.925 ;
        RECT 124.560 97.665 124.820 97.925 ;
        RECT 124.240 95.385 124.500 95.645 ;
        RECT 124.560 95.385 124.820 95.645 ;
        RECT 124.240 93.105 124.500 93.365 ;
        RECT 124.560 93.105 124.820 93.365 ;
        RECT 124.240 90.825 124.500 91.085 ;
        RECT 124.560 90.825 124.820 91.085 ;
        RECT 124.240 88.545 124.500 88.805 ;
        RECT 124.560 88.545 124.820 88.805 ;
        RECT 124.240 86.265 124.500 86.525 ;
        RECT 124.560 86.265 124.820 86.525 ;
        RECT 124.240 83.985 124.500 84.245 ;
        RECT 124.560 83.985 124.820 84.245 ;
        RECT 123.715 83.160 123.975 83.420 ;
        RECT 123.715 82.840 123.975 83.100 ;
        RECT 123.715 82.520 123.975 82.780 ;
        RECT 122.870 81.705 123.130 81.965 ;
        RECT 123.190 81.705 123.450 81.965 ;
        RECT 124.240 81.705 124.500 81.965 ;
        RECT 124.560 81.705 124.820 81.965 ;
        RECT 122.870 79.425 123.130 79.685 ;
        RECT 123.190 79.425 123.450 79.685 ;
        RECT 124.240 79.425 124.500 79.685 ;
        RECT 124.560 79.425 124.820 79.685 ;
        RECT 122.870 77.145 123.130 77.405 ;
        RECT 123.190 77.145 123.450 77.405 ;
        RECT 124.240 77.145 124.500 77.405 ;
        RECT 124.560 77.145 124.820 77.405 ;
        RECT 122.870 76.515 123.130 76.775 ;
        RECT 123.190 76.515 123.450 76.775 ;
        RECT 124.240 76.515 124.500 76.775 ;
        RECT 124.560 76.515 124.820 76.775 ;
        RECT 109.665 62.795 109.925 63.055 ;
        RECT 109.985 62.795 110.245 63.055 ;
        RECT 111.035 62.795 111.295 63.055 ;
        RECT 111.355 62.795 111.615 63.055 ;
        RECT 112.405 62.795 112.665 63.055 ;
        RECT 112.725 62.795 112.985 63.055 ;
        RECT 115.805 70.335 116.065 70.595 ;
        RECT 116.125 70.335 116.385 70.595 ;
        RECT 115.805 69.665 116.065 69.925 ;
        RECT 116.125 69.665 116.385 69.925 ;
        RECT 115.260 69.180 115.520 69.440 ;
        RECT 115.260 68.860 115.520 69.120 ;
        RECT 115.260 68.540 115.520 68.800 ;
        RECT 119.500 70.055 119.760 70.315 ;
        RECT 119.820 70.055 120.080 70.315 ;
        RECT 119.500 69.385 119.760 69.645 ;
        RECT 119.820 69.385 120.080 69.645 ;
        RECT 120.365 69.470 120.625 69.730 ;
        RECT 119.500 68.955 119.760 69.215 ;
        RECT 119.820 68.955 120.080 69.215 ;
        RECT 120.365 69.150 120.625 69.410 ;
        RECT 119.500 68.525 119.760 68.785 ;
        RECT 119.820 68.525 120.080 68.785 ;
        RECT 119.500 68.110 119.760 68.370 ;
        RECT 119.820 68.110 120.080 68.370 ;
        RECT 115.805 67.385 116.065 67.645 ;
        RECT 116.125 67.385 116.385 67.645 ;
        RECT 115.805 65.105 116.065 65.365 ;
        RECT 116.125 65.105 116.385 65.365 ;
        RECT 115.805 62.825 116.065 63.085 ;
        RECT 116.125 62.825 116.385 63.085 ;
        RECT 115.805 60.545 116.065 60.805 ;
        RECT 116.125 60.545 116.385 60.805 ;
        RECT 119.500 67.665 119.760 67.925 ;
        RECT 119.820 67.665 120.080 67.925 ;
        RECT 119.500 67.250 119.760 67.510 ;
        RECT 119.820 67.250 120.080 67.510 ;
        RECT 123.080 69.480 123.340 69.740 ;
        RECT 123.080 69.160 123.340 69.420 ;
        RECT 123.080 68.840 123.340 69.100 ;
        RECT 122.215 68.525 122.475 68.785 ;
        RECT 122.535 68.525 122.795 68.785 ;
        RECT 122.215 68.095 122.475 68.355 ;
        RECT 122.535 68.095 122.795 68.355 ;
        RECT 122.215 67.665 122.475 67.925 ;
        RECT 122.535 67.665 122.795 67.925 ;
        RECT 122.215 67.235 122.475 67.495 ;
        RECT 122.535 67.235 122.795 67.495 ;
        RECT 119.500 66.805 119.760 67.065 ;
        RECT 119.820 66.805 120.080 67.065 ;
        RECT 122.215 66.805 122.475 67.065 ;
        RECT 122.535 66.805 122.795 67.065 ;
        RECT 119.500 66.375 119.760 66.635 ;
        RECT 119.820 66.375 120.080 66.635 ;
        RECT 119.500 65.945 119.760 66.205 ;
        RECT 119.820 65.945 120.080 66.205 ;
        RECT 125.485 70.015 125.745 70.275 ;
        RECT 125.805 70.015 126.065 70.275 ;
        RECT 115.805 59.875 116.065 60.135 ;
        RECT 116.125 59.875 116.385 60.135 ;
        RECT 119.500 64.135 119.760 64.395 ;
        RECT 119.820 64.135 120.080 64.395 ;
        RECT 120.475 64.110 120.735 64.370 ;
        RECT 119.500 63.705 119.760 63.965 ;
        RECT 119.820 63.705 120.080 63.965 ;
        RECT 120.475 63.790 120.735 64.050 ;
        RECT 119.500 63.275 119.760 63.535 ;
        RECT 119.820 63.275 120.080 63.535 ;
        RECT 120.475 63.470 120.735 63.730 ;
        RECT 119.500 62.860 119.760 63.120 ;
        RECT 119.820 62.860 120.080 63.120 ;
        RECT 119.500 62.415 119.760 62.675 ;
        RECT 119.820 62.415 120.080 62.675 ;
        RECT 119.500 62.000 119.760 62.260 ;
        RECT 119.820 62.000 120.080 62.260 ;
        RECT 122.215 63.275 122.475 63.535 ;
        RECT 122.535 63.275 122.795 63.535 ;
        RECT 125.485 69.385 125.745 69.645 ;
        RECT 125.805 69.385 126.065 69.645 ;
        RECT 125.485 68.955 125.745 69.215 ;
        RECT 125.805 68.955 126.065 69.215 ;
        RECT 125.485 68.525 125.745 68.785 ;
        RECT 125.805 68.525 126.065 68.785 ;
        RECT 125.485 68.095 125.745 68.355 ;
        RECT 125.805 68.095 126.065 68.355 ;
        RECT 125.485 67.665 125.745 67.925 ;
        RECT 125.805 67.665 126.065 67.925 ;
        RECT 125.485 67.235 125.745 67.495 ;
        RECT 125.805 67.235 126.065 67.495 ;
        RECT 125.485 66.805 125.745 67.065 ;
        RECT 125.805 66.805 126.065 67.065 ;
        RECT 125.485 66.375 125.745 66.635 ;
        RECT 125.805 66.375 126.065 66.635 ;
        RECT 125.485 65.945 125.745 66.205 ;
        RECT 125.805 65.945 126.065 66.205 ;
        RECT 125.485 65.515 125.745 65.775 ;
        RECT 125.805 65.515 126.065 65.775 ;
        RECT 126.335 65.390 126.595 65.650 ;
        RECT 125.485 65.085 125.745 65.345 ;
        RECT 125.805 65.085 126.065 65.345 ;
        RECT 126.335 65.070 126.595 65.330 ;
        RECT 125.485 64.655 125.745 64.915 ;
        RECT 125.805 64.655 126.065 64.915 ;
        RECT 126.335 64.750 126.595 65.010 ;
        RECT 125.485 64.225 125.745 64.485 ;
        RECT 125.805 64.225 126.065 64.485 ;
        RECT 122.215 62.845 122.475 63.105 ;
        RECT 122.535 62.845 122.795 63.105 ;
        RECT 122.215 62.415 122.475 62.675 ;
        RECT 122.535 62.415 122.795 62.675 ;
        RECT 122.215 61.985 122.475 62.245 ;
        RECT 122.535 61.985 122.795 62.245 ;
        RECT 119.500 61.555 119.760 61.815 ;
        RECT 119.820 61.555 120.080 61.815 ;
        RECT 122.215 61.555 122.475 61.815 ;
        RECT 122.535 61.555 122.795 61.815 ;
        RECT 119.500 61.125 119.760 61.385 ;
        RECT 119.820 61.125 120.080 61.385 ;
        RECT 119.500 60.695 119.760 60.955 ;
        RECT 119.820 60.695 120.080 60.955 ;
        RECT 123.080 61.170 123.340 61.430 ;
        RECT 123.080 60.850 123.340 61.110 ;
        RECT 119.500 60.065 119.760 60.325 ;
        RECT 119.820 60.065 120.080 60.325 ;
        RECT 125.485 63.795 125.745 64.055 ;
        RECT 125.805 63.795 126.065 64.055 ;
        RECT 125.485 63.365 125.745 63.625 ;
        RECT 125.805 63.365 126.065 63.625 ;
        RECT 125.485 62.935 125.745 63.195 ;
        RECT 125.805 62.935 126.065 63.195 ;
        RECT 125.485 62.505 125.745 62.765 ;
        RECT 125.805 62.505 126.065 62.765 ;
        RECT 125.485 62.075 125.745 62.335 ;
        RECT 125.805 62.075 126.065 62.335 ;
        RECT 125.485 61.645 125.745 61.905 ;
        RECT 125.805 61.645 126.065 61.905 ;
        RECT 125.485 61.215 125.745 61.475 ;
        RECT 125.805 61.215 126.065 61.475 ;
        RECT 125.485 60.785 125.745 61.045 ;
        RECT 125.805 60.785 126.065 61.045 ;
        RECT 125.485 60.155 125.745 60.415 ;
        RECT 125.805 60.155 126.065 60.415 ;
      LAYER met2 ;
        RECT 127.375 211.950 144.155 212.280 ;
        RECT 115.355 211.120 158.265 211.450 ;
        RECT 120.335 210.290 147.830 210.620 ;
        RECT 157.665 210.370 158.265 211.120 ;
        RECT 123.680 209.190 157.165 209.790 ;
        RECT 156.565 209.110 157.165 209.190 ;
        RECT 117.715 208.090 142.530 208.690 ;
        RECT 106.100 206.195 118.065 206.795 ;
        RECT 117.695 205.715 118.065 206.195 ;
        RECT 84.950 174.075 85.250 174.645 ;
        RECT 45.995 173.475 85.250 174.075 ;
        RECT 108.195 173.590 109.195 173.880 ;
        RECT 112.045 173.590 113.045 173.880 ;
        RECT 45.995 15.130 46.595 173.475 ;
        RECT 88.630 172.975 88.930 173.545 ;
        RECT 47.095 172.375 88.930 172.975 ;
        RECT 108.195 172.925 109.195 173.205 ;
        RECT 108.195 172.495 109.195 172.775 ;
        RECT 110.205 172.425 110.535 173.195 ;
        RECT 112.045 172.925 113.045 173.205 ;
        RECT 112.045 172.495 113.045 172.775 ;
        RECT 47.095 16.230 47.695 172.375 ;
        RECT 108.195 172.065 109.195 172.345 ;
        RECT 112.045 172.065 113.045 172.345 ;
        RECT 108.195 171.635 113.545 171.915 ;
        RECT 108.195 171.205 109.195 171.485 ;
        RECT 110.205 171.055 110.535 171.635 ;
        RECT 112.045 171.205 113.045 171.485 ;
        RECT 108.195 170.775 113.545 171.055 ;
        RECT 108.195 170.345 109.195 170.625 ;
        RECT 110.205 170.420 110.535 170.775 ;
        RECT 108.195 169.915 109.195 170.195 ;
        RECT 108.195 169.485 109.195 169.765 ;
        RECT 110.195 169.540 110.535 170.420 ;
        RECT 112.045 170.345 113.045 170.625 ;
        RECT 112.045 169.915 113.045 170.195 ;
        RECT 108.195 168.810 109.195 169.100 ;
        RECT 110.195 167.355 110.525 169.540 ;
        RECT 112.045 169.485 113.045 169.765 ;
        RECT 112.045 168.810 113.045 169.100 ;
        RECT 116.785 167.355 117.115 167.775 ;
        RECT 110.195 167.025 117.115 167.355 ;
        RECT 116.785 166.605 117.115 167.025 ;
        RECT 109.605 164.440 110.305 164.730 ;
        RECT 110.975 164.440 111.675 164.730 ;
        RECT 112.345 164.440 113.045 164.730 ;
        RECT 122.810 164.400 123.510 164.690 ;
        RECT 109.605 163.775 110.305 164.055 ;
        RECT 110.975 163.775 111.675 164.055 ;
        RECT 112.345 163.775 113.045 164.055 ;
        RECT 122.810 163.775 123.510 164.055 ;
        RECT 109.605 161.495 110.305 161.775 ;
        RECT 110.975 161.495 111.675 161.775 ;
        RECT 112.345 161.495 113.045 161.775 ;
        RECT 122.810 161.495 123.510 161.775 ;
        RECT 123.680 159.495 124.010 166.330 ;
        RECT 124.180 164.400 124.880 164.690 ;
        RECT 124.180 163.775 124.880 164.055 ;
        RECT 124.180 161.495 124.880 161.775 ;
        RECT 109.605 159.215 110.305 159.495 ;
        RECT 110.975 159.215 111.675 159.495 ;
        RECT 112.345 159.215 113.045 159.495 ;
        RECT 122.810 159.215 124.880 159.495 ;
        RECT 109.605 156.935 113.045 157.215 ;
        RECT 122.810 156.935 123.510 157.215 ;
        RECT 109.605 154.655 110.305 154.935 ;
        RECT 78.045 153.950 106.700 154.550 ;
        RECT 78.045 152.850 106.700 153.450 ;
        RECT 106.100 152.370 106.700 152.850 ;
        RECT 110.475 152.655 110.805 156.935 ;
        RECT 110.975 154.655 111.675 154.935 ;
        RECT 111.845 152.655 112.175 156.935 ;
        RECT 123.680 154.935 124.010 159.215 ;
        RECT 124.180 156.935 124.880 157.215 ;
        RECT 112.345 154.655 113.045 154.935 ;
        RECT 122.810 154.655 124.880 154.935 ;
        RECT 109.605 152.375 113.045 152.655 ;
        RECT 122.810 152.375 123.510 152.655 ;
        RECT 63.150 151.680 71.640 151.960 ;
        RECT 57.150 151.190 58.150 151.480 ;
        RECT 60.740 151.190 61.740 151.480 ;
        RECT 65.405 151.190 65.905 151.480 ;
        RECT 60.740 150.525 61.740 150.805 ;
        RECT 65.405 150.525 65.905 150.805 ;
        RECT 71.310 150.790 71.640 151.680 ;
        RECT 87.150 151.680 95.640 151.960 ;
        RECT 87.150 150.790 87.480 151.680 ;
        RECT 92.885 151.190 93.385 151.480 ;
        RECT 97.050 151.190 98.050 151.480 ;
        RECT 100.640 151.190 101.640 151.480 ;
        RECT 92.885 150.525 93.385 150.805 ;
        RECT 97.050 150.525 98.050 150.805 ;
        RECT 109.605 150.095 110.305 150.375 ;
        RECT 60.740 149.745 61.740 150.025 ;
        RECT 65.405 149.745 65.905 150.025 ;
        RECT 92.885 149.745 93.385 150.025 ;
        RECT 97.050 149.745 98.050 150.025 ;
        RECT 60.740 148.965 61.740 149.245 ;
        RECT 63.170 148.800 63.500 149.680 ;
        RECT 65.405 148.965 65.905 149.245 ;
        RECT 92.885 148.965 93.385 149.245 ;
        RECT 61.930 148.510 63.500 148.800 ;
        RECT 95.290 148.800 95.620 149.680 ;
        RECT 97.050 148.965 98.050 149.245 ;
        RECT 95.290 148.510 96.860 148.800 ;
        RECT 61.930 147.900 62.260 148.510 ;
        RECT 96.530 147.900 96.860 148.510 ;
        RECT 110.475 148.095 110.805 152.375 ;
        RECT 110.975 150.095 111.675 150.375 ;
        RECT 111.845 148.095 112.175 152.375 ;
        RECT 123.680 150.375 124.010 154.655 ;
        RECT 124.180 152.375 124.880 152.655 ;
        RECT 112.345 150.095 113.045 150.375 ;
        RECT 122.810 150.095 124.880 150.375 ;
        RECT 109.605 147.815 113.045 148.095 ;
        RECT 122.810 147.815 123.510 148.095 ;
        RECT 64.885 146.965 65.215 147.275 ;
        RECT 93.575 146.965 93.905 147.275 ;
        RECT 60.740 146.685 63.435 146.965 ;
        RECT 63.765 146.685 65.215 146.965 ;
        RECT 65.405 146.685 72.465 146.965 ;
        RECT 63.765 145.795 64.095 146.685 ;
        RECT 64.885 146.375 65.215 146.685 ;
        RECT 72.135 145.795 72.465 146.685 ;
        RECT 86.325 146.685 93.385 146.965 ;
        RECT 93.575 146.685 95.025 146.965 ;
        RECT 95.355 146.685 98.050 146.965 ;
        RECT 86.325 145.795 86.655 146.685 ;
        RECT 93.575 146.375 93.905 146.685 ;
        RECT 94.695 145.795 95.025 146.685 ;
        RECT 109.605 145.535 110.305 145.815 ;
        RECT 60.740 144.405 61.740 144.685 ;
        RECT 65.405 144.405 65.905 144.685 ;
        RECT 92.885 144.405 93.385 144.685 ;
        RECT 97.050 144.405 98.050 144.685 ;
        RECT 60.740 143.625 61.740 143.905 ;
        RECT 65.405 143.625 65.905 143.905 ;
        RECT 92.885 143.625 93.385 143.905 ;
        RECT 97.050 143.625 98.050 143.905 ;
        RECT 110.475 143.535 110.805 147.815 ;
        RECT 110.975 145.535 111.675 145.815 ;
        RECT 111.845 143.535 112.175 147.815 ;
        RECT 123.680 145.815 124.010 150.095 ;
        RECT 124.180 147.815 124.880 148.095 ;
        RECT 112.345 145.535 113.045 145.815 ;
        RECT 122.810 145.535 124.880 145.815 ;
        RECT 109.605 143.255 113.045 143.535 ;
        RECT 122.810 143.255 123.510 143.535 ;
        RECT 60.740 142.845 61.740 143.125 ;
        RECT 65.405 142.845 65.905 143.125 ;
        RECT 92.885 142.845 93.385 143.125 ;
        RECT 97.050 142.845 98.050 143.125 ;
        RECT 73.560 142.470 74.060 142.760 ;
        RECT 76.300 142.470 76.800 142.760 ;
        RECT 81.990 142.470 82.490 142.760 ;
        RECT 84.730 142.470 85.230 142.760 ;
        RECT 60.740 142.065 61.740 142.345 ;
        RECT 65.405 142.170 65.905 142.460 ;
        RECT 92.885 142.170 93.385 142.460 ;
        RECT 73.560 141.845 74.060 142.125 ;
        RECT 57.150 141.285 58.150 141.565 ;
        RECT 59.255 141.285 61.740 141.565 ;
        RECT 76.300 141.445 76.800 141.725 ;
        RECT 57.150 139.005 58.150 139.285 ;
        RECT 59.255 137.005 59.585 141.285 ;
        RECT 78.045 141.120 78.645 141.895 ;
        RECT 61.930 140.790 78.645 141.120 ;
        RECT 80.145 141.120 80.745 141.895 ;
        RECT 84.730 141.845 85.230 142.125 ;
        RECT 97.050 142.065 98.050 142.345 ;
        RECT 81.990 141.445 82.490 141.725 ;
        RECT 97.050 141.285 99.535 141.565 ;
        RECT 100.640 141.285 101.640 141.565 ;
        RECT 80.145 140.790 96.860 141.120 ;
        RECT 61.930 140.220 62.260 140.790 ;
        RECT 73.040 140.540 73.370 140.790 ;
        RECT 85.420 140.540 85.750 140.790 ;
        RECT 96.530 140.220 96.860 140.790 ;
        RECT 75.035 139.565 75.405 139.765 ;
        RECT 73.560 139.285 75.405 139.565 ;
        RECT 60.740 139.005 63.435 139.285 ;
        RECT 75.035 139.085 75.405 139.285 ;
        RECT 83.385 139.565 83.755 139.765 ;
        RECT 83.385 139.285 85.230 139.565 ;
        RECT 83.385 139.085 83.755 139.285 ;
        RECT 95.355 139.005 98.050 139.285 ;
        RECT 65.405 137.980 65.905 138.270 ;
        RECT 69.160 137.980 70.160 138.270 ;
        RECT 76.300 138.165 76.800 138.445 ;
        RECT 81.990 138.165 82.490 138.445 ;
        RECT 88.630 137.980 89.630 138.270 ;
        RECT 92.885 137.980 93.385 138.270 ;
        RECT 65.405 137.315 65.905 137.595 ;
        RECT 69.160 137.315 70.160 137.595 ;
        RECT 88.630 137.315 89.630 137.595 ;
        RECT 92.885 137.315 93.385 137.595 ;
        RECT 72.135 137.005 74.060 137.285 ;
        RECT 84.730 137.005 86.655 137.285 ;
        RECT 99.205 137.005 99.535 141.285 ;
        RECT 109.605 140.975 110.305 141.255 ;
        RECT 100.640 139.005 101.640 139.285 ;
        RECT 110.475 138.975 110.805 143.255 ;
        RECT 110.975 140.975 111.675 141.255 ;
        RECT 111.845 138.975 112.175 143.255 ;
        RECT 123.680 141.255 124.010 145.535 ;
        RECT 124.180 143.255 124.880 143.535 ;
        RECT 112.345 140.975 113.045 141.255 ;
        RECT 122.810 140.975 124.880 141.255 ;
        RECT 109.605 138.695 113.045 138.975 ;
        RECT 122.810 138.695 123.510 138.975 ;
        RECT 57.150 136.725 58.150 137.005 ;
        RECT 59.255 136.725 61.740 137.005 ;
        RECT 57.150 134.445 58.150 134.725 ;
        RECT 59.255 132.445 59.585 136.725 ;
        RECT 65.405 136.035 65.905 136.315 ;
        RECT 69.160 136.035 70.160 136.315 ;
        RECT 65.405 134.755 65.905 135.035 ;
        RECT 69.160 134.755 70.160 135.035 ;
        RECT 60.740 134.445 65.215 134.725 ;
        RECT 64.885 133.825 65.215 134.445 ;
        RECT 66.095 134.280 66.425 134.590 ;
        RECT 66.095 134.000 68.010 134.280 ;
        RECT 66.095 133.690 66.425 134.000 ;
        RECT 67.680 133.110 68.010 134.000 ;
        RECT 72.135 132.725 72.465 137.005 ;
        RECT 75.035 135.005 75.405 135.205 ;
        RECT 73.560 134.725 75.405 135.005 ;
        RECT 76.300 134.885 76.800 135.165 ;
        RECT 81.990 134.885 82.490 135.165 ;
        RECT 83.385 135.005 83.755 135.205 ;
        RECT 75.035 134.525 75.405 134.725 ;
        RECT 83.385 134.725 85.230 135.005 ;
        RECT 83.385 134.525 83.755 134.725 ;
        RECT 86.325 132.725 86.655 137.005 ;
        RECT 97.050 136.725 99.535 137.005 ;
        RECT 100.640 136.725 101.640 137.005 ;
        RECT 88.630 136.035 89.630 136.315 ;
        RECT 92.885 136.035 93.385 136.315 ;
        RECT 88.630 134.755 89.630 135.035 ;
        RECT 92.885 134.755 93.385 135.035 ;
        RECT 92.365 134.280 92.695 134.590 ;
        RECT 90.780 134.000 92.695 134.280 ;
        RECT 90.780 133.110 91.110 134.000 ;
        RECT 92.365 133.690 92.695 134.000 ;
        RECT 93.575 134.445 98.050 134.725 ;
        RECT 93.575 133.825 93.905 134.445 ;
        RECT 69.160 132.445 74.060 132.725 ;
        RECT 84.730 132.445 89.630 132.725 ;
        RECT 99.205 132.445 99.535 136.725 ;
        RECT 123.680 136.695 124.010 140.975 ;
        RECT 124.180 138.695 124.880 138.975 ;
        RECT 109.605 136.415 110.305 136.695 ;
        RECT 110.975 136.415 111.675 136.695 ;
        RECT 112.345 136.415 113.045 136.695 ;
        RECT 122.810 136.415 124.880 136.695 ;
        RECT 100.640 134.445 101.640 134.725 ;
        RECT 109.605 134.135 114.615 134.415 ;
        RECT 122.810 134.135 123.510 134.415 ;
        RECT 57.150 132.165 58.150 132.445 ;
        RECT 59.255 132.165 61.740 132.445 ;
        RECT 97.050 132.165 99.535 132.445 ;
        RECT 100.640 132.165 101.640 132.445 ;
        RECT 57.150 129.885 58.150 130.165 ;
        RECT 56.100 127.910 56.430 128.750 ;
        RECT 56.630 127.910 56.960 128.195 ;
        RECT 56.100 127.580 56.960 127.910 ;
        RECT 59.255 127.885 59.585 132.165 ;
        RECT 67.000 131.230 67.330 132.120 ;
        RECT 68.640 131.230 68.970 131.540 ;
        RECT 67.000 130.950 68.970 131.230 ;
        RECT 68.640 130.640 68.970 130.950 ;
        RECT 89.820 131.230 90.150 131.540 ;
        RECT 91.460 131.230 91.790 132.120 ;
        RECT 89.820 130.950 91.790 131.230 ;
        RECT 65.405 130.195 65.905 130.475 ;
        RECT 69.160 130.195 70.160 130.475 ;
        RECT 75.035 130.445 75.405 130.645 ;
        RECT 73.560 130.165 75.405 130.445 ;
        RECT 60.740 129.885 63.435 130.165 ;
        RECT 75.035 129.965 75.405 130.165 ;
        RECT 83.385 130.445 83.755 130.645 ;
        RECT 89.820 130.640 90.150 130.950 ;
        RECT 83.385 130.165 85.230 130.445 ;
        RECT 88.630 130.195 89.630 130.475 ;
        RECT 92.885 130.195 93.385 130.475 ;
        RECT 83.385 129.965 83.755 130.165 ;
        RECT 95.355 129.885 98.050 130.165 ;
        RECT 65.405 128.915 65.905 129.195 ;
        RECT 69.160 128.915 70.160 129.195 ;
        RECT 73.560 128.885 74.060 129.165 ;
        RECT 84.730 128.885 85.230 129.165 ;
        RECT 88.630 128.915 89.630 129.195 ;
        RECT 92.885 128.915 93.385 129.195 ;
        RECT 57.150 127.605 61.740 127.885 ;
        RECT 65.405 127.635 65.905 127.915 ;
        RECT 69.160 127.635 70.160 127.915 ;
        RECT 75.055 127.885 75.385 128.330 ;
        RECT 83.405 127.885 83.735 128.330 ;
        RECT 73.560 127.605 74.060 127.885 ;
        RECT 75.055 127.605 76.800 127.885 ;
        RECT 81.990 127.605 83.735 127.885 ;
        RECT 84.730 127.605 85.230 127.885 ;
        RECT 88.630 127.635 89.630 127.915 ;
        RECT 92.885 127.635 93.385 127.915 ;
        RECT 99.205 127.885 99.535 132.165 ;
        RECT 109.605 131.855 110.305 132.135 ;
        RECT 110.975 131.855 111.675 132.135 ;
        RECT 112.345 131.855 113.045 132.135 ;
        RECT 100.640 129.885 101.640 130.165 ;
        RECT 114.285 129.855 114.615 134.135 ;
        RECT 123.680 132.135 124.010 136.415 ;
        RECT 124.180 134.135 124.880 134.415 ;
        RECT 122.810 131.855 124.880 132.135 ;
        RECT 109.605 129.575 114.615 129.855 ;
        RECT 122.810 129.575 123.510 129.855 ;
        RECT 101.830 127.910 102.160 128.195 ;
        RECT 102.360 127.910 102.690 128.750 ;
        RECT 97.050 127.605 101.640 127.885 ;
        RECT 56.630 127.295 56.960 127.580 ;
        RECT 57.150 125.325 58.150 125.605 ;
        RECT 59.255 123.325 59.585 127.605 ;
        RECT 75.055 127.160 75.385 127.605 ;
        RECT 83.405 127.160 83.735 127.605 ;
        RECT 76.990 126.685 77.320 126.795 ;
        RECT 81.470 126.685 81.800 126.795 ;
        RECT 65.405 126.355 65.905 126.635 ;
        RECT 69.160 126.355 70.160 126.635 ;
        RECT 73.560 126.325 74.060 126.605 ;
        RECT 76.990 125.685 77.830 126.685 ;
        RECT 80.960 125.685 81.800 126.685 ;
        RECT 84.730 126.325 85.230 126.605 ;
        RECT 88.630 126.355 89.630 126.635 ;
        RECT 92.885 126.355 93.385 126.635 ;
        RECT 60.740 125.325 63.435 125.605 ;
        RECT 76.990 125.575 77.320 125.685 ;
        RECT 81.470 125.575 81.800 125.685 ;
        RECT 65.405 125.075 65.905 125.355 ;
        RECT 69.160 125.075 70.160 125.355 ;
        RECT 75.035 125.325 75.405 125.525 ;
        RECT 73.560 125.045 75.405 125.325 ;
        RECT 75.035 124.845 75.405 125.045 ;
        RECT 83.385 125.325 83.755 125.525 ;
        RECT 83.385 125.045 85.230 125.325 ;
        RECT 88.630 125.075 89.630 125.355 ;
        RECT 92.885 125.075 93.385 125.355 ;
        RECT 95.355 125.325 98.050 125.605 ;
        RECT 83.385 124.845 83.755 125.045 ;
        RECT 57.150 123.045 58.150 123.325 ;
        RECT 59.255 123.045 61.740 123.325 ;
        RECT 63.085 123.075 63.415 123.520 ;
        RECT 63.765 123.075 64.095 123.965 ;
        RECT 64.880 123.075 65.210 123.385 ;
        RECT 93.580 123.075 93.910 123.385 ;
        RECT 94.695 123.075 95.025 123.965 ;
        RECT 95.375 123.075 95.705 123.520 ;
        RECT 99.205 123.325 99.535 127.605 ;
        RECT 101.830 127.580 102.690 127.910 ;
        RECT 101.830 127.295 102.160 127.580 ;
        RECT 109.605 127.295 110.305 127.575 ;
        RECT 110.975 127.295 111.675 127.575 ;
        RECT 112.345 127.295 113.045 127.575 ;
        RECT 100.640 125.325 101.640 125.605 ;
        RECT 114.285 125.295 114.615 129.575 ;
        RECT 123.680 127.575 124.010 131.855 ;
        RECT 124.180 129.575 124.880 129.855 ;
        RECT 122.810 127.295 124.880 127.575 ;
        RECT 109.605 125.015 114.615 125.295 ;
        RECT 122.810 125.015 123.510 125.295 ;
        RECT 124.180 125.015 124.880 125.295 ;
        RECT 57.150 120.765 58.150 121.045 ;
        RECT 59.255 118.765 59.585 123.045 ;
        RECT 63.085 122.795 65.905 123.075 ;
        RECT 63.085 122.350 63.415 122.795 ;
        RECT 64.880 122.485 65.210 122.795 ;
        RECT 69.160 122.765 74.060 123.045 ;
        RECT 84.730 122.765 89.630 123.045 ;
        RECT 92.885 122.795 95.705 123.075 ;
        RECT 97.050 123.045 99.535 123.325 ;
        RECT 100.640 123.045 101.640 123.325 ;
        RECT 60.740 120.765 63.435 121.045 ;
        RECT 65.405 120.515 65.905 120.795 ;
        RECT 69.160 120.515 70.160 120.795 ;
        RECT 65.405 119.235 65.905 119.515 ;
        RECT 69.160 119.235 70.160 119.515 ;
        RECT 57.150 118.485 58.150 118.765 ;
        RECT 59.255 118.485 61.740 118.765 ;
        RECT 71.310 118.485 71.640 122.765 ;
        RECT 75.035 120.765 75.405 120.965 ;
        RECT 73.560 120.485 75.405 120.765 ;
        RECT 83.385 120.765 83.755 120.965 ;
        RECT 75.035 120.285 75.405 120.485 ;
        RECT 76.300 120.325 76.800 120.605 ;
        RECT 81.990 120.325 82.490 120.605 ;
        RECT 83.385 120.485 85.230 120.765 ;
        RECT 83.385 120.285 83.755 120.485 ;
        RECT 87.150 118.485 87.480 122.765 ;
        RECT 93.580 122.485 93.910 122.795 ;
        RECT 95.375 122.350 95.705 122.795 ;
        RECT 88.630 120.515 89.630 120.795 ;
        RECT 92.885 120.515 93.385 120.795 ;
        RECT 95.355 120.765 98.050 121.045 ;
        RECT 88.630 119.235 89.630 119.515 ;
        RECT 92.885 119.235 93.385 119.515 ;
        RECT 99.205 118.765 99.535 123.045 ;
        RECT 109.605 122.735 110.305 123.015 ;
        RECT 110.975 122.735 111.675 123.015 ;
        RECT 112.345 122.735 113.045 123.015 ;
        RECT 100.640 120.765 101.640 121.045 ;
        RECT 114.285 120.735 114.615 125.015 ;
        RECT 109.605 120.455 114.615 120.735 ;
        RECT 97.050 118.485 99.535 118.765 ;
        RECT 100.640 118.485 101.640 118.765 ;
        RECT 57.150 116.205 58.150 116.485 ;
        RECT 59.255 114.205 59.585 118.485 ;
        RECT 65.405 117.955 65.905 118.235 ;
        RECT 69.160 117.955 70.160 118.235 ;
        RECT 71.310 118.205 74.060 118.485 ;
        RECT 84.730 118.205 87.480 118.485 ;
        RECT 88.630 117.955 89.630 118.235 ;
        RECT 92.885 117.955 93.385 118.235 ;
        RECT 65.405 117.280 65.905 117.570 ;
        RECT 69.160 117.280 70.160 117.570 ;
        RECT 76.300 117.045 76.800 117.325 ;
        RECT 81.990 117.045 82.490 117.325 ;
        RECT 88.630 117.280 89.630 117.570 ;
        RECT 92.885 117.280 93.385 117.570 ;
        RECT 60.740 116.205 63.435 116.485 ;
        RECT 75.035 116.205 75.405 116.405 ;
        RECT 73.560 115.925 75.405 116.205 ;
        RECT 75.035 115.725 75.405 115.925 ;
        RECT 83.385 116.205 83.755 116.405 ;
        RECT 95.355 116.205 98.050 116.485 ;
        RECT 83.385 115.925 85.230 116.205 ;
        RECT 83.385 115.725 83.755 115.925 ;
        RECT 61.930 114.700 62.260 115.270 ;
        RECT 73.040 114.700 73.370 114.950 ;
        RECT 85.420 114.700 85.750 114.950 ;
        RECT 96.530 114.700 96.860 115.270 ;
        RECT 61.930 114.370 96.860 114.700 ;
        RECT 99.205 114.205 99.535 118.485 ;
        RECT 109.605 118.175 110.305 118.455 ;
        RECT 110.975 118.175 111.675 118.455 ;
        RECT 112.345 118.175 113.045 118.455 ;
        RECT 100.640 116.205 101.640 116.485 ;
        RECT 114.285 116.210 114.615 120.455 ;
        RECT 121.785 122.735 124.880 123.015 ;
        RECT 121.785 118.455 122.065 122.735 ;
        RECT 122.810 120.455 123.510 120.735 ;
        RECT 124.180 120.455 124.880 120.735 ;
        RECT 121.785 118.175 124.880 118.455 ;
        RECT 115.375 116.410 115.705 117.180 ;
        RECT 115.895 116.360 118.045 116.640 ;
        RECT 114.285 116.175 116.595 116.210 ;
        RECT 109.605 115.930 116.595 116.175 ;
        RECT 109.605 115.895 114.615 115.930 ;
        RECT 57.150 113.925 58.150 114.205 ;
        RECT 59.255 113.925 61.740 114.205 ;
        RECT 76.300 113.765 76.800 114.045 ;
        RECT 81.990 113.765 82.490 114.045 ;
        RECT 97.050 113.925 99.535 114.205 ;
        RECT 100.640 113.925 101.640 114.205 ;
        RECT 60.740 113.145 61.740 113.425 ;
        RECT 73.560 113.365 74.060 113.645 ;
        RECT 84.730 113.365 85.230 113.645 ;
        RECT 109.605 113.615 110.305 113.895 ;
        RECT 110.975 113.615 111.675 113.895 ;
        RECT 112.345 113.615 113.045 113.895 ;
        RECT 64.315 113.030 65.315 113.320 ;
        RECT 69.115 113.030 69.615 113.320 ;
        RECT 89.175 113.030 89.675 113.320 ;
        RECT 93.475 113.030 94.475 113.320 ;
        RECT 97.050 113.145 98.050 113.425 ;
        RECT 73.560 112.730 74.060 113.020 ;
        RECT 76.300 112.730 76.800 113.020 ;
        RECT 81.990 112.730 82.490 113.020 ;
        RECT 84.730 112.730 85.230 113.020 ;
        RECT 60.740 112.365 61.740 112.645 ;
        RECT 64.315 112.365 65.315 112.645 ;
        RECT 69.115 112.365 69.615 112.645 ;
        RECT 89.175 112.365 89.675 112.645 ;
        RECT 93.475 112.365 94.475 112.645 ;
        RECT 97.050 112.365 98.050 112.645 ;
        RECT 57.150 111.690 58.150 111.980 ;
        RECT 60.740 111.690 61.740 111.980 ;
        RECT 97.050 111.690 98.050 111.980 ;
        RECT 100.640 111.690 101.640 111.980 ;
        RECT 114.285 111.615 114.615 115.895 ;
        RECT 117.715 115.780 118.045 116.360 ;
        RECT 115.895 115.500 118.045 115.780 ;
        RECT 117.715 114.255 118.045 115.500 ;
        RECT 117.715 113.975 120.165 114.255 ;
        RECT 117.715 113.395 118.045 113.975 ;
        RECT 117.715 113.115 120.165 113.395 ;
        RECT 117.715 111.970 118.045 113.115 ;
        RECT 120.355 113.105 120.685 114.275 ;
        RECT 121.785 113.895 122.065 118.175 ;
        RECT 122.810 115.895 123.510 116.175 ;
        RECT 124.180 115.895 124.880 116.175 ;
        RECT 121.785 113.615 124.880 113.895 ;
        RECT 115.895 111.690 118.045 111.970 ;
        RECT 109.605 111.540 114.615 111.615 ;
        RECT 109.605 111.335 116.595 111.540 ;
        RECT 114.285 111.260 116.595 111.335 ;
        RECT 64.315 110.085 65.315 110.365 ;
        RECT 69.115 110.085 69.615 110.365 ;
        RECT 89.175 110.085 89.675 110.365 ;
        RECT 93.475 110.085 94.475 110.365 ;
        RECT 109.605 109.055 110.305 109.335 ;
        RECT 110.975 109.055 111.675 109.335 ;
        RECT 112.345 109.055 113.045 109.335 ;
        RECT 64.315 107.805 65.315 108.085 ;
        RECT 69.115 107.805 69.615 108.085 ;
        RECT 89.175 107.805 89.675 108.085 ;
        RECT 93.475 107.805 94.475 108.085 ;
        RECT 65.505 107.330 65.835 107.640 ;
        RECT 67.000 107.330 67.330 107.775 ;
        RECT 65.505 107.050 67.330 107.330 ;
        RECT 65.505 106.740 65.835 107.050 ;
        RECT 67.000 106.605 67.330 107.050 ;
        RECT 67.680 107.330 68.010 107.775 ;
        RECT 68.595 107.330 68.925 107.640 ;
        RECT 67.680 107.050 68.925 107.330 ;
        RECT 67.680 106.605 68.010 107.050 ;
        RECT 68.595 106.740 68.925 107.050 ;
        RECT 89.865 107.330 90.195 107.640 ;
        RECT 90.780 107.330 91.110 107.775 ;
        RECT 89.865 107.050 91.110 107.330 ;
        RECT 89.865 106.740 90.195 107.050 ;
        RECT 90.780 106.605 91.110 107.050 ;
        RECT 91.460 107.330 91.790 107.775 ;
        RECT 92.955 107.330 93.285 107.640 ;
        RECT 91.460 107.050 93.285 107.330 ;
        RECT 114.285 107.055 114.615 111.260 ;
        RECT 117.715 111.110 118.045 111.690 ;
        RECT 115.895 110.830 118.045 111.110 ;
        RECT 116.785 109.860 117.115 110.630 ;
        RECT 91.460 106.605 91.790 107.050 ;
        RECT 92.955 106.740 93.285 107.050 ;
        RECT 109.605 106.775 114.615 107.055 ;
        RECT 64.315 105.525 69.615 105.805 ;
        RECT 89.175 105.525 94.475 105.805 ;
        RECT 109.605 104.495 110.305 104.775 ;
        RECT 110.975 104.495 111.675 104.775 ;
        RECT 112.345 104.495 113.045 104.775 ;
        RECT 64.315 103.245 65.315 103.525 ;
        RECT 69.115 103.245 69.615 103.525 ;
        RECT 89.175 103.245 89.675 103.525 ;
        RECT 93.475 103.245 94.475 103.525 ;
        RECT 114.285 102.495 114.615 106.775 ;
        RECT 109.605 102.215 114.615 102.495 ;
        RECT 64.315 100.965 69.615 101.245 ;
        RECT 89.175 100.965 94.475 101.245 ;
        RECT 109.605 99.935 110.305 100.215 ;
        RECT 110.975 99.935 111.675 100.215 ;
        RECT 112.345 99.935 113.045 100.215 ;
        RECT 114.285 99.840 114.615 102.215 ;
        RECT 121.785 109.335 122.065 113.615 ;
        RECT 122.810 111.335 123.510 111.615 ;
        RECT 124.180 111.335 124.880 111.615 ;
        RECT 121.785 109.055 124.880 109.335 ;
        RECT 121.785 104.775 122.065 109.055 ;
        RECT 122.810 106.775 123.510 107.055 ;
        RECT 124.180 106.775 124.880 107.055 ;
        RECT 121.785 104.495 124.880 104.775 ;
        RECT 121.785 100.215 122.065 104.495 ;
        RECT 122.810 102.215 123.510 102.495 ;
        RECT 124.180 102.215 124.880 102.495 ;
        RECT 121.785 99.935 124.880 100.215 ;
        RECT 111.845 99.145 112.175 99.505 ;
        RECT 121.785 99.145 122.065 99.935 ;
        RECT 64.315 98.685 65.315 98.965 ;
        RECT 69.115 98.685 69.615 98.965 ;
        RECT 89.175 98.685 89.675 98.965 ;
        RECT 93.475 98.685 94.475 98.965 ;
        RECT 111.845 98.645 122.065 99.145 ;
        RECT 111.845 98.285 112.175 98.645 ;
        RECT 109.605 97.655 114.615 97.935 ;
        RECT 64.315 96.405 69.615 96.685 ;
        RECT 89.175 96.405 94.475 96.685 ;
        RECT 109.605 95.375 110.305 95.655 ;
        RECT 110.975 95.375 111.675 95.655 ;
        RECT 112.345 95.375 113.045 95.655 ;
        RECT 64.315 94.125 65.315 94.405 ;
        RECT 69.115 94.125 69.615 94.405 ;
        RECT 89.175 94.125 89.675 94.405 ;
        RECT 93.475 94.125 94.475 94.405 ;
        RECT 114.285 93.375 114.615 97.655 ;
        RECT 109.605 93.095 114.615 93.375 ;
        RECT 121.785 95.655 122.065 98.645 ;
        RECT 122.810 97.655 123.510 97.935 ;
        RECT 124.180 97.655 124.880 97.935 ;
        RECT 121.785 95.375 124.880 95.655 ;
        RECT 64.315 91.845 65.315 92.125 ;
        RECT 69.115 91.845 69.615 92.125 ;
        RECT 89.175 91.845 89.675 92.125 ;
        RECT 93.475 91.845 94.475 92.125 ;
        RECT 121.785 91.095 122.065 95.375 ;
        RECT 122.810 93.095 123.510 93.375 ;
        RECT 124.180 93.095 124.880 93.375 ;
        RECT 109.605 90.815 110.305 91.095 ;
        RECT 110.975 90.815 111.675 91.095 ;
        RECT 112.345 90.815 113.045 91.095 ;
        RECT 121.785 90.815 124.880 91.095 ;
        RECT 64.315 89.565 65.315 89.845 ;
        RECT 69.115 89.565 69.615 89.845 ;
        RECT 89.175 89.565 89.675 89.845 ;
        RECT 93.475 89.565 94.475 89.845 ;
        RECT 64.315 88.890 65.315 89.180 ;
        RECT 69.115 88.890 69.615 89.180 ;
        RECT 89.175 88.890 89.675 89.180 ;
        RECT 93.475 88.890 94.475 89.180 ;
        RECT 109.605 88.535 114.615 88.815 ;
        RECT 122.810 88.535 123.510 88.815 ;
        RECT 124.180 88.535 124.880 88.815 ;
        RECT 79.165 86.240 104.670 86.840 ;
        RECT 109.605 86.255 110.305 86.535 ;
        RECT 110.975 86.255 111.675 86.535 ;
        RECT 112.345 86.255 113.045 86.535 ;
        RECT 104.070 85.760 104.670 86.240 ;
        RECT 83.780 84.705 88.005 85.035 ;
        RECT 74.410 83.575 87.435 83.905 ;
        RECT 71.925 82.995 78.995 83.275 ;
        RECT 79.565 82.995 86.635 83.275 ;
        RECT 71.925 82.105 72.255 82.995 ;
        RECT 72.595 82.360 73.445 82.650 ;
        RECT 75.820 82.360 76.670 82.650 ;
        RECT 77.395 82.360 78.245 82.650 ;
        RECT 78.585 82.105 78.915 82.995 ;
        RECT 79.645 82.105 79.975 82.995 ;
        RECT 80.315 82.360 81.165 82.650 ;
        RECT 81.890 82.360 82.740 82.650 ;
        RECT 85.115 82.360 85.965 82.650 ;
        RECT 86.305 82.105 86.635 82.995 ;
        RECT 72.595 81.695 73.445 81.975 ;
        RECT 72.595 81.265 73.445 81.545 ;
        RECT 71.905 80.205 72.275 80.885 ;
        RECT 72.595 80.835 73.445 81.115 ;
        RECT 74.430 81.035 74.760 81.895 ;
        RECT 75.820 81.695 76.670 81.975 ;
        RECT 77.395 81.695 78.245 81.975 ;
        RECT 80.315 81.695 81.165 81.975 ;
        RECT 81.890 81.695 82.740 81.975 ;
        RECT 75.820 81.265 76.670 81.545 ;
        RECT 77.395 81.265 78.245 81.545 ;
        RECT 80.315 81.265 81.165 81.545 ;
        RECT 81.890 81.265 82.740 81.545 ;
        RECT 75.745 80.835 77.215 81.115 ;
        RECT 77.395 80.835 78.245 81.115 ;
        RECT 76.925 80.685 77.215 80.835 ;
        RECT 72.445 80.405 76.745 80.685 ;
        RECT 76.925 80.405 78.395 80.685 ;
        RECT 72.595 79.975 73.445 80.255 ;
        RECT 74.430 79.825 74.760 80.405 ;
        RECT 76.925 80.255 77.215 80.405 ;
        RECT 75.745 79.975 77.215 80.255 ;
        RECT 77.395 79.975 78.245 80.255 ;
        RECT 76.925 79.825 77.215 79.975 ;
        RECT 72.445 79.545 76.745 79.825 ;
        RECT 76.925 79.545 78.395 79.825 ;
        RECT 72.595 79.115 73.445 79.395 ;
        RECT 72.595 78.685 73.445 78.965 ;
        RECT 72.595 78.255 73.445 78.535 ;
        RECT 72.595 77.580 73.445 77.885 ;
        RECT 74.430 77.435 74.760 79.545 ;
        RECT 76.925 79.395 77.215 79.545 ;
        RECT 75.745 79.115 77.215 79.395 ;
        RECT 77.395 79.115 78.245 79.395 ;
        RECT 78.585 79.390 78.915 80.840 ;
        RECT 79.645 79.390 79.975 80.840 ;
        RECT 80.315 80.835 81.165 81.115 ;
        RECT 81.345 80.835 82.815 81.115 ;
        RECT 83.800 81.035 84.130 81.895 ;
        RECT 85.115 81.695 85.965 81.975 ;
        RECT 85.115 81.265 85.965 81.545 ;
        RECT 85.115 80.835 85.965 81.115 ;
        RECT 81.345 80.685 81.635 80.835 ;
        RECT 80.165 80.405 81.635 80.685 ;
        RECT 81.815 80.405 86.115 80.685 ;
        RECT 81.345 80.255 81.635 80.405 ;
        RECT 80.315 79.975 81.165 80.255 ;
        RECT 81.345 79.975 82.815 80.255 ;
        RECT 81.345 79.825 81.635 79.975 ;
        RECT 83.800 79.825 84.130 80.405 ;
        RECT 85.115 79.975 85.965 80.255 ;
        RECT 86.285 80.205 86.655 80.885 ;
        RECT 80.165 79.545 81.635 79.825 ;
        RECT 81.815 79.545 86.115 79.825 ;
        RECT 81.345 79.395 81.635 79.545 ;
        RECT 80.315 79.115 81.165 79.395 ;
        RECT 81.345 79.115 82.815 79.395 ;
        RECT 75.820 78.685 76.670 78.965 ;
        RECT 77.395 78.685 78.245 78.965 ;
        RECT 80.315 78.685 81.165 78.965 ;
        RECT 81.890 78.685 82.740 78.965 ;
        RECT 75.820 78.255 76.670 78.535 ;
        RECT 77.395 78.255 78.245 78.535 ;
        RECT 80.315 78.255 81.165 78.535 ;
        RECT 81.890 78.255 82.740 78.535 ;
        RECT 75.820 77.580 76.670 77.885 ;
        RECT 77.395 77.580 78.245 77.885 ;
        RECT 80.315 77.580 81.165 77.885 ;
        RECT 81.890 77.580 82.740 77.885 ;
        RECT 83.800 77.435 84.130 79.545 ;
        RECT 85.115 79.115 85.965 79.395 ;
        RECT 85.115 78.685 85.965 78.965 ;
        RECT 85.115 78.255 85.965 78.535 ;
        RECT 85.115 77.580 85.965 77.885 ;
        RECT 87.085 77.435 87.415 78.275 ;
        RECT 74.430 77.105 79.995 77.435 ;
        RECT 83.800 77.105 87.415 77.435 ;
        RECT 76.360 75.430 76.690 77.105 ;
        RECT 87.675 76.990 88.005 84.705 ;
        RECT 114.285 84.255 114.615 88.535 ;
        RECT 122.810 86.255 123.510 86.535 ;
        RECT 124.180 86.255 124.880 86.535 ;
        RECT 109.605 83.975 114.615 84.255 ;
        RECT 122.810 83.975 123.510 84.255 ;
        RECT 124.180 83.975 124.880 84.255 ;
        RECT 89.110 82.710 90.110 83.000 ;
        RECT 92.960 82.710 93.960 83.000 ;
        RECT 89.110 82.045 90.110 82.325 ;
        RECT 89.110 81.615 90.110 81.895 ;
        RECT 91.120 81.545 91.450 82.315 ;
        RECT 92.960 82.045 93.960 82.325 ;
        RECT 114.285 82.010 114.615 83.975 ;
        RECT 122.330 83.110 122.620 83.450 ;
        RECT 123.680 83.110 124.010 83.420 ;
        RECT 115.375 82.210 115.705 82.980 ;
        RECT 122.330 82.830 124.010 83.110 ;
        RECT 122.330 82.490 122.620 82.830 ;
        RECT 123.680 82.520 124.010 82.830 ;
        RECT 115.895 82.160 118.045 82.440 ;
        RECT 92.960 81.615 93.960 81.895 ;
        RECT 109.605 81.695 110.305 81.975 ;
        RECT 110.975 81.695 111.675 81.975 ;
        RECT 112.345 81.695 113.045 81.975 ;
        RECT 114.285 81.730 116.595 82.010 ;
        RECT 89.110 81.185 90.110 81.465 ;
        RECT 92.960 81.185 93.960 81.465 ;
        RECT 89.110 80.755 94.460 81.035 ;
        RECT 89.110 80.325 90.110 80.605 ;
        RECT 91.120 80.175 91.450 80.755 ;
        RECT 92.960 80.325 93.960 80.605 ;
        RECT 89.110 79.895 94.460 80.175 ;
        RECT 89.110 79.465 90.110 79.745 ;
        RECT 89.110 79.035 90.110 79.315 ;
        RECT 89.110 78.605 90.110 78.885 ;
        RECT 89.110 77.930 90.110 78.220 ;
        RECT 91.120 76.990 91.450 79.895 ;
        RECT 92.960 79.465 93.960 79.745 ;
        RECT 114.285 79.695 114.615 81.730 ;
        RECT 117.715 81.580 118.045 82.160 ;
        RECT 115.895 81.300 118.045 81.580 ;
        RECT 109.605 79.415 114.615 79.695 ;
        RECT 92.960 79.035 93.960 79.315 ;
        RECT 92.960 78.605 93.960 78.885 ;
        RECT 92.960 77.930 93.960 78.220 ;
        RECT 109.605 77.135 110.305 77.415 ;
        RECT 110.975 77.135 111.675 77.415 ;
        RECT 112.345 77.135 113.045 77.415 ;
        RECT 114.285 77.340 114.615 79.415 ;
        RECT 117.715 80.055 118.045 81.300 ;
        RECT 121.155 81.695 123.510 81.975 ;
        RECT 124.180 81.695 124.880 81.975 ;
        RECT 121.155 80.805 121.485 81.695 ;
        RECT 117.715 79.775 120.165 80.055 ;
        RECT 117.715 79.195 118.045 79.775 ;
        RECT 117.715 78.915 120.165 79.195 ;
        RECT 117.715 77.770 118.045 78.915 ;
        RECT 120.355 78.905 120.685 80.075 ;
        RECT 122.810 79.415 123.510 79.695 ;
        RECT 124.180 79.415 124.880 79.695 ;
        RECT 115.895 77.490 118.045 77.770 ;
        RECT 87.675 76.660 91.450 76.990 ;
        RECT 114.285 77.060 116.595 77.340 ;
        RECT 91.120 74.845 95.795 75.175 ;
        RECT 114.285 75.135 114.615 77.060 ;
        RECT 117.715 76.910 118.045 77.490 ;
        RECT 122.810 77.135 123.510 77.415 ;
        RECT 124.180 77.135 124.880 77.415 ;
        RECT 115.895 76.630 118.045 76.910 ;
        RECT 122.810 76.500 123.510 76.790 ;
        RECT 124.180 76.500 124.880 76.790 ;
        RECT 116.785 75.660 117.115 76.430 ;
        RECT 109.605 74.855 114.615 75.135 ;
        RECT 115.745 75.095 116.445 75.385 ;
        RECT 91.120 74.005 91.450 74.845 ;
        RECT 109.605 72.575 110.305 72.855 ;
        RECT 110.975 72.575 111.675 72.855 ;
        RECT 112.345 72.575 113.045 72.855 ;
        RECT 65.330 72.050 66.330 72.340 ;
        RECT 69.180 72.050 70.180 72.340 ;
        RECT 74.350 72.050 75.350 72.340 ;
        RECT 78.200 72.050 79.200 72.340 ;
        RECT 81.290 72.050 82.290 72.340 ;
        RECT 85.140 72.050 86.140 72.340 ;
        RECT 89.110 72.050 90.110 72.340 ;
        RECT 92.960 72.050 93.960 72.340 ;
        RECT 65.330 71.385 66.330 71.665 ;
        RECT 65.330 70.955 66.330 71.235 ;
        RECT 67.340 70.885 67.670 71.655 ;
        RECT 69.180 71.385 70.180 71.665 ;
        RECT 74.350 71.385 75.350 71.665 ;
        RECT 69.180 70.955 70.180 71.235 ;
        RECT 74.350 70.955 75.350 71.235 ;
        RECT 76.360 70.885 76.690 71.655 ;
        RECT 78.200 71.385 79.200 71.665 ;
        RECT 81.290 71.385 82.290 71.665 ;
        RECT 78.200 70.955 79.200 71.235 ;
        RECT 81.290 70.955 82.290 71.235 ;
        RECT 83.800 70.885 84.130 71.655 ;
        RECT 85.140 71.385 86.140 71.665 ;
        RECT 89.110 71.385 90.110 71.665 ;
        RECT 85.140 70.955 86.140 71.235 ;
        RECT 89.110 70.955 90.110 71.235 ;
        RECT 91.120 70.885 91.450 71.655 ;
        RECT 92.960 71.385 93.960 71.665 ;
        RECT 92.960 70.955 93.960 71.235 ;
        RECT 65.330 70.525 66.330 70.805 ;
        RECT 69.180 70.525 70.180 70.805 ;
        RECT 74.350 70.525 75.350 70.805 ;
        RECT 78.200 70.525 79.200 70.805 ;
        RECT 81.290 70.525 82.290 70.805 ;
        RECT 85.140 70.525 86.140 70.805 ;
        RECT 89.110 70.525 90.110 70.805 ;
        RECT 92.960 70.525 93.960 70.805 ;
        RECT 114.285 70.575 114.615 74.855 ;
        RECT 120.330 70.950 124.290 71.280 ;
        RECT 65.330 70.095 70.680 70.375 ;
        RECT 74.350 70.095 79.700 70.375 ;
        RECT 80.790 70.095 86.140 70.375 ;
        RECT 89.110 70.095 94.460 70.375 ;
        RECT 109.605 70.295 114.615 70.575 ;
        RECT 115.745 70.320 116.445 70.610 ;
        RECT 65.330 69.665 66.330 69.945 ;
        RECT 67.340 69.515 67.670 70.095 ;
        RECT 69.180 69.665 70.180 69.945 ;
        RECT 74.350 69.665 75.350 69.945 ;
        RECT 76.360 69.515 76.690 70.095 ;
        RECT 78.200 69.665 79.200 69.945 ;
        RECT 81.290 69.665 82.290 69.945 ;
        RECT 83.800 69.515 84.130 70.095 ;
        RECT 85.140 69.665 86.140 69.945 ;
        RECT 89.110 69.665 90.110 69.945 ;
        RECT 91.120 69.515 91.450 70.095 ;
        RECT 119.440 70.040 120.140 70.330 ;
        RECT 92.960 69.665 93.960 69.945 ;
        RECT 65.330 69.235 70.680 69.515 ;
        RECT 74.350 69.235 79.700 69.515 ;
        RECT 80.790 69.235 86.140 69.515 ;
        RECT 89.110 69.235 94.460 69.515 ;
        RECT 111.845 69.440 112.175 69.750 ;
        RECT 115.745 69.655 116.445 69.935 ;
        RECT 111.845 69.160 115.555 69.440 ;
        RECT 119.440 69.375 120.140 69.655 ;
        RECT 65.330 68.805 66.330 69.085 ;
        RECT 69.180 68.805 70.180 69.085 ;
        RECT 74.350 68.805 75.350 69.085 ;
        RECT 78.200 68.805 79.200 69.085 ;
        RECT 81.290 68.805 82.290 69.085 ;
        RECT 85.140 68.805 86.140 69.085 ;
        RECT 89.110 68.805 90.110 69.085 ;
        RECT 92.960 68.805 93.960 69.085 ;
        RECT 111.845 68.850 112.175 69.160 ;
        RECT 65.330 68.375 70.680 68.655 ;
        RECT 74.350 68.375 79.700 68.655 ;
        RECT 80.790 68.375 86.140 68.655 ;
        RECT 89.110 68.375 94.460 68.655 ;
        RECT 115.225 68.540 115.555 69.160 ;
        RECT 119.440 68.945 120.140 69.225 ;
        RECT 120.330 69.150 120.660 70.950 ;
        RECT 123.960 70.110 124.290 70.950 ;
        RECT 125.425 70.000 126.125 70.290 ;
        RECT 117.715 68.515 120.140 68.795 ;
        RECT 121.155 68.515 122.855 68.795 ;
        RECT 123.045 68.770 123.375 69.805 ;
        RECT 125.425 69.375 126.125 69.655 ;
        RECT 125.425 68.945 126.125 69.225 ;
        RECT 125.425 68.515 126.125 68.795 ;
        RECT 65.330 67.945 66.330 68.225 ;
        RECT 67.340 67.795 67.670 68.375 ;
        RECT 69.180 67.945 70.180 68.225 ;
        RECT 74.350 67.945 75.350 68.225 ;
        RECT 76.360 67.795 76.690 68.375 ;
        RECT 78.200 67.945 79.200 68.225 ;
        RECT 81.290 67.945 82.290 68.225 ;
        RECT 83.800 67.795 84.130 68.375 ;
        RECT 85.140 67.945 86.140 68.225 ;
        RECT 89.110 67.945 90.110 68.225 ;
        RECT 91.120 67.795 91.450 68.375 ;
        RECT 92.960 67.945 93.960 68.225 ;
        RECT 109.605 68.015 110.305 68.295 ;
        RECT 110.975 68.015 111.675 68.295 ;
        RECT 112.345 68.015 113.045 68.295 ;
        RECT 117.715 67.935 118.045 68.515 ;
        RECT 119.440 68.365 120.140 68.370 ;
        RECT 119.440 68.085 124.290 68.365 ;
        RECT 125.425 68.085 126.125 68.365 ;
        RECT 65.330 67.515 70.680 67.795 ;
        RECT 74.350 67.515 79.700 67.795 ;
        RECT 80.790 67.515 86.140 67.795 ;
        RECT 89.110 67.515 94.460 67.795 ;
        RECT 117.715 67.655 120.140 67.935 ;
        RECT 121.155 67.655 122.855 67.935 ;
        RECT 65.330 67.085 66.330 67.365 ;
        RECT 67.340 66.935 67.670 67.515 ;
        RECT 69.180 67.085 70.180 67.365 ;
        RECT 74.350 67.085 75.350 67.365 ;
        RECT 76.360 66.935 76.690 67.515 ;
        RECT 78.200 67.085 79.200 67.365 ;
        RECT 81.290 67.085 82.290 67.365 ;
        RECT 83.800 66.935 84.130 67.515 ;
        RECT 85.140 67.085 86.140 67.365 ;
        RECT 89.110 67.085 90.110 67.365 ;
        RECT 91.120 66.935 91.450 67.515 ;
        RECT 115.745 67.375 116.445 67.655 ;
        RECT 92.960 67.085 93.960 67.365 ;
        RECT 117.715 67.075 118.045 67.655 ;
        RECT 119.440 67.505 120.140 67.510 ;
        RECT 123.960 67.505 124.290 68.085 ;
        RECT 125.425 67.655 126.125 67.935 ;
        RECT 119.440 67.225 124.290 67.505 ;
        RECT 125.425 67.225 126.125 67.505 ;
        RECT 65.330 66.655 70.680 66.935 ;
        RECT 74.350 66.655 79.700 66.935 ;
        RECT 80.790 66.655 86.140 66.935 ;
        RECT 89.110 66.655 94.460 66.935 ;
        RECT 117.715 66.795 120.140 67.075 ;
        RECT 121.155 66.795 122.855 67.075 ;
        RECT 65.330 66.225 66.330 66.505 ;
        RECT 67.340 66.075 67.670 66.655 ;
        RECT 69.180 66.225 70.180 66.505 ;
        RECT 74.350 66.225 75.350 66.505 ;
        RECT 76.360 66.075 76.690 66.655 ;
        RECT 78.200 66.225 79.200 66.505 ;
        RECT 81.290 66.225 82.290 66.505 ;
        RECT 83.800 66.075 84.130 66.655 ;
        RECT 85.140 66.225 86.140 66.505 ;
        RECT 89.110 66.225 90.110 66.505 ;
        RECT 91.120 66.075 91.450 66.655 ;
        RECT 92.960 66.225 93.960 66.505 ;
        RECT 65.330 65.795 70.680 66.075 ;
        RECT 74.350 65.795 79.700 66.075 ;
        RECT 80.790 65.795 86.140 66.075 ;
        RECT 89.110 65.795 94.460 66.075 ;
        RECT 65.330 65.365 66.330 65.645 ;
        RECT 67.340 65.215 67.670 65.795 ;
        RECT 69.180 65.365 70.180 65.645 ;
        RECT 74.350 65.365 75.350 65.645 ;
        RECT 76.360 65.215 76.690 65.795 ;
        RECT 78.200 65.365 79.200 65.645 ;
        RECT 81.290 65.365 82.290 65.645 ;
        RECT 83.800 65.215 84.130 65.795 ;
        RECT 85.140 65.365 86.140 65.645 ;
        RECT 89.110 65.365 90.110 65.645 ;
        RECT 91.120 65.215 91.450 65.795 ;
        RECT 109.605 65.735 110.305 66.015 ;
        RECT 110.975 65.735 111.675 66.015 ;
        RECT 112.345 65.735 113.045 66.015 ;
        RECT 92.960 65.365 93.960 65.645 ;
        RECT 117.715 65.375 118.045 66.795 ;
        RECT 119.440 66.365 120.140 66.645 ;
        RECT 119.440 65.935 120.140 66.215 ;
        RECT 65.330 64.935 70.680 65.215 ;
        RECT 74.350 64.935 79.700 65.215 ;
        RECT 80.790 64.935 86.140 65.215 ;
        RECT 89.110 64.935 94.460 65.215 ;
        RECT 115.745 65.095 118.045 65.375 ;
        RECT 65.330 64.505 66.330 64.785 ;
        RECT 65.330 64.075 66.330 64.355 ;
        RECT 65.330 63.645 66.330 63.925 ;
        RECT 67.340 63.700 67.670 64.935 ;
        RECT 69.180 64.505 70.180 64.785 ;
        RECT 74.350 64.505 75.350 64.785 ;
        RECT 69.180 64.075 70.180 64.355 ;
        RECT 74.350 64.075 75.350 64.355 ;
        RECT 69.180 63.645 70.180 63.925 ;
        RECT 74.350 63.645 75.350 63.925 ;
        RECT 76.360 63.700 76.690 64.935 ;
        RECT 78.200 64.505 79.200 64.785 ;
        RECT 81.290 64.505 82.290 64.785 ;
        RECT 78.200 64.075 79.200 64.355 ;
        RECT 81.290 64.075 82.290 64.355 ;
        RECT 78.200 63.645 79.200 63.925 ;
        RECT 81.290 63.645 82.290 63.925 ;
        RECT 83.800 63.700 84.130 64.935 ;
        RECT 85.140 64.505 86.140 64.785 ;
        RECT 89.110 64.505 90.110 64.785 ;
        RECT 85.140 64.075 86.140 64.355 ;
        RECT 89.110 64.075 90.110 64.355 ;
        RECT 85.140 63.645 86.140 63.925 ;
        RECT 89.110 63.645 90.110 63.925 ;
        RECT 91.120 63.700 91.450 64.935 ;
        RECT 92.960 64.505 93.960 64.785 ;
        RECT 92.960 64.075 93.960 64.355 ;
        RECT 92.960 63.645 93.960 63.925 ;
        RECT 109.605 63.455 110.305 63.735 ;
        RECT 110.975 63.455 111.675 63.735 ;
        RECT 112.345 63.455 113.045 63.735 ;
        RECT 117.715 63.545 118.045 65.095 ;
        RECT 123.960 65.785 124.290 67.225 ;
        RECT 125.425 66.795 126.125 67.075 ;
        RECT 125.425 66.365 126.125 66.645 ;
        RECT 125.425 65.935 126.125 66.215 ;
        RECT 123.960 65.505 126.125 65.785 ;
        RECT 123.960 64.925 124.290 65.505 ;
        RECT 124.640 64.925 125.240 65.505 ;
        RECT 126.305 65.365 126.625 65.650 ;
        RECT 127.395 65.365 127.725 65.785 ;
        RECT 125.425 65.075 126.125 65.355 ;
        RECT 126.305 65.035 127.725 65.365 ;
        RECT 123.960 64.645 126.125 64.925 ;
        RECT 126.305 64.750 126.625 65.035 ;
        RECT 119.440 64.125 120.140 64.405 ;
        RECT 119.440 63.695 120.140 63.975 ;
        RECT 117.715 63.265 120.140 63.545 ;
        RECT 120.440 63.375 120.770 64.465 ;
        RECT 121.155 63.265 122.855 63.545 ;
        RECT 65.330 62.970 66.330 63.260 ;
        RECT 69.180 62.970 70.180 63.260 ;
        RECT 74.350 62.970 75.350 63.260 ;
        RECT 78.200 62.970 79.200 63.260 ;
        RECT 81.290 62.970 82.290 63.260 ;
        RECT 85.140 62.970 86.140 63.260 ;
        RECT 89.110 62.970 90.110 63.260 ;
        RECT 92.960 62.970 93.960 63.260 ;
        RECT 109.605 62.780 110.305 63.070 ;
        RECT 110.975 62.780 111.675 63.070 ;
        RECT 112.345 62.780 113.045 63.070 ;
        RECT 115.745 62.815 116.445 63.095 ;
        RECT 117.715 62.685 118.045 63.265 ;
        RECT 119.440 63.115 120.140 63.120 ;
        RECT 123.960 63.115 124.290 64.645 ;
        RECT 119.440 62.835 124.290 63.115 ;
        RECT 117.715 62.405 120.140 62.685 ;
        RECT 121.155 62.405 122.855 62.685 ;
        RECT 117.715 61.825 118.045 62.405 ;
        RECT 119.440 62.255 120.140 62.260 ;
        RECT 123.960 62.255 124.290 62.835 ;
        RECT 119.440 61.975 124.290 62.255 ;
        RECT 117.715 61.545 120.140 61.825 ;
        RECT 121.135 61.545 122.855 61.825 ;
        RECT 119.440 61.115 120.140 61.395 ;
        RECT 123.045 61.305 123.375 61.430 ;
        RECT 123.940 61.305 124.310 61.480 ;
        RECT 123.045 60.975 124.310 61.305 ;
        RECT 115.745 60.535 116.445 60.815 ;
        RECT 119.440 60.685 120.140 60.965 ;
        RECT 123.045 60.850 123.375 60.975 ;
        RECT 123.940 60.800 124.310 60.975 ;
        RECT 115.745 59.860 116.445 60.150 ;
        RECT 119.440 60.050 120.140 60.340 ;
        RECT 120.420 59.150 123.395 59.480 ;
        RECT 124.640 55.265 125.240 64.645 ;
        RECT 127.395 64.615 127.725 65.035 ;
        RECT 125.425 64.215 126.125 64.495 ;
        RECT 125.425 63.785 126.125 64.065 ;
        RECT 125.425 63.355 126.125 63.635 ;
        RECT 125.425 62.925 126.125 63.205 ;
        RECT 125.425 62.495 126.125 62.775 ;
        RECT 125.425 62.065 126.125 62.345 ;
        RECT 125.425 61.635 126.125 61.915 ;
        RECT 125.425 61.205 126.125 61.485 ;
        RECT 125.425 60.775 126.125 61.055 ;
        RECT 125.425 60.140 126.125 60.430 ;
        RECT 124.640 38.195 142.530 38.795 ;
        RECT 104.070 21.205 104.670 21.710 ;
        RECT 124.640 21.205 125.240 21.445 ;
        RECT 72.280 20.055 72.610 20.895 ;
        RECT 104.070 20.605 125.240 21.205 ;
        RECT 124.640 20.365 125.240 20.605 ;
        RECT 72.280 19.725 124.290 20.055 ;
        RECT 87.515 18.895 123.375 19.225 ;
        RECT 123.960 18.885 124.290 19.725 ;
        RECT 105.170 17.795 118.045 18.395 ;
        RECT 90.985 16.230 91.585 16.710 ;
        RECT 47.095 15.630 91.585 16.230 ;
        RECT 45.995 14.530 84.265 15.130 ;
        RECT 117.715 12.595 142.530 13.195 ;
        RECT 76.225 7.250 113.000 7.850 ;
        RECT 67.205 6.150 90.920 6.750 ;
        RECT 157.665 4.430 158.265 5.310 ;
        RECT 134.480 3.830 158.265 4.430 ;
      LAYER via2 ;
        RECT 127.420 211.975 127.700 212.255 ;
        RECT 127.820 211.975 128.100 212.255 ;
        RECT 128.220 211.975 128.500 212.255 ;
        RECT 143.030 211.975 143.310 212.255 ;
        RECT 143.430 211.975 143.710 212.255 ;
        RECT 143.830 211.975 144.110 212.255 ;
        RECT 115.400 211.145 115.680 211.425 ;
        RECT 115.800 211.145 116.080 211.425 ;
        RECT 116.200 211.145 116.480 211.425 ;
        RECT 157.825 211.170 158.105 211.450 ;
        RECT 157.825 210.770 158.105 211.050 ;
        RECT 120.380 210.315 120.660 210.595 ;
        RECT 120.780 210.315 121.060 210.595 ;
        RECT 121.180 210.315 121.460 210.595 ;
        RECT 146.705 210.315 146.985 210.595 ;
        RECT 147.105 210.315 147.385 210.595 ;
        RECT 147.505 210.315 147.785 210.595 ;
        RECT 157.825 210.370 158.105 210.650 ;
        RECT 123.705 209.350 123.985 209.630 ;
        RECT 124.105 209.350 124.385 209.630 ;
        RECT 156.725 209.510 157.005 209.790 ;
        RECT 156.725 209.110 157.005 209.390 ;
        RECT 117.740 208.250 118.020 208.530 ;
        RECT 118.140 208.250 118.420 208.530 ;
        RECT 118.540 208.250 118.820 208.530 ;
        RECT 140.825 208.250 141.105 208.530 ;
        RECT 141.225 208.250 141.505 208.530 ;
        RECT 141.625 208.250 141.905 208.530 ;
        RECT 142.025 208.250 142.305 208.530 ;
        RECT 106.125 206.355 106.405 206.635 ;
        RECT 106.525 206.355 106.805 206.635 ;
        RECT 106.925 206.355 107.205 206.635 ;
        RECT 117.740 206.515 118.020 206.795 ;
        RECT 117.740 206.115 118.020 206.395 ;
        RECT 117.740 205.715 118.020 205.995 ;
        RECT 84.960 174.320 85.240 174.600 ;
        RECT 84.960 173.920 85.240 174.200 ;
        RECT 84.960 173.520 85.240 173.800 ;
        RECT 108.355 173.595 108.635 173.875 ;
        RECT 108.755 173.595 109.035 173.875 ;
        RECT 112.205 173.595 112.485 173.875 ;
        RECT 112.605 173.595 112.885 173.875 ;
        RECT 88.640 173.220 88.920 173.500 ;
        RECT 88.640 172.820 88.920 173.100 ;
        RECT 108.355 172.925 108.635 173.205 ;
        RECT 108.755 172.925 109.035 173.205 ;
        RECT 110.230 172.870 110.510 173.150 ;
        RECT 112.205 172.925 112.485 173.205 ;
        RECT 112.605 172.925 112.885 173.205 ;
        RECT 88.640 172.420 88.920 172.700 ;
        RECT 108.355 172.495 108.635 172.775 ;
        RECT 108.755 172.495 109.035 172.775 ;
        RECT 110.230 172.470 110.510 172.750 ;
        RECT 112.205 172.495 112.485 172.775 ;
        RECT 112.605 172.495 112.885 172.775 ;
        RECT 108.355 172.065 108.635 172.345 ;
        RECT 108.755 172.065 109.035 172.345 ;
        RECT 112.205 172.065 112.485 172.345 ;
        RECT 112.605 172.065 112.885 172.345 ;
        RECT 108.355 171.205 108.635 171.485 ;
        RECT 108.755 171.205 109.035 171.485 ;
        RECT 112.205 171.205 112.485 171.485 ;
        RECT 112.605 171.205 112.885 171.485 ;
        RECT 108.355 170.345 108.635 170.625 ;
        RECT 108.755 170.345 109.035 170.625 ;
        RECT 112.205 170.345 112.485 170.625 ;
        RECT 112.605 170.345 112.885 170.625 ;
        RECT 108.355 169.915 108.635 170.195 ;
        RECT 108.755 169.915 109.035 170.195 ;
        RECT 110.230 170.035 110.510 170.315 ;
        RECT 112.205 169.915 112.485 170.195 ;
        RECT 112.605 169.915 112.885 170.195 ;
        RECT 108.355 169.485 108.635 169.765 ;
        RECT 108.755 169.485 109.035 169.765 ;
        RECT 110.230 169.635 110.510 169.915 ;
        RECT 108.355 168.815 108.635 169.095 ;
        RECT 108.755 168.815 109.035 169.095 ;
        RECT 112.205 169.485 112.485 169.765 ;
        RECT 112.605 169.485 112.885 169.765 ;
        RECT 112.205 168.815 112.485 169.095 ;
        RECT 112.605 168.815 112.885 169.095 ;
        RECT 116.810 167.450 117.090 167.730 ;
        RECT 116.810 167.050 117.090 167.330 ;
        RECT 116.810 166.650 117.090 166.930 ;
        RECT 123.705 165.930 123.985 166.210 ;
        RECT 123.705 165.530 123.985 165.810 ;
        RECT 123.705 165.130 123.985 165.410 ;
        RECT 109.815 164.445 110.095 164.725 ;
        RECT 111.185 164.445 111.465 164.725 ;
        RECT 112.555 164.445 112.835 164.725 ;
        RECT 123.020 164.405 123.300 164.685 ;
        RECT 109.815 163.775 110.095 164.055 ;
        RECT 111.185 163.775 111.465 164.055 ;
        RECT 112.555 163.775 112.835 164.055 ;
        RECT 123.020 163.775 123.300 164.055 ;
        RECT 109.815 161.495 110.095 161.775 ;
        RECT 111.185 161.495 111.465 161.775 ;
        RECT 112.555 161.495 112.835 161.775 ;
        RECT 123.020 161.495 123.300 161.775 ;
        RECT 124.390 164.405 124.670 164.685 ;
        RECT 124.390 163.775 124.670 164.055 ;
        RECT 124.390 161.495 124.670 161.775 ;
        RECT 109.815 159.215 110.095 159.495 ;
        RECT 111.185 159.215 111.465 159.495 ;
        RECT 112.555 159.215 112.835 159.495 ;
        RECT 123.020 156.935 123.300 157.215 ;
        RECT 109.815 154.655 110.095 154.935 ;
        RECT 78.070 154.110 78.350 154.390 ;
        RECT 78.470 154.110 78.750 154.390 ;
        RECT 78.870 154.110 79.150 154.390 ;
        RECT 104.665 154.110 104.945 154.390 ;
        RECT 105.065 154.110 105.345 154.390 ;
        RECT 105.465 154.110 105.745 154.390 ;
        RECT 80.170 153.010 80.450 153.290 ;
        RECT 80.570 153.010 80.850 153.290 ;
        RECT 80.970 153.010 81.250 153.290 ;
        RECT 106.260 153.170 106.540 153.450 ;
        RECT 106.260 152.770 106.540 153.050 ;
        RECT 111.185 154.655 111.465 154.935 ;
        RECT 124.390 156.935 124.670 157.215 ;
        RECT 112.555 154.655 112.835 154.935 ;
        RECT 106.260 152.370 106.540 152.650 ;
        RECT 123.020 152.375 123.300 152.655 ;
        RECT 63.195 151.680 63.475 151.960 ;
        RECT 63.595 151.680 63.875 151.960 ;
        RECT 63.995 151.680 64.275 151.960 ;
        RECT 71.335 151.635 71.615 151.915 ;
        RECT 57.310 151.195 57.590 151.475 ;
        RECT 57.710 151.195 57.990 151.475 ;
        RECT 60.900 151.195 61.180 151.475 ;
        RECT 61.300 151.195 61.580 151.475 ;
        RECT 65.515 151.195 65.795 151.475 ;
        RECT 71.335 151.235 71.615 151.515 ;
        RECT 71.335 150.835 71.615 151.115 ;
        RECT 60.900 150.525 61.180 150.805 ;
        RECT 61.300 150.525 61.580 150.805 ;
        RECT 65.515 150.525 65.795 150.805 ;
        RECT 87.175 151.635 87.455 151.915 ;
        RECT 94.515 151.680 94.795 151.960 ;
        RECT 94.915 151.680 95.195 151.960 ;
        RECT 95.315 151.680 95.595 151.960 ;
        RECT 87.175 151.235 87.455 151.515 ;
        RECT 92.995 151.195 93.275 151.475 ;
        RECT 97.210 151.195 97.490 151.475 ;
        RECT 97.610 151.195 97.890 151.475 ;
        RECT 100.800 151.195 101.080 151.475 ;
        RECT 101.200 151.195 101.480 151.475 ;
        RECT 87.175 150.835 87.455 151.115 ;
        RECT 92.995 150.525 93.275 150.805 ;
        RECT 97.210 150.525 97.490 150.805 ;
        RECT 97.610 150.525 97.890 150.805 ;
        RECT 109.815 150.095 110.095 150.375 ;
        RECT 60.900 149.745 61.180 150.025 ;
        RECT 61.300 149.745 61.580 150.025 ;
        RECT 65.515 149.745 65.795 150.025 ;
        RECT 92.995 149.745 93.275 150.025 ;
        RECT 97.210 149.745 97.490 150.025 ;
        RECT 97.610 149.745 97.890 150.025 ;
        RECT 63.195 149.355 63.475 149.635 ;
        RECT 60.900 148.965 61.180 149.245 ;
        RECT 61.300 148.965 61.580 149.245 ;
        RECT 95.315 149.355 95.595 149.635 ;
        RECT 63.195 148.955 63.475 149.235 ;
        RECT 65.515 148.965 65.795 149.245 ;
        RECT 92.995 148.965 93.275 149.245 ;
        RECT 63.195 148.555 63.475 148.835 ;
        RECT 95.315 148.955 95.595 149.235 ;
        RECT 97.210 148.965 97.490 149.245 ;
        RECT 97.610 148.965 97.890 149.245 ;
        RECT 95.315 148.555 95.595 148.835 ;
        RECT 111.185 150.095 111.465 150.375 ;
        RECT 124.390 152.375 124.670 152.655 ;
        RECT 112.555 150.095 112.835 150.375 ;
        RECT 123.020 147.815 123.300 148.095 ;
        RECT 62.710 146.685 62.990 146.965 ;
        RECT 63.110 146.685 63.390 146.965 ;
        RECT 63.790 146.640 64.070 146.920 ;
        RECT 63.790 146.240 64.070 146.520 ;
        RECT 72.160 146.640 72.440 146.920 ;
        RECT 63.790 145.840 64.070 146.120 ;
        RECT 72.160 146.240 72.440 146.520 ;
        RECT 72.160 145.840 72.440 146.120 ;
        RECT 86.350 146.640 86.630 146.920 ;
        RECT 86.350 146.240 86.630 146.520 ;
        RECT 94.720 146.640 95.000 146.920 ;
        RECT 95.400 146.685 95.680 146.965 ;
        RECT 95.800 146.685 96.080 146.965 ;
        RECT 86.350 145.840 86.630 146.120 ;
        RECT 94.720 146.240 95.000 146.520 ;
        RECT 94.720 145.840 95.000 146.120 ;
        RECT 109.815 145.535 110.095 145.815 ;
        RECT 60.900 144.405 61.180 144.685 ;
        RECT 61.300 144.405 61.580 144.685 ;
        RECT 65.515 144.405 65.795 144.685 ;
        RECT 92.995 144.405 93.275 144.685 ;
        RECT 97.210 144.405 97.490 144.685 ;
        RECT 97.610 144.405 97.890 144.685 ;
        RECT 60.900 143.625 61.180 143.905 ;
        RECT 61.300 143.625 61.580 143.905 ;
        RECT 65.515 143.625 65.795 143.905 ;
        RECT 92.995 143.625 93.275 143.905 ;
        RECT 97.210 143.625 97.490 143.905 ;
        RECT 97.610 143.625 97.890 143.905 ;
        RECT 111.185 145.535 111.465 145.815 ;
        RECT 124.390 147.815 124.670 148.095 ;
        RECT 112.555 145.535 112.835 145.815 ;
        RECT 123.020 143.255 123.300 143.535 ;
        RECT 60.900 142.845 61.180 143.125 ;
        RECT 61.300 142.845 61.580 143.125 ;
        RECT 65.515 142.845 65.795 143.125 ;
        RECT 92.995 142.845 93.275 143.125 ;
        RECT 97.210 142.845 97.490 143.125 ;
        RECT 97.610 142.845 97.890 143.125 ;
        RECT 73.670 142.475 73.950 142.755 ;
        RECT 76.410 142.475 76.690 142.755 ;
        RECT 82.100 142.475 82.380 142.755 ;
        RECT 84.840 142.475 85.120 142.755 ;
        RECT 60.900 142.065 61.180 142.345 ;
        RECT 61.300 142.065 61.580 142.345 ;
        RECT 65.515 142.175 65.795 142.455 ;
        RECT 92.995 142.175 93.275 142.455 ;
        RECT 73.670 141.845 73.950 142.125 ;
        RECT 57.310 141.285 57.590 141.565 ;
        RECT 57.710 141.285 57.990 141.565 ;
        RECT 76.410 141.445 76.690 141.725 ;
        RECT 78.205 141.615 78.485 141.895 ;
        RECT 57.310 139.005 57.590 139.285 ;
        RECT 57.710 139.005 57.990 139.285 ;
        RECT 78.205 141.215 78.485 141.495 ;
        RECT 78.205 140.815 78.485 141.095 ;
        RECT 80.305 141.615 80.585 141.895 ;
        RECT 84.840 141.845 85.120 142.125 ;
        RECT 97.210 142.065 97.490 142.345 ;
        RECT 97.610 142.065 97.890 142.345 ;
        RECT 80.305 141.215 80.585 141.495 ;
        RECT 82.100 141.445 82.380 141.725 ;
        RECT 100.800 141.285 101.080 141.565 ;
        RECT 101.200 141.285 101.480 141.565 ;
        RECT 80.305 140.815 80.585 141.095 ;
        RECT 75.080 139.485 75.360 139.765 ;
        RECT 62.710 139.005 62.990 139.285 ;
        RECT 63.110 139.005 63.390 139.285 ;
        RECT 75.080 139.085 75.360 139.365 ;
        RECT 83.430 139.485 83.710 139.765 ;
        RECT 83.430 139.085 83.710 139.365 ;
        RECT 95.400 139.005 95.680 139.285 ;
        RECT 95.800 139.005 96.080 139.285 ;
        RECT 65.515 137.985 65.795 138.265 ;
        RECT 69.320 137.985 69.600 138.265 ;
        RECT 69.720 137.985 70.000 138.265 ;
        RECT 76.410 138.165 76.690 138.445 ;
        RECT 82.100 138.165 82.380 138.445 ;
        RECT 88.790 137.985 89.070 138.265 ;
        RECT 89.190 137.985 89.470 138.265 ;
        RECT 92.995 137.985 93.275 138.265 ;
        RECT 65.515 137.315 65.795 137.595 ;
        RECT 69.320 137.315 69.600 137.595 ;
        RECT 69.720 137.315 70.000 137.595 ;
        RECT 88.790 137.315 89.070 137.595 ;
        RECT 89.190 137.315 89.470 137.595 ;
        RECT 92.995 137.315 93.275 137.595 ;
        RECT 57.310 136.725 57.590 137.005 ;
        RECT 57.710 136.725 57.990 137.005 ;
        RECT 72.160 136.960 72.440 137.240 ;
        RECT 57.310 134.445 57.590 134.725 ;
        RECT 57.710 134.445 57.990 134.725 ;
        RECT 72.160 136.560 72.440 136.840 ;
        RECT 65.515 136.035 65.795 136.315 ;
        RECT 69.320 136.035 69.600 136.315 ;
        RECT 69.720 136.035 70.000 136.315 ;
        RECT 72.160 136.160 72.440 136.440 ;
        RECT 65.515 134.755 65.795 135.035 ;
        RECT 69.320 134.755 69.600 135.035 ;
        RECT 69.720 134.755 70.000 135.035 ;
        RECT 62.710 134.445 62.990 134.725 ;
        RECT 63.110 134.445 63.390 134.725 ;
        RECT 67.705 133.955 67.985 134.235 ;
        RECT 67.705 133.555 67.985 133.835 ;
        RECT 67.705 133.155 67.985 133.435 ;
        RECT 86.350 136.960 86.630 137.240 ;
        RECT 109.815 140.975 110.095 141.255 ;
        RECT 100.800 139.005 101.080 139.285 ;
        RECT 101.200 139.005 101.480 139.285 ;
        RECT 111.185 140.975 111.465 141.255 ;
        RECT 124.390 143.255 124.670 143.535 ;
        RECT 112.555 140.975 112.835 141.255 ;
        RECT 123.020 138.695 123.300 138.975 ;
        RECT 86.350 136.560 86.630 136.840 ;
        RECT 100.800 136.725 101.080 137.005 ;
        RECT 101.200 136.725 101.480 137.005 ;
        RECT 86.350 136.160 86.630 136.440 ;
        RECT 75.080 134.925 75.360 135.205 ;
        RECT 76.410 134.885 76.690 135.165 ;
        RECT 82.100 134.885 82.380 135.165 ;
        RECT 83.430 134.925 83.710 135.205 ;
        RECT 75.080 134.525 75.360 134.805 ;
        RECT 83.430 134.525 83.710 134.805 ;
        RECT 88.790 136.035 89.070 136.315 ;
        RECT 89.190 136.035 89.470 136.315 ;
        RECT 92.995 136.035 93.275 136.315 ;
        RECT 88.790 134.755 89.070 135.035 ;
        RECT 89.190 134.755 89.470 135.035 ;
        RECT 92.995 134.755 93.275 135.035 ;
        RECT 90.805 133.955 91.085 134.235 ;
        RECT 90.805 133.555 91.085 133.835 ;
        RECT 95.400 134.445 95.680 134.725 ;
        RECT 95.800 134.445 96.080 134.725 ;
        RECT 90.805 133.155 91.085 133.435 ;
        RECT 124.390 138.695 124.670 138.975 ;
        RECT 109.815 136.415 110.095 136.695 ;
        RECT 111.185 136.415 111.465 136.695 ;
        RECT 112.555 136.415 112.835 136.695 ;
        RECT 100.800 134.445 101.080 134.725 ;
        RECT 101.200 134.445 101.480 134.725 ;
        RECT 123.020 134.135 123.300 134.415 ;
        RECT 57.310 132.165 57.590 132.445 ;
        RECT 57.710 132.165 57.990 132.445 ;
        RECT 100.800 132.165 101.080 132.445 ;
        RECT 101.200 132.165 101.480 132.445 ;
        RECT 57.310 129.885 57.590 130.165 ;
        RECT 57.710 129.885 57.990 130.165 ;
        RECT 56.125 128.425 56.405 128.705 ;
        RECT 56.125 128.025 56.405 128.305 ;
        RECT 56.125 127.625 56.405 127.905 ;
        RECT 67.025 131.795 67.305 132.075 ;
        RECT 67.025 131.395 67.305 131.675 ;
        RECT 91.485 131.795 91.765 132.075 ;
        RECT 67.025 130.995 67.305 131.275 ;
        RECT 91.485 131.395 91.765 131.675 ;
        RECT 91.485 130.995 91.765 131.275 ;
        RECT 65.515 130.195 65.795 130.475 ;
        RECT 69.320 130.195 69.600 130.475 ;
        RECT 69.720 130.195 70.000 130.475 ;
        RECT 75.080 130.365 75.360 130.645 ;
        RECT 62.710 129.885 62.990 130.165 ;
        RECT 63.110 129.885 63.390 130.165 ;
        RECT 75.080 129.965 75.360 130.245 ;
        RECT 83.430 130.365 83.710 130.645 ;
        RECT 83.430 129.965 83.710 130.245 ;
        RECT 88.790 130.195 89.070 130.475 ;
        RECT 89.190 130.195 89.470 130.475 ;
        RECT 92.995 130.195 93.275 130.475 ;
        RECT 95.400 129.885 95.680 130.165 ;
        RECT 95.800 129.885 96.080 130.165 ;
        RECT 65.515 128.915 65.795 129.195 ;
        RECT 69.320 128.915 69.600 129.195 ;
        RECT 69.720 128.915 70.000 129.195 ;
        RECT 73.670 128.885 73.950 129.165 ;
        RECT 84.840 128.885 85.120 129.165 ;
        RECT 88.790 128.915 89.070 129.195 ;
        RECT 89.190 128.915 89.470 129.195 ;
        RECT 92.995 128.915 93.275 129.195 ;
        RECT 75.080 128.005 75.360 128.285 ;
        RECT 65.515 127.635 65.795 127.915 ;
        RECT 69.320 127.635 69.600 127.915 ;
        RECT 69.720 127.635 70.000 127.915 ;
        RECT 83.430 128.005 83.710 128.285 ;
        RECT 73.670 127.605 73.950 127.885 ;
        RECT 75.080 127.605 75.360 127.885 ;
        RECT 83.430 127.605 83.710 127.885 ;
        RECT 84.840 127.605 85.120 127.885 ;
        RECT 88.790 127.635 89.070 127.915 ;
        RECT 89.190 127.635 89.470 127.915 ;
        RECT 92.995 127.635 93.275 127.915 ;
        RECT 109.815 131.855 110.095 132.135 ;
        RECT 111.185 131.855 111.465 132.135 ;
        RECT 112.555 131.855 112.835 132.135 ;
        RECT 100.800 129.885 101.080 130.165 ;
        RECT 101.200 129.885 101.480 130.165 ;
        RECT 124.390 134.135 124.670 134.415 ;
        RECT 123.020 129.575 123.300 129.855 ;
        RECT 102.385 128.425 102.665 128.705 ;
        RECT 102.385 128.025 102.665 128.305 ;
        RECT 102.385 127.625 102.665 127.905 ;
        RECT 57.310 125.325 57.590 125.605 ;
        RECT 57.710 125.325 57.990 125.605 ;
        RECT 75.080 127.205 75.360 127.485 ;
        RECT 83.430 127.205 83.710 127.485 ;
        RECT 65.515 126.355 65.795 126.635 ;
        RECT 69.320 126.355 69.600 126.635 ;
        RECT 69.720 126.355 70.000 126.635 ;
        RECT 73.670 126.325 73.950 126.605 ;
        RECT 77.510 126.245 77.790 126.525 ;
        RECT 77.510 125.845 77.790 126.125 ;
        RECT 81.000 126.245 81.280 126.525 ;
        RECT 84.840 126.325 85.120 126.605 ;
        RECT 88.790 126.355 89.070 126.635 ;
        RECT 89.190 126.355 89.470 126.635 ;
        RECT 92.995 126.355 93.275 126.635 ;
        RECT 81.000 125.845 81.280 126.125 ;
        RECT 62.710 125.325 62.990 125.605 ;
        RECT 63.110 125.325 63.390 125.605 ;
        RECT 65.515 125.075 65.795 125.355 ;
        RECT 69.320 125.075 69.600 125.355 ;
        RECT 69.720 125.075 70.000 125.355 ;
        RECT 75.080 125.245 75.360 125.525 ;
        RECT 75.080 124.845 75.360 125.125 ;
        RECT 83.430 125.245 83.710 125.525 ;
        RECT 83.430 124.845 83.710 125.125 ;
        RECT 88.790 125.075 89.070 125.355 ;
        RECT 89.190 125.075 89.470 125.355 ;
        RECT 92.995 125.075 93.275 125.355 ;
        RECT 95.400 125.325 95.680 125.605 ;
        RECT 95.800 125.325 96.080 125.605 ;
        RECT 63.790 123.640 64.070 123.920 ;
        RECT 57.310 123.045 57.590 123.325 ;
        RECT 57.710 123.045 57.990 123.325 ;
        RECT 63.110 123.195 63.390 123.475 ;
        RECT 63.790 123.240 64.070 123.520 ;
        RECT 94.720 123.640 95.000 123.920 ;
        RECT 57.310 120.765 57.590 121.045 ;
        RECT 57.710 120.765 57.990 121.045 ;
        RECT 63.110 122.795 63.390 123.075 ;
        RECT 63.790 122.840 64.070 123.120 ;
        RECT 94.720 123.240 95.000 123.520 ;
        RECT 63.110 122.395 63.390 122.675 ;
        RECT 71.335 122.640 71.615 122.920 ;
        RECT 71.335 122.240 71.615 122.520 ;
        RECT 71.335 121.840 71.615 122.120 ;
        RECT 71.335 121.440 71.615 121.720 ;
        RECT 62.710 120.765 62.990 121.045 ;
        RECT 63.110 120.765 63.390 121.045 ;
        RECT 65.515 120.515 65.795 120.795 ;
        RECT 69.320 120.515 69.600 120.795 ;
        RECT 69.720 120.515 70.000 120.795 ;
        RECT 65.515 119.235 65.795 119.515 ;
        RECT 69.320 119.235 69.600 119.515 ;
        RECT 69.720 119.235 70.000 119.515 ;
        RECT 57.310 118.485 57.590 118.765 ;
        RECT 57.710 118.485 57.990 118.765 ;
        RECT 87.175 122.640 87.455 122.920 ;
        RECT 94.720 122.840 95.000 123.120 ;
        RECT 95.400 123.195 95.680 123.475 ;
        RECT 109.815 127.295 110.095 127.575 ;
        RECT 111.185 127.295 111.465 127.575 ;
        RECT 112.555 127.295 112.835 127.575 ;
        RECT 100.800 125.325 101.080 125.605 ;
        RECT 101.200 125.325 101.480 125.605 ;
        RECT 124.390 129.575 124.670 129.855 ;
        RECT 123.020 125.015 123.300 125.295 ;
        RECT 124.390 125.015 124.670 125.295 ;
        RECT 95.400 122.795 95.680 123.075 ;
        RECT 100.800 123.045 101.080 123.325 ;
        RECT 101.200 123.045 101.480 123.325 ;
        RECT 87.175 122.240 87.455 122.520 ;
        RECT 95.400 122.395 95.680 122.675 ;
        RECT 87.175 121.840 87.455 122.120 ;
        RECT 87.175 121.440 87.455 121.720 ;
        RECT 75.080 120.685 75.360 120.965 ;
        RECT 83.430 120.685 83.710 120.965 ;
        RECT 75.080 120.285 75.360 120.565 ;
        RECT 76.410 120.325 76.690 120.605 ;
        RECT 82.100 120.325 82.380 120.605 ;
        RECT 83.430 120.285 83.710 120.565 ;
        RECT 88.790 120.515 89.070 120.795 ;
        RECT 89.190 120.515 89.470 120.795 ;
        RECT 92.995 120.515 93.275 120.795 ;
        RECT 95.400 120.765 95.680 121.045 ;
        RECT 95.800 120.765 96.080 121.045 ;
        RECT 88.790 119.235 89.070 119.515 ;
        RECT 89.190 119.235 89.470 119.515 ;
        RECT 92.995 119.235 93.275 119.515 ;
        RECT 109.815 122.735 110.095 123.015 ;
        RECT 111.185 122.735 111.465 123.015 ;
        RECT 112.555 122.735 112.835 123.015 ;
        RECT 100.800 120.765 101.080 121.045 ;
        RECT 101.200 120.765 101.480 121.045 ;
        RECT 100.800 118.485 101.080 118.765 ;
        RECT 101.200 118.485 101.480 118.765 ;
        RECT 57.310 116.205 57.590 116.485 ;
        RECT 57.710 116.205 57.990 116.485 ;
        RECT 65.515 117.955 65.795 118.235 ;
        RECT 69.320 117.955 69.600 118.235 ;
        RECT 69.720 117.955 70.000 118.235 ;
        RECT 88.790 117.955 89.070 118.235 ;
        RECT 89.190 117.955 89.470 118.235 ;
        RECT 92.995 117.955 93.275 118.235 ;
        RECT 65.515 117.285 65.795 117.565 ;
        RECT 69.320 117.285 69.600 117.565 ;
        RECT 69.720 117.285 70.000 117.565 ;
        RECT 76.410 117.045 76.690 117.325 ;
        RECT 82.100 117.045 82.380 117.325 ;
        RECT 88.790 117.285 89.070 117.565 ;
        RECT 89.190 117.285 89.470 117.565 ;
        RECT 92.995 117.285 93.275 117.565 ;
        RECT 62.710 116.205 62.990 116.485 ;
        RECT 63.110 116.205 63.390 116.485 ;
        RECT 75.080 116.125 75.360 116.405 ;
        RECT 75.080 115.725 75.360 116.005 ;
        RECT 83.430 116.125 83.710 116.405 ;
        RECT 95.400 116.205 95.680 116.485 ;
        RECT 95.800 116.205 96.080 116.485 ;
        RECT 83.430 115.725 83.710 116.005 ;
        RECT 78.925 114.395 79.205 114.675 ;
        RECT 79.325 114.395 79.605 114.675 ;
        RECT 79.725 114.395 80.005 114.675 ;
        RECT 109.815 118.175 110.095 118.455 ;
        RECT 111.185 118.175 111.465 118.455 ;
        RECT 112.555 118.175 112.835 118.455 ;
        RECT 100.800 116.205 101.080 116.485 ;
        RECT 101.200 116.205 101.480 116.485 ;
        RECT 123.020 120.455 123.300 120.735 ;
        RECT 124.390 120.455 124.670 120.735 ;
        RECT 115.400 116.855 115.680 117.135 ;
        RECT 115.400 116.455 115.680 116.735 ;
        RECT 117.740 116.195 118.020 116.475 ;
        RECT 57.310 113.925 57.590 114.205 ;
        RECT 57.710 113.925 57.990 114.205 ;
        RECT 76.410 113.765 76.690 114.045 ;
        RECT 82.100 113.765 82.380 114.045 ;
        RECT 100.800 113.925 101.080 114.205 ;
        RECT 101.200 113.925 101.480 114.205 ;
        RECT 60.900 113.145 61.180 113.425 ;
        RECT 61.300 113.145 61.580 113.425 ;
        RECT 73.670 113.365 73.950 113.645 ;
        RECT 84.840 113.365 85.120 113.645 ;
        RECT 109.815 113.615 110.095 113.895 ;
        RECT 111.185 113.615 111.465 113.895 ;
        RECT 112.555 113.615 112.835 113.895 ;
        RECT 64.475 113.035 64.755 113.315 ;
        RECT 64.875 113.035 65.155 113.315 ;
        RECT 69.225 113.035 69.505 113.315 ;
        RECT 89.285 113.035 89.565 113.315 ;
        RECT 93.635 113.035 93.915 113.315 ;
        RECT 94.035 113.035 94.315 113.315 ;
        RECT 97.210 113.145 97.490 113.425 ;
        RECT 97.610 113.145 97.890 113.425 ;
        RECT 73.670 112.735 73.950 113.015 ;
        RECT 76.410 112.735 76.690 113.015 ;
        RECT 82.100 112.735 82.380 113.015 ;
        RECT 84.840 112.735 85.120 113.015 ;
        RECT 60.900 112.365 61.180 112.645 ;
        RECT 61.300 112.365 61.580 112.645 ;
        RECT 64.475 112.365 64.755 112.645 ;
        RECT 64.875 112.365 65.155 112.645 ;
        RECT 69.225 112.365 69.505 112.645 ;
        RECT 89.285 112.365 89.565 112.645 ;
        RECT 93.635 112.365 93.915 112.645 ;
        RECT 94.035 112.365 94.315 112.645 ;
        RECT 97.210 112.365 97.490 112.645 ;
        RECT 97.610 112.365 97.890 112.645 ;
        RECT 57.310 111.695 57.590 111.975 ;
        RECT 57.710 111.695 57.990 111.975 ;
        RECT 60.900 111.695 61.180 111.975 ;
        RECT 61.300 111.695 61.580 111.975 ;
        RECT 97.210 111.695 97.490 111.975 ;
        RECT 97.610 111.695 97.890 111.975 ;
        RECT 100.800 111.695 101.080 111.975 ;
        RECT 101.200 111.695 101.480 111.975 ;
        RECT 117.740 115.795 118.020 116.075 ;
        RECT 117.740 115.395 118.020 115.675 ;
        RECT 117.740 114.995 118.020 115.275 ;
        RECT 117.740 114.595 118.020 114.875 ;
        RECT 117.740 114.195 118.020 114.475 ;
        RECT 117.740 113.795 118.020 114.075 ;
        RECT 117.740 113.395 118.020 113.675 ;
        RECT 120.380 113.950 120.660 114.230 ;
        RECT 120.380 113.550 120.660 113.830 ;
        RECT 117.740 112.995 118.020 113.275 ;
        RECT 120.380 113.150 120.660 113.430 ;
        RECT 123.020 115.895 123.300 116.175 ;
        RECT 124.390 115.895 124.670 116.175 ;
        RECT 117.740 112.595 118.020 112.875 ;
        RECT 117.740 112.195 118.020 112.475 ;
        RECT 117.740 111.795 118.020 112.075 ;
        RECT 117.740 111.395 118.020 111.675 ;
        RECT 64.475 110.085 64.755 110.365 ;
        RECT 64.875 110.085 65.155 110.365 ;
        RECT 69.225 110.085 69.505 110.365 ;
        RECT 89.285 110.085 89.565 110.365 ;
        RECT 93.635 110.085 93.915 110.365 ;
        RECT 94.035 110.085 94.315 110.365 ;
        RECT 109.815 109.055 110.095 109.335 ;
        RECT 111.185 109.055 111.465 109.335 ;
        RECT 112.555 109.055 112.835 109.335 ;
        RECT 64.475 107.805 64.755 108.085 ;
        RECT 64.875 107.805 65.155 108.085 ;
        RECT 69.225 107.805 69.505 108.085 ;
        RECT 89.285 107.805 89.565 108.085 ;
        RECT 93.635 107.805 93.915 108.085 ;
        RECT 94.035 107.805 94.315 108.085 ;
        RECT 67.025 107.450 67.305 107.730 ;
        RECT 67.025 107.050 67.305 107.330 ;
        RECT 67.025 106.650 67.305 106.930 ;
        RECT 67.705 107.450 67.985 107.730 ;
        RECT 67.705 107.050 67.985 107.330 ;
        RECT 67.705 106.650 67.985 106.930 ;
        RECT 90.805 107.450 91.085 107.730 ;
        RECT 90.805 107.050 91.085 107.330 ;
        RECT 90.805 106.650 91.085 106.930 ;
        RECT 91.485 107.450 91.765 107.730 ;
        RECT 91.485 107.050 91.765 107.330 ;
        RECT 117.740 110.995 118.020 111.275 ;
        RECT 116.810 110.305 117.090 110.585 ;
        RECT 116.810 109.905 117.090 110.185 ;
        RECT 91.485 106.650 91.765 106.930 ;
        RECT 109.815 104.495 110.095 104.775 ;
        RECT 111.185 104.495 111.465 104.775 ;
        RECT 112.555 104.495 112.835 104.775 ;
        RECT 64.475 103.245 64.755 103.525 ;
        RECT 64.875 103.245 65.155 103.525 ;
        RECT 69.225 103.245 69.505 103.525 ;
        RECT 89.285 103.245 89.565 103.525 ;
        RECT 93.635 103.245 93.915 103.525 ;
        RECT 94.035 103.245 94.315 103.525 ;
        RECT 114.310 100.695 114.590 100.975 ;
        RECT 114.310 100.295 114.590 100.575 ;
        RECT 109.815 99.935 110.095 100.215 ;
        RECT 111.185 99.935 111.465 100.215 ;
        RECT 112.555 99.935 112.835 100.215 ;
        RECT 114.310 99.895 114.590 100.175 ;
        RECT 123.020 111.335 123.300 111.615 ;
        RECT 124.390 111.335 124.670 111.615 ;
        RECT 123.020 106.775 123.300 107.055 ;
        RECT 124.390 106.775 124.670 107.055 ;
        RECT 123.020 102.215 123.300 102.495 ;
        RECT 124.390 102.215 124.670 102.495 ;
        RECT 64.475 98.685 64.755 98.965 ;
        RECT 64.875 98.685 65.155 98.965 ;
        RECT 69.225 98.685 69.505 98.965 ;
        RECT 89.285 98.685 89.565 98.965 ;
        RECT 93.635 98.685 93.915 98.965 ;
        RECT 94.035 98.685 94.315 98.965 ;
        RECT 114.310 97.525 114.590 97.805 ;
        RECT 114.310 97.125 114.590 97.405 ;
        RECT 114.310 96.725 114.590 97.005 ;
        RECT 66.965 96.405 67.245 96.685 ;
        RECT 67.365 96.405 67.645 96.685 ;
        RECT 67.765 96.405 68.045 96.685 ;
        RECT 90.745 96.405 91.025 96.685 ;
        RECT 91.145 96.405 91.425 96.685 ;
        RECT 91.545 96.405 91.825 96.685 ;
        RECT 109.815 95.375 110.095 95.655 ;
        RECT 111.185 95.375 111.465 95.655 ;
        RECT 112.555 95.375 112.835 95.655 ;
        RECT 64.475 94.125 64.755 94.405 ;
        RECT 64.875 94.125 65.155 94.405 ;
        RECT 69.225 94.125 69.505 94.405 ;
        RECT 89.285 94.125 89.565 94.405 ;
        RECT 93.635 94.125 93.915 94.405 ;
        RECT 94.035 94.125 94.315 94.405 ;
        RECT 123.020 97.655 123.300 97.935 ;
        RECT 124.390 97.655 124.670 97.935 ;
        RECT 64.475 91.845 64.755 92.125 ;
        RECT 64.875 91.845 65.155 92.125 ;
        RECT 69.225 91.845 69.505 92.125 ;
        RECT 89.285 91.845 89.565 92.125 ;
        RECT 93.635 91.845 93.915 92.125 ;
        RECT 94.035 91.845 94.315 92.125 ;
        RECT 123.020 93.095 123.300 93.375 ;
        RECT 124.390 93.095 124.670 93.375 ;
        RECT 109.815 90.815 110.095 91.095 ;
        RECT 111.185 90.815 111.465 91.095 ;
        RECT 112.555 90.815 112.835 91.095 ;
        RECT 64.475 89.565 64.755 89.845 ;
        RECT 64.875 89.565 65.155 89.845 ;
        RECT 69.225 89.565 69.505 89.845 ;
        RECT 89.285 89.565 89.565 89.845 ;
        RECT 93.635 89.565 93.915 89.845 ;
        RECT 94.035 89.565 94.315 89.845 ;
        RECT 64.475 88.895 64.755 89.175 ;
        RECT 64.875 88.895 65.155 89.175 ;
        RECT 69.225 88.895 69.505 89.175 ;
        RECT 89.285 88.895 89.565 89.175 ;
        RECT 93.635 88.895 93.915 89.175 ;
        RECT 94.035 88.895 94.315 89.175 ;
        RECT 123.020 88.535 123.300 88.815 ;
        RECT 124.390 88.535 124.670 88.815 ;
        RECT 79.190 86.400 79.470 86.680 ;
        RECT 79.590 86.400 79.870 86.680 ;
        RECT 79.990 86.400 80.270 86.680 ;
        RECT 104.230 86.560 104.510 86.840 ;
        RECT 104.230 86.160 104.510 86.440 ;
        RECT 109.815 86.255 110.095 86.535 ;
        RECT 111.185 86.255 111.465 86.535 ;
        RECT 112.555 86.255 112.835 86.535 ;
        RECT 104.230 85.760 104.510 86.040 ;
        RECT 83.825 84.730 84.105 85.010 ;
        RECT 84.225 84.730 84.505 85.010 ;
        RECT 74.455 83.600 74.735 83.880 ;
        RECT 74.855 83.600 75.135 83.880 ;
        RECT 75.255 83.600 75.535 83.880 ;
        RECT 86.310 83.600 86.590 83.880 ;
        RECT 86.710 83.600 86.990 83.880 ;
        RECT 87.110 83.600 87.390 83.880 ;
        RECT 71.950 82.950 72.230 83.230 ;
        RECT 71.950 82.550 72.230 82.830 ;
        RECT 78.610 82.950 78.890 83.230 ;
        RECT 71.950 82.150 72.230 82.430 ;
        RECT 72.680 82.365 72.960 82.645 ;
        RECT 73.080 82.365 73.360 82.645 ;
        RECT 75.905 82.365 76.185 82.645 ;
        RECT 76.305 82.365 76.585 82.645 ;
        RECT 77.480 82.365 77.760 82.645 ;
        RECT 77.880 82.365 78.160 82.645 ;
        RECT 78.610 82.550 78.890 82.830 ;
        RECT 78.610 82.150 78.890 82.430 ;
        RECT 79.670 82.950 79.950 83.230 ;
        RECT 79.670 82.550 79.950 82.830 ;
        RECT 86.330 82.950 86.610 83.230 ;
        RECT 79.670 82.150 79.950 82.430 ;
        RECT 80.400 82.365 80.680 82.645 ;
        RECT 80.800 82.365 81.080 82.645 ;
        RECT 81.975 82.365 82.255 82.645 ;
        RECT 82.375 82.365 82.655 82.645 ;
        RECT 85.200 82.365 85.480 82.645 ;
        RECT 85.600 82.365 85.880 82.645 ;
        RECT 86.330 82.550 86.610 82.830 ;
        RECT 86.330 82.150 86.610 82.430 ;
        RECT 72.680 81.695 72.960 81.975 ;
        RECT 73.080 81.695 73.360 81.975 ;
        RECT 72.680 81.265 72.960 81.545 ;
        RECT 73.080 81.265 73.360 81.545 ;
        RECT 74.455 81.525 74.735 81.805 ;
        RECT 75.905 81.695 76.185 81.975 ;
        RECT 76.305 81.695 76.585 81.975 ;
        RECT 77.480 81.695 77.760 81.975 ;
        RECT 77.880 81.695 78.160 81.975 ;
        RECT 80.400 81.695 80.680 81.975 ;
        RECT 80.800 81.695 81.080 81.975 ;
        RECT 81.975 81.695 82.255 81.975 ;
        RECT 82.375 81.695 82.655 81.975 ;
        RECT 74.455 81.125 74.735 81.405 ;
        RECT 75.905 81.265 76.185 81.545 ;
        RECT 76.305 81.265 76.585 81.545 ;
        RECT 77.480 81.265 77.760 81.545 ;
        RECT 77.880 81.265 78.160 81.545 ;
        RECT 80.400 81.265 80.680 81.545 ;
        RECT 80.800 81.265 81.080 81.545 ;
        RECT 81.975 81.265 82.255 81.545 ;
        RECT 82.375 81.265 82.655 81.545 ;
        RECT 83.825 81.525 84.105 81.805 ;
        RECT 85.200 81.695 85.480 81.975 ;
        RECT 85.600 81.695 85.880 81.975 ;
        RECT 71.950 80.605 72.230 80.885 ;
        RECT 72.680 80.835 72.960 81.115 ;
        RECT 73.080 80.835 73.360 81.115 ;
        RECT 83.825 81.125 84.105 81.405 ;
        RECT 85.200 81.265 85.480 81.545 ;
        RECT 85.600 81.265 85.880 81.545 ;
        RECT 77.480 80.835 77.760 81.115 ;
        RECT 77.880 80.835 78.160 81.115 ;
        RECT 71.950 80.205 72.230 80.485 ;
        RECT 72.680 79.975 72.960 80.255 ;
        RECT 73.080 79.975 73.360 80.255 ;
        RECT 78.610 80.375 78.890 80.655 ;
        RECT 77.480 79.975 77.760 80.255 ;
        RECT 77.880 79.975 78.160 80.255 ;
        RECT 78.610 79.975 78.890 80.255 ;
        RECT 78.610 79.575 78.890 79.855 ;
        RECT 72.680 79.115 72.960 79.395 ;
        RECT 73.080 79.115 73.360 79.395 ;
        RECT 72.680 78.685 72.960 78.965 ;
        RECT 73.080 78.685 73.360 78.965 ;
        RECT 74.455 78.905 74.735 79.185 ;
        RECT 77.480 79.115 77.760 79.395 ;
        RECT 77.880 79.115 78.160 79.395 ;
        RECT 80.400 80.835 80.680 81.115 ;
        RECT 80.800 80.835 81.080 81.115 ;
        RECT 85.200 80.835 85.480 81.115 ;
        RECT 85.600 80.835 85.880 81.115 ;
        RECT 79.670 80.375 79.950 80.655 ;
        RECT 86.330 80.605 86.610 80.885 ;
        RECT 79.670 79.975 79.950 80.255 ;
        RECT 80.400 79.975 80.680 80.255 ;
        RECT 80.800 79.975 81.080 80.255 ;
        RECT 79.670 79.575 79.950 79.855 ;
        RECT 85.200 79.975 85.480 80.255 ;
        RECT 85.600 79.975 85.880 80.255 ;
        RECT 86.330 80.205 86.610 80.485 ;
        RECT 80.400 79.115 80.680 79.395 ;
        RECT 80.800 79.115 81.080 79.395 ;
        RECT 72.680 78.255 72.960 78.535 ;
        RECT 73.080 78.255 73.360 78.535 ;
        RECT 74.455 78.505 74.735 78.785 ;
        RECT 75.905 78.685 76.185 78.965 ;
        RECT 76.305 78.685 76.585 78.965 ;
        RECT 77.480 78.685 77.760 78.965 ;
        RECT 77.880 78.685 78.160 78.965 ;
        RECT 80.400 78.685 80.680 78.965 ;
        RECT 80.800 78.685 81.080 78.965 ;
        RECT 81.975 78.685 82.255 78.965 ;
        RECT 82.375 78.685 82.655 78.965 ;
        RECT 83.825 78.905 84.105 79.185 ;
        RECT 85.200 79.115 85.480 79.395 ;
        RECT 85.600 79.115 85.880 79.395 ;
        RECT 75.905 78.255 76.185 78.535 ;
        RECT 76.305 78.255 76.585 78.535 ;
        RECT 77.480 78.255 77.760 78.535 ;
        RECT 77.880 78.255 78.160 78.535 ;
        RECT 80.400 78.255 80.680 78.535 ;
        RECT 80.800 78.255 81.080 78.535 ;
        RECT 81.975 78.255 82.255 78.535 ;
        RECT 82.375 78.255 82.655 78.535 ;
        RECT 83.825 78.505 84.105 78.785 ;
        RECT 85.200 78.685 85.480 78.965 ;
        RECT 85.600 78.685 85.880 78.965 ;
        RECT 74.455 77.950 74.735 78.230 ;
        RECT 72.680 77.605 72.960 77.885 ;
        RECT 73.080 77.605 73.360 77.885 ;
        RECT 85.200 78.255 85.480 78.535 ;
        RECT 85.600 78.255 85.880 78.535 ;
        RECT 83.825 77.950 84.105 78.230 ;
        RECT 74.455 77.550 74.735 77.830 ;
        RECT 75.905 77.605 76.185 77.885 ;
        RECT 76.305 77.605 76.585 77.885 ;
        RECT 77.480 77.605 77.760 77.885 ;
        RECT 77.880 77.605 78.160 77.885 ;
        RECT 80.400 77.605 80.680 77.885 ;
        RECT 80.800 77.605 81.080 77.885 ;
        RECT 81.975 77.605 82.255 77.885 ;
        RECT 82.375 77.605 82.655 77.885 ;
        RECT 87.110 77.950 87.390 78.230 ;
        RECT 83.825 77.550 84.105 77.830 ;
        RECT 85.200 77.605 85.480 77.885 ;
        RECT 85.600 77.605 85.880 77.885 ;
        RECT 87.110 77.550 87.390 77.830 ;
        RECT 74.455 77.150 74.735 77.430 ;
        RECT 78.870 77.130 79.150 77.410 ;
        RECT 79.270 77.130 79.550 77.410 ;
        RECT 79.670 77.130 79.950 77.410 ;
        RECT 83.825 77.150 84.105 77.430 ;
        RECT 87.110 77.150 87.390 77.430 ;
        RECT 123.020 86.255 123.300 86.535 ;
        RECT 124.390 86.255 124.670 86.535 ;
        RECT 123.020 83.975 123.300 84.255 ;
        RECT 124.390 83.975 124.670 84.255 ;
        RECT 89.270 82.715 89.550 82.995 ;
        RECT 89.670 82.715 89.950 82.995 ;
        RECT 93.120 82.715 93.400 82.995 ;
        RECT 93.520 82.715 93.800 82.995 ;
        RECT 89.270 82.045 89.550 82.325 ;
        RECT 89.670 82.045 89.950 82.325 ;
        RECT 91.145 81.990 91.425 82.270 ;
        RECT 93.120 82.045 93.400 82.325 ;
        RECT 93.520 82.045 93.800 82.325 ;
        RECT 89.270 81.615 89.550 81.895 ;
        RECT 89.670 81.615 89.950 81.895 ;
        RECT 115.400 82.655 115.680 82.935 ;
        RECT 115.400 82.255 115.680 82.535 ;
        RECT 91.145 81.590 91.425 81.870 ;
        RECT 93.120 81.615 93.400 81.895 ;
        RECT 93.520 81.615 93.800 81.895 ;
        RECT 109.815 81.695 110.095 81.975 ;
        RECT 111.185 81.695 111.465 81.975 ;
        RECT 112.555 81.695 112.835 81.975 ;
        RECT 117.740 81.995 118.020 82.275 ;
        RECT 89.270 81.185 89.550 81.465 ;
        RECT 89.670 81.185 89.950 81.465 ;
        RECT 93.120 81.185 93.400 81.465 ;
        RECT 93.520 81.185 93.800 81.465 ;
        RECT 89.270 80.325 89.550 80.605 ;
        RECT 89.670 80.325 89.950 80.605 ;
        RECT 93.120 80.325 93.400 80.605 ;
        RECT 93.520 80.325 93.800 80.605 ;
        RECT 89.270 79.465 89.550 79.745 ;
        RECT 89.670 79.465 89.950 79.745 ;
        RECT 93.120 79.465 93.400 79.745 ;
        RECT 93.520 79.465 93.800 79.745 ;
        RECT 117.740 81.595 118.020 81.875 ;
        RECT 89.270 79.035 89.550 79.315 ;
        RECT 89.670 79.035 89.950 79.315 ;
        RECT 91.145 79.155 91.425 79.435 ;
        RECT 93.120 79.035 93.400 79.315 ;
        RECT 93.520 79.035 93.800 79.315 ;
        RECT 89.270 78.605 89.550 78.885 ;
        RECT 89.670 78.605 89.950 78.885 ;
        RECT 91.145 78.755 91.425 79.035 ;
        RECT 89.270 77.935 89.550 78.215 ;
        RECT 89.670 77.935 89.950 78.215 ;
        RECT 93.120 78.605 93.400 78.885 ;
        RECT 93.520 78.605 93.800 78.885 ;
        RECT 93.120 77.935 93.400 78.215 ;
        RECT 93.520 77.935 93.800 78.215 ;
        RECT 109.815 77.135 110.095 77.415 ;
        RECT 111.185 77.135 111.465 77.415 ;
        RECT 112.555 77.135 112.835 77.415 ;
        RECT 117.740 81.195 118.020 81.475 ;
        RECT 117.740 80.795 118.020 81.075 ;
        RECT 121.180 81.650 121.460 81.930 ;
        RECT 124.390 81.695 124.670 81.975 ;
        RECT 121.180 81.250 121.460 81.530 ;
        RECT 121.180 80.850 121.460 81.130 ;
        RECT 117.740 80.395 118.020 80.675 ;
        RECT 117.740 79.995 118.020 80.275 ;
        RECT 117.740 79.595 118.020 79.875 ;
        RECT 117.740 79.195 118.020 79.475 ;
        RECT 120.380 79.750 120.660 80.030 ;
        RECT 120.380 79.350 120.660 79.630 ;
        RECT 123.020 79.415 123.300 79.695 ;
        RECT 124.390 79.415 124.670 79.695 ;
        RECT 117.740 78.795 118.020 79.075 ;
        RECT 120.380 78.950 120.660 79.230 ;
        RECT 117.740 78.395 118.020 78.675 ;
        RECT 117.740 77.995 118.020 78.275 ;
        RECT 117.740 77.595 118.020 77.875 ;
        RECT 117.740 77.195 118.020 77.475 ;
        RECT 123.020 77.135 123.300 77.415 ;
        RECT 124.390 77.135 124.670 77.415 ;
        RECT 76.385 75.920 76.665 76.200 ;
        RECT 76.385 75.520 76.665 75.800 ;
        RECT 91.145 74.850 91.425 75.130 ;
        RECT 94.670 74.870 94.950 75.150 ;
        RECT 95.070 74.870 95.350 75.150 ;
        RECT 95.470 74.870 95.750 75.150 ;
        RECT 117.740 76.795 118.020 77.075 ;
        RECT 123.020 76.505 123.300 76.785 ;
        RECT 124.390 76.505 124.670 76.785 ;
        RECT 116.810 76.105 117.090 76.385 ;
        RECT 116.810 75.705 117.090 75.985 ;
        RECT 115.955 75.100 116.235 75.380 ;
        RECT 91.145 74.450 91.425 74.730 ;
        RECT 91.145 74.050 91.425 74.330 ;
        RECT 109.815 72.575 110.095 72.855 ;
        RECT 111.185 72.575 111.465 72.855 ;
        RECT 112.555 72.575 112.835 72.855 ;
        RECT 65.490 72.055 65.770 72.335 ;
        RECT 65.890 72.055 66.170 72.335 ;
        RECT 69.340 72.055 69.620 72.335 ;
        RECT 69.740 72.055 70.020 72.335 ;
        RECT 74.510 72.055 74.790 72.335 ;
        RECT 74.910 72.055 75.190 72.335 ;
        RECT 78.360 72.055 78.640 72.335 ;
        RECT 78.760 72.055 79.040 72.335 ;
        RECT 81.450 72.055 81.730 72.335 ;
        RECT 81.850 72.055 82.130 72.335 ;
        RECT 85.300 72.055 85.580 72.335 ;
        RECT 85.700 72.055 85.980 72.335 ;
        RECT 89.270 72.055 89.550 72.335 ;
        RECT 89.670 72.055 89.950 72.335 ;
        RECT 93.120 72.055 93.400 72.335 ;
        RECT 93.520 72.055 93.800 72.335 ;
        RECT 65.490 71.385 65.770 71.665 ;
        RECT 65.890 71.385 66.170 71.665 ;
        RECT 67.365 71.330 67.645 71.610 ;
        RECT 69.340 71.385 69.620 71.665 ;
        RECT 69.740 71.385 70.020 71.665 ;
        RECT 74.510 71.385 74.790 71.665 ;
        RECT 74.910 71.385 75.190 71.665 ;
        RECT 65.490 70.955 65.770 71.235 ;
        RECT 65.890 70.955 66.170 71.235 ;
        RECT 76.385 71.330 76.665 71.610 ;
        RECT 78.360 71.385 78.640 71.665 ;
        RECT 78.760 71.385 79.040 71.665 ;
        RECT 81.450 71.385 81.730 71.665 ;
        RECT 81.850 71.385 82.130 71.665 ;
        RECT 67.365 70.930 67.645 71.210 ;
        RECT 69.340 70.955 69.620 71.235 ;
        RECT 69.740 70.955 70.020 71.235 ;
        RECT 74.510 70.955 74.790 71.235 ;
        RECT 74.910 70.955 75.190 71.235 ;
        RECT 83.825 71.330 84.105 71.610 ;
        RECT 85.300 71.385 85.580 71.665 ;
        RECT 85.700 71.385 85.980 71.665 ;
        RECT 89.270 71.385 89.550 71.665 ;
        RECT 89.670 71.385 89.950 71.665 ;
        RECT 76.385 70.930 76.665 71.210 ;
        RECT 78.360 70.955 78.640 71.235 ;
        RECT 78.760 70.955 79.040 71.235 ;
        RECT 81.450 70.955 81.730 71.235 ;
        RECT 81.850 70.955 82.130 71.235 ;
        RECT 91.145 71.330 91.425 71.610 ;
        RECT 93.120 71.385 93.400 71.665 ;
        RECT 93.520 71.385 93.800 71.665 ;
        RECT 83.825 70.930 84.105 71.210 ;
        RECT 85.300 70.955 85.580 71.235 ;
        RECT 85.700 70.955 85.980 71.235 ;
        RECT 89.270 70.955 89.550 71.235 ;
        RECT 89.670 70.955 89.950 71.235 ;
        RECT 91.145 70.930 91.425 71.210 ;
        RECT 93.120 70.955 93.400 71.235 ;
        RECT 93.520 70.955 93.800 71.235 ;
        RECT 65.490 70.525 65.770 70.805 ;
        RECT 65.890 70.525 66.170 70.805 ;
        RECT 69.340 70.525 69.620 70.805 ;
        RECT 69.740 70.525 70.020 70.805 ;
        RECT 74.510 70.525 74.790 70.805 ;
        RECT 74.910 70.525 75.190 70.805 ;
        RECT 78.360 70.525 78.640 70.805 ;
        RECT 78.760 70.525 79.040 70.805 ;
        RECT 81.450 70.525 81.730 70.805 ;
        RECT 81.850 70.525 82.130 70.805 ;
        RECT 85.300 70.525 85.580 70.805 ;
        RECT 85.700 70.525 85.980 70.805 ;
        RECT 89.270 70.525 89.550 70.805 ;
        RECT 89.670 70.525 89.950 70.805 ;
        RECT 93.120 70.525 93.400 70.805 ;
        RECT 93.520 70.525 93.800 70.805 ;
        RECT 123.985 70.955 124.265 71.235 ;
        RECT 115.955 70.325 116.235 70.605 ;
        RECT 65.490 69.665 65.770 69.945 ;
        RECT 65.890 69.665 66.170 69.945 ;
        RECT 69.340 69.665 69.620 69.945 ;
        RECT 69.740 69.665 70.020 69.945 ;
        RECT 74.510 69.665 74.790 69.945 ;
        RECT 74.910 69.665 75.190 69.945 ;
        RECT 78.360 69.665 78.640 69.945 ;
        RECT 78.760 69.665 79.040 69.945 ;
        RECT 81.450 69.665 81.730 69.945 ;
        RECT 81.850 69.665 82.130 69.945 ;
        RECT 85.300 69.665 85.580 69.945 ;
        RECT 85.700 69.665 85.980 69.945 ;
        RECT 89.270 69.665 89.550 69.945 ;
        RECT 89.670 69.665 89.950 69.945 ;
        RECT 119.650 70.045 119.930 70.325 ;
        RECT 93.120 69.665 93.400 69.945 ;
        RECT 93.520 69.665 93.800 69.945 ;
        RECT 115.955 69.655 116.235 69.935 ;
        RECT 119.650 69.375 119.930 69.655 ;
        RECT 65.490 68.805 65.770 69.085 ;
        RECT 65.890 68.805 66.170 69.085 ;
        RECT 69.340 68.805 69.620 69.085 ;
        RECT 69.740 68.805 70.020 69.085 ;
        RECT 74.510 68.805 74.790 69.085 ;
        RECT 74.910 68.805 75.190 69.085 ;
        RECT 78.360 68.805 78.640 69.085 ;
        RECT 78.760 68.805 79.040 69.085 ;
        RECT 81.450 68.805 81.730 69.085 ;
        RECT 81.850 68.805 82.130 69.085 ;
        RECT 85.300 68.805 85.580 69.085 ;
        RECT 85.700 68.805 85.980 69.085 ;
        RECT 89.270 68.805 89.550 69.085 ;
        RECT 89.670 68.805 89.950 69.085 ;
        RECT 93.120 68.805 93.400 69.085 ;
        RECT 93.520 68.805 93.800 69.085 ;
        RECT 119.650 68.945 119.930 69.225 ;
        RECT 123.985 70.555 124.265 70.835 ;
        RECT 123.985 70.155 124.265 70.435 ;
        RECT 125.635 70.005 125.915 70.285 ;
        RECT 123.070 69.350 123.350 69.630 ;
        RECT 125.635 69.375 125.915 69.655 ;
        RECT 123.070 68.950 123.350 69.230 ;
        RECT 121.200 68.515 121.480 68.795 ;
        RECT 121.600 68.515 121.880 68.795 ;
        RECT 125.635 68.945 125.915 69.225 ;
        RECT 125.635 68.515 125.915 68.795 ;
        RECT 65.490 67.945 65.770 68.225 ;
        RECT 65.890 67.945 66.170 68.225 ;
        RECT 69.340 67.945 69.620 68.225 ;
        RECT 69.740 67.945 70.020 68.225 ;
        RECT 74.510 67.945 74.790 68.225 ;
        RECT 74.910 67.945 75.190 68.225 ;
        RECT 78.360 67.945 78.640 68.225 ;
        RECT 78.760 67.945 79.040 68.225 ;
        RECT 81.450 67.945 81.730 68.225 ;
        RECT 81.850 67.945 82.130 68.225 ;
        RECT 85.300 67.945 85.580 68.225 ;
        RECT 85.700 67.945 85.980 68.225 ;
        RECT 89.270 67.945 89.550 68.225 ;
        RECT 89.670 67.945 89.950 68.225 ;
        RECT 93.120 67.945 93.400 68.225 ;
        RECT 93.520 67.945 93.800 68.225 ;
        RECT 109.815 68.015 110.095 68.295 ;
        RECT 111.185 68.015 111.465 68.295 ;
        RECT 112.555 68.015 112.835 68.295 ;
        RECT 125.635 68.085 125.915 68.365 ;
        RECT 121.200 67.655 121.480 67.935 ;
        RECT 121.600 67.655 121.880 67.935 ;
        RECT 65.490 67.085 65.770 67.365 ;
        RECT 65.890 67.085 66.170 67.365 ;
        RECT 69.340 67.085 69.620 67.365 ;
        RECT 69.740 67.085 70.020 67.365 ;
        RECT 74.510 67.085 74.790 67.365 ;
        RECT 74.910 67.085 75.190 67.365 ;
        RECT 78.360 67.085 78.640 67.365 ;
        RECT 78.760 67.085 79.040 67.365 ;
        RECT 81.450 67.085 81.730 67.365 ;
        RECT 81.850 67.085 82.130 67.365 ;
        RECT 85.300 67.085 85.580 67.365 ;
        RECT 85.700 67.085 85.980 67.365 ;
        RECT 89.270 67.085 89.550 67.365 ;
        RECT 89.670 67.085 89.950 67.365 ;
        RECT 115.955 67.375 116.235 67.655 ;
        RECT 93.120 67.085 93.400 67.365 ;
        RECT 93.520 67.085 93.800 67.365 ;
        RECT 125.635 67.655 125.915 67.935 ;
        RECT 125.635 67.225 125.915 67.505 ;
        RECT 121.200 66.795 121.480 67.075 ;
        RECT 121.600 66.795 121.880 67.075 ;
        RECT 65.490 66.225 65.770 66.505 ;
        RECT 65.890 66.225 66.170 66.505 ;
        RECT 69.340 66.225 69.620 66.505 ;
        RECT 69.740 66.225 70.020 66.505 ;
        RECT 74.510 66.225 74.790 66.505 ;
        RECT 74.910 66.225 75.190 66.505 ;
        RECT 78.360 66.225 78.640 66.505 ;
        RECT 78.760 66.225 79.040 66.505 ;
        RECT 81.450 66.225 81.730 66.505 ;
        RECT 81.850 66.225 82.130 66.505 ;
        RECT 85.300 66.225 85.580 66.505 ;
        RECT 85.700 66.225 85.980 66.505 ;
        RECT 89.270 66.225 89.550 66.505 ;
        RECT 89.670 66.225 89.950 66.505 ;
        RECT 93.120 66.225 93.400 66.505 ;
        RECT 93.520 66.225 93.800 66.505 ;
        RECT 65.490 65.365 65.770 65.645 ;
        RECT 65.890 65.365 66.170 65.645 ;
        RECT 69.340 65.365 69.620 65.645 ;
        RECT 69.740 65.365 70.020 65.645 ;
        RECT 74.510 65.365 74.790 65.645 ;
        RECT 74.910 65.365 75.190 65.645 ;
        RECT 78.360 65.365 78.640 65.645 ;
        RECT 78.760 65.365 79.040 65.645 ;
        RECT 81.450 65.365 81.730 65.645 ;
        RECT 81.850 65.365 82.130 65.645 ;
        RECT 85.300 65.365 85.580 65.645 ;
        RECT 85.700 65.365 85.980 65.645 ;
        RECT 89.270 65.365 89.550 65.645 ;
        RECT 89.670 65.365 89.950 65.645 ;
        RECT 109.815 65.735 110.095 66.015 ;
        RECT 111.185 65.735 111.465 66.015 ;
        RECT 112.555 65.735 112.835 66.015 ;
        RECT 93.120 65.365 93.400 65.645 ;
        RECT 93.520 65.365 93.800 65.645 ;
        RECT 119.650 66.365 119.930 66.645 ;
        RECT 119.650 65.935 119.930 66.215 ;
        RECT 65.490 64.505 65.770 64.785 ;
        RECT 65.890 64.505 66.170 64.785 ;
        RECT 69.340 64.505 69.620 64.785 ;
        RECT 69.740 64.505 70.020 64.785 ;
        RECT 74.510 64.505 74.790 64.785 ;
        RECT 74.910 64.505 75.190 64.785 ;
        RECT 65.490 64.075 65.770 64.355 ;
        RECT 65.890 64.075 66.170 64.355 ;
        RECT 67.365 64.195 67.645 64.475 ;
        RECT 78.360 64.505 78.640 64.785 ;
        RECT 78.760 64.505 79.040 64.785 ;
        RECT 81.450 64.505 81.730 64.785 ;
        RECT 81.850 64.505 82.130 64.785 ;
        RECT 69.340 64.075 69.620 64.355 ;
        RECT 69.740 64.075 70.020 64.355 ;
        RECT 74.510 64.075 74.790 64.355 ;
        RECT 74.910 64.075 75.190 64.355 ;
        RECT 76.385 64.195 76.665 64.475 ;
        RECT 85.300 64.505 85.580 64.785 ;
        RECT 85.700 64.505 85.980 64.785 ;
        RECT 89.270 64.505 89.550 64.785 ;
        RECT 89.670 64.505 89.950 64.785 ;
        RECT 78.360 64.075 78.640 64.355 ;
        RECT 78.760 64.075 79.040 64.355 ;
        RECT 81.450 64.075 81.730 64.355 ;
        RECT 81.850 64.075 82.130 64.355 ;
        RECT 83.825 64.195 84.105 64.475 ;
        RECT 93.120 64.505 93.400 64.785 ;
        RECT 93.520 64.505 93.800 64.785 ;
        RECT 85.300 64.075 85.580 64.355 ;
        RECT 85.700 64.075 85.980 64.355 ;
        RECT 89.270 64.075 89.550 64.355 ;
        RECT 89.670 64.075 89.950 64.355 ;
        RECT 91.145 64.195 91.425 64.475 ;
        RECT 93.120 64.075 93.400 64.355 ;
        RECT 93.520 64.075 93.800 64.355 ;
        RECT 65.490 63.645 65.770 63.925 ;
        RECT 65.890 63.645 66.170 63.925 ;
        RECT 67.365 63.795 67.645 64.075 ;
        RECT 69.340 63.645 69.620 63.925 ;
        RECT 69.740 63.645 70.020 63.925 ;
        RECT 74.510 63.645 74.790 63.925 ;
        RECT 74.910 63.645 75.190 63.925 ;
        RECT 76.385 63.795 76.665 64.075 ;
        RECT 78.360 63.645 78.640 63.925 ;
        RECT 78.760 63.645 79.040 63.925 ;
        RECT 81.450 63.645 81.730 63.925 ;
        RECT 81.850 63.645 82.130 63.925 ;
        RECT 83.825 63.795 84.105 64.075 ;
        RECT 85.300 63.645 85.580 63.925 ;
        RECT 85.700 63.645 85.980 63.925 ;
        RECT 89.270 63.645 89.550 63.925 ;
        RECT 89.670 63.645 89.950 63.925 ;
        RECT 91.145 63.795 91.425 64.075 ;
        RECT 93.120 63.645 93.400 63.925 ;
        RECT 93.520 63.645 93.800 63.925 ;
        RECT 109.815 63.455 110.095 63.735 ;
        RECT 111.185 63.455 111.465 63.735 ;
        RECT 112.555 63.455 112.835 63.735 ;
        RECT 125.635 66.795 125.915 67.075 ;
        RECT 125.635 66.365 125.915 66.645 ;
        RECT 125.635 65.935 125.915 66.215 ;
        RECT 127.420 65.460 127.700 65.740 ;
        RECT 125.635 65.075 125.915 65.355 ;
        RECT 127.420 65.060 127.700 65.340 ;
        RECT 127.420 64.660 127.700 64.940 ;
        RECT 119.650 64.125 119.930 64.405 ;
        RECT 120.465 63.980 120.745 64.260 ;
        RECT 119.650 63.695 119.930 63.975 ;
        RECT 120.465 63.580 120.745 63.860 ;
        RECT 121.200 63.265 121.480 63.545 ;
        RECT 121.600 63.265 121.880 63.545 ;
        RECT 65.490 62.975 65.770 63.255 ;
        RECT 65.890 62.975 66.170 63.255 ;
        RECT 69.340 62.975 69.620 63.255 ;
        RECT 69.740 62.975 70.020 63.255 ;
        RECT 74.510 62.975 74.790 63.255 ;
        RECT 74.910 62.975 75.190 63.255 ;
        RECT 78.360 62.975 78.640 63.255 ;
        RECT 78.760 62.975 79.040 63.255 ;
        RECT 81.450 62.975 81.730 63.255 ;
        RECT 81.850 62.975 82.130 63.255 ;
        RECT 85.300 62.975 85.580 63.255 ;
        RECT 85.700 62.975 85.980 63.255 ;
        RECT 89.270 62.975 89.550 63.255 ;
        RECT 89.670 62.975 89.950 63.255 ;
        RECT 93.120 62.975 93.400 63.255 ;
        RECT 93.520 62.975 93.800 63.255 ;
        RECT 109.815 62.785 110.095 63.065 ;
        RECT 111.185 62.785 111.465 63.065 ;
        RECT 112.555 62.785 112.835 63.065 ;
        RECT 115.955 62.815 116.235 63.095 ;
        RECT 121.200 62.405 121.480 62.685 ;
        RECT 121.600 62.405 121.880 62.685 ;
        RECT 121.180 61.545 121.460 61.825 ;
        RECT 121.580 61.545 121.860 61.825 ;
        RECT 119.650 61.115 119.930 61.395 ;
        RECT 123.985 61.200 124.265 61.480 ;
        RECT 115.955 60.535 116.235 60.815 ;
        RECT 119.650 60.685 119.930 60.965 ;
        RECT 123.985 60.800 124.265 61.080 ;
        RECT 115.955 59.865 116.235 60.145 ;
        RECT 119.650 60.055 119.930 60.335 ;
        RECT 120.465 59.175 120.745 59.455 ;
        RECT 120.865 59.175 121.145 59.455 ;
        RECT 122.670 59.175 122.950 59.455 ;
        RECT 123.070 59.175 123.350 59.455 ;
        RECT 125.635 64.215 125.915 64.495 ;
        RECT 125.635 63.785 125.915 64.065 ;
        RECT 125.635 63.355 125.915 63.635 ;
        RECT 125.635 62.925 125.915 63.205 ;
        RECT 125.635 62.495 125.915 62.775 ;
        RECT 125.635 62.065 125.915 62.345 ;
        RECT 125.635 61.635 125.915 61.915 ;
        RECT 125.635 61.205 125.915 61.485 ;
        RECT 125.635 60.775 125.915 61.055 ;
        RECT 125.635 60.145 125.915 60.425 ;
        RECT 124.800 56.950 125.080 57.230 ;
        RECT 124.800 56.550 125.080 56.830 ;
        RECT 124.800 56.150 125.080 56.430 ;
        RECT 124.800 55.750 125.080 56.030 ;
        RECT 124.800 55.350 125.080 55.630 ;
        RECT 124.665 38.355 124.945 38.635 ;
        RECT 125.065 38.355 125.345 38.635 ;
        RECT 125.465 38.355 125.745 38.635 ;
        RECT 140.825 38.355 141.105 38.635 ;
        RECT 141.225 38.355 141.505 38.635 ;
        RECT 141.625 38.355 141.905 38.635 ;
        RECT 142.025 38.355 142.305 38.635 ;
        RECT 104.230 21.430 104.510 21.710 ;
        RECT 104.230 21.030 104.510 21.310 ;
        RECT 124.800 21.165 125.080 21.445 ;
        RECT 72.305 20.570 72.585 20.850 ;
        RECT 104.230 20.630 104.510 20.910 ;
        RECT 124.800 20.765 125.080 21.045 ;
        RECT 72.305 20.170 72.585 20.450 ;
        RECT 124.800 20.365 125.080 20.645 ;
        RECT 72.305 19.770 72.585 20.050 ;
        RECT 123.985 19.730 124.265 20.010 ;
        RECT 123.985 19.330 124.265 19.610 ;
        RECT 87.560 18.920 87.840 19.200 ;
        RECT 87.960 18.920 88.240 19.200 ;
        RECT 88.360 18.920 88.640 19.200 ;
        RECT 122.250 18.920 122.530 19.200 ;
        RECT 122.650 18.920 122.930 19.200 ;
        RECT 123.050 18.920 123.330 19.200 ;
        RECT 123.985 18.930 124.265 19.210 ;
        RECT 105.195 17.955 105.475 18.235 ;
        RECT 105.595 17.955 105.875 18.235 ;
        RECT 105.995 17.955 106.275 18.235 ;
        RECT 116.940 17.955 117.220 18.235 ;
        RECT 117.340 17.955 117.620 18.235 ;
        RECT 117.740 17.955 118.020 18.235 ;
        RECT 91.145 16.430 91.425 16.710 ;
        RECT 91.145 16.030 91.425 16.310 ;
        RECT 91.145 15.630 91.425 15.910 ;
        RECT 83.160 14.690 83.440 14.970 ;
        RECT 83.560 14.690 83.840 14.970 ;
        RECT 83.960 14.690 84.240 14.970 ;
        RECT 117.740 12.755 118.020 13.035 ;
        RECT 118.140 12.755 118.420 13.035 ;
        RECT 118.540 12.755 118.820 13.035 ;
        RECT 140.825 12.755 141.105 13.035 ;
        RECT 141.225 12.755 141.505 13.035 ;
        RECT 141.625 12.755 141.905 13.035 ;
        RECT 142.025 12.755 142.305 13.035 ;
        RECT 76.250 7.410 76.530 7.690 ;
        RECT 76.650 7.410 76.930 7.690 ;
        RECT 77.050 7.410 77.330 7.690 ;
        RECT 112.095 7.410 112.375 7.690 ;
        RECT 112.495 7.410 112.775 7.690 ;
        RECT 67.230 6.310 67.510 6.590 ;
        RECT 67.630 6.310 67.910 6.590 ;
        RECT 68.030 6.310 68.310 6.590 ;
        RECT 90.015 6.310 90.295 6.590 ;
        RECT 90.415 6.310 90.695 6.590 ;
        RECT 157.825 5.030 158.105 5.310 ;
        RECT 157.825 4.630 158.105 4.910 ;
        RECT 134.505 3.990 134.785 4.270 ;
        RECT 134.905 3.990 135.185 4.270 ;
        RECT 135.305 3.990 135.585 4.270 ;
        RECT 135.705 3.990 135.985 4.270 ;
        RECT 157.825 4.230 158.105 4.510 ;
        RECT 157.825 3.830 158.105 4.110 ;
      LAYER met3 ;
        RECT 3.980 219.015 81.585 220.515 ;
        RECT 127.395 211.950 128.525 212.280 ;
        RECT 142.980 211.950 144.160 212.280 ;
        RECT 115.375 211.120 116.505 211.450 ;
        RECT 106.100 206.195 107.230 206.795 ;
        RECT 84.910 173.475 85.290 174.625 ;
        RECT 88.590 172.375 88.970 173.525 ;
        RECT 1.000 168.710 55.500 171.710 ;
        RECT 49.000 64.160 52.000 163.185 ;
        RECT 52.500 59.435 55.500 168.710 ;
        RECT 78.045 153.950 79.175 154.550 ;
        RECT 63.170 151.655 64.300 151.985 ;
        RECT 56.100 127.580 56.430 139.185 ;
        RECT 57.150 89.185 58.150 151.600 ;
        RECT 60.740 111.570 61.740 151.600 ;
        RECT 63.170 148.510 63.500 151.655 ;
        RECT 62.685 146.660 63.415 146.990 ;
        RECT 63.085 139.310 63.415 146.660 ;
        RECT 62.685 138.980 63.415 139.310 ;
        RECT 63.085 134.750 63.415 138.980 ;
        RECT 62.685 134.420 63.415 134.750 ;
        RECT 63.085 130.190 63.415 134.420 ;
        RECT 62.685 129.860 63.415 130.190 ;
        RECT 62.685 125.300 63.415 125.630 ;
        RECT 63.085 121.070 63.415 125.300 ;
        RECT 63.765 122.795 64.095 146.965 ;
        RECT 62.685 120.740 63.415 121.070 ;
        RECT 63.085 116.510 63.415 120.740 ;
        RECT 62.685 116.180 63.415 116.510 ;
        RECT 65.405 114.185 65.905 151.600 ;
        RECT 64.315 88.770 65.315 113.385 ;
        RECT 67.000 106.625 67.330 134.285 ;
        RECT 67.680 106.625 68.010 134.280 ;
        RECT 69.160 117.160 70.160 138.390 ;
        RECT 66.940 96.380 68.070 96.710 ;
        RECT 67.340 83.850 67.670 96.380 ;
        RECT 69.115 88.770 69.615 115.185 ;
        RECT 71.310 111.975 71.640 151.960 ;
        RECT 72.135 136.135 72.465 146.965 ;
        RECT 73.560 91.185 74.060 142.825 ;
        RECT 75.055 115.700 75.385 139.790 ;
        RECT 72.595 89.185 74.060 91.185 ;
        RECT 76.300 89.185 76.800 142.825 ;
        RECT 78.045 140.790 78.645 153.950 ;
        RECT 80.145 153.450 80.745 154.550 ;
        RECT 104.640 153.950 105.770 154.550 ;
        RECT 80.145 152.850 81.275 153.450 ;
        RECT 80.145 140.790 80.745 152.850 ;
        RECT 77.460 125.625 77.840 126.745 ;
        RECT 80.950 125.625 81.330 126.745 ;
        RECT 78.900 114.370 80.030 114.700 ;
        RECT 67.340 83.520 72.255 83.850 ;
        RECT 65.330 62.910 66.330 72.460 ;
        RECT 67.340 70.895 67.670 83.520 ;
        RECT 71.925 80.180 72.255 83.520 ;
        RECT 1.000 56.435 55.500 59.435 ;
        RECT 67.205 6.750 67.805 64.565 ;
        RECT 69.180 62.910 70.180 79.185 ;
        RECT 72.595 77.580 73.445 89.185 ;
        RECT 79.165 86.840 79.765 114.370 ;
        RECT 81.990 89.185 82.490 142.825 ;
        RECT 83.405 115.700 83.735 139.790 ;
        RECT 84.730 91.185 85.230 142.825 ;
        RECT 86.325 136.135 86.655 146.965 ;
        RECT 87.150 111.975 87.480 151.960 ;
        RECT 94.490 151.655 95.620 151.985 ;
        RECT 88.630 117.160 89.630 138.390 ;
        RECT 84.730 89.185 85.965 91.185 ;
        RECT 79.165 86.240 80.295 86.840 ;
        RECT 83.800 84.705 84.530 85.035 ;
        RECT 74.430 83.575 75.560 83.905 ;
        RECT 74.430 81.035 74.760 83.575 ;
        RECT 74.430 77.105 74.760 79.325 ;
        RECT 75.820 77.580 76.670 82.670 ;
        RECT 77.395 77.580 78.245 82.670 ;
        RECT 78.585 79.390 78.915 83.275 ;
        RECT 79.645 77.435 79.975 83.300 ;
        RECT 80.315 79.185 81.165 82.670 ;
        RECT 81.890 79.185 82.740 82.670 ;
        RECT 83.800 81.035 84.130 84.705 ;
        RECT 80.315 77.580 82.740 79.185 ;
        RECT 78.845 77.105 79.975 77.435 ;
        RECT 76.360 74.840 76.690 76.290 ;
        RECT 72.280 74.510 76.690 74.840 ;
        RECT 72.280 19.725 72.610 74.510 ;
        RECT 74.350 62.910 75.350 72.460 ;
        RECT 76.360 70.895 76.690 74.510 ;
        RECT 76.225 7.850 76.825 64.565 ;
        RECT 78.200 62.910 79.200 72.460 ;
        RECT 81.290 62.910 82.290 77.580 ;
        RECT 83.800 74.840 84.130 79.325 ;
        RECT 85.115 77.580 85.965 89.185 ;
        RECT 89.175 88.770 89.675 115.185 ;
        RECT 90.780 106.625 91.110 134.280 ;
        RECT 91.460 106.625 91.790 134.285 ;
        RECT 92.885 114.185 93.385 151.600 ;
        RECT 95.290 148.510 95.620 151.655 ;
        RECT 94.695 122.795 95.025 146.965 ;
        RECT 95.375 146.660 96.105 146.990 ;
        RECT 95.375 139.310 95.705 146.660 ;
        RECT 95.375 138.980 96.105 139.310 ;
        RECT 95.375 134.750 95.705 138.980 ;
        RECT 95.375 134.420 96.105 134.750 ;
        RECT 95.375 130.190 95.705 134.420 ;
        RECT 95.375 129.860 96.105 130.190 ;
        RECT 95.375 125.300 96.105 125.630 ;
        RECT 95.375 121.070 95.705 125.300 ;
        RECT 95.375 120.740 96.105 121.070 ;
        RECT 95.375 116.510 95.705 120.740 ;
        RECT 95.375 116.180 96.105 116.510 ;
        RECT 90.720 96.380 91.850 96.710 ;
        RECT 91.120 84.210 91.450 96.380 ;
        RECT 93.475 88.770 94.475 113.385 ;
        RECT 97.050 111.570 98.050 151.600 ;
        RECT 100.640 89.185 101.640 151.600 ;
        RECT 102.360 127.580 102.690 139.185 ;
        RECT 86.285 83.575 87.415 83.905 ;
        RECT 86.305 80.180 86.635 83.275 ;
        RECT 87.085 77.105 87.415 83.575 ;
        RECT 91.120 83.880 95.775 84.210 ;
        RECT 83.800 74.510 87.845 74.840 ;
        RECT 83.800 70.895 84.130 74.510 ;
        RECT 83.665 15.130 84.265 64.565 ;
        RECT 85.140 62.910 86.140 72.460 ;
        RECT 87.515 19.225 87.845 74.510 ;
        RECT 89.110 62.910 90.110 83.120 ;
        RECT 91.120 81.555 91.450 83.880 ;
        RECT 91.120 78.075 91.450 79.525 ;
        RECT 91.120 70.895 91.450 75.175 ;
        RECT 87.515 18.895 88.665 19.225 ;
        RECT 90.985 15.605 91.585 64.565 ;
        RECT 92.960 62.910 93.960 83.120 ;
        RECT 95.445 75.175 95.775 83.880 ;
        RECT 94.645 74.845 95.775 75.175 ;
        RECT 104.070 20.605 104.670 86.865 ;
        RECT 105.170 18.395 105.770 153.950 ;
        RECT 106.100 18.900 106.700 206.195 ;
        RECT 115.375 175.700 115.705 211.120 ;
        RECT 120.355 210.290 121.485 210.620 ;
        RECT 117.715 208.090 118.845 208.690 ;
        RECT 110.195 175.370 115.705 175.700 ;
        RECT 108.195 168.750 109.195 174.000 ;
        RECT 110.195 173.735 110.525 175.370 ;
        RECT 110.195 173.405 110.535 173.735 ;
        RECT 110.205 172.435 110.535 173.405 ;
        RECT 110.205 168.955 110.535 170.405 ;
        RECT 112.045 168.750 113.045 174.000 ;
        RECT 108.195 167.130 108.895 168.750 ;
        RECT 107.250 166.430 108.895 167.130 ;
        RECT 107.250 161.185 107.950 166.430 ;
        RECT 109.605 62.760 110.305 164.750 ;
        RECT 110.975 62.760 111.675 164.750 ;
        RECT 112.345 62.760 113.045 168.750 ;
        RECT 114.285 96.595 114.615 101.030 ;
        RECT 115.375 76.055 115.705 175.370 ;
        RECT 116.785 75.670 117.115 206.795 ;
        RECT 117.715 110.830 118.045 208.090 ;
        RECT 115.745 59.840 116.445 75.405 ;
        RECT 117.715 18.395 118.045 82.440 ;
        RECT 120.355 78.925 120.685 210.290 ;
        RECT 123.680 209.190 124.410 209.790 ;
        RECT 123.680 165.005 124.010 209.190 ;
        RECT 119.440 65.320 120.140 70.350 ;
        RECT 121.155 68.820 121.485 81.975 ;
        RECT 122.810 76.480 123.510 164.710 ;
        RECT 124.180 73.675 124.880 164.710 ;
        RECT 124.180 72.975 126.125 73.675 ;
        RECT 121.155 68.490 121.905 68.820 ;
        RECT 121.155 67.960 121.485 68.490 ;
        RECT 121.155 67.630 121.905 67.960 ;
        RECT 121.155 67.100 121.485 67.630 ;
        RECT 121.155 66.770 121.905 67.100 ;
        RECT 119.440 60.030 120.140 64.980 ;
        RECT 120.440 59.480 120.770 64.465 ;
        RECT 121.155 63.570 121.485 66.770 ;
        RECT 121.155 63.240 121.905 63.570 ;
        RECT 121.155 62.710 121.485 63.240 ;
        RECT 121.155 62.380 121.905 62.710 ;
        RECT 121.155 61.850 121.485 62.380 ;
        RECT 121.155 61.520 121.885 61.850 ;
        RECT 123.045 59.480 123.375 69.805 ;
        RECT 120.440 59.150 121.170 59.480 ;
        RECT 122.645 59.150 123.375 59.480 ;
        RECT 123.045 19.225 123.375 59.150 ;
        RECT 122.225 18.895 123.375 19.225 ;
        RECT 105.170 17.795 106.300 18.395 ;
        RECT 116.915 17.795 118.045 18.395 ;
        RECT 123.045 17.795 123.375 18.895 ;
        RECT 123.960 17.795 124.290 71.280 ;
        RECT 125.425 60.120 126.125 72.975 ;
        RECT 124.640 38.795 125.240 57.310 ;
        RECT 124.640 38.195 125.770 38.795 ;
        RECT 124.640 17.795 125.240 38.195 ;
        RECT 127.395 17.795 127.725 211.950 ;
        RECT 146.655 210.290 147.835 210.620 ;
        RECT 140.605 208.090 142.530 208.690 ;
        RECT 129.470 184.290 153.530 206.890 ;
        RECT 129.470 158.995 153.530 181.595 ;
        RECT 129.470 135.195 153.530 157.795 ;
        RECT 129.470 111.395 153.530 133.995 ;
        RECT 129.470 87.595 153.530 110.195 ;
        RECT 129.470 63.795 153.530 86.395 ;
        RECT 129.470 39.995 153.530 62.595 ;
        RECT 140.605 38.195 142.530 38.795 ;
        RECT 83.135 14.530 84.265 15.130 ;
        RECT 117.715 13.195 118.045 17.795 ;
        RECT 129.470 14.395 153.530 36.995 ;
        RECT 117.715 12.595 118.845 13.195 ;
        RECT 140.605 12.595 142.530 13.195 ;
        RECT 76.225 7.250 77.355 7.850 ;
        RECT 111.875 7.250 113.000 7.850 ;
        RECT 67.205 6.150 68.335 6.750 ;
        RECT 89.795 6.150 90.920 6.750 ;
        RECT 134.480 3.830 136.010 4.430 ;
        RECT 90.320 1.565 90.920 3.505 ;
        RECT 112.400 1.565 113.000 3.505 ;
        RECT 134.480 1.565 135.080 3.505 ;
        RECT 156.565 1.565 157.165 209.815 ;
        RECT 157.665 3.805 158.265 211.475 ;
      LAYER via3 ;
        RECT 3.980 220.005 4.300 220.325 ;
        RECT 7.660 220.005 7.980 220.325 ;
        RECT 11.340 220.005 11.660 220.325 ;
        RECT 15.020 220.005 15.340 220.325 ;
        RECT 18.700 220.005 19.020 220.325 ;
        RECT 22.380 220.005 22.700 220.325 ;
        RECT 26.060 220.005 26.380 220.325 ;
        RECT 29.740 220.005 30.060 220.325 ;
        RECT 33.420 220.005 33.740 220.325 ;
        RECT 37.100 220.005 37.420 220.325 ;
        RECT 40.780 220.005 41.100 220.325 ;
        RECT 44.460 220.005 44.780 220.325 ;
        RECT 48.140 220.005 48.460 220.325 ;
        RECT 3.980 219.605 4.300 219.925 ;
        RECT 7.660 219.605 7.980 219.925 ;
        RECT 11.340 219.605 11.660 219.925 ;
        RECT 15.020 219.605 15.340 219.925 ;
        RECT 18.700 219.605 19.020 219.925 ;
        RECT 22.380 219.605 22.700 219.925 ;
        RECT 26.060 219.605 26.380 219.925 ;
        RECT 29.740 219.605 30.060 219.925 ;
        RECT 33.420 219.605 33.740 219.925 ;
        RECT 37.100 219.605 37.420 219.925 ;
        RECT 40.780 219.605 41.100 219.925 ;
        RECT 44.460 219.605 44.780 219.925 ;
        RECT 48.140 219.605 48.460 219.925 ;
        RECT 3.980 219.205 4.300 219.525 ;
        RECT 7.660 219.205 7.980 219.525 ;
        RECT 11.340 219.205 11.660 219.525 ;
        RECT 15.020 219.205 15.340 219.525 ;
        RECT 18.700 219.205 19.020 219.525 ;
        RECT 22.380 219.205 22.700 219.525 ;
        RECT 26.060 219.205 26.380 219.525 ;
        RECT 29.740 219.205 30.060 219.525 ;
        RECT 33.420 219.205 33.740 219.525 ;
        RECT 37.100 219.205 37.420 219.525 ;
        RECT 40.780 219.205 41.100 219.525 ;
        RECT 44.460 219.205 44.780 219.525 ;
        RECT 48.140 219.205 48.460 219.525 ;
        RECT 49.190 219.205 50.310 220.325 ;
        RECT 51.820 220.005 52.140 220.325 ;
        RECT 55.500 220.005 55.820 220.325 ;
        RECT 59.180 220.005 59.500 220.325 ;
        RECT 62.860 220.005 63.180 220.325 ;
        RECT 66.540 220.005 66.860 220.325 ;
        RECT 70.220 220.005 70.540 220.325 ;
        RECT 73.900 220.005 74.220 220.325 ;
        RECT 77.580 220.005 77.900 220.325 ;
        RECT 81.260 220.005 81.580 220.325 ;
        RECT 51.820 219.605 52.140 219.925 ;
        RECT 55.500 219.605 55.820 219.925 ;
        RECT 59.180 219.605 59.500 219.925 ;
        RECT 62.860 219.605 63.180 219.925 ;
        RECT 66.540 219.605 66.860 219.925 ;
        RECT 70.220 219.605 70.540 219.925 ;
        RECT 73.900 219.605 74.220 219.925 ;
        RECT 77.580 219.605 77.900 219.925 ;
        RECT 81.260 219.605 81.580 219.925 ;
        RECT 51.820 219.205 52.140 219.525 ;
        RECT 55.500 219.205 55.820 219.525 ;
        RECT 59.180 219.205 59.500 219.525 ;
        RECT 62.860 219.205 63.180 219.525 ;
        RECT 66.540 219.205 66.860 219.525 ;
        RECT 70.220 219.205 70.540 219.525 ;
        RECT 73.900 219.205 74.220 219.525 ;
        RECT 77.580 219.205 77.900 219.525 ;
        RECT 81.260 219.205 81.580 219.525 ;
        RECT 143.010 211.955 143.330 212.275 ;
        RECT 143.410 211.955 143.730 212.275 ;
        RECT 143.810 211.955 144.130 212.275 ;
        RECT 84.940 174.275 85.260 174.595 ;
        RECT 84.940 173.875 85.260 174.195 ;
        RECT 84.940 173.475 85.260 173.795 ;
        RECT 88.620 173.175 88.940 173.495 ;
        RECT 88.620 172.775 88.940 173.095 ;
        RECT 88.620 172.375 88.940 172.695 ;
        RECT 1.190 168.850 2.310 171.570 ;
        RECT 49.140 161.225 51.860 163.145 ;
        RECT 49.190 139.430 50.310 160.950 ;
        RECT 49.140 137.225 51.860 139.145 ;
        RECT 49.190 115.430 50.310 136.950 ;
        RECT 49.140 113.225 51.860 115.145 ;
        RECT 49.190 91.430 50.310 112.950 ;
        RECT 49.140 89.225 51.860 91.145 ;
        RECT 49.190 67.430 50.310 88.950 ;
        RECT 49.140 65.225 51.860 67.145 ;
        RECT 49.190 64.265 50.310 64.985 ;
        RECT 52.640 149.225 55.360 151.145 ;
        RECT 57.290 149.225 58.010 151.145 ;
        RECT 56.105 138.425 56.425 138.745 ;
        RECT 56.105 138.025 56.425 138.345 ;
        RECT 56.105 137.625 56.425 137.945 ;
        RECT 52.640 125.225 55.360 127.145 ;
        RECT 52.640 101.225 55.360 103.145 ;
        RECT 57.290 125.225 58.010 127.145 ;
        RECT 60.880 149.225 61.600 151.145 ;
        RECT 60.880 125.225 61.600 127.145 ;
        RECT 65.495 138.825 65.815 139.145 ;
        RECT 65.495 138.425 65.815 138.745 ;
        RECT 65.495 138.025 65.815 138.345 ;
        RECT 65.495 137.625 65.815 137.945 ;
        RECT 65.495 137.225 65.815 137.545 ;
        RECT 65.495 114.825 65.815 115.145 ;
        RECT 65.495 114.425 65.815 114.745 ;
        RECT 57.290 101.225 58.010 103.145 ;
        RECT 69.300 125.225 70.020 127.145 ;
        RECT 69.205 114.825 69.525 115.145 ;
        RECT 69.205 114.425 69.525 114.745 ;
        RECT 69.205 114.025 69.525 114.345 ;
        RECT 69.205 113.625 69.525 113.945 ;
        RECT 69.205 113.225 69.525 113.545 ;
        RECT 64.455 101.225 65.175 103.145 ;
        RECT 52.640 77.225 55.360 79.145 ;
        RECT 73.650 138.825 73.970 139.145 ;
        RECT 73.650 138.425 73.970 138.745 ;
        RECT 73.650 138.025 73.970 138.345 ;
        RECT 73.650 137.625 73.970 137.945 ;
        RECT 73.650 137.225 73.970 137.545 ;
        RECT 76.390 138.825 76.710 139.145 ;
        RECT 76.390 138.425 76.710 138.745 ;
        RECT 76.390 138.025 76.710 138.345 ;
        RECT 76.390 137.625 76.710 137.945 ;
        RECT 76.390 137.225 76.710 137.545 ;
        RECT 73.650 114.825 73.970 115.145 ;
        RECT 73.650 114.425 73.970 114.745 ;
        RECT 73.650 114.025 73.970 114.345 ;
        RECT 73.650 113.625 73.970 113.945 ;
        RECT 73.650 113.225 73.970 113.545 ;
        RECT 69.205 90.825 69.525 91.145 ;
        RECT 69.205 90.425 69.525 90.745 ;
        RECT 69.205 90.025 69.525 90.345 ;
        RECT 69.205 89.625 69.525 89.945 ;
        RECT 69.205 89.225 69.525 89.545 ;
        RECT 73.650 90.825 73.970 91.145 ;
        RECT 73.650 90.425 73.970 90.745 ;
        RECT 73.650 90.025 73.970 90.345 ;
        RECT 73.650 89.625 73.970 89.945 ;
        RECT 73.650 89.225 73.970 89.545 ;
        RECT 82.080 138.825 82.400 139.145 ;
        RECT 82.080 138.425 82.400 138.745 ;
        RECT 82.080 138.025 82.400 138.345 ;
        RECT 82.080 137.625 82.400 137.945 ;
        RECT 82.080 137.225 82.400 137.545 ;
        RECT 77.490 126.425 77.810 126.745 ;
        RECT 77.490 126.025 77.810 126.345 ;
        RECT 77.490 125.625 77.810 125.945 ;
        RECT 80.980 126.425 81.300 126.745 ;
        RECT 80.980 126.025 81.300 126.345 ;
        RECT 80.980 125.625 81.300 125.945 ;
        RECT 76.390 114.825 76.710 115.145 ;
        RECT 76.390 114.425 76.710 114.745 ;
        RECT 84.820 138.825 85.140 139.145 ;
        RECT 84.820 138.425 85.140 138.745 ;
        RECT 84.820 138.025 85.140 138.345 ;
        RECT 84.820 137.625 85.140 137.945 ;
        RECT 84.820 137.225 85.140 137.545 ;
        RECT 82.080 114.825 82.400 115.145 ;
        RECT 82.080 114.425 82.400 114.745 ;
        RECT 76.390 114.025 76.710 114.345 ;
        RECT 76.390 113.625 76.710 113.945 ;
        RECT 76.390 113.225 76.710 113.545 ;
        RECT 76.390 90.825 76.710 91.145 ;
        RECT 76.390 90.425 76.710 90.745 ;
        RECT 76.390 90.025 76.710 90.345 ;
        RECT 76.390 89.625 76.710 89.945 ;
        RECT 76.390 89.225 76.710 89.545 ;
        RECT 82.080 114.025 82.400 114.345 ;
        RECT 82.080 113.625 82.400 113.945 ;
        RECT 82.080 113.225 82.400 113.545 ;
        RECT 82.080 90.825 82.400 91.145 ;
        RECT 82.080 90.425 82.400 90.745 ;
        RECT 82.080 90.025 82.400 90.345 ;
        RECT 82.080 89.625 82.400 89.945 ;
        RECT 82.080 89.225 82.400 89.545 ;
        RECT 84.820 114.825 85.140 115.145 ;
        RECT 84.820 114.425 85.140 114.745 ;
        RECT 84.820 114.025 85.140 114.345 ;
        RECT 84.820 113.625 85.140 113.945 ;
        RECT 84.820 113.225 85.140 113.545 ;
        RECT 97.190 149.225 97.910 151.145 ;
        RECT 92.975 138.825 93.295 139.145 ;
        RECT 92.975 138.425 93.295 138.745 ;
        RECT 92.975 138.025 93.295 138.345 ;
        RECT 92.975 137.625 93.295 137.945 ;
        RECT 92.975 137.225 93.295 137.545 ;
        RECT 88.770 125.225 89.490 127.145 ;
        RECT 89.265 114.825 89.585 115.145 ;
        RECT 89.265 114.425 89.585 114.745 ;
        RECT 89.265 114.025 89.585 114.345 ;
        RECT 89.265 113.625 89.585 113.945 ;
        RECT 89.265 113.225 89.585 113.545 ;
        RECT 84.820 90.825 85.140 91.145 ;
        RECT 85.460 90.825 85.780 91.145 ;
        RECT 84.820 90.425 85.140 90.745 ;
        RECT 85.460 90.425 85.780 90.745 ;
        RECT 84.820 90.025 85.140 90.345 ;
        RECT 85.460 90.025 85.780 90.345 ;
        RECT 84.820 89.625 85.140 89.945 ;
        RECT 85.460 89.625 85.780 89.945 ;
        RECT 84.820 89.225 85.140 89.545 ;
        RECT 85.460 89.225 85.780 89.545 ;
        RECT 72.660 81.750 73.380 82.470 ;
        RECT 69.320 77.225 70.040 79.145 ;
        RECT 65.470 65.225 66.190 67.145 ;
        RECT 1.190 56.575 2.310 59.295 ;
        RECT 75.885 77.750 76.605 78.470 ;
        RECT 77.460 77.750 78.180 78.470 ;
        RECT 97.190 125.225 97.910 127.145 ;
        RECT 92.975 114.825 93.295 115.145 ;
        RECT 92.975 114.425 93.295 114.745 ;
        RECT 100.780 149.225 101.500 151.145 ;
        RECT 102.365 138.425 102.685 138.745 ;
        RECT 102.365 138.025 102.685 138.345 ;
        RECT 102.365 137.625 102.685 137.945 ;
        RECT 100.780 125.225 101.500 127.145 ;
        RECT 93.615 101.225 94.335 103.145 ;
        RECT 89.265 90.825 89.585 91.145 ;
        RECT 89.265 90.425 89.585 90.745 ;
        RECT 89.265 90.025 89.585 90.345 ;
        RECT 89.265 89.625 89.585 89.945 ;
        RECT 89.265 89.225 89.585 89.545 ;
        RECT 100.780 101.225 101.500 103.145 ;
        RECT 85.180 81.750 85.900 82.470 ;
        RECT 80.380 77.750 81.100 78.470 ;
        RECT 81.955 77.750 82.675 78.470 ;
        RECT 74.490 65.225 75.210 67.145 ;
        RECT 85.280 65.225 86.000 67.145 ;
        RECT 93.100 77.225 93.820 79.145 ;
        RECT 89.250 65.225 89.970 67.145 ;
        RECT 107.440 162.825 107.760 163.145 ;
        RECT 107.440 162.425 107.760 162.745 ;
        RECT 107.440 162.025 107.760 162.345 ;
        RECT 107.440 161.625 107.760 161.945 ;
        RECT 107.440 161.225 107.760 161.545 ;
        RECT 109.795 150.825 110.115 151.145 ;
        RECT 109.795 150.425 110.115 150.745 ;
        RECT 109.795 150.025 110.115 150.345 ;
        RECT 109.795 149.625 110.115 149.945 ;
        RECT 109.795 149.225 110.115 149.545 ;
        RECT 109.795 126.825 110.115 127.145 ;
        RECT 109.795 126.425 110.115 126.745 ;
        RECT 109.795 126.025 110.115 126.345 ;
        RECT 109.795 125.625 110.115 125.945 ;
        RECT 109.795 125.225 110.115 125.545 ;
        RECT 109.795 102.825 110.115 103.145 ;
        RECT 109.795 102.425 110.115 102.745 ;
        RECT 109.795 102.025 110.115 102.345 ;
        RECT 109.795 101.625 110.115 101.945 ;
        RECT 109.795 101.225 110.115 101.545 ;
        RECT 109.795 78.825 110.115 79.145 ;
        RECT 109.795 78.425 110.115 78.745 ;
        RECT 109.795 78.025 110.115 78.345 ;
        RECT 109.795 77.625 110.115 77.945 ;
        RECT 109.795 77.225 110.115 77.545 ;
        RECT 111.165 150.825 111.485 151.145 ;
        RECT 111.165 150.425 111.485 150.745 ;
        RECT 111.165 150.025 111.485 150.345 ;
        RECT 111.165 149.625 111.485 149.945 ;
        RECT 111.165 149.225 111.485 149.545 ;
        RECT 111.165 126.825 111.485 127.145 ;
        RECT 111.165 126.425 111.485 126.745 ;
        RECT 111.165 126.025 111.485 126.345 ;
        RECT 111.165 125.625 111.485 125.945 ;
        RECT 111.165 125.225 111.485 125.545 ;
        RECT 111.165 102.825 111.485 103.145 ;
        RECT 111.165 102.425 111.485 102.745 ;
        RECT 111.165 102.025 111.485 102.345 ;
        RECT 111.165 101.625 111.485 101.945 ;
        RECT 111.165 101.225 111.485 101.545 ;
        RECT 111.165 78.825 111.485 79.145 ;
        RECT 111.165 78.425 111.485 78.745 ;
        RECT 111.165 78.025 111.485 78.345 ;
        RECT 111.165 77.625 111.485 77.945 ;
        RECT 111.165 77.225 111.485 77.545 ;
        RECT 112.535 150.825 112.855 151.145 ;
        RECT 112.535 150.425 112.855 150.745 ;
        RECT 112.535 150.025 112.855 150.345 ;
        RECT 112.535 149.625 112.855 149.945 ;
        RECT 112.535 149.225 112.855 149.545 ;
        RECT 112.535 126.825 112.855 127.145 ;
        RECT 112.535 126.425 112.855 126.745 ;
        RECT 112.535 126.025 112.855 126.345 ;
        RECT 112.535 125.625 112.855 125.945 ;
        RECT 112.535 125.225 112.855 125.545 ;
        RECT 112.535 102.825 112.855 103.145 ;
        RECT 112.535 102.425 112.855 102.745 ;
        RECT 112.535 102.025 112.855 102.345 ;
        RECT 112.535 101.625 112.855 101.945 ;
        RECT 112.535 101.225 112.855 101.545 ;
        RECT 112.535 78.825 112.855 79.145 ;
        RECT 112.535 78.425 112.855 78.745 ;
        RECT 112.535 78.025 112.855 78.345 ;
        RECT 112.535 77.625 112.855 77.945 ;
        RECT 112.535 77.225 112.855 77.545 ;
        RECT 123.000 162.825 123.320 163.145 ;
        RECT 123.000 162.425 123.320 162.745 ;
        RECT 123.000 162.025 123.320 162.345 ;
        RECT 123.000 161.625 123.320 161.945 ;
        RECT 123.000 161.225 123.320 161.545 ;
        RECT 123.000 138.825 123.320 139.145 ;
        RECT 123.000 138.425 123.320 138.745 ;
        RECT 123.000 138.025 123.320 138.345 ;
        RECT 123.000 137.625 123.320 137.945 ;
        RECT 123.000 137.225 123.320 137.545 ;
        RECT 123.000 114.825 123.320 115.145 ;
        RECT 123.000 114.425 123.320 114.745 ;
        RECT 123.000 114.025 123.320 114.345 ;
        RECT 123.000 113.625 123.320 113.945 ;
        RECT 123.000 113.225 123.320 113.545 ;
        RECT 123.000 90.825 123.320 91.145 ;
        RECT 123.000 90.425 123.320 90.745 ;
        RECT 123.000 90.025 123.320 90.345 ;
        RECT 123.000 89.625 123.320 89.945 ;
        RECT 123.000 89.225 123.320 89.545 ;
        RECT 124.370 162.825 124.690 163.145 ;
        RECT 124.370 162.425 124.690 162.745 ;
        RECT 124.370 162.025 124.690 162.345 ;
        RECT 124.370 161.625 124.690 161.945 ;
        RECT 124.370 161.225 124.690 161.545 ;
        RECT 124.370 138.825 124.690 139.145 ;
        RECT 124.370 138.425 124.690 138.745 ;
        RECT 124.370 138.025 124.690 138.345 ;
        RECT 124.370 137.625 124.690 137.945 ;
        RECT 124.370 137.225 124.690 137.545 ;
        RECT 124.370 114.825 124.690 115.145 ;
        RECT 124.370 114.425 124.690 114.745 ;
        RECT 124.370 114.025 124.690 114.345 ;
        RECT 124.370 113.625 124.690 113.945 ;
        RECT 124.370 113.225 124.690 113.545 ;
        RECT 124.370 90.825 124.690 91.145 ;
        RECT 124.370 90.425 124.690 90.745 ;
        RECT 124.370 90.025 124.690 90.345 ;
        RECT 124.370 89.625 124.690 89.945 ;
        RECT 124.370 89.225 124.690 89.545 ;
        RECT 125.615 66.825 125.935 67.145 ;
        RECT 125.615 66.425 125.935 66.745 ;
        RECT 125.615 66.025 125.935 66.345 ;
        RECT 125.615 65.625 125.935 65.945 ;
        RECT 125.615 65.225 125.935 65.545 ;
        RECT 146.685 210.295 147.005 210.615 ;
        RECT 147.085 210.295 147.405 210.615 ;
        RECT 147.485 210.295 147.805 210.615 ;
        RECT 140.605 208.230 140.925 208.550 ;
        RECT 141.005 208.230 141.325 208.550 ;
        RECT 141.405 208.230 141.725 208.550 ;
        RECT 141.805 208.230 142.125 208.550 ;
        RECT 142.205 208.230 142.525 208.550 ;
        RECT 129.570 206.430 129.890 206.750 ;
        RECT 129.570 206.030 129.890 206.350 ;
        RECT 129.570 205.630 129.890 205.950 ;
        RECT 129.570 205.230 129.890 205.550 ;
        RECT 129.570 204.830 129.890 205.150 ;
        RECT 129.570 204.430 129.890 204.750 ;
        RECT 129.570 204.030 129.890 204.350 ;
        RECT 129.570 203.630 129.890 203.950 ;
        RECT 129.570 203.230 129.890 203.550 ;
        RECT 129.570 202.830 129.890 203.150 ;
        RECT 129.570 202.430 129.890 202.750 ;
        RECT 129.570 202.030 129.890 202.350 ;
        RECT 129.570 201.630 129.890 201.950 ;
        RECT 129.570 201.230 129.890 201.550 ;
        RECT 129.570 200.830 129.890 201.150 ;
        RECT 129.570 200.430 129.890 200.750 ;
        RECT 129.570 200.030 129.890 200.350 ;
        RECT 129.570 199.630 129.890 199.950 ;
        RECT 129.570 199.230 129.890 199.550 ;
        RECT 129.570 198.830 129.890 199.150 ;
        RECT 129.570 198.430 129.890 198.750 ;
        RECT 129.570 198.030 129.890 198.350 ;
        RECT 129.570 197.630 129.890 197.950 ;
        RECT 129.570 197.230 129.890 197.550 ;
        RECT 129.570 196.830 129.890 197.150 ;
        RECT 129.570 196.430 129.890 196.750 ;
        RECT 129.570 196.030 129.890 196.350 ;
        RECT 129.570 195.630 129.890 195.950 ;
        RECT 129.570 195.230 129.890 195.550 ;
        RECT 129.570 194.830 129.890 195.150 ;
        RECT 129.570 194.430 129.890 194.750 ;
        RECT 129.570 194.030 129.890 194.350 ;
        RECT 129.570 193.630 129.890 193.950 ;
        RECT 129.570 193.230 129.890 193.550 ;
        RECT 129.570 192.830 129.890 193.150 ;
        RECT 129.570 192.430 129.890 192.750 ;
        RECT 129.570 192.030 129.890 192.350 ;
        RECT 129.570 191.630 129.890 191.950 ;
        RECT 129.570 191.230 129.890 191.550 ;
        RECT 129.570 190.830 129.890 191.150 ;
        RECT 129.570 190.430 129.890 190.750 ;
        RECT 129.570 190.030 129.890 190.350 ;
        RECT 129.570 189.630 129.890 189.950 ;
        RECT 129.570 189.230 129.890 189.550 ;
        RECT 129.570 188.830 129.890 189.150 ;
        RECT 129.570 188.430 129.890 188.750 ;
        RECT 129.570 188.030 129.890 188.350 ;
        RECT 129.570 187.630 129.890 187.950 ;
        RECT 129.570 187.230 129.890 187.550 ;
        RECT 129.570 186.830 129.890 187.150 ;
        RECT 129.570 186.430 129.890 186.750 ;
        RECT 129.570 186.030 129.890 186.350 ;
        RECT 129.570 185.630 129.890 185.950 ;
        RECT 129.570 185.230 129.890 185.550 ;
        RECT 129.570 184.830 129.890 185.150 ;
        RECT 129.570 184.430 129.890 184.750 ;
        RECT 129.570 181.135 129.890 181.455 ;
        RECT 129.570 180.735 129.890 181.055 ;
        RECT 129.570 180.335 129.890 180.655 ;
        RECT 129.570 179.935 129.890 180.255 ;
        RECT 129.570 179.535 129.890 179.855 ;
        RECT 129.570 179.135 129.890 179.455 ;
        RECT 129.570 178.735 129.890 179.055 ;
        RECT 129.570 178.335 129.890 178.655 ;
        RECT 129.570 177.935 129.890 178.255 ;
        RECT 129.570 177.535 129.890 177.855 ;
        RECT 129.570 177.135 129.890 177.455 ;
        RECT 129.570 176.735 129.890 177.055 ;
        RECT 129.570 176.335 129.890 176.655 ;
        RECT 129.570 175.935 129.890 176.255 ;
        RECT 129.570 175.535 129.890 175.855 ;
        RECT 129.570 175.135 129.890 175.455 ;
        RECT 129.570 174.735 129.890 175.055 ;
        RECT 129.570 174.335 129.890 174.655 ;
        RECT 129.570 173.935 129.890 174.255 ;
        RECT 129.570 173.535 129.890 173.855 ;
        RECT 129.570 173.135 129.890 173.455 ;
        RECT 129.570 172.735 129.890 173.055 ;
        RECT 129.570 172.335 129.890 172.655 ;
        RECT 129.570 171.935 129.890 172.255 ;
        RECT 129.570 171.535 129.890 171.855 ;
        RECT 129.570 171.135 129.890 171.455 ;
        RECT 129.570 170.735 129.890 171.055 ;
        RECT 129.570 170.335 129.890 170.655 ;
        RECT 129.570 169.935 129.890 170.255 ;
        RECT 129.570 169.535 129.890 169.855 ;
        RECT 129.570 169.135 129.890 169.455 ;
        RECT 129.570 168.735 129.890 169.055 ;
        RECT 129.570 168.335 129.890 168.655 ;
        RECT 129.570 167.935 129.890 168.255 ;
        RECT 129.570 167.535 129.890 167.855 ;
        RECT 129.570 167.135 129.890 167.455 ;
        RECT 129.570 166.735 129.890 167.055 ;
        RECT 129.570 166.335 129.890 166.655 ;
        RECT 129.570 165.935 129.890 166.255 ;
        RECT 129.570 165.535 129.890 165.855 ;
        RECT 129.570 165.135 129.890 165.455 ;
        RECT 129.570 164.735 129.890 165.055 ;
        RECT 129.570 164.335 129.890 164.655 ;
        RECT 129.570 163.935 129.890 164.255 ;
        RECT 129.570 163.535 129.890 163.855 ;
        RECT 129.570 163.135 129.890 163.455 ;
        RECT 129.570 162.735 129.890 163.055 ;
        RECT 129.570 162.335 129.890 162.655 ;
        RECT 129.570 161.935 129.890 162.255 ;
        RECT 129.570 161.535 129.890 161.855 ;
        RECT 129.570 161.135 129.890 161.455 ;
        RECT 129.570 160.735 129.890 161.055 ;
        RECT 129.570 160.335 129.890 160.655 ;
        RECT 129.570 159.935 129.890 160.255 ;
        RECT 129.570 159.535 129.890 159.855 ;
        RECT 129.570 159.135 129.890 159.455 ;
        RECT 129.570 157.335 129.890 157.655 ;
        RECT 129.570 156.935 129.890 157.255 ;
        RECT 129.570 156.535 129.890 156.855 ;
        RECT 129.570 156.135 129.890 156.455 ;
        RECT 129.570 155.735 129.890 156.055 ;
        RECT 129.570 155.335 129.890 155.655 ;
        RECT 129.570 154.935 129.890 155.255 ;
        RECT 129.570 154.535 129.890 154.855 ;
        RECT 129.570 154.135 129.890 154.455 ;
        RECT 129.570 153.735 129.890 154.055 ;
        RECT 129.570 153.335 129.890 153.655 ;
        RECT 129.570 152.935 129.890 153.255 ;
        RECT 129.570 152.535 129.890 152.855 ;
        RECT 129.570 152.135 129.890 152.455 ;
        RECT 129.570 151.735 129.890 152.055 ;
        RECT 129.570 151.335 129.890 151.655 ;
        RECT 129.570 150.935 129.890 151.255 ;
        RECT 129.570 150.535 129.890 150.855 ;
        RECT 129.570 150.135 129.890 150.455 ;
        RECT 129.570 149.735 129.890 150.055 ;
        RECT 129.570 149.335 129.890 149.655 ;
        RECT 129.570 148.935 129.890 149.255 ;
        RECT 129.570 148.535 129.890 148.855 ;
        RECT 129.570 148.135 129.890 148.455 ;
        RECT 129.570 147.735 129.890 148.055 ;
        RECT 129.570 147.335 129.890 147.655 ;
        RECT 129.570 146.935 129.890 147.255 ;
        RECT 129.570 146.535 129.890 146.855 ;
        RECT 129.570 146.135 129.890 146.455 ;
        RECT 129.570 145.735 129.890 146.055 ;
        RECT 129.570 145.335 129.890 145.655 ;
        RECT 129.570 144.935 129.890 145.255 ;
        RECT 129.570 144.535 129.890 144.855 ;
        RECT 129.570 144.135 129.890 144.455 ;
        RECT 129.570 143.735 129.890 144.055 ;
        RECT 129.570 143.335 129.890 143.655 ;
        RECT 129.570 142.935 129.890 143.255 ;
        RECT 129.570 142.535 129.890 142.855 ;
        RECT 129.570 142.135 129.890 142.455 ;
        RECT 129.570 141.735 129.890 142.055 ;
        RECT 129.570 141.335 129.890 141.655 ;
        RECT 129.570 140.935 129.890 141.255 ;
        RECT 129.570 140.535 129.890 140.855 ;
        RECT 129.570 140.135 129.890 140.455 ;
        RECT 129.570 139.735 129.890 140.055 ;
        RECT 129.570 139.335 129.890 139.655 ;
        RECT 129.570 138.935 129.890 139.255 ;
        RECT 129.570 138.535 129.890 138.855 ;
        RECT 129.570 138.135 129.890 138.455 ;
        RECT 129.570 137.735 129.890 138.055 ;
        RECT 129.570 137.335 129.890 137.655 ;
        RECT 129.570 136.935 129.890 137.255 ;
        RECT 129.570 136.535 129.890 136.855 ;
        RECT 129.570 136.135 129.890 136.455 ;
        RECT 129.570 135.735 129.890 136.055 ;
        RECT 129.570 135.335 129.890 135.655 ;
        RECT 129.570 133.535 129.890 133.855 ;
        RECT 129.570 133.135 129.890 133.455 ;
        RECT 129.570 132.735 129.890 133.055 ;
        RECT 129.570 132.335 129.890 132.655 ;
        RECT 129.570 131.935 129.890 132.255 ;
        RECT 129.570 131.535 129.890 131.855 ;
        RECT 129.570 131.135 129.890 131.455 ;
        RECT 129.570 130.735 129.890 131.055 ;
        RECT 129.570 130.335 129.890 130.655 ;
        RECT 129.570 129.935 129.890 130.255 ;
        RECT 129.570 129.535 129.890 129.855 ;
        RECT 129.570 129.135 129.890 129.455 ;
        RECT 129.570 128.735 129.890 129.055 ;
        RECT 129.570 128.335 129.890 128.655 ;
        RECT 129.570 127.935 129.890 128.255 ;
        RECT 129.570 127.535 129.890 127.855 ;
        RECT 129.570 127.135 129.890 127.455 ;
        RECT 129.570 126.735 129.890 127.055 ;
        RECT 129.570 126.335 129.890 126.655 ;
        RECT 129.570 125.935 129.890 126.255 ;
        RECT 129.570 125.535 129.890 125.855 ;
        RECT 129.570 125.135 129.890 125.455 ;
        RECT 129.570 124.735 129.890 125.055 ;
        RECT 129.570 124.335 129.890 124.655 ;
        RECT 129.570 123.935 129.890 124.255 ;
        RECT 129.570 123.535 129.890 123.855 ;
        RECT 129.570 123.135 129.890 123.455 ;
        RECT 129.570 122.735 129.890 123.055 ;
        RECT 129.570 122.335 129.890 122.655 ;
        RECT 129.570 121.935 129.890 122.255 ;
        RECT 129.570 121.535 129.890 121.855 ;
        RECT 129.570 121.135 129.890 121.455 ;
        RECT 129.570 120.735 129.890 121.055 ;
        RECT 129.570 120.335 129.890 120.655 ;
        RECT 129.570 119.935 129.890 120.255 ;
        RECT 129.570 119.535 129.890 119.855 ;
        RECT 129.570 119.135 129.890 119.455 ;
        RECT 129.570 118.735 129.890 119.055 ;
        RECT 129.570 118.335 129.890 118.655 ;
        RECT 129.570 117.935 129.890 118.255 ;
        RECT 129.570 117.535 129.890 117.855 ;
        RECT 129.570 117.135 129.890 117.455 ;
        RECT 129.570 116.735 129.890 117.055 ;
        RECT 129.570 116.335 129.890 116.655 ;
        RECT 129.570 115.935 129.890 116.255 ;
        RECT 129.570 115.535 129.890 115.855 ;
        RECT 129.570 115.135 129.890 115.455 ;
        RECT 129.570 114.735 129.890 115.055 ;
        RECT 129.570 114.335 129.890 114.655 ;
        RECT 129.570 113.935 129.890 114.255 ;
        RECT 129.570 113.535 129.890 113.855 ;
        RECT 129.570 113.135 129.890 113.455 ;
        RECT 129.570 112.735 129.890 113.055 ;
        RECT 129.570 112.335 129.890 112.655 ;
        RECT 129.570 111.935 129.890 112.255 ;
        RECT 129.570 111.535 129.890 111.855 ;
        RECT 129.570 109.735 129.890 110.055 ;
        RECT 129.570 109.335 129.890 109.655 ;
        RECT 129.570 108.935 129.890 109.255 ;
        RECT 129.570 108.535 129.890 108.855 ;
        RECT 129.570 108.135 129.890 108.455 ;
        RECT 129.570 107.735 129.890 108.055 ;
        RECT 129.570 107.335 129.890 107.655 ;
        RECT 129.570 106.935 129.890 107.255 ;
        RECT 129.570 106.535 129.890 106.855 ;
        RECT 129.570 106.135 129.890 106.455 ;
        RECT 129.570 105.735 129.890 106.055 ;
        RECT 129.570 105.335 129.890 105.655 ;
        RECT 129.570 104.935 129.890 105.255 ;
        RECT 129.570 104.535 129.890 104.855 ;
        RECT 129.570 104.135 129.890 104.455 ;
        RECT 129.570 103.735 129.890 104.055 ;
        RECT 129.570 103.335 129.890 103.655 ;
        RECT 129.570 102.935 129.890 103.255 ;
        RECT 129.570 102.535 129.890 102.855 ;
        RECT 129.570 102.135 129.890 102.455 ;
        RECT 129.570 101.735 129.890 102.055 ;
        RECT 129.570 101.335 129.890 101.655 ;
        RECT 129.570 100.935 129.890 101.255 ;
        RECT 129.570 100.535 129.890 100.855 ;
        RECT 129.570 100.135 129.890 100.455 ;
        RECT 129.570 99.735 129.890 100.055 ;
        RECT 129.570 99.335 129.890 99.655 ;
        RECT 129.570 98.935 129.890 99.255 ;
        RECT 129.570 98.535 129.890 98.855 ;
        RECT 129.570 98.135 129.890 98.455 ;
        RECT 129.570 97.735 129.890 98.055 ;
        RECT 129.570 97.335 129.890 97.655 ;
        RECT 129.570 96.935 129.890 97.255 ;
        RECT 129.570 96.535 129.890 96.855 ;
        RECT 129.570 96.135 129.890 96.455 ;
        RECT 129.570 95.735 129.890 96.055 ;
        RECT 129.570 95.335 129.890 95.655 ;
        RECT 129.570 94.935 129.890 95.255 ;
        RECT 129.570 94.535 129.890 94.855 ;
        RECT 129.570 94.135 129.890 94.455 ;
        RECT 129.570 93.735 129.890 94.055 ;
        RECT 129.570 93.335 129.890 93.655 ;
        RECT 129.570 92.935 129.890 93.255 ;
        RECT 129.570 92.535 129.890 92.855 ;
        RECT 129.570 92.135 129.890 92.455 ;
        RECT 129.570 91.735 129.890 92.055 ;
        RECT 129.570 91.335 129.890 91.655 ;
        RECT 129.570 90.935 129.890 91.255 ;
        RECT 129.570 90.535 129.890 90.855 ;
        RECT 129.570 90.135 129.890 90.455 ;
        RECT 129.570 89.735 129.890 90.055 ;
        RECT 129.570 89.335 129.890 89.655 ;
        RECT 129.570 88.935 129.890 89.255 ;
        RECT 129.570 88.535 129.890 88.855 ;
        RECT 129.570 88.135 129.890 88.455 ;
        RECT 129.570 87.735 129.890 88.055 ;
        RECT 129.570 85.935 129.890 86.255 ;
        RECT 129.570 85.535 129.890 85.855 ;
        RECT 129.570 85.135 129.890 85.455 ;
        RECT 129.570 84.735 129.890 85.055 ;
        RECT 129.570 84.335 129.890 84.655 ;
        RECT 129.570 83.935 129.890 84.255 ;
        RECT 129.570 83.535 129.890 83.855 ;
        RECT 129.570 83.135 129.890 83.455 ;
        RECT 129.570 82.735 129.890 83.055 ;
        RECT 129.570 82.335 129.890 82.655 ;
        RECT 129.570 81.935 129.890 82.255 ;
        RECT 129.570 81.535 129.890 81.855 ;
        RECT 129.570 81.135 129.890 81.455 ;
        RECT 129.570 80.735 129.890 81.055 ;
        RECT 129.570 80.335 129.890 80.655 ;
        RECT 129.570 79.935 129.890 80.255 ;
        RECT 129.570 79.535 129.890 79.855 ;
        RECT 129.570 79.135 129.890 79.455 ;
        RECT 129.570 78.735 129.890 79.055 ;
        RECT 129.570 78.335 129.890 78.655 ;
        RECT 129.570 77.935 129.890 78.255 ;
        RECT 129.570 77.535 129.890 77.855 ;
        RECT 129.570 77.135 129.890 77.455 ;
        RECT 129.570 76.735 129.890 77.055 ;
        RECT 129.570 76.335 129.890 76.655 ;
        RECT 129.570 75.935 129.890 76.255 ;
        RECT 129.570 75.535 129.890 75.855 ;
        RECT 129.570 75.135 129.890 75.455 ;
        RECT 129.570 74.735 129.890 75.055 ;
        RECT 129.570 74.335 129.890 74.655 ;
        RECT 129.570 73.935 129.890 74.255 ;
        RECT 129.570 73.535 129.890 73.855 ;
        RECT 129.570 73.135 129.890 73.455 ;
        RECT 129.570 72.735 129.890 73.055 ;
        RECT 129.570 72.335 129.890 72.655 ;
        RECT 129.570 71.935 129.890 72.255 ;
        RECT 129.570 71.535 129.890 71.855 ;
        RECT 129.570 71.135 129.890 71.455 ;
        RECT 129.570 70.735 129.890 71.055 ;
        RECT 129.570 70.335 129.890 70.655 ;
        RECT 129.570 69.935 129.890 70.255 ;
        RECT 129.570 69.535 129.890 69.855 ;
        RECT 129.570 69.135 129.890 69.455 ;
        RECT 129.570 68.735 129.890 69.055 ;
        RECT 129.570 68.335 129.890 68.655 ;
        RECT 129.570 67.935 129.890 68.255 ;
        RECT 129.570 67.535 129.890 67.855 ;
        RECT 129.570 67.135 129.890 67.455 ;
        RECT 129.570 66.735 129.890 67.055 ;
        RECT 129.570 66.335 129.890 66.655 ;
        RECT 129.570 65.935 129.890 66.255 ;
        RECT 129.570 65.535 129.890 65.855 ;
        RECT 129.570 65.135 129.890 65.455 ;
        RECT 129.570 64.735 129.890 65.055 ;
        RECT 129.570 64.335 129.890 64.655 ;
        RECT 129.570 63.935 129.890 64.255 ;
        RECT 129.570 62.135 129.890 62.455 ;
        RECT 129.570 61.735 129.890 62.055 ;
        RECT 129.570 61.335 129.890 61.655 ;
        RECT 129.570 60.935 129.890 61.255 ;
        RECT 129.570 60.535 129.890 60.855 ;
        RECT 129.570 60.135 129.890 60.455 ;
        RECT 129.570 59.735 129.890 60.055 ;
        RECT 129.570 59.335 129.890 59.655 ;
        RECT 129.570 58.935 129.890 59.255 ;
        RECT 129.570 58.535 129.890 58.855 ;
        RECT 129.570 58.135 129.890 58.455 ;
        RECT 129.570 57.735 129.890 58.055 ;
        RECT 129.570 57.335 129.890 57.655 ;
        RECT 129.570 56.935 129.890 57.255 ;
        RECT 129.570 56.535 129.890 56.855 ;
        RECT 129.570 56.135 129.890 56.455 ;
        RECT 129.570 55.735 129.890 56.055 ;
        RECT 129.570 55.335 129.890 55.655 ;
        RECT 129.570 54.935 129.890 55.255 ;
        RECT 129.570 54.535 129.890 54.855 ;
        RECT 129.570 54.135 129.890 54.455 ;
        RECT 129.570 53.735 129.890 54.055 ;
        RECT 129.570 53.335 129.890 53.655 ;
        RECT 129.570 52.935 129.890 53.255 ;
        RECT 129.570 52.535 129.890 52.855 ;
        RECT 129.570 52.135 129.890 52.455 ;
        RECT 129.570 51.735 129.890 52.055 ;
        RECT 129.570 51.335 129.890 51.655 ;
        RECT 129.570 50.935 129.890 51.255 ;
        RECT 129.570 50.535 129.890 50.855 ;
        RECT 129.570 50.135 129.890 50.455 ;
        RECT 129.570 49.735 129.890 50.055 ;
        RECT 129.570 49.335 129.890 49.655 ;
        RECT 129.570 48.935 129.890 49.255 ;
        RECT 129.570 48.535 129.890 48.855 ;
        RECT 129.570 48.135 129.890 48.455 ;
        RECT 129.570 47.735 129.890 48.055 ;
        RECT 129.570 47.335 129.890 47.655 ;
        RECT 129.570 46.935 129.890 47.255 ;
        RECT 129.570 46.535 129.890 46.855 ;
        RECT 129.570 46.135 129.890 46.455 ;
        RECT 129.570 45.735 129.890 46.055 ;
        RECT 129.570 45.335 129.890 45.655 ;
        RECT 129.570 44.935 129.890 45.255 ;
        RECT 129.570 44.535 129.890 44.855 ;
        RECT 129.570 44.135 129.890 44.455 ;
        RECT 129.570 43.735 129.890 44.055 ;
        RECT 129.570 43.335 129.890 43.655 ;
        RECT 129.570 42.935 129.890 43.255 ;
        RECT 129.570 42.535 129.890 42.855 ;
        RECT 129.570 42.135 129.890 42.455 ;
        RECT 129.570 41.735 129.890 42.055 ;
        RECT 129.570 41.335 129.890 41.655 ;
        RECT 129.570 40.935 129.890 41.255 ;
        RECT 129.570 40.535 129.890 40.855 ;
        RECT 129.570 40.135 129.890 40.455 ;
        RECT 140.605 38.335 140.925 38.655 ;
        RECT 141.005 38.335 141.325 38.655 ;
        RECT 141.405 38.335 141.725 38.655 ;
        RECT 141.805 38.335 142.125 38.655 ;
        RECT 142.205 38.335 142.525 38.655 ;
        RECT 129.570 36.535 129.890 36.855 ;
        RECT 129.570 36.135 129.890 36.455 ;
        RECT 129.570 35.735 129.890 36.055 ;
        RECT 129.570 35.335 129.890 35.655 ;
        RECT 129.570 34.935 129.890 35.255 ;
        RECT 129.570 34.535 129.890 34.855 ;
        RECT 129.570 34.135 129.890 34.455 ;
        RECT 129.570 33.735 129.890 34.055 ;
        RECT 129.570 33.335 129.890 33.655 ;
        RECT 129.570 32.935 129.890 33.255 ;
        RECT 129.570 32.535 129.890 32.855 ;
        RECT 129.570 32.135 129.890 32.455 ;
        RECT 129.570 31.735 129.890 32.055 ;
        RECT 129.570 31.335 129.890 31.655 ;
        RECT 129.570 30.935 129.890 31.255 ;
        RECT 129.570 30.535 129.890 30.855 ;
        RECT 129.570 30.135 129.890 30.455 ;
        RECT 129.570 29.735 129.890 30.055 ;
        RECT 129.570 29.335 129.890 29.655 ;
        RECT 129.570 28.935 129.890 29.255 ;
        RECT 129.570 28.535 129.890 28.855 ;
        RECT 129.570 28.135 129.890 28.455 ;
        RECT 129.570 27.735 129.890 28.055 ;
        RECT 129.570 27.335 129.890 27.655 ;
        RECT 129.570 26.935 129.890 27.255 ;
        RECT 129.570 26.535 129.890 26.855 ;
        RECT 129.570 26.135 129.890 26.455 ;
        RECT 129.570 25.735 129.890 26.055 ;
        RECT 129.570 25.335 129.890 25.655 ;
        RECT 129.570 24.935 129.890 25.255 ;
        RECT 129.570 24.535 129.890 24.855 ;
        RECT 129.570 24.135 129.890 24.455 ;
        RECT 129.570 23.735 129.890 24.055 ;
        RECT 129.570 23.335 129.890 23.655 ;
        RECT 129.570 22.935 129.890 23.255 ;
        RECT 129.570 22.535 129.890 22.855 ;
        RECT 129.570 22.135 129.890 22.455 ;
        RECT 129.570 21.735 129.890 22.055 ;
        RECT 129.570 21.335 129.890 21.655 ;
        RECT 129.570 20.935 129.890 21.255 ;
        RECT 129.570 20.535 129.890 20.855 ;
        RECT 129.570 20.135 129.890 20.455 ;
        RECT 129.570 19.735 129.890 20.055 ;
        RECT 129.570 19.335 129.890 19.655 ;
        RECT 129.570 18.935 129.890 19.255 ;
        RECT 129.570 18.535 129.890 18.855 ;
        RECT 129.570 18.135 129.890 18.455 ;
        RECT 129.570 17.735 129.890 18.055 ;
        RECT 129.570 17.335 129.890 17.655 ;
        RECT 129.570 16.935 129.890 17.255 ;
        RECT 129.570 16.535 129.890 16.855 ;
        RECT 129.570 16.135 129.890 16.455 ;
        RECT 129.570 15.735 129.890 16.055 ;
        RECT 129.570 15.335 129.890 15.655 ;
        RECT 129.570 14.935 129.890 15.255 ;
        RECT 129.570 14.535 129.890 14.855 ;
        RECT 140.605 12.735 140.925 13.055 ;
        RECT 141.005 12.735 141.325 13.055 ;
        RECT 141.405 12.735 141.725 13.055 ;
        RECT 141.805 12.735 142.125 13.055 ;
        RECT 142.205 12.735 142.525 13.055 ;
        RECT 111.875 7.390 112.195 7.710 ;
        RECT 112.275 7.390 112.595 7.710 ;
        RECT 112.675 7.390 112.995 7.710 ;
        RECT 89.795 6.290 90.115 6.610 ;
        RECT 90.195 6.290 90.515 6.610 ;
        RECT 90.595 6.290 90.915 6.610 ;
        RECT 134.485 3.970 134.805 4.290 ;
        RECT 134.885 3.970 135.205 4.290 ;
        RECT 135.285 3.970 135.605 4.290 ;
        RECT 135.685 3.970 136.005 4.290 ;
        RECT 90.460 3.175 90.780 3.495 ;
        RECT 90.460 2.775 90.780 3.095 ;
        RECT 90.460 2.375 90.780 2.695 ;
        RECT 90.460 1.975 90.780 2.295 ;
        RECT 90.460 1.575 90.780 1.895 ;
        RECT 112.540 3.175 112.860 3.495 ;
        RECT 112.540 2.775 112.860 3.095 ;
        RECT 112.540 2.375 112.860 2.695 ;
        RECT 112.540 1.975 112.860 2.295 ;
        RECT 112.540 1.575 112.860 1.895 ;
        RECT 134.620 3.175 134.940 3.495 ;
        RECT 134.620 2.775 134.940 3.095 ;
        RECT 134.620 2.375 134.940 2.695 ;
        RECT 134.620 1.975 134.940 2.295 ;
        RECT 134.620 1.575 134.940 1.895 ;
        RECT 156.705 3.175 157.025 3.495 ;
        RECT 156.705 2.775 157.025 3.095 ;
        RECT 156.705 2.375 157.025 2.695 ;
        RECT 156.705 1.975 157.025 2.295 ;
        RECT 156.705 1.575 157.025 1.895 ;
      LAYER met4 ;
        RECT 144.130 224.760 144.135 225.405 ;
        RECT 3.990 220.515 4.290 224.760 ;
        RECT 7.670 220.515 7.970 224.760 ;
        RECT 11.350 220.515 11.650 224.760 ;
        RECT 15.030 220.515 15.330 224.760 ;
        RECT 18.710 220.515 19.010 224.760 ;
        RECT 22.390 220.515 22.690 224.760 ;
        RECT 26.070 220.515 26.370 224.760 ;
        RECT 29.750 220.515 30.050 224.760 ;
        RECT 33.430 220.515 33.730 224.760 ;
        RECT 37.110 220.515 37.410 224.760 ;
        RECT 40.790 220.515 41.090 224.760 ;
        RECT 44.470 220.515 44.770 224.760 ;
        RECT 48.150 220.515 48.450 224.760 ;
        RECT 51.830 220.515 52.130 224.760 ;
        RECT 55.510 220.515 55.810 224.760 ;
        RECT 59.190 220.515 59.490 224.760 ;
        RECT 62.870 220.515 63.170 224.760 ;
        RECT 66.550 220.515 66.850 224.760 ;
        RECT 70.230 220.515 70.530 224.760 ;
        RECT 73.910 220.515 74.210 224.760 ;
        RECT 77.590 220.515 77.890 224.760 ;
        RECT 81.270 220.515 81.570 224.760 ;
        RECT 3.975 219.015 4.305 220.515 ;
        RECT 7.655 219.015 7.985 220.515 ;
        RECT 11.335 219.015 11.665 220.515 ;
        RECT 15.015 219.015 15.345 220.515 ;
        RECT 18.695 219.015 19.025 220.515 ;
        RECT 22.375 219.015 22.705 220.515 ;
        RECT 26.055 219.015 26.385 220.515 ;
        RECT 29.735 219.015 30.065 220.515 ;
        RECT 33.415 219.015 33.745 220.515 ;
        RECT 37.095 219.015 37.425 220.515 ;
        RECT 40.775 219.015 41.105 220.515 ;
        RECT 44.455 219.015 44.785 220.515 ;
        RECT 48.135 219.015 48.465 220.515 ;
        RECT 51.815 219.015 52.145 220.515 ;
        RECT 55.495 219.015 55.825 220.515 ;
        RECT 59.175 219.015 59.505 220.515 ;
        RECT 62.855 219.015 63.185 220.515 ;
        RECT 66.535 219.015 66.865 220.515 ;
        RECT 70.215 219.015 70.545 220.515 ;
        RECT 73.895 219.015 74.225 220.515 ;
        RECT 77.575 219.015 77.905 220.515 ;
        RECT 81.255 219.015 81.585 220.515 ;
        RECT 84.950 174.600 85.250 224.760 ;
        RECT 84.935 173.470 85.265 174.600 ;
        RECT 88.630 173.500 88.930 224.760 ;
        RECT 143.835 212.280 144.135 224.760 ;
        RECT 143.005 211.950 144.135 212.280 ;
        RECT 147.510 210.620 147.810 224.760 ;
        RECT 146.680 210.290 147.810 210.620 ;
        RECT 140.600 208.090 142.530 208.690 ;
        RECT 129.490 206.810 129.970 206.830 ;
        RECT 88.615 172.370 88.945 173.500 ;
        RECT 129.470 163.185 130.070 206.810 ;
        RECT 141.930 206.495 142.530 208.090 ;
        RECT 131.325 184.685 153.135 206.495 ;
        RECT 141.930 184.525 142.530 184.685 ;
        RECT 141.930 181.200 142.530 181.270 ;
        RECT 50.500 161.185 130.070 163.185 ;
        RECT 52.500 149.185 127.725 151.185 ;
        RECT 129.470 139.185 130.070 161.185 ;
        RECT 131.325 159.390 153.135 181.200 ;
        RECT 141.930 157.400 142.530 159.390 ;
        RECT 50.500 137.185 130.070 139.185 ;
        RECT 52.500 125.185 127.725 127.185 ;
        RECT 129.470 115.185 130.070 137.185 ;
        RECT 131.325 135.590 153.135 157.400 ;
        RECT 141.930 133.600 142.530 135.590 ;
        RECT 50.500 113.185 130.070 115.185 ;
        RECT 52.500 101.185 127.725 103.185 ;
        RECT 129.470 91.185 130.070 113.185 ;
        RECT 131.325 111.790 153.135 133.600 ;
        RECT 141.930 109.800 142.530 111.790 ;
        RECT 50.500 89.185 130.070 91.185 ;
        RECT 71.350 81.610 87.210 82.610 ;
        RECT 52.500 77.185 127.725 79.185 ;
        RECT 129.470 67.185 130.070 89.185 ;
        RECT 131.325 87.990 153.135 109.800 ;
        RECT 141.930 86.000 142.530 87.990 ;
        RECT 50.500 65.185 130.070 67.185 ;
        RECT 129.470 14.395 130.070 65.185 ;
        RECT 131.325 64.190 153.135 86.000 ;
        RECT 141.930 62.200 142.530 64.190 ;
        RECT 131.325 40.390 153.135 62.200 ;
        RECT 141.930 38.795 142.530 40.390 ;
        RECT 140.600 38.195 142.530 38.795 ;
        RECT 141.930 36.600 142.530 36.795 ;
        RECT 131.325 14.790 153.135 36.600 ;
        RECT 141.930 13.195 142.530 14.790 ;
        RECT 140.600 12.595 142.530 13.195 ;
        RECT 111.870 7.250 113.000 7.850 ;
        RECT 89.790 6.150 90.920 6.750 ;
        RECT 90.320 1.000 90.920 6.150 ;
        RECT 112.400 1.000 113.000 7.250 ;
        RECT 134.480 3.830 136.010 4.430 ;
        RECT 134.480 1.000 135.080 3.830 ;
        RECT 156.565 1.000 157.165 3.505 ;
  END
END tt_um_lcasimon_tdc
END LIBRARY

