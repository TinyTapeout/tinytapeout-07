VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_twin_tee_opamp_osc
  CLASS BLOCK ;
  FOREIGN tt_um_twin_tee_opamp_osc ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.060000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 32.495098 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 130.110 94.370 142.570 99.700 ;
        RECT 111.250 88.080 123.710 93.410 ;
        RECT 113.870 48.000 142.850 50.010 ;
        RECT 114.200 15.650 116.210 41.630 ;
        RECT 118.250 15.850 120.260 41.830 ;
        RECT 126.150 34.000 128.160 42.880 ;
        RECT 125.600 22.350 128.700 33.180 ;
      LAYER nwell ;
        RECT 130.200 28.400 133.390 43.810 ;
        RECT 136.550 28.400 139.740 43.810 ;
      LAYER pwell ;
        RECT 130.350 25.550 139.550 28.010 ;
      LAYER nwell ;
        RECT 141.150 26.600 144.340 44.070 ;
      LAYER pwell ;
        RECT 137.150 25.500 137.700 25.550 ;
        RECT 129.650 22.400 140.480 25.500 ;
        RECT 145.150 22.400 148.250 40.100 ;
      LAYER li1 ;
        RECT 130.290 99.350 142.390 99.520 ;
        RECT 130.290 94.720 130.460 99.350 ;
        RECT 130.940 98.520 133.100 98.870 ;
        RECT 139.580 95.200 141.740 95.550 ;
        RECT 142.220 94.720 142.390 99.350 ;
        RECT 130.290 94.550 142.390 94.720 ;
        RECT 111.430 93.060 123.530 93.230 ;
        RECT 111.430 88.430 111.600 93.060 ;
        RECT 112.080 92.230 114.240 92.580 ;
        RECT 120.720 88.910 122.880 89.260 ;
        RECT 123.360 88.430 123.530 93.060 ;
        RECT 111.430 88.260 123.530 88.430 ;
        RECT 105.310 83.690 107.600 86.540 ;
        RECT 114.050 49.660 142.670 49.830 ;
        RECT 114.050 48.350 114.220 49.660 ;
        RECT 114.700 48.830 116.860 49.180 ;
        RECT 139.860 48.830 142.020 49.180 ;
        RECT 142.500 48.350 142.670 49.660 ;
        RECT 114.050 48.180 142.670 48.350 ;
        RECT 141.330 43.720 144.160 43.890 ;
        RECT 130.380 43.460 133.210 43.630 ;
        RECT 130.380 43.100 130.550 43.460 ;
        RECT 126.330 42.530 127.980 42.700 ;
        RECT 126.330 42.400 126.500 42.530 ;
        RECT 118.430 41.480 120.080 41.650 ;
        RECT 114.380 41.280 116.030 41.450 ;
        RECT 114.380 16.000 114.550 41.280 ;
        RECT 115.030 38.640 115.380 40.800 ;
        RECT 115.030 16.480 115.380 18.640 ;
        RECT 115.860 16.000 116.030 41.280 ;
        RECT 118.430 16.200 118.600 41.480 ;
        RECT 119.080 38.840 119.430 41.000 ;
        RECT 119.080 16.680 119.430 18.840 ;
        RECT 119.910 16.200 120.080 41.480 ;
        RECT 124.500 34.350 126.500 42.400 ;
        RECT 126.980 39.890 127.330 42.050 ;
        RECT 126.980 34.830 127.330 36.990 ;
        RECT 127.810 34.350 127.980 42.530 ;
        RECT 124.500 34.180 127.980 34.350 ;
        RECT 124.500 33.000 127.650 34.180 ;
        RECT 124.500 32.830 128.520 33.000 ;
        RECT 124.500 22.700 125.950 32.830 ;
        RECT 126.630 32.260 127.670 32.430 ;
        RECT 126.290 30.200 126.460 32.200 ;
        RECT 127.840 30.200 128.010 32.200 ;
        RECT 126.630 29.970 127.670 30.140 ;
        RECT 126.290 27.910 126.460 29.910 ;
        RECT 127.840 27.910 128.010 29.910 ;
        RECT 126.630 27.680 127.670 27.850 ;
        RECT 126.290 25.620 126.460 27.620 ;
        RECT 127.840 25.620 128.010 27.620 ;
        RECT 126.630 25.390 127.670 25.560 ;
        RECT 126.290 23.330 126.460 25.330 ;
        RECT 127.840 23.330 128.010 25.330 ;
        RECT 128.350 25.000 128.520 32.830 ;
        RECT 130.250 31.200 130.550 43.100 ;
        RECT 131.275 42.890 132.315 43.060 ;
        RECT 130.890 40.830 131.060 42.830 ;
        RECT 132.530 40.830 132.700 42.830 ;
        RECT 131.275 40.600 132.315 40.770 ;
        RECT 130.890 38.540 131.060 40.540 ;
        RECT 132.530 38.540 132.700 40.540 ;
        RECT 131.275 38.310 132.315 38.480 ;
        RECT 130.890 36.250 131.060 38.250 ;
        RECT 132.530 36.250 132.700 38.250 ;
        RECT 131.275 36.020 132.315 36.190 ;
        RECT 130.890 33.960 131.060 35.960 ;
        RECT 132.530 33.960 132.700 35.960 ;
        RECT 131.275 33.730 132.315 33.900 ;
        RECT 130.890 31.670 131.060 33.670 ;
        RECT 132.530 31.670 132.700 33.670 ;
        RECT 131.275 31.440 132.315 31.610 ;
        RECT 130.380 28.750 130.550 31.200 ;
        RECT 130.890 29.380 131.060 31.380 ;
        RECT 132.530 29.380 132.700 31.380 ;
        RECT 131.275 29.150 132.315 29.320 ;
        RECT 133.040 28.750 133.210 43.460 ;
        RECT 130.380 28.580 133.210 28.750 ;
        RECT 136.730 43.460 139.560 43.630 ;
        RECT 136.730 28.750 136.900 43.460 ;
        RECT 139.390 43.100 139.560 43.460 ;
        RECT 141.330 43.350 141.500 43.720 ;
        RECT 137.625 42.890 138.665 43.060 ;
        RECT 137.240 40.830 137.410 42.830 ;
        RECT 138.880 40.830 139.050 42.830 ;
        RECT 137.625 40.600 138.665 40.770 ;
        RECT 137.240 38.540 137.410 40.540 ;
        RECT 138.880 38.540 139.050 40.540 ;
        RECT 137.625 38.310 138.665 38.480 ;
        RECT 137.240 36.250 137.410 38.250 ;
        RECT 138.880 36.250 139.050 38.250 ;
        RECT 137.625 36.020 138.665 36.190 ;
        RECT 137.240 33.960 137.410 35.960 ;
        RECT 138.880 33.960 139.050 35.960 ;
        RECT 137.625 33.730 138.665 33.900 ;
        RECT 137.240 31.670 137.410 33.670 ;
        RECT 138.880 31.670 139.050 33.670 ;
        RECT 137.625 31.440 138.665 31.610 ;
        RECT 137.240 29.380 137.410 31.380 ;
        RECT 138.880 29.380 139.050 31.380 ;
        RECT 139.390 31.200 139.700 43.100 ;
        RECT 137.625 29.150 138.665 29.320 ;
        RECT 139.390 28.750 139.560 31.200 ;
        RECT 136.730 28.580 139.560 28.750 ;
        RECT 130.530 27.660 134.770 27.830 ;
        RECT 130.530 25.900 130.700 27.660 ;
        RECT 131.380 27.090 133.920 27.260 ;
        RECT 131.040 26.530 131.210 27.030 ;
        RECT 134.090 26.530 134.260 27.030 ;
        RECT 131.380 26.300 133.920 26.470 ;
        RECT 134.600 25.900 134.770 27.660 ;
        RECT 130.530 25.730 134.770 25.900 ;
        RECT 135.130 27.660 139.370 27.830 ;
        RECT 141.300 27.800 141.500 43.350 ;
        RECT 142.225 43.150 143.265 43.320 ;
        RECT 141.840 42.590 142.010 43.090 ;
        RECT 143.480 42.590 143.650 43.090 ;
        RECT 142.225 42.360 143.265 42.530 ;
        RECT 141.840 41.800 142.010 42.300 ;
        RECT 143.480 41.800 143.650 42.300 ;
        RECT 142.225 41.570 143.265 41.740 ;
        RECT 141.840 41.010 142.010 41.510 ;
        RECT 143.480 41.010 143.650 41.510 ;
        RECT 142.225 40.780 143.265 40.950 ;
        RECT 141.840 40.220 142.010 40.720 ;
        RECT 143.480 40.220 143.650 40.720 ;
        RECT 142.225 39.990 143.265 40.160 ;
        RECT 141.840 39.430 142.010 39.930 ;
        RECT 143.480 39.430 143.650 39.930 ;
        RECT 142.225 39.200 143.265 39.370 ;
        RECT 141.840 38.640 142.010 39.140 ;
        RECT 143.480 38.640 143.650 39.140 ;
        RECT 142.225 38.410 143.265 38.580 ;
        RECT 141.840 37.850 142.010 38.350 ;
        RECT 143.480 37.850 143.650 38.350 ;
        RECT 142.225 37.620 143.265 37.790 ;
        RECT 141.840 37.060 142.010 37.560 ;
        RECT 143.480 37.060 143.650 37.560 ;
        RECT 142.225 36.830 143.265 37.000 ;
        RECT 141.840 36.270 142.010 36.770 ;
        RECT 143.480 36.270 143.650 36.770 ;
        RECT 142.225 36.040 143.265 36.210 ;
        RECT 141.840 35.480 142.010 35.980 ;
        RECT 143.480 35.480 143.650 35.980 ;
        RECT 142.225 35.250 143.265 35.420 ;
        RECT 141.840 34.690 142.010 35.190 ;
        RECT 143.480 34.690 143.650 35.190 ;
        RECT 142.225 34.460 143.265 34.630 ;
        RECT 141.840 33.900 142.010 34.400 ;
        RECT 143.480 33.900 143.650 34.400 ;
        RECT 142.225 33.670 143.265 33.840 ;
        RECT 141.840 33.110 142.010 33.610 ;
        RECT 143.480 33.110 143.650 33.610 ;
        RECT 142.225 32.880 143.265 33.050 ;
        RECT 141.840 32.320 142.010 32.820 ;
        RECT 143.480 32.320 143.650 32.820 ;
        RECT 142.225 32.090 143.265 32.260 ;
        RECT 141.840 31.530 142.010 32.030 ;
        RECT 143.480 31.530 143.650 32.030 ;
        RECT 142.225 31.300 143.265 31.470 ;
        RECT 141.840 30.740 142.010 31.240 ;
        RECT 143.480 30.740 143.650 31.240 ;
        RECT 142.225 30.510 143.265 30.680 ;
        RECT 141.840 29.950 142.010 30.450 ;
        RECT 143.480 29.950 143.650 30.450 ;
        RECT 142.225 29.720 143.265 29.890 ;
        RECT 141.840 29.160 142.010 29.660 ;
        RECT 143.480 29.160 143.650 29.660 ;
        RECT 142.225 28.930 143.265 29.100 ;
        RECT 141.840 28.370 142.010 28.870 ;
        RECT 143.480 28.370 143.650 28.870 ;
        RECT 142.225 28.140 143.265 28.310 ;
        RECT 135.130 25.900 135.300 27.660 ;
        RECT 135.980 27.090 138.520 27.260 ;
        RECT 135.640 26.530 135.810 27.030 ;
        RECT 138.690 26.530 138.860 27.030 ;
        RECT 135.980 26.300 138.520 26.470 ;
        RECT 139.200 25.900 139.370 27.660 ;
        RECT 141.330 26.950 141.500 27.800 ;
        RECT 141.840 27.580 142.010 28.080 ;
        RECT 143.480 27.580 143.650 28.080 ;
        RECT 142.225 27.350 143.265 27.520 ;
        RECT 143.990 26.950 144.160 43.720 ;
        RECT 141.330 26.780 144.160 26.950 ;
        RECT 145.330 39.750 148.070 39.920 ;
        RECT 135.130 25.730 139.500 25.900 ;
        RECT 130.550 25.700 131.350 25.730 ;
        RECT 138.700 25.700 139.500 25.730 ;
        RECT 129.830 25.250 140.300 25.320 ;
        RECT 145.330 25.250 145.500 39.750 ;
        RECT 146.180 39.180 147.220 39.350 ;
        RECT 145.840 37.120 146.010 39.120 ;
        RECT 147.390 37.120 147.560 39.120 ;
        RECT 146.180 36.890 147.220 37.060 ;
        RECT 147.900 37.050 148.070 39.750 ;
        RECT 145.840 34.830 146.010 36.830 ;
        RECT 147.390 34.830 147.560 36.830 ;
        RECT 146.180 34.600 147.220 34.770 ;
        RECT 145.840 32.540 146.010 34.540 ;
        RECT 147.390 32.540 147.560 34.540 ;
        RECT 146.180 32.310 147.220 32.480 ;
        RECT 145.840 30.250 146.010 32.250 ;
        RECT 147.390 30.250 147.560 32.250 ;
        RECT 146.180 30.020 147.220 30.190 ;
        RECT 145.840 27.960 146.010 29.960 ;
        RECT 147.390 27.960 147.560 29.960 ;
        RECT 146.180 27.730 147.220 27.900 ;
        RECT 145.840 25.670 146.010 27.670 ;
        RECT 147.390 25.670 147.560 27.670 ;
        RECT 146.180 25.440 147.220 25.610 ;
        RECT 129.830 25.150 145.500 25.250 ;
        RECT 129.830 25.000 130.000 25.150 ;
        RECT 126.630 23.100 127.670 23.270 ;
        RECT 128.350 22.750 130.000 25.000 ;
        RECT 130.630 24.640 132.630 24.810 ;
        RECT 132.920 24.640 134.920 24.810 ;
        RECT 135.210 24.640 137.210 24.810 ;
        RECT 137.500 24.640 139.500 24.810 ;
        RECT 140.130 24.650 145.500 25.150 ;
        RECT 130.400 23.430 130.570 24.470 ;
        RECT 132.690 23.430 132.860 24.470 ;
        RECT 134.980 23.430 135.150 24.470 ;
        RECT 137.270 23.430 137.440 24.470 ;
        RECT 139.560 23.430 139.730 24.470 ;
        RECT 130.630 23.090 132.630 23.260 ;
        RECT 132.920 23.090 134.920 23.260 ;
        RECT 135.210 23.090 137.210 23.260 ;
        RECT 137.500 23.090 139.500 23.260 ;
        RECT 140.100 23.050 145.500 24.650 ;
        RECT 145.840 23.380 146.010 25.380 ;
        RECT 147.390 23.380 147.560 25.380 ;
        RECT 146.180 23.150 147.220 23.320 ;
        RECT 140.130 22.750 145.500 23.050 ;
        RECT 147.900 22.750 148.650 37.050 ;
        RECT 126.200 22.700 128.100 22.750 ;
        RECT 128.350 22.700 148.650 22.750 ;
        RECT 124.500 20.500 148.650 22.700 ;
        RECT 118.430 16.030 120.080 16.200 ;
        RECT 114.380 15.830 116.030 16.000 ;
      LAYER mcon ;
        RECT 105.310 84.070 107.600 86.060 ;
        RECT 114.790 48.910 116.775 49.100 ;
        RECT 139.945 48.910 141.930 49.100 ;
        RECT 115.110 38.725 115.300 40.710 ;
        RECT 115.110 16.570 115.300 18.555 ;
        RECT 119.160 38.925 119.350 40.910 ;
        RECT 119.160 16.770 119.350 18.755 ;
        RECT 125.000 38.100 125.850 41.800 ;
        RECT 126.250 34.800 126.500 41.950 ;
        RECT 127.060 39.975 127.250 41.960 ;
        RECT 127.060 34.920 127.250 36.905 ;
        RECT 125.700 23.550 125.950 32.900 ;
        RECT 126.710 32.260 127.590 32.430 ;
        RECT 126.290 30.280 126.460 32.120 ;
        RECT 127.840 30.280 128.010 32.120 ;
        RECT 126.710 29.970 127.590 30.140 ;
        RECT 126.290 27.990 126.460 29.830 ;
        RECT 127.840 27.990 128.010 29.830 ;
        RECT 126.710 27.680 127.590 27.850 ;
        RECT 126.290 25.700 126.460 27.540 ;
        RECT 127.840 25.700 128.010 27.540 ;
        RECT 126.710 25.390 127.590 25.560 ;
        RECT 126.290 23.410 126.460 25.250 ;
        RECT 127.840 23.410 128.010 25.250 ;
        RECT 130.250 31.200 130.550 43.100 ;
        RECT 131.355 42.890 132.235 43.060 ;
        RECT 130.890 40.910 131.060 42.750 ;
        RECT 132.530 40.910 132.700 42.750 ;
        RECT 131.355 40.600 132.235 40.770 ;
        RECT 130.890 38.620 131.060 40.460 ;
        RECT 132.530 38.620 132.700 40.460 ;
        RECT 131.355 38.310 132.235 38.480 ;
        RECT 130.890 36.330 131.060 38.170 ;
        RECT 132.530 36.330 132.700 38.170 ;
        RECT 131.355 36.020 132.235 36.190 ;
        RECT 130.890 34.040 131.060 35.880 ;
        RECT 132.530 34.040 132.700 35.880 ;
        RECT 131.355 33.730 132.235 33.900 ;
        RECT 130.890 31.750 131.060 33.590 ;
        RECT 132.530 31.750 132.700 33.590 ;
        RECT 131.355 31.440 132.235 31.610 ;
        RECT 130.890 29.460 131.060 31.300 ;
        RECT 132.530 29.460 132.700 31.300 ;
        RECT 131.355 29.150 132.235 29.320 ;
        RECT 137.705 42.890 138.585 43.060 ;
        RECT 137.240 40.910 137.410 42.750 ;
        RECT 138.880 40.910 139.050 42.750 ;
        RECT 137.705 40.600 138.585 40.770 ;
        RECT 137.240 38.620 137.410 40.460 ;
        RECT 138.880 38.620 139.050 40.460 ;
        RECT 137.705 38.310 138.585 38.480 ;
        RECT 137.240 36.330 137.410 38.170 ;
        RECT 138.880 36.330 139.050 38.170 ;
        RECT 137.705 36.020 138.585 36.190 ;
        RECT 137.240 34.040 137.410 35.880 ;
        RECT 138.880 34.040 139.050 35.880 ;
        RECT 137.705 33.730 138.585 33.900 ;
        RECT 137.240 31.750 137.410 33.590 ;
        RECT 138.880 31.750 139.050 33.590 ;
        RECT 137.705 31.440 138.585 31.610 ;
        RECT 137.240 29.460 137.410 31.300 ;
        RECT 138.880 29.460 139.050 31.300 ;
        RECT 139.400 31.200 139.700 43.100 ;
        RECT 137.705 29.150 138.585 29.320 ;
        RECT 131.460 27.090 133.840 27.260 ;
        RECT 131.040 26.610 131.210 26.950 ;
        RECT 134.090 26.610 134.260 26.950 ;
        RECT 131.460 26.300 133.840 26.470 ;
        RECT 141.300 27.800 141.500 43.350 ;
        RECT 142.305 43.150 143.185 43.320 ;
        RECT 141.840 42.670 142.010 43.010 ;
        RECT 143.480 42.670 143.650 43.010 ;
        RECT 142.305 42.360 143.185 42.530 ;
        RECT 141.840 41.880 142.010 42.220 ;
        RECT 143.480 41.880 143.650 42.220 ;
        RECT 142.305 41.570 143.185 41.740 ;
        RECT 141.840 41.090 142.010 41.430 ;
        RECT 143.480 41.090 143.650 41.430 ;
        RECT 142.305 40.780 143.185 40.950 ;
        RECT 141.840 40.300 142.010 40.640 ;
        RECT 143.480 40.300 143.650 40.640 ;
        RECT 142.305 39.990 143.185 40.160 ;
        RECT 141.840 39.510 142.010 39.850 ;
        RECT 143.480 39.510 143.650 39.850 ;
        RECT 142.305 39.200 143.185 39.370 ;
        RECT 141.840 38.720 142.010 39.060 ;
        RECT 143.480 38.720 143.650 39.060 ;
        RECT 142.305 38.410 143.185 38.580 ;
        RECT 141.840 37.930 142.010 38.270 ;
        RECT 143.480 37.930 143.650 38.270 ;
        RECT 142.305 37.620 143.185 37.790 ;
        RECT 141.840 37.140 142.010 37.480 ;
        RECT 143.480 37.140 143.650 37.480 ;
        RECT 142.305 36.830 143.185 37.000 ;
        RECT 141.840 36.350 142.010 36.690 ;
        RECT 143.480 36.350 143.650 36.690 ;
        RECT 142.305 36.040 143.185 36.210 ;
        RECT 141.840 35.560 142.010 35.900 ;
        RECT 143.480 35.560 143.650 35.900 ;
        RECT 142.305 35.250 143.185 35.420 ;
        RECT 141.840 34.770 142.010 35.110 ;
        RECT 143.480 34.770 143.650 35.110 ;
        RECT 142.305 34.460 143.185 34.630 ;
        RECT 141.840 33.980 142.010 34.320 ;
        RECT 143.480 33.980 143.650 34.320 ;
        RECT 142.305 33.670 143.185 33.840 ;
        RECT 141.840 33.190 142.010 33.530 ;
        RECT 143.480 33.190 143.650 33.530 ;
        RECT 142.305 32.880 143.185 33.050 ;
        RECT 141.840 32.400 142.010 32.740 ;
        RECT 143.480 32.400 143.650 32.740 ;
        RECT 142.305 32.090 143.185 32.260 ;
        RECT 141.840 31.610 142.010 31.950 ;
        RECT 143.480 31.610 143.650 31.950 ;
        RECT 142.305 31.300 143.185 31.470 ;
        RECT 141.840 30.820 142.010 31.160 ;
        RECT 143.480 30.820 143.650 31.160 ;
        RECT 142.305 30.510 143.185 30.680 ;
        RECT 141.840 30.030 142.010 30.370 ;
        RECT 143.480 30.030 143.650 30.370 ;
        RECT 142.305 29.720 143.185 29.890 ;
        RECT 141.840 29.240 142.010 29.580 ;
        RECT 143.480 29.240 143.650 29.580 ;
        RECT 142.305 28.930 143.185 29.100 ;
        RECT 141.840 28.450 142.010 28.790 ;
        RECT 143.480 28.450 143.650 28.790 ;
        RECT 142.305 28.140 143.185 28.310 ;
        RECT 136.060 27.090 138.440 27.260 ;
        RECT 135.640 26.610 135.810 26.950 ;
        RECT 138.690 26.610 138.860 26.950 ;
        RECT 136.060 26.300 138.440 26.470 ;
        RECT 141.840 27.660 142.010 28.000 ;
        RECT 143.480 27.660 143.650 28.000 ;
        RECT 142.305 27.350 143.185 27.520 ;
        RECT 146.260 39.180 147.140 39.350 ;
        RECT 145.840 37.200 146.010 39.040 ;
        RECT 147.390 37.200 147.560 39.040 ;
        RECT 146.260 36.890 147.140 37.060 ;
        RECT 145.840 34.910 146.010 36.750 ;
        RECT 147.390 34.910 147.560 36.750 ;
        RECT 146.260 34.600 147.140 34.770 ;
        RECT 145.840 32.620 146.010 34.460 ;
        RECT 147.390 32.620 147.560 34.460 ;
        RECT 146.260 32.310 147.140 32.480 ;
        RECT 145.840 30.330 146.010 32.170 ;
        RECT 147.390 30.330 147.560 32.170 ;
        RECT 146.260 30.020 147.140 30.190 ;
        RECT 145.840 28.040 146.010 29.880 ;
        RECT 147.390 28.040 147.560 29.880 ;
        RECT 146.260 27.730 147.140 27.900 ;
        RECT 145.840 25.750 146.010 27.590 ;
        RECT 147.390 25.750 147.560 27.590 ;
        RECT 146.260 25.440 147.140 25.610 ;
        RECT 126.710 23.100 127.590 23.270 ;
        RECT 130.710 24.640 132.550 24.810 ;
        RECT 133.000 24.640 134.840 24.810 ;
        RECT 135.290 24.640 137.130 24.810 ;
        RECT 137.580 24.640 139.420 24.810 ;
        RECT 130.400 23.510 130.570 24.390 ;
        RECT 132.690 23.510 132.860 24.390 ;
        RECT 134.980 23.510 135.150 24.390 ;
        RECT 137.270 23.510 137.440 24.390 ;
        RECT 139.560 23.510 139.730 24.390 ;
        RECT 130.710 23.090 132.550 23.260 ;
        RECT 133.000 23.090 134.840 23.260 ;
        RECT 135.290 23.090 137.130 23.260 ;
        RECT 137.580 23.090 139.420 23.260 ;
        RECT 145.250 23.050 145.500 24.200 ;
        RECT 145.840 23.460 146.010 25.300 ;
        RECT 147.390 23.460 147.560 25.300 ;
        RECT 146.260 23.150 147.140 23.320 ;
        RECT 147.900 23.050 148.150 24.200 ;
        RECT 126.200 22.450 128.100 22.750 ;
        RECT 130.300 22.500 139.850 22.750 ;
        RECT 145.600 22.550 147.800 22.750 ;
        RECT 127.800 20.800 146.750 21.350 ;
      LAYER met1 ;
        RECT 130.800 98.900 133.230 98.950 ;
        RECT 129.080 98.220 133.230 98.900 ;
        RECT 103.750 92.910 106.020 93.680 ;
        RECT 102.090 92.770 106.020 92.910 ;
        RECT 129.080 92.800 129.760 98.220 ;
        RECT 130.800 98.200 133.230 98.220 ;
        RECT 138.715 95.030 144.130 95.765 ;
        RECT 143.395 92.805 144.130 95.030 ;
        RECT 146.620 94.300 148.890 94.360 ;
        RECT 146.620 93.005 152.400 94.300 ;
        RECT 146.440 92.805 152.400 93.005 ;
        RECT 102.090 92.030 114.890 92.770 ;
        RECT 124.840 92.120 129.860 92.800 ;
        RECT 102.090 91.885 106.020 92.030 ;
        RECT 102.090 91.360 103.115 91.885 ;
        RECT 102.060 90.335 103.145 91.360 ;
        RECT 103.750 91.170 106.020 91.885 ;
        RECT 109.470 86.880 110.210 92.030 ;
        RECT 124.840 89.370 125.520 92.120 ;
        RECT 143.380 92.045 152.400 92.805 ;
        RECT 146.480 92.000 152.400 92.045 ;
        RECT 146.480 91.900 149.400 92.000 ;
        RECT 146.480 91.850 148.890 91.900 ;
        RECT 120.110 88.690 127.130 89.370 ;
        RECT 146.480 86.950 147.425 91.850 ;
        RECT 105.160 83.400 107.800 86.460 ;
        RECT 109.470 86.140 117.530 86.880 ;
        RECT 93.750 83.250 95.250 83.280 ;
        RECT 104.290 83.250 107.800 83.400 ;
        RECT 93.750 81.750 107.800 83.250 ;
        RECT 93.750 81.720 95.250 81.750 ;
        RECT 104.290 80.990 107.800 81.750 ;
        RECT 104.290 80.890 106.560 80.990 ;
        RECT 104.780 69.235 105.970 80.890 ;
        RECT 104.780 68.045 112.295 69.235 ;
        RECT 104.780 49.410 105.970 68.045 ;
        RECT 106.510 68.040 109.590 68.045 ;
        RECT 116.800 67.720 117.520 86.140 ;
        RECT 146.400 83.110 147.500 86.950 ;
        RECT 146.370 82.010 147.530 83.110 ;
        RECT 111.770 67.000 117.520 67.720 ;
        RECT 144.090 49.490 145.010 49.520 ;
        RECT 104.780 48.655 117.005 49.410 ;
        RECT 142.840 49.370 145.010 49.490 ;
        RECT 104.780 40.645 105.970 48.655 ;
        RECT 139.690 48.590 145.010 49.370 ;
        RECT 142.840 48.570 145.010 48.590 ;
        RECT 144.090 48.540 145.010 48.570 ;
        RECT 110.750 45.250 112.250 45.280 ;
        RECT 124.400 45.250 148.650 45.900 ;
        RECT 110.750 43.750 148.650 45.250 ;
        RECT 110.750 43.720 112.250 43.750 ;
        RECT 115.080 40.645 115.330 40.770 ;
        RECT 104.780 39.455 115.595 40.645 ;
        RECT 104.780 21.595 105.970 39.455 ;
        RECT 115.080 38.665 115.330 39.455 ;
        RECT 118.850 38.700 119.550 43.750 ;
        RECT 124.400 43.550 148.650 43.750 ;
        RECT 124.400 34.650 126.600 42.400 ;
        RECT 126.750 39.650 127.700 43.550 ;
        RECT 127.030 36.950 127.280 36.965 ;
        RECT 124.400 22.800 126.050 34.650 ;
        RECT 126.900 34.450 128.750 36.950 ;
        RECT 126.650 32.200 127.650 32.550 ;
        RECT 126.260 31.750 126.490 32.180 ;
        RECT 127.800 31.750 128.750 34.450 ;
        RECT 126.250 30.600 128.750 31.750 ;
        RECT 128.900 31.050 130.650 43.550 ;
        RECT 131.250 42.850 136.600 43.200 ;
        RECT 137.600 42.850 138.700 43.150 ;
        RECT 130.860 42.450 131.090 42.810 ;
        RECT 132.450 42.800 136.600 42.850 ;
        RECT 132.450 42.450 136.950 42.800 ;
        RECT 137.210 42.450 137.440 42.810 ;
        RECT 138.850 42.450 139.080 42.810 ;
        RECT 130.850 41.650 139.080 42.450 ;
        RECT 130.850 41.250 134.450 41.650 ;
        RECT 130.860 40.850 131.090 41.250 ;
        RECT 132.450 41.200 134.450 41.250 ;
        RECT 132.500 40.850 134.450 41.200 ;
        RECT 131.300 40.800 132.300 40.850 ;
        RECT 131.295 40.570 132.300 40.800 ;
        RECT 131.300 40.550 132.300 40.570 ;
        RECT 132.550 40.520 134.450 40.850 ;
        RECT 130.860 40.100 131.090 40.520 ;
        RECT 132.500 40.100 134.450 40.520 ;
        RECT 130.850 38.850 134.450 40.100 ;
        RECT 130.860 38.560 131.090 38.850 ;
        RECT 132.450 38.550 134.450 38.850 ;
        RECT 131.250 38.250 134.450 38.550 ;
        RECT 130.860 37.950 131.090 38.230 ;
        RECT 132.450 37.950 134.450 38.250 ;
        RECT 130.850 36.750 134.450 37.950 ;
        RECT 130.860 36.270 131.090 36.750 ;
        RECT 131.300 36.220 132.300 36.250 ;
        RECT 131.295 35.990 132.300 36.220 ;
        RECT 131.300 35.950 132.300 35.990 ;
        RECT 130.860 35.650 131.090 35.940 ;
        RECT 132.450 35.650 134.450 36.750 ;
        RECT 130.850 34.450 134.450 35.650 ;
        RECT 130.860 33.980 131.090 34.450 ;
        RECT 132.450 33.950 134.450 34.450 ;
        RECT 131.250 33.700 134.450 33.950 ;
        RECT 130.860 33.250 131.090 33.650 ;
        RECT 132.450 33.250 134.450 33.700 ;
        RECT 130.850 32.050 134.450 33.250 ;
        RECT 130.860 31.690 131.090 32.050 ;
        RECT 131.300 31.640 132.300 31.700 ;
        RECT 131.295 31.410 132.300 31.640 ;
        RECT 131.300 31.400 132.300 31.410 ;
        RECT 130.860 31.000 131.090 31.360 ;
        RECT 132.450 31.000 134.450 32.050 ;
        RECT 126.260 30.220 126.490 30.600 ;
        RECT 127.800 30.200 128.750 30.600 ;
        RECT 126.650 29.900 128.750 30.200 ;
        RECT 126.260 29.500 126.490 29.890 ;
        RECT 127.800 29.500 128.750 29.900 ;
        RECT 130.850 29.800 134.450 31.000 ;
        RECT 126.250 28.350 128.750 29.500 ;
        RECT 130.860 29.400 131.090 29.800 ;
        RECT 132.450 29.350 134.450 29.800 ;
        RECT 131.250 29.150 134.450 29.350 ;
        RECT 135.450 41.250 139.080 41.650 ;
        RECT 135.450 40.050 136.950 41.250 ;
        RECT 137.210 40.850 137.440 41.250 ;
        RECT 138.850 40.850 139.080 41.250 ;
        RECT 137.650 40.800 138.700 40.850 ;
        RECT 137.645 40.570 138.700 40.800 ;
        RECT 137.650 40.550 138.700 40.570 ;
        RECT 137.210 40.050 137.440 40.520 ;
        RECT 138.850 40.050 139.080 40.520 ;
        RECT 135.450 38.850 139.080 40.050 ;
        RECT 135.450 37.950 136.950 38.850 ;
        RECT 137.210 38.560 137.440 38.850 ;
        RECT 138.850 38.560 139.080 38.850 ;
        RECT 137.600 38.250 138.700 38.550 ;
        RECT 137.210 37.950 137.440 38.230 ;
        RECT 138.850 37.950 139.080 38.230 ;
        RECT 135.450 36.750 139.080 37.950 ;
        RECT 135.450 35.650 136.950 36.750 ;
        RECT 137.210 36.270 137.440 36.750 ;
        RECT 138.850 36.270 139.080 36.750 ;
        RECT 137.650 36.220 138.700 36.250 ;
        RECT 137.645 35.990 138.700 36.220 ;
        RECT 137.650 35.950 138.700 35.990 ;
        RECT 137.210 35.650 137.440 35.940 ;
        RECT 138.850 35.650 139.080 35.940 ;
        RECT 135.450 34.450 139.080 35.650 ;
        RECT 135.450 33.250 136.950 34.450 ;
        RECT 137.210 33.980 137.440 34.450 ;
        RECT 138.850 33.980 139.080 34.450 ;
        RECT 137.600 33.650 138.700 33.950 ;
        RECT 137.210 33.250 137.440 33.650 ;
        RECT 138.850 33.250 139.080 33.650 ;
        RECT 135.450 32.050 139.080 33.250 ;
        RECT 135.450 31.000 136.950 32.050 ;
        RECT 137.210 31.690 137.440 32.050 ;
        RECT 137.650 31.640 138.700 31.700 ;
        RECT 138.850 31.690 139.080 32.050 ;
        RECT 137.645 31.410 138.700 31.640 ;
        RECT 137.650 31.400 138.700 31.410 ;
        RECT 137.210 31.000 137.440 31.360 ;
        RECT 138.850 31.000 139.080 31.360 ;
        RECT 139.250 31.050 141.550 43.550 ;
        RECT 142.200 43.100 143.250 43.400 ;
        RECT 135.450 29.800 139.080 31.000 ;
        RECT 135.450 29.150 136.950 29.800 ;
        RECT 137.210 29.400 137.440 29.800 ;
        RECT 138.850 29.400 139.080 29.800 ;
        RECT 137.925 29.350 138.475 29.380 ;
        RECT 131.250 29.100 136.950 29.150 ;
        RECT 126.260 27.930 126.490 28.350 ;
        RECT 126.650 27.600 127.650 27.950 ;
        RECT 126.260 27.200 126.490 27.600 ;
        RECT 127.800 27.200 128.750 28.350 ;
        RECT 132.450 28.200 136.950 29.100 ;
        RECT 137.600 29.050 138.700 29.350 ;
        RECT 137.700 28.800 138.650 29.050 ;
        RECT 137.925 28.770 138.475 28.800 ;
        RECT 132.450 27.400 134.800 28.200 ;
        RECT 137.650 27.700 138.650 28.100 ;
        RECT 131.550 27.290 134.800 27.400 ;
        RECT 136.100 27.450 138.650 27.700 ;
        RECT 136.100 27.290 138.500 27.450 ;
        RECT 139.700 27.400 141.550 31.050 ;
        RECT 141.700 30.300 142.050 43.100 ;
        RECT 143.450 42.610 143.680 43.070 ;
        RECT 142.250 42.560 143.300 42.600 ;
        RECT 142.245 42.330 143.300 42.560 ;
        RECT 142.250 42.300 143.300 42.330 ;
        RECT 144.050 42.500 148.650 42.650 ;
        RECT 150.100 42.500 152.400 92.000 ;
        RECT 143.450 41.820 143.680 42.280 ;
        RECT 142.200 41.500 143.250 41.800 ;
        RECT 144.050 41.700 155.700 42.500 ;
        RECT 143.450 41.030 143.680 41.490 ;
        RECT 142.250 40.980 143.300 41.000 ;
        RECT 142.245 40.750 143.300 40.980 ;
        RECT 142.250 40.700 143.300 40.750 ;
        RECT 144.050 40.800 157.310 41.700 ;
        RECT 142.200 39.950 143.250 40.250 ;
        RECT 143.450 40.240 143.680 40.700 ;
        RECT 144.050 40.200 155.700 40.800 ;
        RECT 156.410 40.600 157.310 40.800 ;
        RECT 143.450 39.450 143.680 39.910 ;
        RECT 144.050 39.450 148.650 40.200 ;
        RECT 156.380 39.700 157.340 40.600 ;
        RECT 142.250 39.400 143.300 39.450 ;
        RECT 142.245 39.170 143.300 39.400 ;
        RECT 142.250 39.150 143.300 39.170 ;
        RECT 144.050 39.400 147.400 39.450 ;
        RECT 143.450 38.660 143.680 39.120 ;
        RECT 142.200 38.350 143.250 38.650 ;
        RECT 143.450 37.870 143.680 38.330 ;
        RECT 142.250 37.820 143.300 37.850 ;
        RECT 142.245 37.590 143.300 37.820 ;
        RECT 142.250 37.550 143.300 37.590 ;
        RECT 143.450 37.080 143.680 37.540 ;
        RECT 142.200 36.750 143.250 37.050 ;
        RECT 143.450 36.290 143.680 36.750 ;
        RECT 142.250 36.240 143.300 36.250 ;
        RECT 142.245 36.010 143.300 36.240 ;
        RECT 142.250 35.950 143.300 36.010 ;
        RECT 143.450 35.500 143.680 35.960 ;
        RECT 142.200 35.200 143.250 35.500 ;
        RECT 143.450 34.710 143.680 35.170 ;
        RECT 142.250 34.660 143.300 34.700 ;
        RECT 142.245 34.430 143.300 34.660 ;
        RECT 142.250 34.400 143.300 34.430 ;
        RECT 143.450 33.920 143.680 34.380 ;
        RECT 142.200 33.600 143.250 33.900 ;
        RECT 142.250 33.080 143.300 33.150 ;
        RECT 143.450 33.130 143.680 33.590 ;
        RECT 142.245 32.850 143.300 33.080 ;
        RECT 142.200 32.050 143.250 32.350 ;
        RECT 143.450 32.340 143.680 32.800 ;
        RECT 143.450 31.550 143.680 32.010 ;
        RECT 142.250 31.500 143.300 31.550 ;
        RECT 142.245 31.270 143.300 31.500 ;
        RECT 142.250 31.250 143.300 31.270 ;
        RECT 143.450 30.760 143.680 31.220 ;
        RECT 142.200 30.450 143.250 30.750 ;
        RECT 141.700 29.400 142.100 30.300 ;
        RECT 143.450 29.970 143.680 30.430 ;
        RECT 142.250 29.920 143.300 29.950 ;
        RECT 142.245 29.690 143.300 29.920 ;
        RECT 142.250 29.650 143.300 29.690 ;
        RECT 141.700 27.550 142.050 29.400 ;
        RECT 143.450 29.180 143.680 29.640 ;
        RECT 142.200 28.850 143.250 29.150 ;
        RECT 142.250 28.340 143.300 28.400 ;
        RECT 143.450 28.390 143.680 28.850 ;
        RECT 142.245 28.110 143.300 28.340 ;
        RECT 142.250 28.100 143.300 28.110 ;
        RECT 143.450 27.600 143.680 28.060 ;
        RECT 142.200 27.300 143.250 27.600 ;
        RECT 126.250 26.050 128.750 27.200 ;
        RECT 129.550 26.860 130.550 27.250 ;
        RECT 131.400 27.150 134.800 27.290 ;
        RECT 131.400 27.060 133.900 27.150 ;
        RECT 136.000 27.060 138.500 27.290 ;
        RECT 131.550 27.050 133.850 27.060 ;
        RECT 131.010 26.950 131.240 27.010 ;
        RECT 134.060 26.950 134.290 27.010 ;
        RECT 135.610 26.950 135.840 27.010 ;
        RECT 138.660 26.950 138.890 27.010 ;
        RECT 130.900 26.860 131.300 26.950 ;
        RECT 134.000 26.860 134.400 26.950 ;
        RECT 129.550 26.645 134.400 26.860 ;
        RECT 129.550 26.250 130.550 26.645 ;
        RECT 130.900 26.600 131.300 26.645 ;
        RECT 134.000 26.600 134.400 26.645 ;
        RECT 135.500 26.875 135.900 26.950 ;
        RECT 138.600 26.875 139.000 26.950 ;
        RECT 139.400 26.875 140.400 27.250 ;
        RECT 135.500 26.650 140.400 26.875 ;
        RECT 135.500 26.600 135.900 26.650 ;
        RECT 138.600 26.630 140.400 26.650 ;
        RECT 138.600 26.600 139.000 26.630 ;
        RECT 131.010 26.550 131.240 26.600 ;
        RECT 134.060 26.550 134.290 26.600 ;
        RECT 135.610 26.550 135.840 26.600 ;
        RECT 138.660 26.550 138.890 26.600 ;
        RECT 131.400 26.400 133.900 26.500 ;
        RECT 136.000 26.400 138.500 26.500 ;
        RECT 131.400 26.270 138.500 26.400 ;
        RECT 131.600 26.050 138.250 26.270 ;
        RECT 139.400 26.250 140.400 26.630 ;
        RECT 144.050 26.600 145.350 39.400 ;
        RECT 146.150 39.250 147.200 39.400 ;
        RECT 146.200 39.150 147.200 39.250 ;
        RECT 145.810 38.750 146.040 39.100 ;
        RECT 145.700 38.550 146.050 38.750 ;
        RECT 147.360 38.550 147.590 39.100 ;
        RECT 145.700 37.600 147.590 38.550 ;
        RECT 145.700 36.300 146.050 37.600 ;
        RECT 146.200 36.850 147.200 37.150 ;
        RECT 147.360 37.140 147.590 37.600 ;
        RECT 147.360 36.300 147.590 36.810 ;
        RECT 145.700 35.350 147.590 36.300 ;
        RECT 145.700 33.950 146.050 35.350 ;
        RECT 147.360 34.850 147.590 35.350 ;
        RECT 146.200 34.550 147.200 34.850 ;
        RECT 147.360 33.950 147.590 34.520 ;
        RECT 145.700 33.000 147.590 33.950 ;
        RECT 145.700 31.800 146.050 33.000 ;
        RECT 147.360 32.560 147.590 33.000 ;
        RECT 146.200 32.250 147.200 32.550 ;
        RECT 147.360 31.800 147.590 32.230 ;
        RECT 145.700 30.850 147.590 31.800 ;
        RECT 145.700 29.500 146.050 30.850 ;
        RECT 146.200 29.950 147.200 30.300 ;
        RECT 147.360 30.270 147.590 30.850 ;
        RECT 147.360 29.500 147.590 29.940 ;
        RECT 145.700 28.550 147.590 29.500 ;
        RECT 145.700 27.250 146.050 28.550 ;
        RECT 146.200 27.650 147.200 28.000 ;
        RECT 147.360 27.980 147.590 28.550 ;
        RECT 147.360 27.250 147.590 27.650 ;
        RECT 145.700 26.300 147.590 27.250 ;
        RECT 126.260 25.640 126.490 26.050 ;
        RECT 127.800 25.800 128.750 26.050 ;
        RECT 127.800 25.650 129.130 25.800 ;
        RECT 130.450 25.650 131.450 25.950 ;
        RECT 126.650 25.350 129.130 25.650 ;
        RECT 126.260 24.950 126.490 25.310 ;
        RECT 127.800 25.150 129.130 25.350 ;
        RECT 127.800 24.950 128.750 25.150 ;
        RECT 132.450 25.100 137.700 26.050 ;
        RECT 138.600 25.650 139.600 25.950 ;
        RECT 143.555 25.920 144.445 25.950 ;
        RECT 145.700 25.920 146.050 26.300 ;
        RECT 143.555 25.030 146.050 25.920 ;
        RECT 147.360 25.690 147.590 26.300 ;
        RECT 146.300 25.640 147.200 25.650 ;
        RECT 146.200 25.410 147.200 25.640 ;
        RECT 146.300 25.350 147.200 25.410 ;
        RECT 143.555 25.000 144.445 25.030 ;
        RECT 126.250 23.800 128.750 24.950 ;
        RECT 145.700 24.900 146.050 25.030 ;
        RECT 147.360 24.900 147.590 25.360 ;
        RECT 130.650 24.610 132.610 24.840 ;
        RECT 132.940 24.610 134.900 24.840 ;
        RECT 135.230 24.610 137.190 24.840 ;
        RECT 137.520 24.610 139.480 24.840 ;
        RECT 130.370 24.400 130.600 24.450 ;
        RECT 126.260 23.350 126.490 23.800 ;
        RECT 127.800 23.350 128.750 23.800 ;
        RECT 130.250 23.500 130.650 24.400 ;
        RECT 130.370 23.450 130.600 23.500 ;
        RECT 127.850 23.300 128.750 23.350 ;
        RECT 131.100 23.300 132.000 24.610 ;
        RECT 132.660 24.300 132.890 24.450 ;
        RECT 132.550 23.600 133.000 24.300 ;
        RECT 132.660 23.450 132.890 23.600 ;
        RECT 133.500 23.300 134.400 24.610 ;
        RECT 134.950 24.300 135.180 24.450 ;
        RECT 134.850 23.600 135.300 24.300 ;
        RECT 134.950 23.450 135.180 23.600 ;
        RECT 135.800 23.300 136.700 24.610 ;
        RECT 137.240 24.300 137.470 24.450 ;
        RECT 137.150 23.600 137.600 24.300 ;
        RECT 137.240 23.450 137.470 23.600 ;
        RECT 138.050 23.300 138.950 24.610 ;
        RECT 139.530 24.400 139.760 24.450 ;
        RECT 139.450 23.500 139.850 24.400 ;
        RECT 139.530 23.450 139.760 23.500 ;
        RECT 126.650 22.950 127.650 23.300 ;
        RECT 127.850 23.290 139.450 23.300 ;
        RECT 127.850 23.060 139.480 23.290 ;
        RECT 127.850 23.000 139.450 23.060 ;
        RECT 140.050 22.800 141.400 24.850 ;
        RECT 143.850 22.800 145.550 24.300 ;
        RECT 145.700 23.950 147.650 24.900 ;
        RECT 147.900 24.300 148.650 37.250 ;
        RECT 145.700 23.450 146.050 23.950 ;
        RECT 145.810 23.400 146.040 23.450 ;
        RECT 147.360 23.400 147.590 23.950 ;
        RECT 146.200 23.050 147.200 23.400 ;
        RECT 147.800 22.800 148.650 24.300 ;
        RECT 124.450 21.595 148.650 22.800 ;
        RECT 104.780 20.450 148.650 21.595 ;
        RECT 104.780 20.405 117.950 20.450 ;
        RECT 121.950 20.405 129.595 20.450 ;
        RECT 114.850 20.400 115.600 20.405 ;
        RECT 115.080 18.300 115.330 18.615 ;
        RECT 119.130 18.300 119.380 18.815 ;
        RECT 114.850 17.100 119.650 18.300 ;
        RECT 115.080 16.510 115.330 17.100 ;
        RECT 116.650 14.850 117.850 17.100 ;
        RECT 119.130 16.710 119.380 17.100 ;
        RECT 150.250 14.850 151.450 14.880 ;
        RECT 116.650 13.650 151.450 14.850 ;
        RECT 150.250 13.620 151.450 13.650 ;
      LAYER via ;
        RECT 102.090 90.335 103.115 91.360 ;
        RECT 126.420 88.690 127.100 89.370 ;
        RECT 111.075 68.045 112.265 69.235 ;
        RECT 146.400 82.010 147.500 83.110 ;
        RECT 111.800 67.000 112.520 67.720 ;
        RECT 144.090 48.570 145.010 49.490 ;
        RECT 137.650 42.850 138.650 43.150 ;
        RECT 129.200 40.850 130.050 41.200 ;
        RECT 129.100 40.550 130.050 40.850 ;
        RECT 124.600 22.900 125.400 32.700 ;
        RECT 126.700 32.200 127.600 32.550 ;
        RECT 129.200 36.250 130.050 40.550 ;
        RECT 129.100 35.950 130.050 36.250 ;
        RECT 129.200 31.700 130.050 35.950 ;
        RECT 129.100 31.400 130.050 31.700 ;
        RECT 129.200 31.250 130.050 31.400 ;
        RECT 131.350 40.550 132.250 40.850 ;
        RECT 131.350 35.950 132.250 36.250 ;
        RECT 131.350 31.400 132.250 31.700 ;
        RECT 137.750 40.550 138.650 40.850 ;
        RECT 137.650 38.250 138.650 38.550 ;
        RECT 137.750 35.950 138.650 36.250 ;
        RECT 137.650 33.650 138.650 33.950 ;
        RECT 137.750 31.400 138.650 31.700 ;
        RECT 139.950 33.950 140.800 43.600 ;
        RECT 142.250 43.100 143.200 43.400 ;
        RECT 139.950 33.550 140.850 33.950 ;
        RECT 139.950 32.400 140.800 33.550 ;
        RECT 139.950 32.000 140.850 32.400 ;
        RECT 126.700 27.600 127.600 27.950 ;
        RECT 137.650 29.050 138.650 29.350 ;
        RECT 137.925 28.800 138.475 29.050 ;
        RECT 137.700 27.450 138.550 28.100 ;
        RECT 139.950 30.800 140.800 32.000 ;
        RECT 139.950 27.800 140.850 30.800 ;
        RECT 139.950 27.450 141.200 27.800 ;
        RECT 140.050 27.400 141.200 27.450 ;
        RECT 142.300 42.300 143.250 42.600 ;
        RECT 142.250 41.500 143.200 41.800 ;
        RECT 142.300 40.700 143.250 41.000 ;
        RECT 142.250 39.950 143.200 40.250 ;
        RECT 142.300 39.150 143.250 39.450 ;
        RECT 142.250 38.350 143.200 38.650 ;
        RECT 142.300 37.550 143.250 37.850 ;
        RECT 142.250 36.750 143.200 37.050 ;
        RECT 142.300 35.950 143.250 36.250 ;
        RECT 142.250 35.200 143.200 35.500 ;
        RECT 142.300 34.400 143.250 34.700 ;
        RECT 142.250 33.600 143.200 33.900 ;
        RECT 142.300 32.850 143.250 33.150 ;
        RECT 142.250 32.050 143.200 32.350 ;
        RECT 142.300 31.250 143.250 31.550 ;
        RECT 142.250 30.450 143.200 30.750 ;
        RECT 141.750 29.600 142.050 30.000 ;
        RECT 142.300 29.650 143.250 29.950 ;
        RECT 142.250 28.850 143.200 29.150 ;
        RECT 142.300 28.100 143.250 28.400 ;
        RECT 142.250 27.300 143.200 27.600 ;
        RECT 129.650 27.030 130.350 27.050 ;
        RECT 129.625 26.475 130.350 27.030 ;
        RECT 129.650 26.450 130.350 26.475 ;
        RECT 130.950 26.600 131.250 26.950 ;
        RECT 134.050 26.600 134.350 26.950 ;
        RECT 135.550 26.600 135.850 26.950 ;
        RECT 138.650 26.600 138.950 26.950 ;
        RECT 139.675 26.480 140.225 27.030 ;
        RECT 144.400 26.600 145.000 42.450 ;
        RECT 148.100 39.750 148.500 42.450 ;
        RECT 156.410 39.700 157.310 40.600 ;
        RECT 146.200 39.250 147.150 39.550 ;
        RECT 146.350 39.150 147.100 39.250 ;
        RECT 146.250 36.850 147.150 37.150 ;
        RECT 146.250 34.550 147.150 34.850 ;
        RECT 146.250 32.250 147.150 32.550 ;
        RECT 146.250 29.950 147.150 30.300 ;
        RECT 146.250 27.650 147.150 28.000 ;
        RECT 128.450 25.150 129.100 25.800 ;
        RECT 130.500 25.650 131.400 25.950 ;
        RECT 132.600 25.400 133.000 26.100 ;
        RECT 137.150 25.400 137.550 26.100 ;
        RECT 138.650 25.650 139.550 25.950 ;
        RECT 146.350 25.350 147.150 25.650 ;
        RECT 130.300 23.500 130.600 24.400 ;
        RECT 132.600 23.600 132.950 24.300 ;
        RECT 134.900 23.600 135.250 24.300 ;
        RECT 137.200 23.600 137.550 24.300 ;
        RECT 139.500 23.500 139.800 24.400 ;
        RECT 126.700 22.950 127.600 23.300 ;
        RECT 148.050 24.600 148.450 37.100 ;
        RECT 146.250 23.050 147.150 23.400 ;
        RECT 130.150 22.250 130.650 22.350 ;
        RECT 134.900 22.250 135.250 22.350 ;
        RECT 139.300 22.250 139.800 22.350 ;
        RECT 130.150 21.900 139.800 22.250 ;
        RECT 130.150 21.600 139.750 21.900 ;
        RECT 150.250 13.650 151.450 14.850 ;
      LAYER met2 ;
        RECT 102.090 89.435 103.115 91.390 ;
        RECT 102.070 88.460 103.135 89.435 ;
        RECT 102.090 88.435 103.115 88.460 ;
        RECT 126.420 87.565 127.100 89.400 ;
        RECT 90.275 83.250 91.725 83.270 ;
        RECT 90.250 81.750 95.280 83.250 ;
        RECT 90.275 81.730 91.725 81.750 ;
        RECT 146.400 79.595 147.500 83.140 ;
        RECT 146.380 78.545 147.520 79.595 ;
        RECT 146.400 78.520 147.500 78.545 ;
        RECT 111.075 69.235 112.265 69.265 ;
        RECT 111.075 68.045 114.150 69.235 ;
        RECT 111.075 68.015 112.265 68.045 ;
        RECT 107.070 67.720 107.790 67.765 ;
        RECT 111.800 67.720 112.520 67.750 ;
        RECT 107.070 67.000 112.520 67.720 ;
        RECT 107.070 66.955 107.790 67.000 ;
        RECT 111.800 66.970 112.520 67.000 ;
        RECT 144.060 49.465 145.780 49.490 ;
        RECT 144.060 48.595 145.800 49.465 ;
        RECT 144.060 48.570 145.780 48.595 ;
        RECT 66.775 45.250 68.225 45.270 ;
        RECT 66.750 43.750 112.280 45.250 ;
        RECT 66.775 43.730 68.225 43.750 ;
        RECT 139.950 43.450 140.800 43.650 ;
        RECT 134.060 43.400 135.840 43.440 ;
        RECT 134.050 43.150 138.700 43.400 ;
        RECT 134.060 42.850 138.700 43.150 ;
        RECT 139.950 43.050 143.250 43.450 ;
        RECT 134.060 42.810 138.650 42.850 ;
        RECT 129.200 40.900 130.050 41.250 ;
        RECT 129.100 40.850 130.050 40.900 ;
        RECT 131.350 40.850 132.250 40.900 ;
        RECT 129.050 40.550 132.500 40.850 ;
        RECT 129.100 40.500 130.050 40.550 ;
        RECT 131.350 40.500 132.250 40.550 ;
        RECT 129.200 36.300 130.050 40.500 ;
        RECT 134.060 38.590 135.840 42.810 ;
        RECT 137.650 42.800 138.650 42.810 ;
        RECT 139.950 41.850 140.800 43.050 ;
        RECT 142.250 42.250 148.650 42.650 ;
        RECT 139.950 41.450 143.250 41.850 ;
        RECT 139.950 40.900 140.800 41.450 ;
        RECT 144.050 41.000 148.650 42.250 ;
        RECT 137.750 40.550 140.800 40.900 ;
        RECT 142.250 40.700 148.650 41.000 ;
        RECT 137.750 40.500 138.650 40.550 ;
        RECT 139.950 40.300 140.800 40.550 ;
        RECT 139.950 39.900 143.250 40.300 ;
        RECT 139.950 38.700 140.800 39.900 ;
        RECT 144.100 39.450 148.650 40.700 ;
        RECT 142.250 39.150 147.350 39.450 ;
        RECT 144.050 39.000 147.350 39.150 ;
        RECT 137.650 38.590 138.650 38.600 ;
        RECT 134.060 38.210 138.700 38.590 ;
        RECT 139.950 38.300 143.250 38.700 ;
        RECT 129.100 36.250 130.050 36.300 ;
        RECT 131.350 36.250 132.250 36.300 ;
        RECT 129.050 35.950 132.500 36.250 ;
        RECT 129.100 35.900 130.050 35.950 ;
        RECT 131.350 35.900 132.250 35.950 ;
        RECT 124.600 32.700 125.400 32.750 ;
        RECT 124.600 32.050 127.750 32.700 ;
        RECT 124.600 28.150 125.400 32.050 ;
        RECT 129.200 31.750 130.050 35.900 ;
        RECT 134.060 33.990 135.840 38.210 ;
        RECT 137.650 38.200 138.650 38.210 ;
        RECT 139.950 37.100 140.800 38.300 ;
        RECT 144.050 37.850 145.350 39.000 ;
        RECT 142.250 37.550 145.350 37.850 ;
        RECT 139.950 36.700 143.200 37.100 ;
        RECT 139.950 36.350 140.800 36.700 ;
        RECT 137.750 35.950 140.800 36.350 ;
        RECT 144.050 36.300 145.350 37.550 ;
        RECT 146.200 36.700 148.650 37.250 ;
        RECT 142.250 35.950 145.350 36.300 ;
        RECT 137.750 35.900 138.650 35.950 ;
        RECT 139.950 35.550 140.800 35.950 ;
        RECT 139.950 35.150 143.200 35.550 ;
        RECT 137.650 33.990 138.650 34.000 ;
        RECT 134.060 33.610 138.650 33.990 ;
        RECT 129.100 31.700 130.050 31.750 ;
        RECT 131.350 31.700 132.250 31.750 ;
        RECT 129.050 31.400 132.500 31.700 ;
        RECT 129.100 31.350 130.050 31.400 ;
        RECT 131.350 31.350 132.250 31.400 ;
        RECT 129.200 31.200 130.050 31.350 ;
        RECT 134.060 30.110 135.840 33.610 ;
        RECT 137.650 33.600 138.650 33.610 ;
        RECT 139.950 33.950 140.800 35.150 ;
        RECT 144.050 34.950 145.350 35.950 ;
        RECT 144.050 34.700 147.350 34.950 ;
        RECT 142.250 34.400 147.350 34.700 ;
        RECT 142.250 34.350 145.350 34.400 ;
        RECT 139.950 33.550 143.250 33.950 ;
        RECT 139.950 32.400 140.800 33.550 ;
        RECT 144.050 33.150 145.350 34.350 ;
        RECT 142.250 32.800 145.350 33.150 ;
        RECT 139.950 32.000 143.250 32.400 ;
        RECT 139.950 31.750 140.800 32.000 ;
        RECT 137.750 31.400 140.800 31.750 ;
        RECT 144.050 31.550 145.350 32.800 ;
        RECT 147.900 32.700 148.650 36.700 ;
        RECT 156.410 34.925 157.310 40.630 ;
        RECT 156.390 34.075 157.330 34.925 ;
        RECT 156.410 34.050 157.310 34.075 ;
        RECT 146.200 32.150 148.650 32.700 ;
        RECT 137.750 31.350 138.650 31.400 ;
        RECT 139.950 30.800 140.800 31.400 ;
        RECT 142.250 31.200 145.350 31.550 ;
        RECT 139.950 30.400 143.250 30.800 ;
        RECT 134.070 28.870 135.830 30.110 ;
        RECT 137.925 29.400 138.475 29.970 ;
        RECT 124.600 27.500 127.750 28.150 ;
        RECT 137.650 27.850 138.650 29.400 ;
        RECT 139.950 29.200 140.850 30.400 ;
        RECT 144.050 30.350 145.350 31.200 ;
        RECT 141.050 29.550 142.050 30.050 ;
        RECT 144.050 30.000 147.350 30.350 ;
        RECT 142.250 29.800 147.350 30.000 ;
        RECT 142.250 29.600 145.350 29.800 ;
        RECT 141.050 29.500 141.750 29.550 ;
        RECT 139.950 28.800 143.200 29.200 ;
        RECT 139.950 27.850 140.850 28.800 ;
        RECT 144.050 28.450 145.350 29.600 ;
        RECT 142.250 28.050 145.350 28.450 ;
        RECT 147.900 28.100 148.650 32.150 ;
        RECT 124.600 23.550 125.400 27.500 ;
        RECT 129.250 27.030 130.450 27.750 ;
        RECT 137.700 27.400 138.550 27.850 ;
        RECT 139.950 27.700 141.200 27.850 ;
        RECT 139.950 27.400 143.200 27.700 ;
        RECT 141.100 27.250 143.200 27.400 ;
        RECT 139.600 27.030 140.900 27.250 ;
        RECT 129.250 27.000 134.325 27.030 ;
        RECT 135.575 27.000 140.900 27.030 ;
        RECT 129.250 26.550 134.350 27.000 ;
        RECT 135.550 26.550 140.900 27.000 ;
        RECT 144.050 27.200 145.350 28.050 ;
        RECT 146.200 27.550 148.650 28.100 ;
        RECT 144.050 26.600 147.150 27.200 ;
        RECT 129.250 26.475 134.325 26.550 ;
        RECT 135.575 26.480 140.900 26.550 ;
        RECT 129.250 26.300 130.450 26.475 ;
        RECT 139.600 26.250 140.900 26.480 ;
        RECT 128.450 25.800 129.100 25.830 ;
        RECT 128.450 25.150 129.820 25.800 ;
        RECT 130.100 25.550 131.450 26.000 ;
        RECT 128.450 25.120 129.100 25.150 ;
        RECT 124.600 22.900 127.750 23.550 ;
        RECT 124.600 22.850 125.400 22.900 ;
        RECT 130.100 22.350 130.750 25.550 ;
        RECT 132.500 23.450 133.100 26.200 ;
        RECT 134.800 22.350 135.350 24.450 ;
        RECT 137.050 23.450 137.650 26.200 ;
        RECT 138.550 25.550 139.900 26.000 ;
        RECT 142.535 25.920 143.375 26.095 ;
        RECT 139.250 22.350 139.900 25.550 ;
        RECT 142.510 25.030 144.475 25.920 ;
        RECT 146.350 25.300 147.150 26.600 ;
        RECT 142.535 24.855 143.375 25.030 ;
        RECT 147.900 23.550 148.650 27.550 ;
        RECT 146.200 23.000 148.650 23.550 ;
        RECT 130.100 21.450 139.900 22.350 ;
        RECT 150.250 14.850 151.450 22.145 ;
        RECT 150.220 13.650 151.480 14.850 ;
      LAYER via2 ;
        RECT 102.115 88.460 103.090 89.435 ;
        RECT 126.420 87.610 127.100 88.290 ;
        RECT 90.275 81.775 91.725 83.225 ;
        RECT 146.425 78.545 147.475 79.595 ;
        RECT 112.915 68.045 114.105 69.235 ;
        RECT 144.885 48.595 145.755 49.465 ;
        RECT 66.775 43.775 68.225 45.225 ;
        RECT 156.435 34.075 157.285 34.925 ;
        RECT 134.300 29.350 135.750 30.150 ;
        RECT 137.925 29.375 138.475 29.925 ;
        RECT 129.350 27.100 129.950 27.650 ;
        RECT 140.200 26.450 140.800 27.150 ;
        RECT 129.125 25.150 129.775 25.800 ;
        RECT 142.535 24.900 143.375 26.050 ;
        RECT 150.250 20.900 151.450 22.100 ;
      LAYER met3 ;
        RECT 87.255 83.250 88.745 83.275 ;
        RECT 87.250 81.750 91.750 83.250 ;
        RECT 87.255 81.725 88.745 81.750 ;
        RECT 28.255 45.250 29.745 45.275 ;
        RECT 28.250 43.750 68.250 45.250 ;
        RECT 28.255 43.725 29.745 43.750 ;
        RECT 102.090 27.500 103.115 89.460 ;
        RECT 126.395 87.585 127.125 88.315 ;
        RECT 126.420 86.790 127.100 87.585 ;
        RECT 109.380 70.450 126.240 85.850 ;
        RECT 128.080 69.740 144.940 85.140 ;
        RECT 112.890 69.235 114.130 69.260 ;
        RECT 112.890 68.045 115.675 69.235 ;
        RECT 112.890 68.020 114.130 68.045 ;
        RECT 146.400 67.985 147.500 79.620 ;
        RECT 107.045 66.975 107.815 67.745 ;
        RECT 107.070 63.140 107.790 66.975 ;
        RECT 109.290 51.330 126.150 66.730 ;
        RECT 128.250 51.530 145.110 66.930 ;
        RECT 146.375 66.895 147.525 67.985 ;
        RECT 146.400 66.890 147.500 66.895 ;
        RECT 144.860 50.055 145.780 50.060 ;
        RECT 144.835 49.145 145.805 50.055 ;
        RECT 144.860 48.570 145.780 49.145 ;
        RECT 134.200 30.165 141.150 30.200 ;
        RECT 134.200 29.975 141.715 30.165 ;
        RECT 134.200 29.525 141.750 29.975 ;
        RECT 134.200 29.340 141.715 29.525 ;
        RECT 134.200 29.250 141.150 29.340 ;
        RECT 136.500 28.750 139.350 29.250 ;
        RECT 123.300 27.500 130.150 27.850 ;
        RECT 102.090 26.950 130.150 27.500 ;
        RECT 140.150 27.300 150.000 27.400 ;
        RECT 102.090 26.500 123.950 26.950 ;
        RECT 140.150 26.600 151.450 27.300 ;
        RECT 102.090 26.490 103.115 26.500 ;
        RECT 140.150 26.400 140.950 26.600 ;
        RECT 149.150 26.100 151.450 26.600 ;
        RECT 128.850 24.875 143.400 26.075 ;
        RECT 150.250 22.125 151.450 26.100 ;
        RECT 150.225 20.875 151.475 22.125 ;
        RECT 156.410 8.645 157.310 34.950 ;
        RECT 156.385 7.755 157.335 8.645 ;
        RECT 156.410 7.750 157.310 7.755 ;
      LAYER via3 ;
        RECT 87.255 81.755 88.745 83.245 ;
        RECT 28.255 43.755 29.745 45.245 ;
        RECT 126.420 86.820 127.100 87.500 ;
        RECT 125.820 70.590 126.140 85.710 ;
        RECT 144.520 69.880 144.840 85.000 ;
        RECT 114.455 68.045 115.645 69.235 ;
        RECT 146.405 66.895 147.495 67.985 ;
        RECT 107.070 63.170 107.790 63.890 ;
        RECT 125.730 51.470 126.050 66.590 ;
        RECT 144.690 51.670 145.010 66.790 ;
        RECT 144.865 49.145 145.775 50.055 ;
        RECT 156.415 7.755 157.305 8.645 ;
      LAYER met4 ;
        RECT 3.990 223.800 4.290 224.760 ;
        RECT 7.670 223.800 7.970 224.760 ;
        RECT 11.350 223.800 11.650 224.760 ;
        RECT 15.030 223.800 15.330 224.760 ;
        RECT 18.710 223.800 19.010 224.760 ;
        RECT 22.390 223.800 22.690 224.760 ;
        RECT 26.070 223.800 26.370 224.760 ;
        RECT 29.750 223.800 30.050 224.760 ;
        RECT 33.430 223.800 33.730 224.760 ;
        RECT 37.110 223.800 37.410 224.760 ;
        RECT 40.790 223.800 41.090 224.760 ;
        RECT 44.470 223.800 44.770 224.760 ;
        RECT 48.150 223.800 48.450 224.760 ;
        RECT 51.830 223.800 52.130 224.760 ;
        RECT 55.510 223.800 55.810 224.760 ;
        RECT 59.190 223.800 59.490 224.760 ;
        RECT 62.870 223.800 63.170 224.760 ;
        RECT 66.550 223.800 66.850 224.760 ;
        RECT 70.230 223.800 70.530 224.760 ;
        RECT 73.910 223.800 74.210 224.760 ;
        RECT 77.590 223.800 77.890 224.760 ;
        RECT 81.270 223.800 81.570 224.760 ;
        RECT 84.950 223.800 85.250 224.760 ;
        RECT 88.630 223.800 88.930 224.760 ;
        RECT 3.200 223.500 88.930 223.800 ;
        RECT 49.000 220.760 50.500 223.500 ;
        RECT 66.550 223.450 66.850 223.500 ;
        RECT 84.950 223.450 85.250 223.500 ;
        RECT 126.415 87.010 127.105 87.505 ;
        RECT 125.300 85.830 145.270 87.010 ;
        RECT 50.500 81.750 88.750 83.250 ;
        RECT 109.775 70.845 124.385 85.455 ;
        RECT 125.300 79.990 126.480 85.830 ;
        RECT 116.170 69.275 117.300 70.845 ;
        RECT 125.740 70.510 126.220 79.990 ;
        RECT 128.475 70.135 143.085 84.745 ;
        RECT 144.090 79.430 145.270 85.830 ;
        RECT 136.165 69.275 137.295 70.135 ;
        RECT 144.440 69.800 144.920 79.430 ;
        RECT 114.450 69.235 115.650 69.240 ;
        RECT 116.170 69.235 137.295 69.275 ;
        RECT 114.450 68.145 137.295 69.235 ;
        RECT 114.450 68.045 117.095 68.145 ;
        RECT 114.450 68.040 115.650 68.045 ;
        RECT 144.260 66.890 147.500 67.990 ;
        RECT 107.065 63.890 107.795 63.895 ;
        RECT 109.685 63.890 124.295 66.335 ;
        RECT 125.650 66.210 126.130 66.670 ;
        RECT 128.645 66.210 143.255 66.535 ;
        RECT 107.065 63.170 124.295 63.890 ;
        RECT 107.065 63.165 107.795 63.170 ;
        RECT 109.685 51.725 124.295 63.170 ;
        RECT 125.410 61.400 143.255 66.210 ;
        RECT 144.260 62.050 145.360 66.890 ;
        RECT 125.650 51.390 126.130 61.400 ;
        RECT 126.690 50.780 127.610 61.400 ;
        RECT 128.645 51.925 143.255 61.400 ;
        RECT 144.610 51.590 145.090 62.050 ;
        RECT 126.690 49.860 145.780 50.780 ;
        RECT 144.860 49.140 145.780 49.860 ;
        RECT 2.500 43.750 29.750 45.250 ;
        RECT 156.410 1.000 157.310 8.650 ;
  END
END tt_um_twin_tee_opamp_osc
END LIBRARY

