VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_analog_rf_readout_circuit
  CLASS BLOCK ;
  FOREIGN tt_um_analog_rf_readout_circuit ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.000000 ;
    ANTENNADIFFAREA 56.617199 ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 22.000000 ;
    ANTENNADIFFAREA 56.617199 ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 103.665 45.850 107.785 47.470 ;
        RECT 124.660 47.425 129.890 48.360 ;
        RECT 123.175 47.415 129.890 47.425 ;
        RECT 120.445 43.100 129.890 47.415 ;
        RECT 120.450 43.085 129.890 43.100 ;
        RECT 124.660 41.740 129.890 43.085 ;
        RECT 135.950 47.390 137.390 54.395 ;
        RECT 135.950 47.385 139.730 47.390 ;
        RECT 135.950 43.065 142.920 47.385 ;
        RECT 135.950 33.775 137.390 43.065 ;
        RECT 139.670 43.055 142.920 43.065 ;
        RECT 111.955 6.105 113.485 6.520 ;
        RECT 90.150 5.735 91.240 5.995 ;
        RECT 89.260 5.660 91.240 5.735 ;
        RECT 89.260 4.875 92.195 5.660 ;
        RECT 111.955 5.165 114.415 6.105 ;
        RECT 134.000 6.095 135.530 6.515 ;
        RECT 111.955 4.900 113.485 5.165 ;
        RECT 134.000 5.155 136.455 6.095 ;
        RECT 156.100 5.830 157.630 6.515 ;
        RECT 134.000 4.895 135.530 5.155 ;
        RECT 154.130 4.895 157.630 5.830 ;
        RECT 154.130 4.890 155.100 4.895 ;
        RECT 90.150 4.720 92.195 4.875 ;
        RECT 90.150 4.375 91.240 4.720 ;
      LAYER li1 ;
        RECT 121.435 56.235 122.505 56.440 ;
        RECT 98.005 51.200 98.355 53.360 ;
        RECT 98.005 48.540 98.355 50.700 ;
        RECT 105.435 47.650 105.605 56.155 ;
        RECT 104.150 47.480 107.105 47.650 ;
        RECT 104.150 47.240 104.320 47.480 ;
        RECT 103.945 46.080 104.645 47.240 ;
        RECT 105.035 45.880 105.205 47.180 ;
        RECT 105.475 46.140 105.645 47.480 ;
        RECT 105.915 46.320 106.085 47.180 ;
        RECT 104.795 45.520 105.295 45.880 ;
        RECT 104.795 44.100 104.965 45.520 ;
        RECT 105.235 44.350 105.405 45.140 ;
        RECT 103.960 43.730 104.130 44.060 ;
        RECT 105.225 43.640 105.405 44.350 ;
        RECT 104.505 42.330 105.405 43.640 ;
        RECT 105.895 43.000 106.095 46.320 ;
        RECT 106.495 45.880 106.665 47.180 ;
        RECT 106.935 46.140 107.105 47.480 ;
        RECT 106.415 45.520 106.755 45.880 ;
        RECT 107.375 45.840 107.555 47.180 ;
        RECT 121.425 47.115 122.505 56.235 ;
        RECT 129.480 54.575 136.855 54.745 ;
        RECT 124.950 49.135 125.665 49.160 ;
        RECT 124.900 48.595 125.665 49.135 ;
        RECT 107.365 45.745 107.555 45.840 ;
        RECT 109.720 45.745 110.320 45.780 ;
        RECT 106.485 44.970 106.665 45.520 ;
        RECT 107.365 45.210 110.320 45.745 ;
        RECT 106.485 44.120 106.655 44.970 ;
        RECT 106.925 43.260 107.095 45.160 ;
        RECT 107.365 45.010 107.555 45.210 ;
        RECT 109.720 45.180 110.320 45.210 ;
        RECT 107.365 44.120 107.535 45.010 ;
        RECT 106.785 43.080 107.095 43.260 ;
        RECT 107.800 43.095 107.970 43.425 ;
        RECT 120.735 43.355 123.095 47.115 ;
        RECT 108.585 43.130 108.915 43.300 ;
        RECT 104.770 42.170 105.060 42.330 ;
        RECT 105.905 42.010 106.075 43.000 ;
        RECT 105.885 41.400 106.075 42.010 ;
        RECT 106.345 41.830 106.515 43.010 ;
        RECT 106.785 41.970 106.955 43.080 ;
        RECT 106.315 41.570 106.575 41.830 ;
        RECT 105.885 41.060 106.285 41.400 ;
        RECT 124.900 41.370 125.070 48.595 ;
        RECT 127.190 42.030 127.360 48.070 ;
        RECT 129.480 41.370 129.650 54.575 ;
        RECT 136.495 54.310 136.855 54.575 ;
        RECT 134.795 53.870 135.120 53.875 ;
        RECT 131.170 51.555 135.120 53.870 ;
        RECT 130.800 51.385 135.120 51.555 ;
        RECT 130.800 41.640 130.970 51.385 ;
        RECT 131.170 50.900 135.120 51.385 ;
        RECT 131.170 50.885 135.115 50.900 ;
        RECT 131.405 49.380 133.545 50.220 ;
        RECT 134.255 49.255 135.115 50.885 ;
        RECT 133.090 48.670 133.260 48.680 ;
        RECT 136.190 48.670 136.360 54.105 ;
        RECT 133.085 41.635 136.360 48.670 ;
        RECT 124.900 41.200 126.585 41.370 ;
        RECT 98.010 37.010 98.360 39.170 ;
        RECT 126.415 38.345 126.585 41.200 ;
        RECT 127.995 41.200 129.650 41.370 ;
        RECT 127.205 38.360 127.375 40.885 ;
        RECT 127.200 37.995 127.375 38.360 ;
        RECT 127.995 38.345 128.165 41.200 ;
        RECT 128.655 40.320 133.715 40.490 ;
        RECT 128.655 40.315 129.695 40.320 ;
        RECT 128.655 37.995 128.830 40.315 ;
        RECT 129.675 38.045 133.715 38.200 ;
        RECT 129.675 38.030 133.720 38.045 ;
        RECT 125.200 37.430 125.590 37.825 ;
        RECT 127.200 37.820 128.830 37.995 ;
        RECT 130.205 37.280 133.720 38.030 ;
        RECT 130.205 37.270 133.890 37.280 ;
        RECT 127.540 37.115 127.790 37.155 ;
        RECT 127.500 36.945 127.830 37.115 ;
        RECT 127.540 36.905 127.790 36.945 ;
        RECT 98.010 34.350 98.360 36.510 ;
        RECT 128.470 35.915 128.640 35.955 ;
        RECT 128.435 35.670 128.680 35.915 ;
        RECT 128.470 35.625 128.640 35.670 ;
        RECT 130.210 34.295 133.890 37.270 ;
        RECT 130.210 34.270 133.125 34.295 ;
        RECT 131.080 31.500 133.125 34.270 ;
        RECT 135.415 34.065 136.360 41.635 ;
        RECT 136.980 47.080 137.150 54.105 ;
        RECT 137.750 47.080 138.920 56.265 ;
        RECT 139.955 47.080 142.315 47.085 ;
        RECT 136.980 43.325 142.315 47.080 ;
        RECT 136.980 34.065 137.150 43.325 ;
        RECT 135.415 30.125 136.195 34.065 ;
        RECT 135.355 29.215 136.260 30.125 ;
        RECT 111.870 6.505 112.040 10.020 ;
        RECT 112.285 7.110 112.615 7.280 ;
        RECT 111.870 6.335 112.365 6.505 ;
        RECT 90.390 5.685 90.560 5.705 ;
        RECT 87.310 4.690 90.560 5.685 ;
        RECT 90.390 4.665 90.560 4.690 ;
        RECT 90.390 4.000 90.560 4.035 ;
        RECT 84.775 3.005 90.560 4.000 ;
        RECT 90.390 2.995 90.560 3.005 ;
        RECT 90.830 2.995 91.000 5.705 ;
        RECT 91.415 4.910 91.915 5.885 ;
        RECT 92.295 3.320 92.725 4.350 ;
        RECT 112.195 3.240 112.365 6.335 ;
        RECT 90.430 1.680 90.970 2.200 ;
        RECT 112.635 1.700 112.805 6.230 ;
        RECT 113.075 3.240 113.245 10.005 ;
        RECT 133.775 6.655 133.945 9.920 ;
        RECT 134.265 7.460 134.595 7.630 ;
        RECT 133.775 6.485 134.410 6.655 ;
        RECT 113.635 5.735 114.140 6.280 ;
        RECT 113.635 5.355 114.135 5.735 ;
        RECT 114.515 3.765 114.945 4.620 ;
        RECT 134.240 3.235 134.410 6.485 ;
        RECT 113.135 2.980 113.305 3.000 ;
        RECT 113.075 2.690 113.365 2.980 ;
        RECT 113.135 2.670 113.305 2.690 ;
        RECT 112.460 1.220 112.970 1.700 ;
        RECT 134.680 1.695 134.850 6.225 ;
        RECT 135.120 3.235 135.290 9.930 ;
        RECT 155.790 6.695 155.960 10.265 ;
        RECT 156.870 8.665 157.590 9.385 ;
        RECT 156.285 7.440 156.615 7.610 ;
        RECT 155.790 6.525 156.510 6.695 ;
        RECT 135.675 5.345 136.175 6.320 ;
        RECT 154.320 5.080 154.820 6.245 ;
        RECT 136.555 3.755 136.985 4.835 ;
        RECT 155.200 3.950 155.635 4.450 ;
        RECT 155.200 3.570 155.630 3.950 ;
        RECT 156.340 3.235 156.510 6.525 ;
        RECT 135.180 2.930 135.350 2.950 ;
        RECT 135.120 2.640 135.410 2.930 ;
        RECT 135.180 2.620 135.350 2.640 ;
        RECT 156.780 1.695 156.950 6.225 ;
        RECT 157.220 3.235 157.390 8.665 ;
        RECT 157.280 2.930 157.450 2.950 ;
        RECT 157.220 2.640 157.510 2.930 ;
        RECT 157.280 2.620 157.450 2.640 ;
        RECT 134.505 1.215 135.015 1.695 ;
        RECT 156.605 1.215 157.115 1.695 ;
      LAYER mcon ;
        RECT 105.435 55.985 105.605 56.155 ;
        RECT 98.085 51.285 98.275 53.270 ;
        RECT 98.085 48.630 98.275 50.615 ;
        RECT 121.585 55.595 122.325 56.145 ;
        RECT 105.035 46.220 105.205 47.100 ;
        RECT 105.475 46.220 105.645 47.100 ;
        RECT 105.915 46.220 106.085 47.100 ;
        RECT 104.795 44.180 104.965 45.060 ;
        RECT 105.235 44.180 105.405 45.060 ;
        RECT 103.960 43.810 104.130 43.980 ;
        RECT 106.495 46.220 106.665 47.100 ;
        RECT 106.935 46.220 107.105 47.100 ;
        RECT 137.890 55.450 138.745 55.995 ;
        RECT 107.375 46.220 107.545 47.100 ;
        RECT 109.780 45.240 110.255 45.715 ;
        RECT 106.485 44.200 106.655 45.080 ;
        RECT 106.925 44.200 107.095 45.080 ;
        RECT 107.365 44.200 107.535 45.080 ;
        RECT 107.800 43.175 107.970 43.345 ;
        RECT 108.665 43.130 108.835 43.300 ;
        RECT 104.830 42.200 105.000 42.370 ;
        RECT 105.905 42.050 106.075 42.930 ;
        RECT 106.345 42.050 106.515 42.930 ;
        RECT 106.785 42.050 106.955 42.930 ;
        RECT 124.900 42.110 125.070 47.990 ;
        RECT 106.345 41.600 106.515 41.770 ;
        RECT 127.190 42.110 127.360 47.990 ;
        RECT 129.480 42.110 129.650 47.990 ;
        RECT 132.945 49.555 133.405 50.030 ;
        RECT 134.425 49.370 134.960 49.910 ;
        RECT 130.800 41.720 130.970 48.600 ;
        RECT 133.090 41.720 133.260 48.600 ;
        RECT 98.090 37.095 98.280 39.080 ;
        RECT 126.415 38.425 126.585 40.805 ;
        RECT 127.205 38.425 127.375 40.805 ;
        RECT 127.995 38.425 128.165 40.805 ;
        RECT 129.755 40.320 133.635 40.490 ;
        RECT 129.755 38.030 133.635 38.200 ;
        RECT 125.270 37.500 125.520 37.750 ;
        RECT 98.090 34.440 98.280 36.425 ;
        RECT 131.495 31.685 132.590 32.465 ;
        RECT 136.190 34.145 136.360 54.025 ;
        RECT 136.980 34.145 137.150 54.025 ;
        RECT 135.415 29.280 136.195 30.060 ;
        RECT 155.790 10.095 155.960 10.265 ;
        RECT 111.870 9.845 112.040 10.015 ;
        RECT 113.075 9.835 113.245 10.005 ;
        RECT 112.365 7.110 112.535 7.280 ;
        RECT 87.340 4.690 88.335 5.685 ;
        RECT 90.390 4.745 90.560 5.625 ;
        RECT 90.830 4.745 91.000 5.625 ;
        RECT 91.415 5.385 91.915 5.885 ;
        RECT 112.195 5.270 112.365 6.150 ;
        RECT 84.805 3.035 85.740 3.970 ;
        RECT 90.390 3.075 90.560 3.955 ;
        RECT 90.830 3.075 91.000 3.955 ;
        RECT 92.295 3.920 92.725 4.350 ;
        RECT 112.195 3.320 112.365 4.200 ;
        RECT 112.635 5.270 112.805 6.150 ;
        RECT 112.635 3.320 112.805 4.200 ;
        RECT 90.610 1.860 90.780 2.030 ;
        RECT 133.775 9.750 133.945 9.920 ;
        RECT 135.120 9.760 135.290 9.930 ;
        RECT 134.345 7.460 134.515 7.630 ;
        RECT 113.075 5.270 113.245 6.150 ;
        RECT 113.635 5.775 114.140 6.280 ;
        RECT 134.240 5.265 134.410 6.145 ;
        RECT 113.075 3.320 113.245 4.200 ;
        RECT 114.515 4.190 114.945 4.620 ;
        RECT 134.240 3.315 134.410 4.195 ;
        RECT 134.680 5.265 134.850 6.145 ;
        RECT 134.680 3.315 134.850 4.195 ;
        RECT 113.135 2.750 113.305 2.920 ;
        RECT 156.365 7.440 156.535 7.610 ;
        RECT 135.120 5.265 135.290 6.145 ;
        RECT 135.675 5.820 136.175 6.320 ;
        RECT 154.320 5.745 154.820 6.245 ;
        RECT 156.340 5.265 156.510 6.145 ;
        RECT 135.120 3.315 135.290 4.195 ;
        RECT 136.555 4.405 136.985 4.835 ;
        RECT 155.200 4.015 155.635 4.450 ;
        RECT 156.340 3.315 156.510 4.195 ;
        RECT 156.780 5.265 156.950 6.145 ;
        RECT 156.780 3.315 156.950 4.195 ;
        RECT 135.180 2.700 135.350 2.870 ;
        RECT 157.220 5.265 157.390 6.145 ;
        RECT 157.220 3.315 157.390 4.195 ;
        RECT 157.280 2.700 157.450 2.870 ;
        RECT 112.635 1.365 112.805 1.535 ;
        RECT 134.680 1.360 134.850 1.530 ;
        RECT 156.780 1.360 156.950 1.530 ;
      LAYER met1 ;
        RECT 98.525 142.685 100.525 172.685 ;
        RECT 99.805 56.725 101.390 56.775 ;
        RECT 98.005 56.670 98.355 56.675 ;
        RECT 97.680 56.555 98.795 56.670 ;
        RECT 97.640 55.315 98.845 56.555 ;
        RECT 98.005 53.360 98.355 55.315 ;
        RECT 99.805 55.245 139.210 56.725 ;
        RECT 99.805 55.240 121.115 55.245 ;
        RECT 99.805 55.190 101.390 55.240 ;
        RECT 98.055 51.225 98.305 53.360 ;
        RECT 98.055 48.625 98.305 50.675 ;
        RECT 98.010 43.980 98.360 48.625 ;
        RECT 105.005 46.160 105.235 47.160 ;
        RECT 105.445 46.160 105.675 47.160 ;
        RECT 105.885 46.160 106.115 47.160 ;
        RECT 106.465 46.160 106.695 47.160 ;
        RECT 106.905 46.160 107.135 47.160 ;
        RECT 107.345 46.160 107.575 47.160 ;
        RECT 109.720 45.180 110.320 45.780 ;
        RECT 104.765 44.120 104.995 45.120 ;
        RECT 105.205 44.120 105.435 45.120 ;
        RECT 106.455 44.140 106.685 45.140 ;
        RECT 106.895 44.140 107.125 45.140 ;
        RECT 107.335 44.140 107.565 45.140 ;
        RECT 103.875 43.980 104.210 44.065 ;
        RECT 98.010 43.810 104.210 43.980 ;
        RECT 98.010 39.170 98.360 43.810 ;
        RECT 103.875 43.730 104.210 43.810 ;
        RECT 107.720 43.100 108.055 43.430 ;
        RECT 108.585 43.050 108.920 43.380 ;
        RECT 104.770 42.370 105.060 42.400 ;
        RECT 104.770 42.200 105.720 42.370 ;
        RECT 104.770 42.170 105.060 42.200 ;
        RECT 105.515 41.770 105.720 42.200 ;
        RECT 105.875 41.990 106.105 42.990 ;
        RECT 106.315 41.990 106.545 42.990 ;
        RECT 106.755 41.990 106.985 42.990 ;
        RECT 106.315 41.770 106.575 41.830 ;
        RECT 105.515 41.600 106.575 41.770 ;
        RECT 98.060 37.035 98.310 39.170 ;
        RECT 98.060 34.350 98.310 36.485 ;
        RECT 98.010 32.350 98.360 34.350 ;
        RECT 99.810 32.650 101.395 32.710 ;
        RECT 105.515 32.650 105.685 41.600 ;
        RECT 106.315 41.570 106.575 41.600 ;
        RECT 123.620 35.915 123.865 55.245 ;
        RECT 124.870 42.050 125.100 48.050 ;
        RECT 126.860 41.705 127.675 55.245 ;
        RECT 132.865 49.380 133.585 55.245 ;
        RECT 129.450 42.050 129.680 48.050 ;
        RECT 130.770 41.660 131.000 48.660 ;
        RECT 133.060 41.660 133.290 48.660 ;
        RECT 126.385 38.365 126.615 40.865 ;
        RECT 127.175 38.365 127.405 40.865 ;
        RECT 127.965 38.365 128.195 40.865 ;
        RECT 129.695 40.290 133.695 40.520 ;
        RECT 129.695 38.000 133.695 38.230 ;
        RECT 125.200 37.430 125.590 37.825 ;
        RECT 127.465 36.845 127.870 37.235 ;
        RECT 128.405 35.915 128.710 35.975 ;
        RECT 123.620 35.670 128.710 35.915 ;
        RECT 128.405 35.610 128.710 35.670 ;
        RECT 131.495 32.650 132.815 32.680 ;
        RECT 134.255 32.650 135.110 50.130 ;
        RECT 136.160 34.085 136.390 54.085 ;
        RECT 136.950 34.085 137.180 54.085 ;
        RECT 97.660 31.230 98.800 32.350 ;
        RECT 99.810 31.170 139.345 32.650 ;
        RECT 99.810 31.165 124.195 31.170 ;
        RECT 99.810 31.115 101.395 31.165 ;
        RECT 135.355 29.215 136.260 30.125 ;
        RECT 113.000 25.965 113.320 26.010 ;
        RECT 125.255 25.965 125.515 26.040 ;
        RECT 113.000 25.795 125.515 25.965 ;
        RECT 113.000 25.750 113.320 25.795 ;
        RECT 125.255 25.720 125.515 25.795 ;
        RECT 114.440 24.295 114.720 24.380 ;
        RECT 133.700 24.295 134.020 24.340 ;
        RECT 114.440 24.125 134.020 24.295 ;
        RECT 114.440 24.040 114.720 24.125 ;
        RECT 133.700 24.080 134.020 24.125 ;
        RECT 117.325 21.825 117.585 21.900 ;
        RECT 155.745 21.825 156.005 21.900 ;
        RECT 117.325 21.655 156.005 21.825 ;
        RECT 117.325 21.580 117.585 21.655 ;
        RECT 155.745 21.580 156.005 21.655 ;
        RECT 155.760 10.310 155.990 10.325 ;
        RECT 111.795 9.770 112.115 10.090 ;
        RECT 113.000 9.760 113.320 10.080 ;
        RECT 155.715 10.050 156.035 10.310 ;
        RECT 155.760 10.035 155.990 10.050 ;
        RECT 133.700 9.675 134.020 9.995 ;
        RECT 135.045 9.685 135.365 10.005 ;
        RECT 156.810 8.635 157.650 9.415 ;
        RECT 90.800 8.245 156.535 8.475 ;
        RECT 87.265 4.615 88.430 5.765 ;
        RECT 90.360 4.685 90.590 5.685 ;
        RECT 90.800 4.685 91.030 8.245 ;
        RECT 112.365 7.360 112.535 8.245 ;
        RECT 134.345 7.710 134.515 8.245 ;
        RECT 134.265 7.380 134.595 7.710 ;
        RECT 156.365 7.690 156.535 8.245 ;
        RECT 156.285 7.360 156.615 7.690 ;
        RECT 112.285 7.030 112.615 7.360 ;
        RECT 91.355 5.325 91.980 5.960 ;
        RECT 112.165 5.210 112.395 6.210 ;
        RECT 112.605 5.210 112.835 6.210 ;
        RECT 113.045 5.210 113.275 6.210 ;
        RECT 113.560 5.700 114.215 6.360 ;
        RECT 134.210 5.205 134.440 6.205 ;
        RECT 134.650 5.205 134.880 6.205 ;
        RECT 135.090 5.205 135.320 6.205 ;
        RECT 135.600 5.745 136.250 6.395 ;
        RECT 154.245 5.670 154.895 6.320 ;
        RECT 156.310 5.205 156.540 6.205 ;
        RECT 156.750 5.205 156.980 6.205 ;
        RECT 157.190 5.205 157.420 6.205 ;
        RECT 84.745 2.975 85.805 4.035 ;
        RECT 90.360 3.015 90.590 4.015 ;
        RECT 90.800 3.015 91.030 4.015 ;
        RECT 92.220 3.840 92.800 4.435 ;
        RECT 112.165 3.260 112.395 4.260 ;
        RECT 112.605 3.260 112.835 4.260 ;
        RECT 113.045 3.260 113.275 4.260 ;
        RECT 114.440 4.115 115.020 4.705 ;
        RECT 136.470 4.320 137.070 4.920 ;
        RECT 134.210 3.255 134.440 4.255 ;
        RECT 134.650 3.255 134.880 4.255 ;
        RECT 135.090 3.255 135.320 4.255 ;
        RECT 155.110 3.930 155.720 4.535 ;
        RECT 156.310 3.255 156.540 4.255 ;
        RECT 156.750 3.255 156.980 4.255 ;
        RECT 157.190 3.255 157.420 4.255 ;
        RECT 113.075 2.575 113.365 2.980 ;
        RECT 135.120 2.575 135.410 2.930 ;
        RECT 157.220 2.575 157.510 2.930 ;
        RECT 90.430 2.285 157.510 2.575 ;
        RECT 90.430 1.680 90.970 2.285 ;
        RECT 112.460 1.220 112.970 1.700 ;
        RECT 134.505 1.215 135.015 1.695 ;
        RECT 156.605 1.215 157.115 1.695 ;
      LAYER via ;
        RECT 99.030 171.105 100.005 172.170 ;
        RECT 99.050 143.170 100.025 144.235 ;
        RECT 97.680 55.375 98.795 56.490 ;
        RECT 99.860 55.240 101.345 56.725 ;
        RECT 109.750 45.210 110.285 45.745 ;
        RECT 107.755 43.130 108.015 43.390 ;
        RECT 108.620 43.085 108.880 43.345 ;
        RECT 125.240 37.470 125.550 37.780 ;
        RECT 127.510 36.875 127.820 37.185 ;
        RECT 97.730 31.280 98.750 32.300 ;
        RECT 99.860 31.165 101.345 32.650 ;
        RECT 135.385 29.250 136.225 30.090 ;
        RECT 113.030 25.750 113.290 26.010 ;
        RECT 125.255 25.750 125.515 26.010 ;
        RECT 114.440 24.070 114.720 24.350 ;
        RECT 133.730 24.080 133.990 24.340 ;
        RECT 117.325 21.610 117.585 21.870 ;
        RECT 155.745 21.610 156.005 21.870 ;
        RECT 111.825 9.800 112.085 10.060 ;
        RECT 155.745 10.050 156.005 10.310 ;
        RECT 113.030 9.790 113.290 10.050 ;
        RECT 133.730 9.705 133.990 9.965 ;
        RECT 135.075 9.715 135.335 9.975 ;
        RECT 156.840 8.635 157.620 9.415 ;
        RECT 87.310 4.660 88.365 5.715 ;
        RECT 91.385 5.355 91.945 5.915 ;
        RECT 113.605 5.745 114.170 6.310 ;
        RECT 135.645 5.790 136.205 6.350 ;
        RECT 154.290 5.715 154.850 6.275 ;
        RECT 84.775 3.005 85.770 4.000 ;
        RECT 92.265 3.890 92.755 4.380 ;
        RECT 114.485 4.160 114.975 4.650 ;
        RECT 136.525 4.375 137.015 4.865 ;
        RECT 155.170 3.985 155.665 4.480 ;
        RECT 90.565 1.815 90.825 2.075 ;
        RECT 112.590 1.320 112.850 1.580 ;
        RECT 134.635 1.315 134.895 1.575 ;
        RECT 156.735 1.315 156.995 1.575 ;
      LAYER met2 ;
        RECT 98.525 170.685 100.525 172.685 ;
        RECT 98.525 142.685 100.525 144.685 ;
        RECT 97.640 55.315 98.845 56.555 ;
        RECT 99.805 55.190 101.390 56.775 ;
        RECT 109.720 45.180 110.320 45.780 ;
        RECT 103.190 38.430 103.830 39.055 ;
        RECT 97.660 31.230 98.800 32.350 ;
        RECT 99.810 31.115 101.395 32.710 ;
        RECT 103.230 26.020 103.765 38.430 ;
        RECT 107.720 27.300 108.055 43.430 ;
        RECT 108.590 30.325 108.915 43.380 ;
        RECT 108.590 29.970 117.540 30.325 ;
        RECT 107.720 27.020 114.720 27.300 ;
        RECT 103.230 25.745 112.045 26.020 ;
        RECT 111.870 10.090 112.040 25.745 ;
        RECT 113.030 25.720 113.290 26.040 ;
        RECT 111.795 9.770 112.115 10.090 ;
        RECT 113.075 10.080 113.245 25.720 ;
        RECT 114.440 24.350 114.720 27.020 ;
        RECT 114.410 24.070 114.750 24.350 ;
        RECT 117.295 21.870 117.540 29.970 ;
        RECT 125.090 29.835 125.700 37.930 ;
        RECT 125.225 25.720 125.550 29.835 ;
        RECT 127.465 25.255 127.870 37.235 ;
        RECT 135.355 30.060 136.260 30.125 ;
        RECT 135.355 29.280 157.620 30.060 ;
        RECT 135.355 29.215 136.260 29.280 ;
        RECT 127.465 24.895 135.345 25.255 ;
        RECT 127.465 24.890 127.830 24.895 ;
        RECT 133.730 24.050 133.990 24.370 ;
        RECT 117.295 21.610 117.615 21.870 ;
        RECT 113.000 9.760 113.320 10.080 ;
        RECT 133.775 9.995 133.945 24.050 ;
        RECT 135.065 10.005 135.345 24.895 ;
        RECT 155.715 21.610 156.035 21.870 ;
        RECT 155.790 10.340 155.960 21.610 ;
        RECT 155.745 10.020 156.005 10.340 ;
        RECT 133.700 9.675 134.020 9.995 ;
        RECT 135.045 9.685 135.365 10.005 ;
        RECT 156.840 8.605 157.620 29.280 ;
        RECT 87.265 4.615 88.430 5.765 ;
        RECT 91.355 5.325 91.980 5.960 ;
        RECT 113.560 5.700 114.215 6.360 ;
        RECT 135.600 5.745 136.250 6.395 ;
        RECT 154.245 5.670 154.895 6.320 ;
        RECT 84.745 2.975 85.805 4.035 ;
        RECT 92.220 3.840 92.800 4.435 ;
        RECT 114.440 4.115 115.020 4.705 ;
        RECT 136.470 4.320 137.070 4.920 ;
        RECT 155.110 3.930 155.720 4.535 ;
        RECT 90.430 1.680 90.970 2.200 ;
        RECT 112.460 1.220 112.970 1.700 ;
        RECT 134.505 1.215 135.015 1.695 ;
        RECT 156.605 1.215 157.115 1.695 ;
      LAYER via2 ;
        RECT 99.030 171.105 100.005 172.170 ;
        RECT 99.050 143.170 100.025 144.235 ;
        RECT 97.680 55.375 98.795 56.490 ;
        RECT 99.860 55.240 101.345 56.725 ;
        RECT 109.775 45.235 110.260 45.720 ;
        RECT 103.230 38.465 103.765 39.000 ;
        RECT 97.730 31.280 98.750 32.300 ;
        RECT 99.860 31.165 101.345 32.650 ;
        RECT 87.310 4.660 88.365 5.715 ;
        RECT 91.385 5.415 91.945 5.915 ;
        RECT 113.605 5.745 114.170 6.310 ;
        RECT 135.645 5.790 136.205 6.350 ;
        RECT 154.290 5.715 154.850 6.275 ;
        RECT 84.800 3.030 85.745 3.975 ;
        RECT 92.265 3.890 92.755 4.380 ;
        RECT 114.485 4.160 114.975 4.650 ;
        RECT 136.525 4.375 137.015 4.865 ;
        RECT 155.170 3.985 155.665 4.480 ;
        RECT 90.545 1.795 90.845 2.095 ;
        RECT 112.570 1.300 112.870 1.600 ;
        RECT 134.615 1.295 134.915 1.595 ;
        RECT 156.715 1.295 157.015 1.595 ;
      LAYER met3 ;
        RECT 98.525 170.685 100.525 172.685 ;
        RECT 98.525 142.685 100.525 144.685 ;
        RECT 48.970 135.650 100.525 135.655 ;
        RECT 48.970 133.660 100.550 135.650 ;
        RECT 48.970 133.655 100.525 133.660 ;
        RECT 99.835 56.725 101.370 56.750 ;
        RECT 49.005 55.240 101.370 56.725 ;
        RECT 99.835 55.215 101.370 55.240 ;
        RECT 19.220 46.145 21.760 46.815 ;
        RECT 19.220 45.505 50.265 46.145 ;
        RECT 19.220 44.765 21.760 45.505 ;
        RECT 103.205 39.000 103.790 39.025 ;
        RECT 109.750 39.000 110.285 45.745 ;
        RECT 103.205 38.465 110.285 39.000 ;
        RECT 103.205 38.440 103.790 38.465 ;
        RECT 99.835 32.650 101.370 32.675 ;
        RECT 48.970 31.165 101.370 32.650 ;
        RECT 99.835 31.140 101.370 31.165 ;
        RECT 19.220 18.715 21.770 19.365 ;
        RECT 19.220 18.710 43.660 18.715 ;
        RECT 19.220 17.820 43.685 18.710 ;
        RECT 19.220 17.815 43.660 17.820 ;
        RECT 19.220 17.305 21.770 17.815 ;
        RECT 1.000 8.230 155.640 9.350 ;
        RECT 49.000 6.360 85.770 7.355 ;
        RECT 84.775 3.005 85.770 6.360 ;
        RECT 87.310 5.740 88.430 8.230 ;
        RECT 91.415 5.960 91.915 8.230 ;
        RECT 113.635 6.335 114.140 8.230 ;
        RECT 135.675 6.375 136.175 8.230 ;
        RECT 87.285 4.690 88.430 5.740 ;
        RECT 91.355 5.325 91.980 5.960 ;
        RECT 113.580 5.720 114.195 6.335 ;
        RECT 135.620 5.765 136.230 6.375 ;
        RECT 154.320 6.300 154.820 8.230 ;
        RECT 154.265 5.690 154.875 6.300 ;
        RECT 87.285 4.635 88.390 4.690 ;
        RECT 92.220 3.840 92.800 4.435 ;
        RECT 114.460 4.135 115.000 4.705 ;
        RECT 136.470 4.320 137.070 4.920 ;
        RECT 155.110 3.930 155.720 4.535 ;
        RECT 90.430 1.680 90.970 2.200 ;
        RECT 112.460 1.220 112.970 1.700 ;
        RECT 134.505 1.215 135.015 1.695 ;
        RECT 156.605 1.215 157.115 1.695 ;
      LAYER via3 ;
        RECT 99.030 171.105 100.005 172.170 ;
        RECT 99.050 143.170 100.025 144.235 ;
        RECT 49.000 133.655 51.000 135.655 ;
        RECT 98.530 133.660 100.520 135.650 ;
        RECT 49.035 55.240 50.520 56.725 ;
        RECT 19.840 45.255 21.120 46.425 ;
        RECT 49.595 45.505 50.235 46.145 ;
        RECT 49.000 31.165 50.485 32.650 ;
        RECT 19.860 17.735 21.140 18.905 ;
        RECT 42.765 17.820 43.655 18.710 ;
        RECT 1.215 8.260 2.275 9.320 ;
        RECT 49.300 6.440 50.025 7.230 ;
        RECT 84.705 6.360 85.710 7.355 ;
        RECT 92.240 3.975 92.780 4.405 ;
        RECT 114.460 4.245 115.000 4.675 ;
        RECT 136.500 4.350 137.040 4.890 ;
        RECT 155.145 3.960 155.690 4.505 ;
        RECT 90.520 1.770 90.870 2.120 ;
        RECT 112.545 1.275 112.895 1.625 ;
        RECT 134.590 1.270 134.940 1.620 ;
        RECT 156.690 1.270 157.040 1.620 ;
      LAYER met4 ;
        RECT 73.525 214.685 139.525 216.685 ;
        RECT 73.525 144.685 75.525 214.685 ;
        RECT 80.525 207.685 132.525 209.685 ;
        RECT 80.525 151.685 82.525 207.685 ;
        RECT 87.525 199.685 125.525 201.685 ;
        RECT 87.525 158.685 89.525 199.685 ;
        RECT 94.525 192.685 118.525 194.685 ;
        RECT 94.525 165.685 96.525 192.685 ;
        RECT 100.525 172.685 100.945 172.690 ;
        RECT 116.525 172.685 118.525 192.685 ;
        RECT 98.525 170.685 118.525 172.685 ;
        RECT 123.525 165.685 125.525 199.685 ;
        RECT 94.525 163.685 125.525 165.685 ;
        RECT 130.525 158.685 132.525 207.685 ;
        RECT 87.525 156.685 132.525 158.685 ;
        RECT 137.515 151.685 139.525 214.685 ;
        RECT 80.525 149.685 139.525 151.685 ;
        RECT 73.525 142.685 96.525 144.685 ;
        RECT 48.995 133.650 49.000 135.660 ;
        RECT 50.500 133.650 51.005 135.660 ;
        RECT 94.525 129.775 96.525 142.685 ;
        RECT 98.525 133.655 100.525 144.685 ;
        RECT 57.690 127.775 96.525 129.775 ;
        RECT 50.500 55.235 50.525 56.730 ;
        RECT 19.220 19.365 21.760 46.815 ;
        RECT 48.995 31.160 49.000 32.655 ;
        RECT 19.220 17.305 21.770 19.365 ;
        RECT 42.760 1.000 43.660 18.715 ;
        RECT 57.690 5.250 59.690 127.775 ;
        RECT 84.700 7.355 85.715 7.360 ;
        RECT 84.700 6.360 155.635 7.355 ;
        RECT 84.700 6.355 85.715 6.360 ;
        RECT 57.690 3.250 68.990 5.250 ;
        RECT 92.295 4.435 92.725 6.360 ;
        RECT 114.515 4.680 114.945 6.360 ;
        RECT 136.555 4.895 136.985 6.360 ;
        RECT 92.220 3.840 92.800 4.435 ;
        RECT 114.455 4.240 115.005 4.680 ;
        RECT 136.495 4.345 137.045 4.895 ;
        RECT 155.200 4.510 155.635 6.360 ;
        RECT 155.140 3.955 155.695 4.510 ;
        RECT 68.090 1.000 68.990 3.250 ;
        RECT 90.430 1.680 90.970 2.200 ;
        RECT 90.545 1.000 90.845 1.680 ;
        RECT 112.460 1.000 112.970 1.700 ;
        RECT 134.505 1.000 135.015 1.695 ;
        RECT 156.605 1.000 157.115 1.695 ;
        RECT 42.760 0.100 46.010 1.000 ;
  END
END tt_um_analog_rf_readout_circuit
END LIBRARY

