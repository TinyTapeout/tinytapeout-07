VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_mux
  CLASS BLOCK ;
  FOREIGN tt_mux ;
  ORIGIN 0.000 0.000 ;
  SIZE 1359.760 BY 54.400 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 402.280 2.480 403.880 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 555.880 2.480 557.480 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 709.480 2.480 711.080 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.080 2.480 864.680 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1016.680 2.480 1018.280 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1170.280 2.480 1171.880 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1323.880 2.480 1325.480 51.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 479.080 2.480 480.680 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.680 2.480 634.280 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.280 2.480 787.880 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 939.880 2.480 941.480 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1093.480 2.480 1095.080 51.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1247.080 2.480 1248.680 51.920 ;
    END
  END VPWR
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 47.110 1359.760 47.410 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 46.430 1359.760 46.730 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 45.750 1359.760 46.050 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 45.070 1359.760 45.370 ;
    END
  END addr[3]
  PIN k_one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1358.760 44.390 1359.760 44.690 ;
    END
  END k_one
  PIN k_zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1358.760 43.710 1359.760 44.010 ;
    END
  END k_zero
  PIN spine_iw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 43.030 1359.760 43.330 ;
    END
  END spine_iw[0]
  PIN spine_iw[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 36.230 1359.760 36.530 ;
    END
  END spine_iw[10]
  PIN spine_iw[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 35.550 1359.760 35.850 ;
    END
  END spine_iw[11]
  PIN spine_iw[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 34.870 1359.760 35.170 ;
    END
  END spine_iw[12]
  PIN spine_iw[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 34.190 1359.760 34.490 ;
    END
  END spine_iw[13]
  PIN spine_iw[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 33.510 1359.760 33.810 ;
    END
  END spine_iw[14]
  PIN spine_iw[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 32.830 1359.760 33.130 ;
    END
  END spine_iw[15]
  PIN spine_iw[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 32.150 1359.760 32.450 ;
    END
  END spine_iw[16]
  PIN spine_iw[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 31.470 1359.760 31.770 ;
    END
  END spine_iw[17]
  PIN spine_iw[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 30.790 1359.760 31.090 ;
    END
  END spine_iw[18]
  PIN spine_iw[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 30.110 1359.760 30.410 ;
    END
  END spine_iw[19]
  PIN spine_iw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 42.350 1359.760 42.650 ;
    END
  END spine_iw[1]
  PIN spine_iw[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 29.430 1359.760 29.730 ;
    END
  END spine_iw[20]
  PIN spine_iw[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 28.750 1359.760 29.050 ;
    END
  END spine_iw[21]
  PIN spine_iw[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 28.070 1359.760 28.370 ;
    END
  END spine_iw[22]
  PIN spine_iw[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 27.390 1359.760 27.690 ;
    END
  END spine_iw[23]
  PIN spine_iw[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 26.710 1359.760 27.010 ;
    END
  END spine_iw[24]
  PIN spine_iw[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 26.030 1359.760 26.330 ;
    END
  END spine_iw[25]
  PIN spine_iw[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 25.350 1359.760 25.650 ;
    END
  END spine_iw[26]
  PIN spine_iw[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 24.670 1359.760 24.970 ;
    END
  END spine_iw[27]
  PIN spine_iw[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 23.990 1359.760 24.290 ;
    END
  END spine_iw[28]
  PIN spine_iw[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 23.310 1359.760 23.610 ;
    END
  END spine_iw[29]
  PIN spine_iw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 41.670 1359.760 41.970 ;
    END
  END spine_iw[2]
  PIN spine_iw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 40.990 1359.760 41.290 ;
    END
  END spine_iw[3]
  PIN spine_iw[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 40.310 1359.760 40.610 ;
    END
  END spine_iw[4]
  PIN spine_iw[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 39.630 1359.760 39.930 ;
    END
  END spine_iw[5]
  PIN spine_iw[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 38.950 1359.760 39.250 ;
    END
  END spine_iw[6]
  PIN spine_iw[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 38.270 1359.760 38.570 ;
    END
  END spine_iw[7]
  PIN spine_iw[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 37.590 1359.760 37.890 ;
    END
  END spine_iw[8]
  PIN spine_iw[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 36.910 1359.760 37.210 ;
    END
  END spine_iw[9]
  PIN spine_ow[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1358.760 22.630 1359.760 22.930 ;
    END
  END spine_ow[0]
  PIN spine_ow[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 15.830 1359.760 16.130 ;
    END
  END spine_ow[10]
  PIN spine_ow[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 15.150 1359.760 15.450 ;
    END
  END spine_ow[11]
  PIN spine_ow[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 14.470 1359.760 14.770 ;
    END
  END spine_ow[12]
  PIN spine_ow[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 13.790 1359.760 14.090 ;
    END
  END spine_ow[13]
  PIN spine_ow[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 13.110 1359.760 13.410 ;
    END
  END spine_ow[14]
  PIN spine_ow[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 12.430 1359.760 12.730 ;
    END
  END spine_ow[15]
  PIN spine_ow[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 11.750 1359.760 12.050 ;
    END
  END spine_ow[16]
  PIN spine_ow[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 11.070 1359.760 11.370 ;
    END
  END spine_ow[17]
  PIN spine_ow[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 10.390 1359.760 10.690 ;
    END
  END spine_ow[18]
  PIN spine_ow[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 9.710 1359.760 10.010 ;
    END
  END spine_ow[19]
  PIN spine_ow[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 21.950 1359.760 22.250 ;
    END
  END spine_ow[1]
  PIN spine_ow[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 9.030 1359.760 9.330 ;
    END
  END spine_ow[20]
  PIN spine_ow[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 8.350 1359.760 8.650 ;
    END
  END spine_ow[21]
  PIN spine_ow[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 7.670 1359.760 7.970 ;
    END
  END spine_ow[22]
  PIN spine_ow[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 6.990 1359.760 7.290 ;
    END
  END spine_ow[23]
  PIN spine_ow[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 6.310 1359.760 6.610 ;
    END
  END spine_ow[24]
  PIN spine_ow[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1358.760 5.630 1359.760 5.930 ;
    END
  END spine_ow[25]
  PIN spine_ow[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 21.270 1359.760 21.570 ;
    END
  END spine_ow[2]
  PIN spine_ow[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 20.590 1359.760 20.890 ;
    END
  END spine_ow[3]
  PIN spine_ow[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 19.910 1359.760 20.210 ;
    END
  END spine_ow[4]
  PIN spine_ow[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 19.230 1359.760 19.530 ;
    END
  END spine_ow[5]
  PIN spine_ow[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 18.550 1359.760 18.850 ;
    END
  END spine_ow[6]
  PIN spine_ow[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 17.870 1359.760 18.170 ;
    END
  END spine_ow[7]
  PIN spine_ow[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 17.190 1359.760 17.490 ;
    END
  END spine_ow[8]
  PIN spine_ow[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 1358.760 16.510 1359.760 16.810 ;
    END
  END spine_ow[9]
  PIN um_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1339.830 53.400 1340.130 54.400 ;
    END
  END um_ena[0]
  PIN um_ena[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 488.830 53.400 489.130 54.400 ;
    END
  END um_ena[10]
  PIN um_ena[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 488.830 0.000 489.130 1.000 ;
    END
  END um_ena[11]
  PIN um_ena[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 318.630 53.400 318.930 54.400 ;
    END
  END um_ena[12]
  PIN um_ena[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 318.630 0.000 318.930 1.000 ;
    END
  END um_ena[13]
  PIN um_ena[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 148.430 53.400 148.730 54.400 ;
    END
  END um_ena[14]
  PIN um_ena[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 148.430 0.000 148.730 1.000 ;
    END
  END um_ena[15]
  PIN um_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1339.830 0.000 1340.130 1.000 ;
    END
  END um_ena[1]
  PIN um_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1169.630 53.400 1169.930 54.400 ;
    END
  END um_ena[2]
  PIN um_ena[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1169.630 0.000 1169.930 1.000 ;
    END
  END um_ena[3]
  PIN um_ena[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 999.430 53.400 999.730 54.400 ;
    END
  END um_ena[4]
  PIN um_ena[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 999.430 0.000 999.730 1.000 ;
    END
  END um_ena[5]
  PIN um_ena[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 829.230 53.400 829.530 54.400 ;
    END
  END um_ena[6]
  PIN um_ena[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 829.230 0.000 829.530 1.000 ;
    END
  END um_ena[7]
  PIN um_ena[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 659.030 53.400 659.330 54.400 ;
    END
  END um_ena[8]
  PIN um_ena[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 659.030 0.000 659.330 1.000 ;
    END
  END um_ena[9]
  PIN um_iw[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1337.070 53.400 1337.370 54.400 ;
    END
  END um_iw[0]
  PIN um_iw[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 969.070 0.000 969.370 1.000 ;
    END
  END um_iw[100]
  PIN um_iw[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 966.310 0.000 966.610 1.000 ;
    END
  END um_iw[101]
  PIN um_iw[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 963.550 0.000 963.850 1.000 ;
    END
  END um_iw[102]
  PIN um_iw[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 960.790 0.000 961.090 1.000 ;
    END
  END um_iw[103]
  PIN um_iw[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 958.030 0.000 958.330 1.000 ;
    END
  END um_iw[104]
  PIN um_iw[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 955.270 0.000 955.570 1.000 ;
    END
  END um_iw[105]
  PIN um_iw[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 952.510 0.000 952.810 1.000 ;
    END
  END um_iw[106]
  PIN um_iw[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 949.750 0.000 950.050 1.000 ;
    END
  END um_iw[107]
  PIN um_iw[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 826.470 53.400 826.770 54.400 ;
    END
  END um_iw[108]
  PIN um_iw[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 823.710 53.400 824.010 54.400 ;
    END
  END um_iw[109]
  PIN um_iw[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1309.470 53.400 1309.770 54.400 ;
    END
  END um_iw[10]
  PIN um_iw[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 820.950 53.400 821.250 54.400 ;
    END
  END um_iw[110]
  PIN um_iw[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 818.190 53.400 818.490 54.400 ;
    END
  END um_iw[111]
  PIN um_iw[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 815.430 53.400 815.730 54.400 ;
    END
  END um_iw[112]
  PIN um_iw[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 812.670 53.400 812.970 54.400 ;
    END
  END um_iw[113]
  PIN um_iw[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 809.910 53.400 810.210 54.400 ;
    END
  END um_iw[114]
  PIN um_iw[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 807.150 53.400 807.450 54.400 ;
    END
  END um_iw[115]
  PIN um_iw[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 804.390 53.400 804.690 54.400 ;
    END
  END um_iw[116]
  PIN um_iw[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 801.630 53.400 801.930 54.400 ;
    END
  END um_iw[117]
  PIN um_iw[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 798.870 53.400 799.170 54.400 ;
    END
  END um_iw[118]
  PIN um_iw[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 796.110 53.400 796.410 54.400 ;
    END
  END um_iw[119]
  PIN um_iw[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1306.710 53.400 1307.010 54.400 ;
    END
  END um_iw[11]
  PIN um_iw[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 793.350 53.400 793.650 54.400 ;
    END
  END um_iw[120]
  PIN um_iw[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 790.590 53.400 790.890 54.400 ;
    END
  END um_iw[121]
  PIN um_iw[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 787.830 53.400 788.130 54.400 ;
    END
  END um_iw[122]
  PIN um_iw[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 785.070 53.400 785.370 54.400 ;
    END
  END um_iw[123]
  PIN um_iw[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 782.310 53.400 782.610 54.400 ;
    END
  END um_iw[124]
  PIN um_iw[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 779.550 53.400 779.850 54.400 ;
    END
  END um_iw[125]
  PIN um_iw[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 826.470 0.000 826.770 1.000 ;
    END
  END um_iw[126]
  PIN um_iw[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 823.710 0.000 824.010 1.000 ;
    END
  END um_iw[127]
  PIN um_iw[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 820.950 0.000 821.250 1.000 ;
    END
  END um_iw[128]
  PIN um_iw[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 818.190 0.000 818.490 1.000 ;
    END
  END um_iw[129]
  PIN um_iw[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1303.950 53.400 1304.250 54.400 ;
    END
  END um_iw[12]
  PIN um_iw[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 815.430 0.000 815.730 1.000 ;
    END
  END um_iw[130]
  PIN um_iw[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 812.670 0.000 812.970 1.000 ;
    END
  END um_iw[131]
  PIN um_iw[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 809.910 0.000 810.210 1.000 ;
    END
  END um_iw[132]
  PIN um_iw[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 807.150 0.000 807.450 1.000 ;
    END
  END um_iw[133]
  PIN um_iw[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 804.390 0.000 804.690 1.000 ;
    END
  END um_iw[134]
  PIN um_iw[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 801.630 0.000 801.930 1.000 ;
    END
  END um_iw[135]
  PIN um_iw[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 798.870 0.000 799.170 1.000 ;
    END
  END um_iw[136]
  PIN um_iw[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 796.110 0.000 796.410 1.000 ;
    END
  END um_iw[137]
  PIN um_iw[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 793.350 0.000 793.650 1.000 ;
    END
  END um_iw[138]
  PIN um_iw[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 790.590 0.000 790.890 1.000 ;
    END
  END um_iw[139]
  PIN um_iw[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1301.190 53.400 1301.490 54.400 ;
    END
  END um_iw[13]
  PIN um_iw[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 787.830 0.000 788.130 1.000 ;
    END
  END um_iw[140]
  PIN um_iw[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 785.070 0.000 785.370 1.000 ;
    END
  END um_iw[141]
  PIN um_iw[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 782.310 0.000 782.610 1.000 ;
    END
  END um_iw[142]
  PIN um_iw[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 779.550 0.000 779.850 1.000 ;
    END
  END um_iw[143]
  PIN um_iw[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 656.270 53.400 656.570 54.400 ;
    END
  END um_iw[144]
  PIN um_iw[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 653.510 53.400 653.810 54.400 ;
    END
  END um_iw[145]
  PIN um_iw[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 650.750 53.400 651.050 54.400 ;
    END
  END um_iw[146]
  PIN um_iw[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 647.990 53.400 648.290 54.400 ;
    END
  END um_iw[147]
  PIN um_iw[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 645.230 53.400 645.530 54.400 ;
    END
  END um_iw[148]
  PIN um_iw[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 642.470 53.400 642.770 54.400 ;
    END
  END um_iw[149]
  PIN um_iw[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1298.430 53.400 1298.730 54.400 ;
    END
  END um_iw[14]
  PIN um_iw[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 639.710 53.400 640.010 54.400 ;
    END
  END um_iw[150]
  PIN um_iw[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 636.950 53.400 637.250 54.400 ;
    END
  END um_iw[151]
  PIN um_iw[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 634.190 53.400 634.490 54.400 ;
    END
  END um_iw[152]
  PIN um_iw[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 631.430 53.400 631.730 54.400 ;
    END
  END um_iw[153]
  PIN um_iw[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 628.670 53.400 628.970 54.400 ;
    END
  END um_iw[154]
  PIN um_iw[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 625.910 53.400 626.210 54.400 ;
    END
  END um_iw[155]
  PIN um_iw[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 623.150 53.400 623.450 54.400 ;
    END
  END um_iw[156]
  PIN um_iw[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 620.390 53.400 620.690 54.400 ;
    END
  END um_iw[157]
  PIN um_iw[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 617.630 53.400 617.930 54.400 ;
    END
  END um_iw[158]
  PIN um_iw[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 614.870 53.400 615.170 54.400 ;
    END
  END um_iw[159]
  PIN um_iw[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1295.670 53.400 1295.970 54.400 ;
    END
  END um_iw[15]
  PIN um_iw[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 612.110 53.400 612.410 54.400 ;
    END
  END um_iw[160]
  PIN um_iw[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 609.350 53.400 609.650 54.400 ;
    END
  END um_iw[161]
  PIN um_iw[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 656.270 0.000 656.570 1.000 ;
    END
  END um_iw[162]
  PIN um_iw[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 653.510 0.000 653.810 1.000 ;
    END
  END um_iw[163]
  PIN um_iw[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 650.750 0.000 651.050 1.000 ;
    END
  END um_iw[164]
  PIN um_iw[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 647.990 0.000 648.290 1.000 ;
    END
  END um_iw[165]
  PIN um_iw[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 645.230 0.000 645.530 1.000 ;
    END
  END um_iw[166]
  PIN um_iw[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 642.470 0.000 642.770 1.000 ;
    END
  END um_iw[167]
  PIN um_iw[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 639.710 0.000 640.010 1.000 ;
    END
  END um_iw[168]
  PIN um_iw[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 636.950 0.000 637.250 1.000 ;
    END
  END um_iw[169]
  PIN um_iw[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1292.910 53.400 1293.210 54.400 ;
    END
  END um_iw[16]
  PIN um_iw[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 634.190 0.000 634.490 1.000 ;
    END
  END um_iw[170]
  PIN um_iw[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 631.430 0.000 631.730 1.000 ;
    END
  END um_iw[171]
  PIN um_iw[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 628.670 0.000 628.970 1.000 ;
    END
  END um_iw[172]
  PIN um_iw[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 625.910 0.000 626.210 1.000 ;
    END
  END um_iw[173]
  PIN um_iw[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 623.150 0.000 623.450 1.000 ;
    END
  END um_iw[174]
  PIN um_iw[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 620.390 0.000 620.690 1.000 ;
    END
  END um_iw[175]
  PIN um_iw[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 617.630 0.000 617.930 1.000 ;
    END
  END um_iw[176]
  PIN um_iw[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 614.870 0.000 615.170 1.000 ;
    END
  END um_iw[177]
  PIN um_iw[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 612.110 0.000 612.410 1.000 ;
    END
  END um_iw[178]
  PIN um_iw[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 609.350 0.000 609.650 1.000 ;
    END
  END um_iw[179]
  PIN um_iw[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1290.150 53.400 1290.450 54.400 ;
    END
  END um_iw[17]
  PIN um_iw[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 486.070 53.400 486.370 54.400 ;
    END
  END um_iw[180]
  PIN um_iw[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 483.310 53.400 483.610 54.400 ;
    END
  END um_iw[181]
  PIN um_iw[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 480.550 53.400 480.850 54.400 ;
    END
  END um_iw[182]
  PIN um_iw[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 477.790 53.400 478.090 54.400 ;
    END
  END um_iw[183]
  PIN um_iw[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 475.030 53.400 475.330 54.400 ;
    END
  END um_iw[184]
  PIN um_iw[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 472.270 53.400 472.570 54.400 ;
    END
  END um_iw[185]
  PIN um_iw[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 469.510 53.400 469.810 54.400 ;
    END
  END um_iw[186]
  PIN um_iw[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 466.750 53.400 467.050 54.400 ;
    END
  END um_iw[187]
  PIN um_iw[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 463.990 53.400 464.290 54.400 ;
    END
  END um_iw[188]
  PIN um_iw[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 461.230 53.400 461.530 54.400 ;
    END
  END um_iw[189]
  PIN um_iw[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1337.070 0.000 1337.370 1.000 ;
    END
  END um_iw[18]
  PIN um_iw[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 458.470 53.400 458.770 54.400 ;
    END
  END um_iw[190]
  PIN um_iw[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 455.710 53.400 456.010 54.400 ;
    END
  END um_iw[191]
  PIN um_iw[192]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 452.950 53.400 453.250 54.400 ;
    END
  END um_iw[192]
  PIN um_iw[193]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 450.190 53.400 450.490 54.400 ;
    END
  END um_iw[193]
  PIN um_iw[194]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 447.430 53.400 447.730 54.400 ;
    END
  END um_iw[194]
  PIN um_iw[195]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 444.670 53.400 444.970 54.400 ;
    END
  END um_iw[195]
  PIN um_iw[196]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 441.910 53.400 442.210 54.400 ;
    END
  END um_iw[196]
  PIN um_iw[197]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 439.150 53.400 439.450 54.400 ;
    END
  END um_iw[197]
  PIN um_iw[198]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 486.070 0.000 486.370 1.000 ;
    END
  END um_iw[198]
  PIN um_iw[199]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 483.310 0.000 483.610 1.000 ;
    END
  END um_iw[199]
  PIN um_iw[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1334.310 0.000 1334.610 1.000 ;
    END
  END um_iw[19]
  PIN um_iw[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1334.310 53.400 1334.610 54.400 ;
    END
  END um_iw[1]
  PIN um_iw[200]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 480.550 0.000 480.850 1.000 ;
    END
  END um_iw[200]
  PIN um_iw[201]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 477.790 0.000 478.090 1.000 ;
    END
  END um_iw[201]
  PIN um_iw[202]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 475.030 0.000 475.330 1.000 ;
    END
  END um_iw[202]
  PIN um_iw[203]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 472.270 0.000 472.570 1.000 ;
    END
  END um_iw[203]
  PIN um_iw[204]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 469.510 0.000 469.810 1.000 ;
    END
  END um_iw[204]
  PIN um_iw[205]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 466.750 0.000 467.050 1.000 ;
    END
  END um_iw[205]
  PIN um_iw[206]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 463.990 0.000 464.290 1.000 ;
    END
  END um_iw[206]
  PIN um_iw[207]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 461.230 0.000 461.530 1.000 ;
    END
  END um_iw[207]
  PIN um_iw[208]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 458.470 0.000 458.770 1.000 ;
    END
  END um_iw[208]
  PIN um_iw[209]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 455.710 0.000 456.010 1.000 ;
    END
  END um_iw[209]
  PIN um_iw[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1331.550 0.000 1331.850 1.000 ;
    END
  END um_iw[20]
  PIN um_iw[210]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 452.950 0.000 453.250 1.000 ;
    END
  END um_iw[210]
  PIN um_iw[211]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 450.190 0.000 450.490 1.000 ;
    END
  END um_iw[211]
  PIN um_iw[212]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 447.430 0.000 447.730 1.000 ;
    END
  END um_iw[212]
  PIN um_iw[213]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 444.670 0.000 444.970 1.000 ;
    END
  END um_iw[213]
  PIN um_iw[214]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 441.910 0.000 442.210 1.000 ;
    END
  END um_iw[214]
  PIN um_iw[215]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 439.150 0.000 439.450 1.000 ;
    END
  END um_iw[215]
  PIN um_iw[216]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 315.870 53.400 316.170 54.400 ;
    END
  END um_iw[216]
  PIN um_iw[217]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 313.110 53.400 313.410 54.400 ;
    END
  END um_iw[217]
  PIN um_iw[218]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 310.350 53.400 310.650 54.400 ;
    END
  END um_iw[218]
  PIN um_iw[219]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 307.590 53.400 307.890 54.400 ;
    END
  END um_iw[219]
  PIN um_iw[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1328.790 0.000 1329.090 1.000 ;
    END
  END um_iw[21]
  PIN um_iw[220]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 304.830 53.400 305.130 54.400 ;
    END
  END um_iw[220]
  PIN um_iw[221]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 302.070 53.400 302.370 54.400 ;
    END
  END um_iw[221]
  PIN um_iw[222]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 299.310 53.400 299.610 54.400 ;
    END
  END um_iw[222]
  PIN um_iw[223]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 296.550 53.400 296.850 54.400 ;
    END
  END um_iw[223]
  PIN um_iw[224]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 293.790 53.400 294.090 54.400 ;
    END
  END um_iw[224]
  PIN um_iw[225]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 291.030 53.400 291.330 54.400 ;
    END
  END um_iw[225]
  PIN um_iw[226]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 288.270 53.400 288.570 54.400 ;
    END
  END um_iw[226]
  PIN um_iw[227]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 285.510 53.400 285.810 54.400 ;
    END
  END um_iw[227]
  PIN um_iw[228]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 282.750 53.400 283.050 54.400 ;
    END
  END um_iw[228]
  PIN um_iw[229]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 279.990 53.400 280.290 54.400 ;
    END
  END um_iw[229]
  PIN um_iw[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1326.030 0.000 1326.330 1.000 ;
    END
  END um_iw[22]
  PIN um_iw[230]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 277.230 53.400 277.530 54.400 ;
    END
  END um_iw[230]
  PIN um_iw[231]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 274.470 53.400 274.770 54.400 ;
    END
  END um_iw[231]
  PIN um_iw[232]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 271.710 53.400 272.010 54.400 ;
    END
  END um_iw[232]
  PIN um_iw[233]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 268.950 53.400 269.250 54.400 ;
    END
  END um_iw[233]
  PIN um_iw[234]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 315.870 0.000 316.170 1.000 ;
    END
  END um_iw[234]
  PIN um_iw[235]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 313.110 0.000 313.410 1.000 ;
    END
  END um_iw[235]
  PIN um_iw[236]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 310.350 0.000 310.650 1.000 ;
    END
  END um_iw[236]
  PIN um_iw[237]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 307.590 0.000 307.890 1.000 ;
    END
  END um_iw[237]
  PIN um_iw[238]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 304.830 0.000 305.130 1.000 ;
    END
  END um_iw[238]
  PIN um_iw[239]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 302.070 0.000 302.370 1.000 ;
    END
  END um_iw[239]
  PIN um_iw[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1323.270 0.000 1323.570 1.000 ;
    END
  END um_iw[23]
  PIN um_iw[240]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 299.310 0.000 299.610 1.000 ;
    END
  END um_iw[240]
  PIN um_iw[241]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 296.550 0.000 296.850 1.000 ;
    END
  END um_iw[241]
  PIN um_iw[242]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 293.790 0.000 294.090 1.000 ;
    END
  END um_iw[242]
  PIN um_iw[243]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 291.030 0.000 291.330 1.000 ;
    END
  END um_iw[243]
  PIN um_iw[244]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 288.270 0.000 288.570 1.000 ;
    END
  END um_iw[244]
  PIN um_iw[245]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 285.510 0.000 285.810 1.000 ;
    END
  END um_iw[245]
  PIN um_iw[246]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 282.750 0.000 283.050 1.000 ;
    END
  END um_iw[246]
  PIN um_iw[247]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 279.990 0.000 280.290 1.000 ;
    END
  END um_iw[247]
  PIN um_iw[248]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 277.230 0.000 277.530 1.000 ;
    END
  END um_iw[248]
  PIN um_iw[249]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 274.470 0.000 274.770 1.000 ;
    END
  END um_iw[249]
  PIN um_iw[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1320.510 0.000 1320.810 1.000 ;
    END
  END um_iw[24]
  PIN um_iw[250]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 271.710 0.000 272.010 1.000 ;
    END
  END um_iw[250]
  PIN um_iw[251]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 268.950 0.000 269.250 1.000 ;
    END
  END um_iw[251]
  PIN um_iw[252]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 145.670 53.400 145.970 54.400 ;
    END
  END um_iw[252]
  PIN um_iw[253]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 142.910 53.400 143.210 54.400 ;
    END
  END um_iw[253]
  PIN um_iw[254]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 53.400 140.450 54.400 ;
    END
  END um_iw[254]
  PIN um_iw[255]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 137.390 53.400 137.690 54.400 ;
    END
  END um_iw[255]
  PIN um_iw[256]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 134.630 53.400 134.930 54.400 ;
    END
  END um_iw[256]
  PIN um_iw[257]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 131.870 53.400 132.170 54.400 ;
    END
  END um_iw[257]
  PIN um_iw[258]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 53.400 129.410 54.400 ;
    END
  END um_iw[258]
  PIN um_iw[259]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 126.350 53.400 126.650 54.400 ;
    END
  END um_iw[259]
  PIN um_iw[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1317.750 0.000 1318.050 1.000 ;
    END
  END um_iw[25]
  PIN um_iw[260]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 123.590 53.400 123.890 54.400 ;
    END
  END um_iw[260]
  PIN um_iw[261]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 120.830 53.400 121.130 54.400 ;
    END
  END um_iw[261]
  PIN um_iw[262]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 118.070 53.400 118.370 54.400 ;
    END
  END um_iw[262]
  PIN um_iw[263]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 115.310 53.400 115.610 54.400 ;
    END
  END um_iw[263]
  PIN um_iw[264]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 112.550 53.400 112.850 54.400 ;
    END
  END um_iw[264]
  PIN um_iw[265]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 109.790 53.400 110.090 54.400 ;
    END
  END um_iw[265]
  PIN um_iw[266]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 107.030 53.400 107.330 54.400 ;
    END
  END um_iw[266]
  PIN um_iw[267]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 104.270 53.400 104.570 54.400 ;
    END
  END um_iw[267]
  PIN um_iw[268]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 101.510 53.400 101.810 54.400 ;
    END
  END um_iw[268]
  PIN um_iw[269]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 98.750 53.400 99.050 54.400 ;
    END
  END um_iw[269]
  PIN um_iw[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1314.990 0.000 1315.290 1.000 ;
    END
  END um_iw[26]
  PIN um_iw[270]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 145.670 0.000 145.970 1.000 ;
    END
  END um_iw[270]
  PIN um_iw[271]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 142.910 0.000 143.210 1.000 ;
    END
  END um_iw[271]
  PIN um_iw[272]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 0.000 140.450 1.000 ;
    END
  END um_iw[272]
  PIN um_iw[273]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 137.390 0.000 137.690 1.000 ;
    END
  END um_iw[273]
  PIN um_iw[274]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 134.630 0.000 134.930 1.000 ;
    END
  END um_iw[274]
  PIN um_iw[275]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 131.870 0.000 132.170 1.000 ;
    END
  END um_iw[275]
  PIN um_iw[276]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 0.000 129.410 1.000 ;
    END
  END um_iw[276]
  PIN um_iw[277]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 126.350 0.000 126.650 1.000 ;
    END
  END um_iw[277]
  PIN um_iw[278]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 123.590 0.000 123.890 1.000 ;
    END
  END um_iw[278]
  PIN um_iw[279]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 120.830 0.000 121.130 1.000 ;
    END
  END um_iw[279]
  PIN um_iw[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1312.230 0.000 1312.530 1.000 ;
    END
  END um_iw[27]
  PIN um_iw[280]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 118.070 0.000 118.370 1.000 ;
    END
  END um_iw[280]
  PIN um_iw[281]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 115.310 0.000 115.610 1.000 ;
    END
  END um_iw[281]
  PIN um_iw[282]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 112.550 0.000 112.850 1.000 ;
    END
  END um_iw[282]
  PIN um_iw[283]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 109.790 0.000 110.090 1.000 ;
    END
  END um_iw[283]
  PIN um_iw[284]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 107.030 0.000 107.330 1.000 ;
    END
  END um_iw[284]
  PIN um_iw[285]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 104.270 0.000 104.570 1.000 ;
    END
  END um_iw[285]
  PIN um_iw[286]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 101.510 0.000 101.810 1.000 ;
    END
  END um_iw[286]
  PIN um_iw[287]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 98.750 0.000 99.050 1.000 ;
    END
  END um_iw[287]
  PIN um_iw[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1309.470 0.000 1309.770 1.000 ;
    END
  END um_iw[28]
  PIN um_iw[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1306.710 0.000 1307.010 1.000 ;
    END
  END um_iw[29]
  PIN um_iw[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1331.550 53.400 1331.850 54.400 ;
    END
  END um_iw[2]
  PIN um_iw[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1303.950 0.000 1304.250 1.000 ;
    END
  END um_iw[30]
  PIN um_iw[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1301.190 0.000 1301.490 1.000 ;
    END
  END um_iw[31]
  PIN um_iw[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1298.430 0.000 1298.730 1.000 ;
    END
  END um_iw[32]
  PIN um_iw[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1295.670 0.000 1295.970 1.000 ;
    END
  END um_iw[33]
  PIN um_iw[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1292.910 0.000 1293.210 1.000 ;
    END
  END um_iw[34]
  PIN um_iw[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1290.150 0.000 1290.450 1.000 ;
    END
  END um_iw[35]
  PIN um_iw[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1166.870 53.400 1167.170 54.400 ;
    END
  END um_iw[36]
  PIN um_iw[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1164.110 53.400 1164.410 54.400 ;
    END
  END um_iw[37]
  PIN um_iw[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1161.350 53.400 1161.650 54.400 ;
    END
  END um_iw[38]
  PIN um_iw[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1158.590 53.400 1158.890 54.400 ;
    END
  END um_iw[39]
  PIN um_iw[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1328.790 53.400 1329.090 54.400 ;
    END
  END um_iw[3]
  PIN um_iw[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1155.830 53.400 1156.130 54.400 ;
    END
  END um_iw[40]
  PIN um_iw[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1153.070 53.400 1153.370 54.400 ;
    END
  END um_iw[41]
  PIN um_iw[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1150.310 53.400 1150.610 54.400 ;
    END
  END um_iw[42]
  PIN um_iw[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1147.550 53.400 1147.850 54.400 ;
    END
  END um_iw[43]
  PIN um_iw[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1144.790 53.400 1145.090 54.400 ;
    END
  END um_iw[44]
  PIN um_iw[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1142.030 53.400 1142.330 54.400 ;
    END
  END um_iw[45]
  PIN um_iw[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1139.270 53.400 1139.570 54.400 ;
    END
  END um_iw[46]
  PIN um_iw[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1136.510 53.400 1136.810 54.400 ;
    END
  END um_iw[47]
  PIN um_iw[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1133.750 53.400 1134.050 54.400 ;
    END
  END um_iw[48]
  PIN um_iw[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1130.990 53.400 1131.290 54.400 ;
    END
  END um_iw[49]
  PIN um_iw[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1326.030 53.400 1326.330 54.400 ;
    END
  END um_iw[4]
  PIN um_iw[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1128.230 53.400 1128.530 54.400 ;
    END
  END um_iw[50]
  PIN um_iw[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1125.470 53.400 1125.770 54.400 ;
    END
  END um_iw[51]
  PIN um_iw[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1122.710 53.400 1123.010 54.400 ;
    END
  END um_iw[52]
  PIN um_iw[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1119.950 53.400 1120.250 54.400 ;
    END
  END um_iw[53]
  PIN um_iw[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1166.870 0.000 1167.170 1.000 ;
    END
  END um_iw[54]
  PIN um_iw[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1164.110 0.000 1164.410 1.000 ;
    END
  END um_iw[55]
  PIN um_iw[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1161.350 0.000 1161.650 1.000 ;
    END
  END um_iw[56]
  PIN um_iw[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1158.590 0.000 1158.890 1.000 ;
    END
  END um_iw[57]
  PIN um_iw[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1155.830 0.000 1156.130 1.000 ;
    END
  END um_iw[58]
  PIN um_iw[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1153.070 0.000 1153.370 1.000 ;
    END
  END um_iw[59]
  PIN um_iw[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1323.270 53.400 1323.570 54.400 ;
    END
  END um_iw[5]
  PIN um_iw[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1150.310 0.000 1150.610 1.000 ;
    END
  END um_iw[60]
  PIN um_iw[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1147.550 0.000 1147.850 1.000 ;
    END
  END um_iw[61]
  PIN um_iw[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1144.790 0.000 1145.090 1.000 ;
    END
  END um_iw[62]
  PIN um_iw[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1142.030 0.000 1142.330 1.000 ;
    END
  END um_iw[63]
  PIN um_iw[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1139.270 0.000 1139.570 1.000 ;
    END
  END um_iw[64]
  PIN um_iw[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1136.510 0.000 1136.810 1.000 ;
    END
  END um_iw[65]
  PIN um_iw[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1133.750 0.000 1134.050 1.000 ;
    END
  END um_iw[66]
  PIN um_iw[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1130.990 0.000 1131.290 1.000 ;
    END
  END um_iw[67]
  PIN um_iw[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1128.230 0.000 1128.530 1.000 ;
    END
  END um_iw[68]
  PIN um_iw[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1125.470 0.000 1125.770 1.000 ;
    END
  END um_iw[69]
  PIN um_iw[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1320.510 53.400 1320.810 54.400 ;
    END
  END um_iw[6]
  PIN um_iw[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1122.710 0.000 1123.010 1.000 ;
    END
  END um_iw[70]
  PIN um_iw[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1119.950 0.000 1120.250 1.000 ;
    END
  END um_iw[71]
  PIN um_iw[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 996.670 53.400 996.970 54.400 ;
    END
  END um_iw[72]
  PIN um_iw[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 993.910 53.400 994.210 54.400 ;
    END
  END um_iw[73]
  PIN um_iw[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 991.150 53.400 991.450 54.400 ;
    END
  END um_iw[74]
  PIN um_iw[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 988.390 53.400 988.690 54.400 ;
    END
  END um_iw[75]
  PIN um_iw[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 985.630 53.400 985.930 54.400 ;
    END
  END um_iw[76]
  PIN um_iw[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 982.870 53.400 983.170 54.400 ;
    END
  END um_iw[77]
  PIN um_iw[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 980.110 53.400 980.410 54.400 ;
    END
  END um_iw[78]
  PIN um_iw[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 977.350 53.400 977.650 54.400 ;
    END
  END um_iw[79]
  PIN um_iw[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1317.750 53.400 1318.050 54.400 ;
    END
  END um_iw[7]
  PIN um_iw[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 974.590 53.400 974.890 54.400 ;
    END
  END um_iw[80]
  PIN um_iw[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 971.830 53.400 972.130 54.400 ;
    END
  END um_iw[81]
  PIN um_iw[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 969.070 53.400 969.370 54.400 ;
    END
  END um_iw[82]
  PIN um_iw[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 966.310 53.400 966.610 54.400 ;
    END
  END um_iw[83]
  PIN um_iw[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 963.550 53.400 963.850 54.400 ;
    END
  END um_iw[84]
  PIN um_iw[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 960.790 53.400 961.090 54.400 ;
    END
  END um_iw[85]
  PIN um_iw[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 958.030 53.400 958.330 54.400 ;
    END
  END um_iw[86]
  PIN um_iw[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 955.270 53.400 955.570 54.400 ;
    END
  END um_iw[87]
  PIN um_iw[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 952.510 53.400 952.810 54.400 ;
    END
  END um_iw[88]
  PIN um_iw[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 949.750 53.400 950.050 54.400 ;
    END
  END um_iw[89]
  PIN um_iw[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1314.990 53.400 1315.290 54.400 ;
    END
  END um_iw[8]
  PIN um_iw[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 996.670 0.000 996.970 1.000 ;
    END
  END um_iw[90]
  PIN um_iw[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 993.910 0.000 994.210 1.000 ;
    END
  END um_iw[91]
  PIN um_iw[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 991.150 0.000 991.450 1.000 ;
    END
  END um_iw[92]
  PIN um_iw[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 988.390 0.000 988.690 1.000 ;
    END
  END um_iw[93]
  PIN um_iw[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 985.630 0.000 985.930 1.000 ;
    END
  END um_iw[94]
  PIN um_iw[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 982.870 0.000 983.170 1.000 ;
    END
  END um_iw[95]
  PIN um_iw[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 980.110 0.000 980.410 1.000 ;
    END
  END um_iw[96]
  PIN um_iw[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 977.350 0.000 977.650 1.000 ;
    END
  END um_iw[97]
  PIN um_iw[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 974.590 0.000 974.890 1.000 ;
    END
  END um_iw[98]
  PIN um_iw[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 971.830 0.000 972.130 1.000 ;
    END
  END um_iw[99]
  PIN um_iw[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER met4 ;
        RECT 1312.230 53.400 1312.530 54.400 ;
    END
  END um_iw[9]
  PIN um_k_zero[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1221.150 53.400 1221.450 54.400 ;
    END
  END um_k_zero[0]
  PIN um_k_zero[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 370.150 53.400 370.450 54.400 ;
    END
  END um_k_zero[10]
  PIN um_k_zero[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 370.150 0.000 370.450 1.000 ;
    END
  END um_k_zero[11]
  PIN um_k_zero[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 199.950 53.400 200.250 54.400 ;
    END
  END um_k_zero[12]
  PIN um_k_zero[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 199.950 0.000 200.250 1.000 ;
    END
  END um_k_zero[13]
  PIN um_k_zero[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 53.400 30.050 54.400 ;
    END
  END um_k_zero[14]
  PIN um_k_zero[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 0.000 30.050 1.000 ;
    END
  END um_k_zero[15]
  PIN um_k_zero[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1221.150 0.000 1221.450 1.000 ;
    END
  END um_k_zero[1]
  PIN um_k_zero[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1050.950 53.400 1051.250 54.400 ;
    END
  END um_k_zero[2]
  PIN um_k_zero[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1050.950 0.000 1051.250 1.000 ;
    END
  END um_k_zero[3]
  PIN um_k_zero[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 880.750 53.400 881.050 54.400 ;
    END
  END um_k_zero[4]
  PIN um_k_zero[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 880.750 0.000 881.050 1.000 ;
    END
  END um_k_zero[5]
  PIN um_k_zero[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 710.550 53.400 710.850 54.400 ;
    END
  END um_k_zero[6]
  PIN um_k_zero[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 710.550 0.000 710.850 1.000 ;
    END
  END um_k_zero[7]
  PIN um_k_zero[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 540.350 53.400 540.650 54.400 ;
    END
  END um_k_zero[8]
  PIN um_k_zero[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 540.350 0.000 540.650 1.000 ;
    END
  END um_k_zero[9]
  PIN um_ow[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1287.390 53.400 1287.690 54.400 ;
    END
  END um_ow[0]
  PIN um_ow[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 935.950 53.400 936.250 54.400 ;
    END
  END um_ow[100]
  PIN um_ow[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 933.190 53.400 933.490 54.400 ;
    END
  END um_ow[101]
  PIN um_ow[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 930.430 53.400 930.730 54.400 ;
    END
  END um_ow[102]
  PIN um_ow[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 927.670 53.400 927.970 54.400 ;
    END
  END um_ow[103]
  PIN um_ow[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 924.910 53.400 925.210 54.400 ;
    END
  END um_ow[104]
  PIN um_ow[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 922.150 53.400 922.450 54.400 ;
    END
  END um_ow[105]
  PIN um_ow[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 919.390 53.400 919.690 54.400 ;
    END
  END um_ow[106]
  PIN um_ow[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 916.630 53.400 916.930 54.400 ;
    END
  END um_ow[107]
  PIN um_ow[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 913.870 53.400 914.170 54.400 ;
    END
  END um_ow[108]
  PIN um_ow[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 911.110 53.400 911.410 54.400 ;
    END
  END um_ow[109]
  PIN um_ow[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1259.790 53.400 1260.090 54.400 ;
    END
  END um_ow[10]
  PIN um_ow[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 908.350 53.400 908.650 54.400 ;
    END
  END um_ow[110]
  PIN um_ow[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 905.590 53.400 905.890 54.400 ;
    END
  END um_ow[111]
  PIN um_ow[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 902.830 53.400 903.130 54.400 ;
    END
  END um_ow[112]
  PIN um_ow[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 900.070 53.400 900.370 54.400 ;
    END
  END um_ow[113]
  PIN um_ow[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met4 ;
        RECT 897.310 53.400 897.610 54.400 ;
    END
  END um_ow[114]
  PIN um_ow[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 894.550 53.400 894.850 54.400 ;
    END
  END um_ow[115]
  PIN um_ow[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 891.790 53.400 892.090 54.400 ;
    END
  END um_ow[116]
  PIN um_ow[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 889.030 53.400 889.330 54.400 ;
    END
  END um_ow[117]
  PIN um_ow[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met4 ;
        RECT 886.270 53.400 886.570 54.400 ;
    END
  END um_ow[118]
  PIN um_ow[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met4 ;
        RECT 883.510 53.400 883.810 54.400 ;
    END
  END um_ow[119]
  PIN um_ow[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1257.030 53.400 1257.330 54.400 ;
    END
  END um_ow[11]
  PIN um_ow[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 946.990 0.000 947.290 1.000 ;
    END
  END um_ow[120]
  PIN um_ow[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 944.230 0.000 944.530 1.000 ;
    END
  END um_ow[121]
  PIN um_ow[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 941.470 0.000 941.770 1.000 ;
    END
  END um_ow[122]
  PIN um_ow[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 938.710 0.000 939.010 1.000 ;
    END
  END um_ow[123]
  PIN um_ow[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 935.950 0.000 936.250 1.000 ;
    END
  END um_ow[124]
  PIN um_ow[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 933.190 0.000 933.490 1.000 ;
    END
  END um_ow[125]
  PIN um_ow[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 930.430 0.000 930.730 1.000 ;
    END
  END um_ow[126]
  PIN um_ow[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 927.670 0.000 927.970 1.000 ;
    END
  END um_ow[127]
  PIN um_ow[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 924.910 0.000 925.210 1.000 ;
    END
  END um_ow[128]
  PIN um_ow[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 922.150 0.000 922.450 1.000 ;
    END
  END um_ow[129]
  PIN um_ow[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1254.270 53.400 1254.570 54.400 ;
    END
  END um_ow[12]
  PIN um_ow[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 919.390 0.000 919.690 1.000 ;
    END
  END um_ow[130]
  PIN um_ow[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 916.630 0.000 916.930 1.000 ;
    END
  END um_ow[131]
  PIN um_ow[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 913.870 0.000 914.170 1.000 ;
    END
  END um_ow[132]
  PIN um_ow[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 911.110 0.000 911.410 1.000 ;
    END
  END um_ow[133]
  PIN um_ow[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 908.350 0.000 908.650 1.000 ;
    END
  END um_ow[134]
  PIN um_ow[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 905.590 0.000 905.890 1.000 ;
    END
  END um_ow[135]
  PIN um_ow[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 902.830 0.000 903.130 1.000 ;
    END
  END um_ow[136]
  PIN um_ow[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 900.070 0.000 900.370 1.000 ;
    END
  END um_ow[137]
  PIN um_ow[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 897.310 0.000 897.610 1.000 ;
    END
  END um_ow[138]
  PIN um_ow[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met4 ;
        RECT 894.550 0.000 894.850 1.000 ;
    END
  END um_ow[139]
  PIN um_ow[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1251.510 53.400 1251.810 54.400 ;
    END
  END um_ow[13]
  PIN um_ow[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met4 ;
        RECT 891.790 0.000 892.090 1.000 ;
    END
  END um_ow[140]
  PIN um_ow[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 889.030 0.000 889.330 1.000 ;
    END
  END um_ow[141]
  PIN um_ow[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 886.270 0.000 886.570 1.000 ;
    END
  END um_ow[142]
  PIN um_ow[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 883.510 0.000 883.810 1.000 ;
    END
  END um_ow[143]
  PIN um_ow[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 776.790 53.400 777.090 54.400 ;
    END
  END um_ow[144]
  PIN um_ow[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 774.030 53.400 774.330 54.400 ;
    END
  END um_ow[145]
  PIN um_ow[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 771.270 53.400 771.570 54.400 ;
    END
  END um_ow[146]
  PIN um_ow[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 768.510 53.400 768.810 54.400 ;
    END
  END um_ow[147]
  PIN um_ow[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 765.750 53.400 766.050 54.400 ;
    END
  END um_ow[148]
  PIN um_ow[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 762.990 53.400 763.290 54.400 ;
    END
  END um_ow[149]
  PIN um_ow[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1248.750 53.400 1249.050 54.400 ;
    END
  END um_ow[14]
  PIN um_ow[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 760.230 53.400 760.530 54.400 ;
    END
  END um_ow[150]
  PIN um_ow[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 757.470 53.400 757.770 54.400 ;
    END
  END um_ow[151]
  PIN um_ow[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 754.710 53.400 755.010 54.400 ;
    END
  END um_ow[152]
  PIN um_ow[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 751.950 53.400 752.250 54.400 ;
    END
  END um_ow[153]
  PIN um_ow[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 749.190 53.400 749.490 54.400 ;
    END
  END um_ow[154]
  PIN um_ow[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 746.430 53.400 746.730 54.400 ;
    END
  END um_ow[155]
  PIN um_ow[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 743.670 53.400 743.970 54.400 ;
    END
  END um_ow[156]
  PIN um_ow[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 740.910 53.400 741.210 54.400 ;
    END
  END um_ow[157]
  PIN um_ow[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 738.150 53.400 738.450 54.400 ;
    END
  END um_ow[158]
  PIN um_ow[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 735.390 53.400 735.690 54.400 ;
    END
  END um_ow[159]
  PIN um_ow[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1245.990 53.400 1246.290 54.400 ;
    END
  END um_ow[15]
  PIN um_ow[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 732.630 53.400 732.930 54.400 ;
    END
  END um_ow[160]
  PIN um_ow[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 729.870 53.400 730.170 54.400 ;
    END
  END um_ow[161]
  PIN um_ow[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 727.110 53.400 727.410 54.400 ;
    END
  END um_ow[162]
  PIN um_ow[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 724.350 53.400 724.650 54.400 ;
    END
  END um_ow[163]
  PIN um_ow[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 721.590 53.400 721.890 54.400 ;
    END
  END um_ow[164]
  PIN um_ow[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 718.830 53.400 719.130 54.400 ;
    END
  END um_ow[165]
  PIN um_ow[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 716.070 53.400 716.370 54.400 ;
    END
  END um_ow[166]
  PIN um_ow[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 713.310 53.400 713.610 54.400 ;
    END
  END um_ow[167]
  PIN um_ow[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 776.790 0.000 777.090 1.000 ;
    END
  END um_ow[168]
  PIN um_ow[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 774.030 0.000 774.330 1.000 ;
    END
  END um_ow[169]
  PIN um_ow[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1243.230 53.400 1243.530 54.400 ;
    END
  END um_ow[16]
  PIN um_ow[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 771.270 0.000 771.570 1.000 ;
    END
  END um_ow[170]
  PIN um_ow[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 768.510 0.000 768.810 1.000 ;
    END
  END um_ow[171]
  PIN um_ow[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 765.750 0.000 766.050 1.000 ;
    END
  END um_ow[172]
  PIN um_ow[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 762.990 0.000 763.290 1.000 ;
    END
  END um_ow[173]
  PIN um_ow[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 760.230 0.000 760.530 1.000 ;
    END
  END um_ow[174]
  PIN um_ow[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 757.470 0.000 757.770 1.000 ;
    END
  END um_ow[175]
  PIN um_ow[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 754.710 0.000 755.010 1.000 ;
    END
  END um_ow[176]
  PIN um_ow[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 751.950 0.000 752.250 1.000 ;
    END
  END um_ow[177]
  PIN um_ow[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 749.190 0.000 749.490 1.000 ;
    END
  END um_ow[178]
  PIN um_ow[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 746.430 0.000 746.730 1.000 ;
    END
  END um_ow[179]
  PIN um_ow[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1240.470 53.400 1240.770 54.400 ;
    END
  END um_ow[17]
  PIN um_ow[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 743.670 0.000 743.970 1.000 ;
    END
  END um_ow[180]
  PIN um_ow[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 740.910 0.000 741.210 1.000 ;
    END
  END um_ow[181]
  PIN um_ow[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 738.150 0.000 738.450 1.000 ;
    END
  END um_ow[182]
  PIN um_ow[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 735.390 0.000 735.690 1.000 ;
    END
  END um_ow[183]
  PIN um_ow[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 732.630 0.000 732.930 1.000 ;
    END
  END um_ow[184]
  PIN um_ow[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 729.870 0.000 730.170 1.000 ;
    END
  END um_ow[185]
  PIN um_ow[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 727.110 0.000 727.410 1.000 ;
    END
  END um_ow[186]
  PIN um_ow[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 724.350 0.000 724.650 1.000 ;
    END
  END um_ow[187]
  PIN um_ow[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 721.590 0.000 721.890 1.000 ;
    END
  END um_ow[188]
  PIN um_ow[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 718.830 0.000 719.130 1.000 ;
    END
  END um_ow[189]
  PIN um_ow[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1237.710 53.400 1238.010 54.400 ;
    END
  END um_ow[18]
  PIN um_ow[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 716.070 0.000 716.370 1.000 ;
    END
  END um_ow[190]
  PIN um_ow[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 713.310 0.000 713.610 1.000 ;
    END
  END um_ow[191]
  PIN um_ow[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 606.590 53.400 606.890 54.400 ;
    END
  END um_ow[192]
  PIN um_ow[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 603.830 53.400 604.130 54.400 ;
    END
  END um_ow[193]
  PIN um_ow[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 601.070 53.400 601.370 54.400 ;
    END
  END um_ow[194]
  PIN um_ow[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 598.310 53.400 598.610 54.400 ;
    END
  END um_ow[195]
  PIN um_ow[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 595.550 53.400 595.850 54.400 ;
    END
  END um_ow[196]
  PIN um_ow[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 592.790 53.400 593.090 54.400 ;
    END
  END um_ow[197]
  PIN um_ow[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 590.030 53.400 590.330 54.400 ;
    END
  END um_ow[198]
  PIN um_ow[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 587.270 53.400 587.570 54.400 ;
    END
  END um_ow[199]
  PIN um_ow[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1234.950 53.400 1235.250 54.400 ;
    END
  END um_ow[19]
  PIN um_ow[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met4 ;
        RECT 1284.630 53.400 1284.930 54.400 ;
    END
  END um_ow[1]
  PIN um_ow[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 584.510 53.400 584.810 54.400 ;
    END
  END um_ow[200]
  PIN um_ow[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 581.750 53.400 582.050 54.400 ;
    END
  END um_ow[201]
  PIN um_ow[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 578.990 53.400 579.290 54.400 ;
    END
  END um_ow[202]
  PIN um_ow[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 576.230 53.400 576.530 54.400 ;
    END
  END um_ow[203]
  PIN um_ow[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 573.470 53.400 573.770 54.400 ;
    END
  END um_ow[204]
  PIN um_ow[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 570.710 53.400 571.010 54.400 ;
    END
  END um_ow[205]
  PIN um_ow[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 567.950 53.400 568.250 54.400 ;
    END
  END um_ow[206]
  PIN um_ow[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 565.190 53.400 565.490 54.400 ;
    END
  END um_ow[207]
  PIN um_ow[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 562.430 53.400 562.730 54.400 ;
    END
  END um_ow[208]
  PIN um_ow[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 559.670 53.400 559.970 54.400 ;
    END
  END um_ow[209]
  PIN um_ow[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1232.190 53.400 1232.490 54.400 ;
    END
  END um_ow[20]
  PIN um_ow[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 556.910 53.400 557.210 54.400 ;
    END
  END um_ow[210]
  PIN um_ow[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 554.150 53.400 554.450 54.400 ;
    END
  END um_ow[211]
  PIN um_ow[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 551.390 53.400 551.690 54.400 ;
    END
  END um_ow[212]
  PIN um_ow[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 548.630 53.400 548.930 54.400 ;
    END
  END um_ow[213]
  PIN um_ow[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 545.870 53.400 546.170 54.400 ;
    END
  END um_ow[214]
  PIN um_ow[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 543.110 53.400 543.410 54.400 ;
    END
  END um_ow[215]
  PIN um_ow[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 606.590 0.000 606.890 1.000 ;
    END
  END um_ow[216]
  PIN um_ow[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 603.830 0.000 604.130 1.000 ;
    END
  END um_ow[217]
  PIN um_ow[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 601.070 0.000 601.370 1.000 ;
    END
  END um_ow[218]
  PIN um_ow[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 598.310 0.000 598.610 1.000 ;
    END
  END um_ow[219]
  PIN um_ow[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met4 ;
        RECT 1229.430 53.400 1229.730 54.400 ;
    END
  END um_ow[21]
  PIN um_ow[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 595.550 0.000 595.850 1.000 ;
    END
  END um_ow[220]
  PIN um_ow[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 592.790 0.000 593.090 1.000 ;
    END
  END um_ow[221]
  PIN um_ow[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 590.030 0.000 590.330 1.000 ;
    END
  END um_ow[222]
  PIN um_ow[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 587.270 0.000 587.570 1.000 ;
    END
  END um_ow[223]
  PIN um_ow[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 584.510 0.000 584.810 1.000 ;
    END
  END um_ow[224]
  PIN um_ow[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 581.750 0.000 582.050 1.000 ;
    END
  END um_ow[225]
  PIN um_ow[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 578.990 0.000 579.290 1.000 ;
    END
  END um_ow[226]
  PIN um_ow[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 576.230 0.000 576.530 1.000 ;
    END
  END um_ow[227]
  PIN um_ow[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 573.470 0.000 573.770 1.000 ;
    END
  END um_ow[228]
  PIN um_ow[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 570.710 0.000 571.010 1.000 ;
    END
  END um_ow[229]
  PIN um_ow[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1226.670 53.400 1226.970 54.400 ;
    END
  END um_ow[22]
  PIN um_ow[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 567.950 0.000 568.250 1.000 ;
    END
  END um_ow[230]
  PIN um_ow[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 565.190 0.000 565.490 1.000 ;
    END
  END um_ow[231]
  PIN um_ow[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 562.430 0.000 562.730 1.000 ;
    END
  END um_ow[232]
  PIN um_ow[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 559.670 0.000 559.970 1.000 ;
    END
  END um_ow[233]
  PIN um_ow[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 556.910 0.000 557.210 1.000 ;
    END
  END um_ow[234]
  PIN um_ow[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 554.150 0.000 554.450 1.000 ;
    END
  END um_ow[235]
  PIN um_ow[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 551.390 0.000 551.690 1.000 ;
    END
  END um_ow[236]
  PIN um_ow[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 548.630 0.000 548.930 1.000 ;
    END
  END um_ow[237]
  PIN um_ow[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 545.870 0.000 546.170 1.000 ;
    END
  END um_ow[238]
  PIN um_ow[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 543.110 0.000 543.410 1.000 ;
    END
  END um_ow[239]
  PIN um_ow[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met4 ;
        RECT 1223.910 53.400 1224.210 54.400 ;
    END
  END um_ow[23]
  PIN um_ow[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 436.390 53.400 436.690 54.400 ;
    END
  END um_ow[240]
  PIN um_ow[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 433.630 53.400 433.930 54.400 ;
    END
  END um_ow[241]
  PIN um_ow[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 430.870 53.400 431.170 54.400 ;
    END
  END um_ow[242]
  PIN um_ow[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 428.110 53.400 428.410 54.400 ;
    END
  END um_ow[243]
  PIN um_ow[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 425.350 53.400 425.650 54.400 ;
    END
  END um_ow[244]
  PIN um_ow[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 422.590 53.400 422.890 54.400 ;
    END
  END um_ow[245]
  PIN um_ow[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 419.830 53.400 420.130 54.400 ;
    END
  END um_ow[246]
  PIN um_ow[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 417.070 53.400 417.370 54.400 ;
    END
  END um_ow[247]
  PIN um_ow[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 414.310 53.400 414.610 54.400 ;
    END
  END um_ow[248]
  PIN um_ow[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 411.550 53.400 411.850 54.400 ;
    END
  END um_ow[249]
  PIN um_ow[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1287.390 0.000 1287.690 1.000 ;
    END
  END um_ow[24]
  PIN um_ow[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 408.790 53.400 409.090 54.400 ;
    END
  END um_ow[250]
  PIN um_ow[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 406.030 53.400 406.330 54.400 ;
    END
  END um_ow[251]
  PIN um_ow[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 403.270 53.400 403.570 54.400 ;
    END
  END um_ow[252]
  PIN um_ow[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 400.510 53.400 400.810 54.400 ;
    END
  END um_ow[253]
  PIN um_ow[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 397.750 53.400 398.050 54.400 ;
    END
  END um_ow[254]
  PIN um_ow[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 394.990 53.400 395.290 54.400 ;
    END
  END um_ow[255]
  PIN um_ow[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 392.230 53.400 392.530 54.400 ;
    END
  END um_ow[256]
  PIN um_ow[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 389.470 53.400 389.770 54.400 ;
    END
  END um_ow[257]
  PIN um_ow[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 386.710 53.400 387.010 54.400 ;
    END
  END um_ow[258]
  PIN um_ow[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 383.950 53.400 384.250 54.400 ;
    END
  END um_ow[259]
  PIN um_ow[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1284.630 0.000 1284.930 1.000 ;
    END
  END um_ow[25]
  PIN um_ow[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 381.190 53.400 381.490 54.400 ;
    END
  END um_ow[260]
  PIN um_ow[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 378.430 53.400 378.730 54.400 ;
    END
  END um_ow[261]
  PIN um_ow[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 375.670 53.400 375.970 54.400 ;
    END
  END um_ow[262]
  PIN um_ow[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 372.910 53.400 373.210 54.400 ;
    END
  END um_ow[263]
  PIN um_ow[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 436.390 0.000 436.690 1.000 ;
    END
  END um_ow[264]
  PIN um_ow[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 433.630 0.000 433.930 1.000 ;
    END
  END um_ow[265]
  PIN um_ow[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 430.870 0.000 431.170 1.000 ;
    END
  END um_ow[266]
  PIN um_ow[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 428.110 0.000 428.410 1.000 ;
    END
  END um_ow[267]
  PIN um_ow[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 425.350 0.000 425.650 1.000 ;
    END
  END um_ow[268]
  PIN um_ow[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 422.590 0.000 422.890 1.000 ;
    END
  END um_ow[269]
  PIN um_ow[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1281.870 0.000 1282.170 1.000 ;
    END
  END um_ow[26]
  PIN um_ow[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 419.830 0.000 420.130 1.000 ;
    END
  END um_ow[270]
  PIN um_ow[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 417.070 0.000 417.370 1.000 ;
    END
  END um_ow[271]
  PIN um_ow[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 414.310 0.000 414.610 1.000 ;
    END
  END um_ow[272]
  PIN um_ow[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 411.550 0.000 411.850 1.000 ;
    END
  END um_ow[273]
  PIN um_ow[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 408.790 0.000 409.090 1.000 ;
    END
  END um_ow[274]
  PIN um_ow[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 406.030 0.000 406.330 1.000 ;
    END
  END um_ow[275]
  PIN um_ow[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 403.270 0.000 403.570 1.000 ;
    END
  END um_ow[276]
  PIN um_ow[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 400.510 0.000 400.810 1.000 ;
    END
  END um_ow[277]
  PIN um_ow[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 397.750 0.000 398.050 1.000 ;
    END
  END um_ow[278]
  PIN um_ow[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 394.990 0.000 395.290 1.000 ;
    END
  END um_ow[279]
  PIN um_ow[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1279.110 0.000 1279.410 1.000 ;
    END
  END um_ow[27]
  PIN um_ow[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 392.230 0.000 392.530 1.000 ;
    END
  END um_ow[280]
  PIN um_ow[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 389.470 0.000 389.770 1.000 ;
    END
  END um_ow[281]
  PIN um_ow[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 386.710 0.000 387.010 1.000 ;
    END
  END um_ow[282]
  PIN um_ow[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 383.950 0.000 384.250 1.000 ;
    END
  END um_ow[283]
  PIN um_ow[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 381.190 0.000 381.490 1.000 ;
    END
  END um_ow[284]
  PIN um_ow[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 378.430 0.000 378.730 1.000 ;
    END
  END um_ow[285]
  PIN um_ow[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 375.670 0.000 375.970 1.000 ;
    END
  END um_ow[286]
  PIN um_ow[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 372.910 0.000 373.210 1.000 ;
    END
  END um_ow[287]
  PIN um_ow[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 266.190 53.400 266.490 54.400 ;
    END
  END um_ow[288]
  PIN um_ow[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 263.430 53.400 263.730 54.400 ;
    END
  END um_ow[289]
  PIN um_ow[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1276.350 0.000 1276.650 1.000 ;
    END
  END um_ow[28]
  PIN um_ow[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 260.670 53.400 260.970 54.400 ;
    END
  END um_ow[290]
  PIN um_ow[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 257.910 53.400 258.210 54.400 ;
    END
  END um_ow[291]
  PIN um_ow[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 255.150 53.400 255.450 54.400 ;
    END
  END um_ow[292]
  PIN um_ow[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 252.390 53.400 252.690 54.400 ;
    END
  END um_ow[293]
  PIN um_ow[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 249.630 53.400 249.930 54.400 ;
    END
  END um_ow[294]
  PIN um_ow[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 246.870 53.400 247.170 54.400 ;
    END
  END um_ow[295]
  PIN um_ow[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 244.110 53.400 244.410 54.400 ;
    END
  END um_ow[296]
  PIN um_ow[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 241.350 53.400 241.650 54.400 ;
    END
  END um_ow[297]
  PIN um_ow[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 238.590 53.400 238.890 54.400 ;
    END
  END um_ow[298]
  PIN um_ow[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 235.830 53.400 236.130 54.400 ;
    END
  END um_ow[299]
  PIN um_ow[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1273.590 0.000 1273.890 1.000 ;
    END
  END um_ow[29]
  PIN um_ow[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1281.870 53.400 1282.170 54.400 ;
    END
  END um_ow[2]
  PIN um_ow[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 233.070 53.400 233.370 54.400 ;
    END
  END um_ow[300]
  PIN um_ow[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 230.310 53.400 230.610 54.400 ;
    END
  END um_ow[301]
  PIN um_ow[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 227.550 53.400 227.850 54.400 ;
    END
  END um_ow[302]
  PIN um_ow[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 224.790 53.400 225.090 54.400 ;
    END
  END um_ow[303]
  PIN um_ow[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 222.030 53.400 222.330 54.400 ;
    END
  END um_ow[304]
  PIN um_ow[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 219.270 53.400 219.570 54.400 ;
    END
  END um_ow[305]
  PIN um_ow[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 216.510 53.400 216.810 54.400 ;
    END
  END um_ow[306]
  PIN um_ow[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 213.750 53.400 214.050 54.400 ;
    END
  END um_ow[307]
  PIN um_ow[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 210.990 53.400 211.290 54.400 ;
    END
  END um_ow[308]
  PIN um_ow[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 208.230 53.400 208.530 54.400 ;
    END
  END um_ow[309]
  PIN um_ow[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1270.830 0.000 1271.130 1.000 ;
    END
  END um_ow[30]
  PIN um_ow[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 205.470 53.400 205.770 54.400 ;
    END
  END um_ow[310]
  PIN um_ow[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 202.710 53.400 203.010 54.400 ;
    END
  END um_ow[311]
  PIN um_ow[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 266.190 0.000 266.490 1.000 ;
    END
  END um_ow[312]
  PIN um_ow[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 263.430 0.000 263.730 1.000 ;
    END
  END um_ow[313]
  PIN um_ow[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 260.670 0.000 260.970 1.000 ;
    END
  END um_ow[314]
  PIN um_ow[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 257.910 0.000 258.210 1.000 ;
    END
  END um_ow[315]
  PIN um_ow[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 255.150 0.000 255.450 1.000 ;
    END
  END um_ow[316]
  PIN um_ow[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 252.390 0.000 252.690 1.000 ;
    END
  END um_ow[317]
  PIN um_ow[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 249.630 0.000 249.930 1.000 ;
    END
  END um_ow[318]
  PIN um_ow[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 246.870 0.000 247.170 1.000 ;
    END
  END um_ow[319]
  PIN um_ow[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1268.070 0.000 1268.370 1.000 ;
    END
  END um_ow[31]
  PIN um_ow[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 244.110 0.000 244.410 1.000 ;
    END
  END um_ow[320]
  PIN um_ow[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 241.350 0.000 241.650 1.000 ;
    END
  END um_ow[321]
  PIN um_ow[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 238.590 0.000 238.890 1.000 ;
    END
  END um_ow[322]
  PIN um_ow[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 235.830 0.000 236.130 1.000 ;
    END
  END um_ow[323]
  PIN um_ow[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 233.070 0.000 233.370 1.000 ;
    END
  END um_ow[324]
  PIN um_ow[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 230.310 0.000 230.610 1.000 ;
    END
  END um_ow[325]
  PIN um_ow[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 227.550 0.000 227.850 1.000 ;
    END
  END um_ow[326]
  PIN um_ow[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 224.790 0.000 225.090 1.000 ;
    END
  END um_ow[327]
  PIN um_ow[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 222.030 0.000 222.330 1.000 ;
    END
  END um_ow[328]
  PIN um_ow[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 219.270 0.000 219.570 1.000 ;
    END
  END um_ow[329]
  PIN um_ow[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1265.310 0.000 1265.610 1.000 ;
    END
  END um_ow[32]
  PIN um_ow[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 216.510 0.000 216.810 1.000 ;
    END
  END um_ow[330]
  PIN um_ow[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 213.750 0.000 214.050 1.000 ;
    END
  END um_ow[331]
  PIN um_ow[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 210.990 0.000 211.290 1.000 ;
    END
  END um_ow[332]
  PIN um_ow[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 208.230 0.000 208.530 1.000 ;
    END
  END um_ow[333]
  PIN um_ow[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 205.470 0.000 205.770 1.000 ;
    END
  END um_ow[334]
  PIN um_ow[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 202.710 0.000 203.010 1.000 ;
    END
  END um_ow[335]
  PIN um_ow[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 95.990 53.400 96.290 54.400 ;
    END
  END um_ow[336]
  PIN um_ow[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 93.230 53.400 93.530 54.400 ;
    END
  END um_ow[337]
  PIN um_ow[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 90.470 53.400 90.770 54.400 ;
    END
  END um_ow[338]
  PIN um_ow[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 87.710 53.400 88.010 54.400 ;
    END
  END um_ow[339]
  PIN um_ow[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met4 ;
        RECT 1262.550 0.000 1262.850 1.000 ;
    END
  END um_ow[33]
  PIN um_ow[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 84.950 53.400 85.250 54.400 ;
    END
  END um_ow[340]
  PIN um_ow[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 82.190 53.400 82.490 54.400 ;
    END
  END um_ow[341]
  PIN um_ow[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 79.430 53.400 79.730 54.400 ;
    END
  END um_ow[342]
  PIN um_ow[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 76.670 53.400 76.970 54.400 ;
    END
  END um_ow[343]
  PIN um_ow[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 73.910 53.400 74.210 54.400 ;
    END
  END um_ow[344]
  PIN um_ow[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 71.150 53.400 71.450 54.400 ;
    END
  END um_ow[345]
  PIN um_ow[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 68.390 53.400 68.690 54.400 ;
    END
  END um_ow[346]
  PIN um_ow[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 65.630 53.400 65.930 54.400 ;
    END
  END um_ow[347]
  PIN um_ow[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 62.870 53.400 63.170 54.400 ;
    END
  END um_ow[348]
  PIN um_ow[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 60.110 53.400 60.410 54.400 ;
    END
  END um_ow[349]
  PIN um_ow[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1259.790 0.000 1260.090 1.000 ;
    END
  END um_ow[34]
  PIN um_ow[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 57.350 53.400 57.650 54.400 ;
    END
  END um_ow[350]
  PIN um_ow[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 54.590 53.400 54.890 54.400 ;
    END
  END um_ow[351]
  PIN um_ow[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 51.830 53.400 52.130 54.400 ;
    END
  END um_ow[352]
  PIN um_ow[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 49.070 53.400 49.370 54.400 ;
    END
  END um_ow[353]
  PIN um_ow[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 46.310 53.400 46.610 54.400 ;
    END
  END um_ow[354]
  PIN um_ow[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 43.550 53.400 43.850 54.400 ;
    END
  END um_ow[355]
  PIN um_ow[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 40.790 53.400 41.090 54.400 ;
    END
  END um_ow[356]
  PIN um_ow[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 38.030 53.400 38.330 54.400 ;
    END
  END um_ow[357]
  PIN um_ow[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 35.270 53.400 35.570 54.400 ;
    END
  END um_ow[358]
  PIN um_ow[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 32.510 53.400 32.810 54.400 ;
    END
  END um_ow[359]
  PIN um_ow[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1257.030 0.000 1257.330 1.000 ;
    END
  END um_ow[35]
  PIN um_ow[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 95.990 0.000 96.290 1.000 ;
    END
  END um_ow[360]
  PIN um_ow[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 93.230 0.000 93.530 1.000 ;
    END
  END um_ow[361]
  PIN um_ow[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 90.470 0.000 90.770 1.000 ;
    END
  END um_ow[362]
  PIN um_ow[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 87.710 0.000 88.010 1.000 ;
    END
  END um_ow[363]
  PIN um_ow[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 84.950 0.000 85.250 1.000 ;
    END
  END um_ow[364]
  PIN um_ow[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 82.190 0.000 82.490 1.000 ;
    END
  END um_ow[365]
  PIN um_ow[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 79.430 0.000 79.730 1.000 ;
    END
  END um_ow[366]
  PIN um_ow[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 76.670 0.000 76.970 1.000 ;
    END
  END um_ow[367]
  PIN um_ow[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 73.910 0.000 74.210 1.000 ;
    END
  END um_ow[368]
  PIN um_ow[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 71.150 0.000 71.450 1.000 ;
    END
  END um_ow[369]
  PIN um_ow[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1254.270 0.000 1254.570 1.000 ;
    END
  END um_ow[36]
  PIN um_ow[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 68.390 0.000 68.690 1.000 ;
    END
  END um_ow[370]
  PIN um_ow[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 65.630 0.000 65.930 1.000 ;
    END
  END um_ow[371]
  PIN um_ow[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 62.870 0.000 63.170 1.000 ;
    END
  END um_ow[372]
  PIN um_ow[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 60.110 0.000 60.410 1.000 ;
    END
  END um_ow[373]
  PIN um_ow[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 57.350 0.000 57.650 1.000 ;
    END
  END um_ow[374]
  PIN um_ow[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 54.590 0.000 54.890 1.000 ;
    END
  END um_ow[375]
  PIN um_ow[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 51.830 0.000 52.130 1.000 ;
    END
  END um_ow[376]
  PIN um_ow[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 49.070 0.000 49.370 1.000 ;
    END
  END um_ow[377]
  PIN um_ow[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 46.310 0.000 46.610 1.000 ;
    END
  END um_ow[378]
  PIN um_ow[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 43.550 0.000 43.850 1.000 ;
    END
  END um_ow[379]
  PIN um_ow[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1251.510 0.000 1251.810 1.000 ;
    END
  END um_ow[37]
  PIN um_ow[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 40.790 0.000 41.090 1.000 ;
    END
  END um_ow[380]
  PIN um_ow[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 38.030 0.000 38.330 1.000 ;
    END
  END um_ow[381]
  PIN um_ow[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 35.270 0.000 35.570 1.000 ;
    END
  END um_ow[382]
  PIN um_ow[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 32.510 0.000 32.810 1.000 ;
    END
  END um_ow[383]
  PIN um_ow[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1248.750 0.000 1249.050 1.000 ;
    END
  END um_ow[38]
  PIN um_ow[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1245.990 0.000 1246.290 1.000 ;
    END
  END um_ow[39]
  PIN um_ow[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1279.110 53.400 1279.410 54.400 ;
    END
  END um_ow[3]
  PIN um_ow[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1243.230 0.000 1243.530 1.000 ;
    END
  END um_ow[40]
  PIN um_ow[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1240.470 0.000 1240.770 1.000 ;
    END
  END um_ow[41]
  PIN um_ow[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met4 ;
        RECT 1237.710 0.000 1238.010 1.000 ;
    END
  END um_ow[42]
  PIN um_ow[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1234.950 0.000 1235.250 1.000 ;
    END
  END um_ow[43]
  PIN um_ow[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1232.190 0.000 1232.490 1.000 ;
    END
  END um_ow[44]
  PIN um_ow[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1229.430 0.000 1229.730 1.000 ;
    END
  END um_ow[45]
  PIN um_ow[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1226.670 0.000 1226.970 1.000 ;
    END
  END um_ow[46]
  PIN um_ow[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1223.910 0.000 1224.210 1.000 ;
    END
  END um_ow[47]
  PIN um_ow[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1117.190 53.400 1117.490 54.400 ;
    END
  END um_ow[48]
  PIN um_ow[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1114.430 53.400 1114.730 54.400 ;
    END
  END um_ow[49]
  PIN um_ow[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1276.350 53.400 1276.650 54.400 ;
    END
  END um_ow[4]
  PIN um_ow[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1111.670 53.400 1111.970 54.400 ;
    END
  END um_ow[50]
  PIN um_ow[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1108.910 53.400 1109.210 54.400 ;
    END
  END um_ow[51]
  PIN um_ow[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1106.150 53.400 1106.450 54.400 ;
    END
  END um_ow[52]
  PIN um_ow[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1103.390 53.400 1103.690 54.400 ;
    END
  END um_ow[53]
  PIN um_ow[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1100.630 53.400 1100.930 54.400 ;
    END
  END um_ow[54]
  PIN um_ow[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1097.870 53.400 1098.170 54.400 ;
    END
  END um_ow[55]
  PIN um_ow[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1095.110 53.400 1095.410 54.400 ;
    END
  END um_ow[56]
  PIN um_ow[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1092.350 53.400 1092.650 54.400 ;
    END
  END um_ow[57]
  PIN um_ow[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1089.590 53.400 1089.890 54.400 ;
    END
  END um_ow[58]
  PIN um_ow[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1086.830 53.400 1087.130 54.400 ;
    END
  END um_ow[59]
  PIN um_ow[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1273.590 53.400 1273.890 54.400 ;
    END
  END um_ow[5]
  PIN um_ow[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1084.070 53.400 1084.370 54.400 ;
    END
  END um_ow[60]
  PIN um_ow[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1081.310 53.400 1081.610 54.400 ;
    END
  END um_ow[61]
  PIN um_ow[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1078.550 53.400 1078.850 54.400 ;
    END
  END um_ow[62]
  PIN um_ow[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1075.790 53.400 1076.090 54.400 ;
    END
  END um_ow[63]
  PIN um_ow[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1073.030 53.400 1073.330 54.400 ;
    END
  END um_ow[64]
  PIN um_ow[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1070.270 53.400 1070.570 54.400 ;
    END
  END um_ow[65]
  PIN um_ow[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1067.510 53.400 1067.810 54.400 ;
    END
  END um_ow[66]
  PIN um_ow[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1064.750 53.400 1065.050 54.400 ;
    END
  END um_ow[67]
  PIN um_ow[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1061.990 53.400 1062.290 54.400 ;
    END
  END um_ow[68]
  PIN um_ow[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1059.230 53.400 1059.530 54.400 ;
    END
  END um_ow[69]
  PIN um_ow[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1270.830 53.400 1271.130 54.400 ;
    END
  END um_ow[6]
  PIN um_ow[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1056.470 53.400 1056.770 54.400 ;
    END
  END um_ow[70]
  PIN um_ow[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1053.710 53.400 1054.010 54.400 ;
    END
  END um_ow[71]
  PIN um_ow[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1117.190 0.000 1117.490 1.000 ;
    END
  END um_ow[72]
  PIN um_ow[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1114.430 0.000 1114.730 1.000 ;
    END
  END um_ow[73]
  PIN um_ow[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1111.670 0.000 1111.970 1.000 ;
    END
  END um_ow[74]
  PIN um_ow[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1108.910 0.000 1109.210 1.000 ;
    END
  END um_ow[75]
  PIN um_ow[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1106.150 0.000 1106.450 1.000 ;
    END
  END um_ow[76]
  PIN um_ow[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1103.390 0.000 1103.690 1.000 ;
    END
  END um_ow[77]
  PIN um_ow[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1100.630 0.000 1100.930 1.000 ;
    END
  END um_ow[78]
  PIN um_ow[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1097.870 0.000 1098.170 1.000 ;
    END
  END um_ow[79]
  PIN um_ow[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1268.070 53.400 1268.370 54.400 ;
    END
  END um_ow[7]
  PIN um_ow[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1095.110 0.000 1095.410 1.000 ;
    END
  END um_ow[80]
  PIN um_ow[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1092.350 0.000 1092.650 1.000 ;
    END
  END um_ow[81]
  PIN um_ow[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1089.590 0.000 1089.890 1.000 ;
    END
  END um_ow[82]
  PIN um_ow[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1086.830 0.000 1087.130 1.000 ;
    END
  END um_ow[83]
  PIN um_ow[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1084.070 0.000 1084.370 1.000 ;
    END
  END um_ow[84]
  PIN um_ow[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1081.310 0.000 1081.610 1.000 ;
    END
  END um_ow[85]
  PIN um_ow[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1078.550 0.000 1078.850 1.000 ;
    END
  END um_ow[86]
  PIN um_ow[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1075.790 0.000 1076.090 1.000 ;
    END
  END um_ow[87]
  PIN um_ow[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1073.030 0.000 1073.330 1.000 ;
    END
  END um_ow[88]
  PIN um_ow[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1070.270 0.000 1070.570 1.000 ;
    END
  END um_ow[89]
  PIN um_ow[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1265.310 53.400 1265.610 54.400 ;
    END
  END um_ow[8]
  PIN um_ow[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1067.510 0.000 1067.810 1.000 ;
    END
  END um_ow[90]
  PIN um_ow[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1064.750 0.000 1065.050 1.000 ;
    END
  END um_ow[91]
  PIN um_ow[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1061.990 0.000 1062.290 1.000 ;
    END
  END um_ow[92]
  PIN um_ow[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1059.230 0.000 1059.530 1.000 ;
    END
  END um_ow[93]
  PIN um_ow[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1056.470 0.000 1056.770 1.000 ;
    END
  END um_ow[94]
  PIN um_ow[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1053.710 0.000 1054.010 1.000 ;
    END
  END um_ow[95]
  PIN um_ow[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 946.990 53.400 947.290 54.400 ;
    END
  END um_ow[96]
  PIN um_ow[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 944.230 53.400 944.530 54.400 ;
    END
  END um_ow[97]
  PIN um_ow[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 941.470 53.400 941.770 54.400 ;
    END
  END um_ow[98]
  PIN um_ow[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 938.710 53.400 939.010 54.400 ;
    END
  END um_ow[99]
  PIN um_ow[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 1262.550 53.400 1262.850 54.400 ;
    END
  END um_ow[9]
  PIN um_pg_vdd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 1195.390 53.400 1195.690 54.400 ;
    END
  END um_pg_vdd[0]
  PIN um_pg_vdd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 344.390 53.400 344.690 54.400 ;
    END
  END um_pg_vdd[10]
  PIN um_pg_vdd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 344.390 0.000 344.690 1.000 ;
    END
  END um_pg_vdd[11]
  PIN um_pg_vdd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 174.190 53.400 174.490 54.400 ;
    END
  END um_pg_vdd[12]
  PIN um_pg_vdd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 174.190 0.000 174.490 1.000 ;
    END
  END um_pg_vdd[13]
  PIN um_pg_vdd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 3.990 53.400 4.290 54.400 ;
    END
  END um_pg_vdd[14]
  PIN um_pg_vdd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 3.990 0.000 4.290 1.000 ;
    END
  END um_pg_vdd[15]
  PIN um_pg_vdd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 1195.390 0.000 1195.690 1.000 ;
    END
  END um_pg_vdd[1]
  PIN um_pg_vdd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 1025.190 53.400 1025.490 54.400 ;
    END
  END um_pg_vdd[2]
  PIN um_pg_vdd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 1025.190 0.000 1025.490 1.000 ;
    END
  END um_pg_vdd[3]
  PIN um_pg_vdd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 854.990 53.400 855.290 54.400 ;
    END
  END um_pg_vdd[4]
  PIN um_pg_vdd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 854.990 0.000 855.290 1.000 ;
    END
  END um_pg_vdd[5]
  PIN um_pg_vdd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 684.790 53.400 685.090 54.400 ;
    END
  END um_pg_vdd[6]
  PIN um_pg_vdd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 684.790 0.000 685.090 1.000 ;
    END
  END um_pg_vdd[7]
  PIN um_pg_vdd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 514.590 53.400 514.890 54.400 ;
    END
  END um_pg_vdd[8]
  PIN um_pg_vdd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 514.590 0.000 514.890 1.000 ;
    END
  END um_pg_vdd[9]
  OBS
      LAYER nwell ;
        RECT 2.570 47.545 1357.190 50.375 ;
        RECT 2.570 42.105 1357.190 44.935 ;
        RECT 2.570 36.665 1357.190 39.495 ;
        RECT 2.570 31.225 1357.190 34.055 ;
        RECT 2.570 25.785 1357.190 28.615 ;
        RECT 2.570 20.345 1357.190 23.175 ;
        RECT 2.570 14.905 1357.190 17.735 ;
        RECT 2.570 9.465 1357.190 12.295 ;
        RECT 2.570 4.025 1357.190 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 1357.000 51.765 ;
      LAYER met1 ;
        RECT 2.760 0.040 1357.000 54.360 ;
      LAYER met2 ;
        RECT 6.530 0.010 1356.450 54.390 ;
      LAYER met3 ;
        RECT 3.950 47.810 1358.760 53.545 ;
        RECT 3.950 5.230 1358.360 47.810 ;
        RECT 3.950 0.175 1358.760 5.230 ;
      LAYER met4 ;
        RECT 4.690 53.000 29.350 53.545 ;
        RECT 30.450 53.000 32.110 53.545 ;
        RECT 33.210 53.000 34.870 53.545 ;
        RECT 35.970 53.000 37.630 53.545 ;
        RECT 38.730 53.000 40.390 53.545 ;
        RECT 41.490 53.000 43.150 53.545 ;
        RECT 44.250 53.000 45.910 53.545 ;
        RECT 47.010 53.000 48.670 53.545 ;
        RECT 49.770 53.000 51.430 53.545 ;
        RECT 52.530 53.000 54.190 53.545 ;
        RECT 55.290 53.000 56.950 53.545 ;
        RECT 58.050 53.000 59.710 53.545 ;
        RECT 60.810 53.000 62.470 53.545 ;
        RECT 63.570 53.000 65.230 53.545 ;
        RECT 66.330 53.000 67.990 53.545 ;
        RECT 69.090 53.000 70.750 53.545 ;
        RECT 71.850 53.000 73.510 53.545 ;
        RECT 74.610 53.000 76.270 53.545 ;
        RECT 77.370 53.000 79.030 53.545 ;
        RECT 80.130 53.000 81.790 53.545 ;
        RECT 82.890 53.000 84.550 53.545 ;
        RECT 85.650 53.000 87.310 53.545 ;
        RECT 88.410 53.000 90.070 53.545 ;
        RECT 91.170 53.000 92.830 53.545 ;
        RECT 93.930 53.000 95.590 53.545 ;
        RECT 96.690 53.000 98.350 53.545 ;
        RECT 99.450 53.000 101.110 53.545 ;
        RECT 102.210 53.000 103.870 53.545 ;
        RECT 104.970 53.000 106.630 53.545 ;
        RECT 107.730 53.000 109.390 53.545 ;
        RECT 110.490 53.000 112.150 53.545 ;
        RECT 113.250 53.000 114.910 53.545 ;
        RECT 116.010 53.000 117.670 53.545 ;
        RECT 118.770 53.000 120.430 53.545 ;
        RECT 121.530 53.000 123.190 53.545 ;
        RECT 124.290 53.000 125.950 53.545 ;
        RECT 127.050 53.000 128.710 53.545 ;
        RECT 129.810 53.000 131.470 53.545 ;
        RECT 132.570 53.000 134.230 53.545 ;
        RECT 135.330 53.000 136.990 53.545 ;
        RECT 138.090 53.000 139.750 53.545 ;
        RECT 140.850 53.000 142.510 53.545 ;
        RECT 143.610 53.000 145.270 53.545 ;
        RECT 146.370 53.000 148.030 53.545 ;
        RECT 149.130 53.000 173.790 53.545 ;
        RECT 174.890 53.000 199.550 53.545 ;
        RECT 200.650 53.000 202.310 53.545 ;
        RECT 203.410 53.000 205.070 53.545 ;
        RECT 206.170 53.000 207.830 53.545 ;
        RECT 208.930 53.000 210.590 53.545 ;
        RECT 211.690 53.000 213.350 53.545 ;
        RECT 214.450 53.000 216.110 53.545 ;
        RECT 217.210 53.000 218.870 53.545 ;
        RECT 219.970 53.000 221.630 53.545 ;
        RECT 222.730 53.000 224.390 53.545 ;
        RECT 225.490 53.000 227.150 53.545 ;
        RECT 228.250 53.000 229.910 53.545 ;
        RECT 231.010 53.000 232.670 53.545 ;
        RECT 233.770 53.000 235.430 53.545 ;
        RECT 236.530 53.000 238.190 53.545 ;
        RECT 239.290 53.000 240.950 53.545 ;
        RECT 242.050 53.000 243.710 53.545 ;
        RECT 244.810 53.000 246.470 53.545 ;
        RECT 247.570 53.000 249.230 53.545 ;
        RECT 250.330 53.000 251.990 53.545 ;
        RECT 253.090 53.000 254.750 53.545 ;
        RECT 255.850 53.000 257.510 53.545 ;
        RECT 258.610 53.000 260.270 53.545 ;
        RECT 261.370 53.000 263.030 53.545 ;
        RECT 264.130 53.000 265.790 53.545 ;
        RECT 266.890 53.000 268.550 53.545 ;
        RECT 269.650 53.000 271.310 53.545 ;
        RECT 272.410 53.000 274.070 53.545 ;
        RECT 275.170 53.000 276.830 53.545 ;
        RECT 277.930 53.000 279.590 53.545 ;
        RECT 280.690 53.000 282.350 53.545 ;
        RECT 283.450 53.000 285.110 53.545 ;
        RECT 286.210 53.000 287.870 53.545 ;
        RECT 288.970 53.000 290.630 53.545 ;
        RECT 291.730 53.000 293.390 53.545 ;
        RECT 294.490 53.000 296.150 53.545 ;
        RECT 297.250 53.000 298.910 53.545 ;
        RECT 300.010 53.000 301.670 53.545 ;
        RECT 302.770 53.000 304.430 53.545 ;
        RECT 305.530 53.000 307.190 53.545 ;
        RECT 308.290 53.000 309.950 53.545 ;
        RECT 311.050 53.000 312.710 53.545 ;
        RECT 313.810 53.000 315.470 53.545 ;
        RECT 316.570 53.000 318.230 53.545 ;
        RECT 319.330 53.000 343.990 53.545 ;
        RECT 345.090 53.000 369.750 53.545 ;
        RECT 370.850 53.000 372.510 53.545 ;
        RECT 373.610 53.000 375.270 53.545 ;
        RECT 376.370 53.000 378.030 53.545 ;
        RECT 379.130 53.000 380.790 53.545 ;
        RECT 381.890 53.000 383.550 53.545 ;
        RECT 384.650 53.000 386.310 53.545 ;
        RECT 387.410 53.000 389.070 53.545 ;
        RECT 390.170 53.000 391.830 53.545 ;
        RECT 392.930 53.000 394.590 53.545 ;
        RECT 395.690 53.000 397.350 53.545 ;
        RECT 398.450 53.000 400.110 53.545 ;
        RECT 401.210 53.000 402.870 53.545 ;
        RECT 403.970 53.000 405.630 53.545 ;
        RECT 406.730 53.000 408.390 53.545 ;
        RECT 409.490 53.000 411.150 53.545 ;
        RECT 412.250 53.000 413.910 53.545 ;
        RECT 415.010 53.000 416.670 53.545 ;
        RECT 417.770 53.000 419.430 53.545 ;
        RECT 420.530 53.000 422.190 53.545 ;
        RECT 423.290 53.000 424.950 53.545 ;
        RECT 426.050 53.000 427.710 53.545 ;
        RECT 428.810 53.000 430.470 53.545 ;
        RECT 431.570 53.000 433.230 53.545 ;
        RECT 434.330 53.000 435.990 53.545 ;
        RECT 437.090 53.000 438.750 53.545 ;
        RECT 439.850 53.000 441.510 53.545 ;
        RECT 442.610 53.000 444.270 53.545 ;
        RECT 445.370 53.000 447.030 53.545 ;
        RECT 448.130 53.000 449.790 53.545 ;
        RECT 450.890 53.000 452.550 53.545 ;
        RECT 453.650 53.000 455.310 53.545 ;
        RECT 456.410 53.000 458.070 53.545 ;
        RECT 459.170 53.000 460.830 53.545 ;
        RECT 461.930 53.000 463.590 53.545 ;
        RECT 464.690 53.000 466.350 53.545 ;
        RECT 467.450 53.000 469.110 53.545 ;
        RECT 470.210 53.000 471.870 53.545 ;
        RECT 472.970 53.000 474.630 53.545 ;
        RECT 475.730 53.000 477.390 53.545 ;
        RECT 478.490 53.000 480.150 53.545 ;
        RECT 481.250 53.000 482.910 53.545 ;
        RECT 484.010 53.000 485.670 53.545 ;
        RECT 486.770 53.000 488.430 53.545 ;
        RECT 489.530 53.000 514.190 53.545 ;
        RECT 515.290 53.000 539.950 53.545 ;
        RECT 541.050 53.000 542.710 53.545 ;
        RECT 543.810 53.000 545.470 53.545 ;
        RECT 546.570 53.000 548.230 53.545 ;
        RECT 549.330 53.000 550.990 53.545 ;
        RECT 552.090 53.000 553.750 53.545 ;
        RECT 554.850 53.000 556.510 53.545 ;
        RECT 557.610 53.000 559.270 53.545 ;
        RECT 560.370 53.000 562.030 53.545 ;
        RECT 563.130 53.000 564.790 53.545 ;
        RECT 565.890 53.000 567.550 53.545 ;
        RECT 568.650 53.000 570.310 53.545 ;
        RECT 571.410 53.000 573.070 53.545 ;
        RECT 574.170 53.000 575.830 53.545 ;
        RECT 576.930 53.000 578.590 53.545 ;
        RECT 579.690 53.000 581.350 53.545 ;
        RECT 582.450 53.000 584.110 53.545 ;
        RECT 585.210 53.000 586.870 53.545 ;
        RECT 587.970 53.000 589.630 53.545 ;
        RECT 590.730 53.000 592.390 53.545 ;
        RECT 593.490 53.000 595.150 53.545 ;
        RECT 596.250 53.000 597.910 53.545 ;
        RECT 599.010 53.000 600.670 53.545 ;
        RECT 601.770 53.000 603.430 53.545 ;
        RECT 604.530 53.000 606.190 53.545 ;
        RECT 607.290 53.000 608.950 53.545 ;
        RECT 610.050 53.000 611.710 53.545 ;
        RECT 612.810 53.000 614.470 53.545 ;
        RECT 615.570 53.000 617.230 53.545 ;
        RECT 618.330 53.000 619.990 53.545 ;
        RECT 621.090 53.000 622.750 53.545 ;
        RECT 623.850 53.000 625.510 53.545 ;
        RECT 626.610 53.000 628.270 53.545 ;
        RECT 629.370 53.000 631.030 53.545 ;
        RECT 632.130 53.000 633.790 53.545 ;
        RECT 634.890 53.000 636.550 53.545 ;
        RECT 637.650 53.000 639.310 53.545 ;
        RECT 640.410 53.000 642.070 53.545 ;
        RECT 643.170 53.000 644.830 53.545 ;
        RECT 645.930 53.000 647.590 53.545 ;
        RECT 648.690 53.000 650.350 53.545 ;
        RECT 651.450 53.000 653.110 53.545 ;
        RECT 654.210 53.000 655.870 53.545 ;
        RECT 656.970 53.000 658.630 53.545 ;
        RECT 659.730 53.000 684.390 53.545 ;
        RECT 685.490 53.000 710.150 53.545 ;
        RECT 711.250 53.000 712.910 53.545 ;
        RECT 714.010 53.000 715.670 53.545 ;
        RECT 716.770 53.000 718.430 53.545 ;
        RECT 719.530 53.000 721.190 53.545 ;
        RECT 722.290 53.000 723.950 53.545 ;
        RECT 725.050 53.000 726.710 53.545 ;
        RECT 727.810 53.000 729.470 53.545 ;
        RECT 730.570 53.000 732.230 53.545 ;
        RECT 733.330 53.000 734.990 53.545 ;
        RECT 736.090 53.000 737.750 53.545 ;
        RECT 738.850 53.000 740.510 53.545 ;
        RECT 741.610 53.000 743.270 53.545 ;
        RECT 744.370 53.000 746.030 53.545 ;
        RECT 747.130 53.000 748.790 53.545 ;
        RECT 749.890 53.000 751.550 53.545 ;
        RECT 752.650 53.000 754.310 53.545 ;
        RECT 755.410 53.000 757.070 53.545 ;
        RECT 758.170 53.000 759.830 53.545 ;
        RECT 760.930 53.000 762.590 53.545 ;
        RECT 763.690 53.000 765.350 53.545 ;
        RECT 766.450 53.000 768.110 53.545 ;
        RECT 769.210 53.000 770.870 53.545 ;
        RECT 771.970 53.000 773.630 53.545 ;
        RECT 774.730 53.000 776.390 53.545 ;
        RECT 777.490 53.000 779.150 53.545 ;
        RECT 780.250 53.000 781.910 53.545 ;
        RECT 783.010 53.000 784.670 53.545 ;
        RECT 785.770 53.000 787.430 53.545 ;
        RECT 788.530 53.000 790.190 53.545 ;
        RECT 791.290 53.000 792.950 53.545 ;
        RECT 794.050 53.000 795.710 53.545 ;
        RECT 796.810 53.000 798.470 53.545 ;
        RECT 799.570 53.000 801.230 53.545 ;
        RECT 802.330 53.000 803.990 53.545 ;
        RECT 805.090 53.000 806.750 53.545 ;
        RECT 807.850 53.000 809.510 53.545 ;
        RECT 810.610 53.000 812.270 53.545 ;
        RECT 813.370 53.000 815.030 53.545 ;
        RECT 816.130 53.000 817.790 53.545 ;
        RECT 818.890 53.000 820.550 53.545 ;
        RECT 821.650 53.000 823.310 53.545 ;
        RECT 824.410 53.000 826.070 53.545 ;
        RECT 827.170 53.000 828.830 53.545 ;
        RECT 829.930 53.000 854.590 53.545 ;
        RECT 855.690 53.000 880.350 53.545 ;
        RECT 881.450 53.000 883.110 53.545 ;
        RECT 884.210 53.000 885.870 53.545 ;
        RECT 886.970 53.000 888.630 53.545 ;
        RECT 889.730 53.000 891.390 53.545 ;
        RECT 892.490 53.000 894.150 53.545 ;
        RECT 895.250 53.000 896.910 53.545 ;
        RECT 898.010 53.000 899.670 53.545 ;
        RECT 900.770 53.000 902.430 53.545 ;
        RECT 903.530 53.000 905.190 53.545 ;
        RECT 906.290 53.000 907.950 53.545 ;
        RECT 909.050 53.000 910.710 53.545 ;
        RECT 911.810 53.000 913.470 53.545 ;
        RECT 914.570 53.000 916.230 53.545 ;
        RECT 917.330 53.000 918.990 53.545 ;
        RECT 920.090 53.000 921.750 53.545 ;
        RECT 922.850 53.000 924.510 53.545 ;
        RECT 925.610 53.000 927.270 53.545 ;
        RECT 928.370 53.000 930.030 53.545 ;
        RECT 931.130 53.000 932.790 53.545 ;
        RECT 933.890 53.000 935.550 53.545 ;
        RECT 936.650 53.000 938.310 53.545 ;
        RECT 939.410 53.000 941.070 53.545 ;
        RECT 942.170 53.000 943.830 53.545 ;
        RECT 944.930 53.000 946.590 53.545 ;
        RECT 947.690 53.000 949.350 53.545 ;
        RECT 950.450 53.000 952.110 53.545 ;
        RECT 953.210 53.000 954.870 53.545 ;
        RECT 955.970 53.000 957.630 53.545 ;
        RECT 958.730 53.000 960.390 53.545 ;
        RECT 961.490 53.000 963.150 53.545 ;
        RECT 964.250 53.000 965.910 53.545 ;
        RECT 967.010 53.000 968.670 53.545 ;
        RECT 969.770 53.000 971.430 53.545 ;
        RECT 972.530 53.000 974.190 53.545 ;
        RECT 975.290 53.000 976.950 53.545 ;
        RECT 978.050 53.000 979.710 53.545 ;
        RECT 980.810 53.000 982.470 53.545 ;
        RECT 983.570 53.000 985.230 53.545 ;
        RECT 986.330 53.000 987.990 53.545 ;
        RECT 989.090 53.000 990.750 53.545 ;
        RECT 991.850 53.000 993.510 53.545 ;
        RECT 994.610 53.000 996.270 53.545 ;
        RECT 997.370 53.000 999.030 53.545 ;
        RECT 1000.130 53.000 1024.790 53.545 ;
        RECT 1025.890 53.000 1050.550 53.545 ;
        RECT 1051.650 53.000 1053.310 53.545 ;
        RECT 1054.410 53.000 1056.070 53.545 ;
        RECT 1057.170 53.000 1058.830 53.545 ;
        RECT 1059.930 53.000 1061.590 53.545 ;
        RECT 1062.690 53.000 1064.350 53.545 ;
        RECT 1065.450 53.000 1067.110 53.545 ;
        RECT 1068.210 53.000 1069.870 53.545 ;
        RECT 1070.970 53.000 1072.630 53.545 ;
        RECT 1073.730 53.000 1075.390 53.545 ;
        RECT 1076.490 53.000 1078.150 53.545 ;
        RECT 1079.250 53.000 1080.910 53.545 ;
        RECT 1082.010 53.000 1083.670 53.545 ;
        RECT 1084.770 53.000 1086.430 53.545 ;
        RECT 1087.530 53.000 1089.190 53.545 ;
        RECT 1090.290 53.000 1091.950 53.545 ;
        RECT 1093.050 53.000 1094.710 53.545 ;
        RECT 1095.810 53.000 1097.470 53.545 ;
        RECT 1098.570 53.000 1100.230 53.545 ;
        RECT 1101.330 53.000 1102.990 53.545 ;
        RECT 1104.090 53.000 1105.750 53.545 ;
        RECT 1106.850 53.000 1108.510 53.545 ;
        RECT 1109.610 53.000 1111.270 53.545 ;
        RECT 1112.370 53.000 1114.030 53.545 ;
        RECT 1115.130 53.000 1116.790 53.545 ;
        RECT 1117.890 53.000 1119.550 53.545 ;
        RECT 1120.650 53.000 1122.310 53.545 ;
        RECT 1123.410 53.000 1125.070 53.545 ;
        RECT 1126.170 53.000 1127.830 53.545 ;
        RECT 1128.930 53.000 1130.590 53.545 ;
        RECT 1131.690 53.000 1133.350 53.545 ;
        RECT 1134.450 53.000 1136.110 53.545 ;
        RECT 1137.210 53.000 1138.870 53.545 ;
        RECT 1139.970 53.000 1141.630 53.545 ;
        RECT 1142.730 53.000 1144.390 53.545 ;
        RECT 1145.490 53.000 1147.150 53.545 ;
        RECT 1148.250 53.000 1149.910 53.545 ;
        RECT 1151.010 53.000 1152.670 53.545 ;
        RECT 1153.770 53.000 1155.430 53.545 ;
        RECT 1156.530 53.000 1158.190 53.545 ;
        RECT 1159.290 53.000 1160.950 53.545 ;
        RECT 1162.050 53.000 1163.710 53.545 ;
        RECT 1164.810 53.000 1166.470 53.545 ;
        RECT 1167.570 53.000 1169.230 53.545 ;
        RECT 1170.330 53.000 1194.990 53.545 ;
        RECT 1196.090 53.000 1220.750 53.545 ;
        RECT 1221.850 53.000 1223.510 53.545 ;
        RECT 1224.610 53.000 1226.270 53.545 ;
        RECT 1227.370 53.000 1229.030 53.545 ;
        RECT 1230.130 53.000 1231.790 53.545 ;
        RECT 1232.890 53.000 1234.550 53.545 ;
        RECT 1235.650 53.000 1237.310 53.545 ;
        RECT 1238.410 53.000 1240.070 53.545 ;
        RECT 1241.170 53.000 1242.830 53.545 ;
        RECT 1243.930 53.000 1245.590 53.545 ;
        RECT 1246.690 53.000 1248.350 53.545 ;
        RECT 1249.450 53.000 1251.110 53.545 ;
        RECT 1252.210 53.000 1253.870 53.545 ;
        RECT 1254.970 53.000 1256.630 53.545 ;
        RECT 1257.730 53.000 1259.390 53.545 ;
        RECT 1260.490 53.000 1262.150 53.545 ;
        RECT 1263.250 53.000 1264.910 53.545 ;
        RECT 1266.010 53.000 1267.670 53.545 ;
        RECT 1268.770 53.000 1270.430 53.545 ;
        RECT 1271.530 53.000 1273.190 53.545 ;
        RECT 1274.290 53.000 1275.950 53.545 ;
        RECT 1277.050 53.000 1278.710 53.545 ;
        RECT 1279.810 53.000 1281.470 53.545 ;
        RECT 1282.570 53.000 1284.230 53.545 ;
        RECT 1285.330 53.000 1286.990 53.545 ;
        RECT 1288.090 53.000 1289.750 53.545 ;
        RECT 1290.850 53.000 1292.510 53.545 ;
        RECT 1293.610 53.000 1295.270 53.545 ;
        RECT 1296.370 53.000 1298.030 53.545 ;
        RECT 1299.130 53.000 1300.790 53.545 ;
        RECT 1301.890 53.000 1303.550 53.545 ;
        RECT 1304.650 53.000 1306.310 53.545 ;
        RECT 1307.410 53.000 1309.070 53.545 ;
        RECT 1310.170 53.000 1311.830 53.545 ;
        RECT 1312.930 53.000 1314.590 53.545 ;
        RECT 1315.690 53.000 1317.350 53.545 ;
        RECT 1318.450 53.000 1320.110 53.545 ;
        RECT 1321.210 53.000 1322.870 53.545 ;
        RECT 1323.970 53.000 1325.630 53.545 ;
        RECT 1326.730 53.000 1328.390 53.545 ;
        RECT 1329.490 53.000 1331.150 53.545 ;
        RECT 1332.250 53.000 1333.910 53.545 ;
        RECT 1335.010 53.000 1336.670 53.545 ;
        RECT 1337.770 53.000 1339.430 53.545 ;
        RECT 3.975 52.320 1340.145 53.000 ;
        RECT 3.975 2.080 17.880 52.320 ;
        RECT 20.280 2.080 94.680 52.320 ;
        RECT 97.080 2.080 171.480 52.320 ;
        RECT 173.880 2.080 248.280 52.320 ;
        RECT 250.680 2.080 325.080 52.320 ;
        RECT 327.480 2.080 401.880 52.320 ;
        RECT 404.280 2.080 478.680 52.320 ;
        RECT 481.080 2.080 555.480 52.320 ;
        RECT 557.880 2.080 632.280 52.320 ;
        RECT 634.680 2.080 709.080 52.320 ;
        RECT 711.480 2.080 785.880 52.320 ;
        RECT 788.280 2.080 862.680 52.320 ;
        RECT 865.080 2.080 939.480 52.320 ;
        RECT 941.880 2.080 1016.280 52.320 ;
        RECT 1018.680 2.080 1093.080 52.320 ;
        RECT 1095.480 2.080 1169.880 52.320 ;
        RECT 1172.280 2.080 1246.680 52.320 ;
        RECT 1249.080 2.080 1323.480 52.320 ;
        RECT 1325.880 2.080 1340.145 52.320 ;
        RECT 3.975 1.400 1340.145 2.080 ;
        RECT 4.690 0.855 29.350 1.400 ;
        RECT 30.450 0.855 32.110 1.400 ;
        RECT 33.210 0.855 34.870 1.400 ;
        RECT 35.970 0.855 37.630 1.400 ;
        RECT 38.730 0.855 40.390 1.400 ;
        RECT 41.490 0.855 43.150 1.400 ;
        RECT 44.250 0.855 45.910 1.400 ;
        RECT 47.010 0.855 48.670 1.400 ;
        RECT 49.770 0.855 51.430 1.400 ;
        RECT 52.530 0.855 54.190 1.400 ;
        RECT 55.290 0.855 56.950 1.400 ;
        RECT 58.050 0.855 59.710 1.400 ;
        RECT 60.810 0.855 62.470 1.400 ;
        RECT 63.570 0.855 65.230 1.400 ;
        RECT 66.330 0.855 67.990 1.400 ;
        RECT 69.090 0.855 70.750 1.400 ;
        RECT 71.850 0.855 73.510 1.400 ;
        RECT 74.610 0.855 76.270 1.400 ;
        RECT 77.370 0.855 79.030 1.400 ;
        RECT 80.130 0.855 81.790 1.400 ;
        RECT 82.890 0.855 84.550 1.400 ;
        RECT 85.650 0.855 87.310 1.400 ;
        RECT 88.410 0.855 90.070 1.400 ;
        RECT 91.170 0.855 92.830 1.400 ;
        RECT 93.930 0.855 95.590 1.400 ;
        RECT 96.690 0.855 98.350 1.400 ;
        RECT 99.450 0.855 101.110 1.400 ;
        RECT 102.210 0.855 103.870 1.400 ;
        RECT 104.970 0.855 106.630 1.400 ;
        RECT 107.730 0.855 109.390 1.400 ;
        RECT 110.490 0.855 112.150 1.400 ;
        RECT 113.250 0.855 114.910 1.400 ;
        RECT 116.010 0.855 117.670 1.400 ;
        RECT 118.770 0.855 120.430 1.400 ;
        RECT 121.530 0.855 123.190 1.400 ;
        RECT 124.290 0.855 125.950 1.400 ;
        RECT 127.050 0.855 128.710 1.400 ;
        RECT 129.810 0.855 131.470 1.400 ;
        RECT 132.570 0.855 134.230 1.400 ;
        RECT 135.330 0.855 136.990 1.400 ;
        RECT 138.090 0.855 139.750 1.400 ;
        RECT 140.850 0.855 142.510 1.400 ;
        RECT 143.610 0.855 145.270 1.400 ;
        RECT 146.370 0.855 148.030 1.400 ;
        RECT 149.130 0.855 173.790 1.400 ;
        RECT 174.890 0.855 199.550 1.400 ;
        RECT 200.650 0.855 202.310 1.400 ;
        RECT 203.410 0.855 205.070 1.400 ;
        RECT 206.170 0.855 207.830 1.400 ;
        RECT 208.930 0.855 210.590 1.400 ;
        RECT 211.690 0.855 213.350 1.400 ;
        RECT 214.450 0.855 216.110 1.400 ;
        RECT 217.210 0.855 218.870 1.400 ;
        RECT 219.970 0.855 221.630 1.400 ;
        RECT 222.730 0.855 224.390 1.400 ;
        RECT 225.490 0.855 227.150 1.400 ;
        RECT 228.250 0.855 229.910 1.400 ;
        RECT 231.010 0.855 232.670 1.400 ;
        RECT 233.770 0.855 235.430 1.400 ;
        RECT 236.530 0.855 238.190 1.400 ;
        RECT 239.290 0.855 240.950 1.400 ;
        RECT 242.050 0.855 243.710 1.400 ;
        RECT 244.810 0.855 246.470 1.400 ;
        RECT 247.570 0.855 249.230 1.400 ;
        RECT 250.330 0.855 251.990 1.400 ;
        RECT 253.090 0.855 254.750 1.400 ;
        RECT 255.850 0.855 257.510 1.400 ;
        RECT 258.610 0.855 260.270 1.400 ;
        RECT 261.370 0.855 263.030 1.400 ;
        RECT 264.130 0.855 265.790 1.400 ;
        RECT 266.890 0.855 268.550 1.400 ;
        RECT 269.650 0.855 271.310 1.400 ;
        RECT 272.410 0.855 274.070 1.400 ;
        RECT 275.170 0.855 276.830 1.400 ;
        RECT 277.930 0.855 279.590 1.400 ;
        RECT 280.690 0.855 282.350 1.400 ;
        RECT 283.450 0.855 285.110 1.400 ;
        RECT 286.210 0.855 287.870 1.400 ;
        RECT 288.970 0.855 290.630 1.400 ;
        RECT 291.730 0.855 293.390 1.400 ;
        RECT 294.490 0.855 296.150 1.400 ;
        RECT 297.250 0.855 298.910 1.400 ;
        RECT 300.010 0.855 301.670 1.400 ;
        RECT 302.770 0.855 304.430 1.400 ;
        RECT 305.530 0.855 307.190 1.400 ;
        RECT 308.290 0.855 309.950 1.400 ;
        RECT 311.050 0.855 312.710 1.400 ;
        RECT 313.810 0.855 315.470 1.400 ;
        RECT 316.570 0.855 318.230 1.400 ;
        RECT 319.330 0.855 343.990 1.400 ;
        RECT 345.090 0.855 369.750 1.400 ;
        RECT 370.850 0.855 372.510 1.400 ;
        RECT 373.610 0.855 375.270 1.400 ;
        RECT 376.370 0.855 378.030 1.400 ;
        RECT 379.130 0.855 380.790 1.400 ;
        RECT 381.890 0.855 383.550 1.400 ;
        RECT 384.650 0.855 386.310 1.400 ;
        RECT 387.410 0.855 389.070 1.400 ;
        RECT 390.170 0.855 391.830 1.400 ;
        RECT 392.930 0.855 394.590 1.400 ;
        RECT 395.690 0.855 397.350 1.400 ;
        RECT 398.450 0.855 400.110 1.400 ;
        RECT 401.210 0.855 402.870 1.400 ;
        RECT 403.970 0.855 405.630 1.400 ;
        RECT 406.730 0.855 408.390 1.400 ;
        RECT 409.490 0.855 411.150 1.400 ;
        RECT 412.250 0.855 413.910 1.400 ;
        RECT 415.010 0.855 416.670 1.400 ;
        RECT 417.770 0.855 419.430 1.400 ;
        RECT 420.530 0.855 422.190 1.400 ;
        RECT 423.290 0.855 424.950 1.400 ;
        RECT 426.050 0.855 427.710 1.400 ;
        RECT 428.810 0.855 430.470 1.400 ;
        RECT 431.570 0.855 433.230 1.400 ;
        RECT 434.330 0.855 435.990 1.400 ;
        RECT 437.090 0.855 438.750 1.400 ;
        RECT 439.850 0.855 441.510 1.400 ;
        RECT 442.610 0.855 444.270 1.400 ;
        RECT 445.370 0.855 447.030 1.400 ;
        RECT 448.130 0.855 449.790 1.400 ;
        RECT 450.890 0.855 452.550 1.400 ;
        RECT 453.650 0.855 455.310 1.400 ;
        RECT 456.410 0.855 458.070 1.400 ;
        RECT 459.170 0.855 460.830 1.400 ;
        RECT 461.930 0.855 463.590 1.400 ;
        RECT 464.690 0.855 466.350 1.400 ;
        RECT 467.450 0.855 469.110 1.400 ;
        RECT 470.210 0.855 471.870 1.400 ;
        RECT 472.970 0.855 474.630 1.400 ;
        RECT 475.730 0.855 477.390 1.400 ;
        RECT 478.490 0.855 480.150 1.400 ;
        RECT 481.250 0.855 482.910 1.400 ;
        RECT 484.010 0.855 485.670 1.400 ;
        RECT 486.770 0.855 488.430 1.400 ;
        RECT 489.530 0.855 514.190 1.400 ;
        RECT 515.290 0.855 539.950 1.400 ;
        RECT 541.050 0.855 542.710 1.400 ;
        RECT 543.810 0.855 545.470 1.400 ;
        RECT 546.570 0.855 548.230 1.400 ;
        RECT 549.330 0.855 550.990 1.400 ;
        RECT 552.090 0.855 553.750 1.400 ;
        RECT 554.850 0.855 556.510 1.400 ;
        RECT 557.610 0.855 559.270 1.400 ;
        RECT 560.370 0.855 562.030 1.400 ;
        RECT 563.130 0.855 564.790 1.400 ;
        RECT 565.890 0.855 567.550 1.400 ;
        RECT 568.650 0.855 570.310 1.400 ;
        RECT 571.410 0.855 573.070 1.400 ;
        RECT 574.170 0.855 575.830 1.400 ;
        RECT 576.930 0.855 578.590 1.400 ;
        RECT 579.690 0.855 581.350 1.400 ;
        RECT 582.450 0.855 584.110 1.400 ;
        RECT 585.210 0.855 586.870 1.400 ;
        RECT 587.970 0.855 589.630 1.400 ;
        RECT 590.730 0.855 592.390 1.400 ;
        RECT 593.490 0.855 595.150 1.400 ;
        RECT 596.250 0.855 597.910 1.400 ;
        RECT 599.010 0.855 600.670 1.400 ;
        RECT 601.770 0.855 603.430 1.400 ;
        RECT 604.530 0.855 606.190 1.400 ;
        RECT 607.290 0.855 608.950 1.400 ;
        RECT 610.050 0.855 611.710 1.400 ;
        RECT 612.810 0.855 614.470 1.400 ;
        RECT 615.570 0.855 617.230 1.400 ;
        RECT 618.330 0.855 619.990 1.400 ;
        RECT 621.090 0.855 622.750 1.400 ;
        RECT 623.850 0.855 625.510 1.400 ;
        RECT 626.610 0.855 628.270 1.400 ;
        RECT 629.370 0.855 631.030 1.400 ;
        RECT 632.130 0.855 633.790 1.400 ;
        RECT 634.890 0.855 636.550 1.400 ;
        RECT 637.650 0.855 639.310 1.400 ;
        RECT 640.410 0.855 642.070 1.400 ;
        RECT 643.170 0.855 644.830 1.400 ;
        RECT 645.930 0.855 647.590 1.400 ;
        RECT 648.690 0.855 650.350 1.400 ;
        RECT 651.450 0.855 653.110 1.400 ;
        RECT 654.210 0.855 655.870 1.400 ;
        RECT 656.970 0.855 658.630 1.400 ;
        RECT 659.730 0.855 684.390 1.400 ;
        RECT 685.490 0.855 710.150 1.400 ;
        RECT 711.250 0.855 712.910 1.400 ;
        RECT 714.010 0.855 715.670 1.400 ;
        RECT 716.770 0.855 718.430 1.400 ;
        RECT 719.530 0.855 721.190 1.400 ;
        RECT 722.290 0.855 723.950 1.400 ;
        RECT 725.050 0.855 726.710 1.400 ;
        RECT 727.810 0.855 729.470 1.400 ;
        RECT 730.570 0.855 732.230 1.400 ;
        RECT 733.330 0.855 734.990 1.400 ;
        RECT 736.090 0.855 737.750 1.400 ;
        RECT 738.850 0.855 740.510 1.400 ;
        RECT 741.610 0.855 743.270 1.400 ;
        RECT 744.370 0.855 746.030 1.400 ;
        RECT 747.130 0.855 748.790 1.400 ;
        RECT 749.890 0.855 751.550 1.400 ;
        RECT 752.650 0.855 754.310 1.400 ;
        RECT 755.410 0.855 757.070 1.400 ;
        RECT 758.170 0.855 759.830 1.400 ;
        RECT 760.930 0.855 762.590 1.400 ;
        RECT 763.690 0.855 765.350 1.400 ;
        RECT 766.450 0.855 768.110 1.400 ;
        RECT 769.210 0.855 770.870 1.400 ;
        RECT 771.970 0.855 773.630 1.400 ;
        RECT 774.730 0.855 776.390 1.400 ;
        RECT 777.490 0.855 779.150 1.400 ;
        RECT 780.250 0.855 781.910 1.400 ;
        RECT 783.010 0.855 784.670 1.400 ;
        RECT 785.770 0.855 787.430 1.400 ;
        RECT 788.530 0.855 790.190 1.400 ;
        RECT 791.290 0.855 792.950 1.400 ;
        RECT 794.050 0.855 795.710 1.400 ;
        RECT 796.810 0.855 798.470 1.400 ;
        RECT 799.570 0.855 801.230 1.400 ;
        RECT 802.330 0.855 803.990 1.400 ;
        RECT 805.090 0.855 806.750 1.400 ;
        RECT 807.850 0.855 809.510 1.400 ;
        RECT 810.610 0.855 812.270 1.400 ;
        RECT 813.370 0.855 815.030 1.400 ;
        RECT 816.130 0.855 817.790 1.400 ;
        RECT 818.890 0.855 820.550 1.400 ;
        RECT 821.650 0.855 823.310 1.400 ;
        RECT 824.410 0.855 826.070 1.400 ;
        RECT 827.170 0.855 828.830 1.400 ;
        RECT 829.930 0.855 854.590 1.400 ;
        RECT 855.690 0.855 880.350 1.400 ;
        RECT 881.450 0.855 883.110 1.400 ;
        RECT 884.210 0.855 885.870 1.400 ;
        RECT 886.970 0.855 888.630 1.400 ;
        RECT 889.730 0.855 891.390 1.400 ;
        RECT 892.490 0.855 894.150 1.400 ;
        RECT 895.250 0.855 896.910 1.400 ;
        RECT 898.010 0.855 899.670 1.400 ;
        RECT 900.770 0.855 902.430 1.400 ;
        RECT 903.530 0.855 905.190 1.400 ;
        RECT 906.290 0.855 907.950 1.400 ;
        RECT 909.050 0.855 910.710 1.400 ;
        RECT 911.810 0.855 913.470 1.400 ;
        RECT 914.570 0.855 916.230 1.400 ;
        RECT 917.330 0.855 918.990 1.400 ;
        RECT 920.090 0.855 921.750 1.400 ;
        RECT 922.850 0.855 924.510 1.400 ;
        RECT 925.610 0.855 927.270 1.400 ;
        RECT 928.370 0.855 930.030 1.400 ;
        RECT 931.130 0.855 932.790 1.400 ;
        RECT 933.890 0.855 935.550 1.400 ;
        RECT 936.650 0.855 938.310 1.400 ;
        RECT 939.410 0.855 941.070 1.400 ;
        RECT 942.170 0.855 943.830 1.400 ;
        RECT 944.930 0.855 946.590 1.400 ;
        RECT 947.690 0.855 949.350 1.400 ;
        RECT 950.450 0.855 952.110 1.400 ;
        RECT 953.210 0.855 954.870 1.400 ;
        RECT 955.970 0.855 957.630 1.400 ;
        RECT 958.730 0.855 960.390 1.400 ;
        RECT 961.490 0.855 963.150 1.400 ;
        RECT 964.250 0.855 965.910 1.400 ;
        RECT 967.010 0.855 968.670 1.400 ;
        RECT 969.770 0.855 971.430 1.400 ;
        RECT 972.530 0.855 974.190 1.400 ;
        RECT 975.290 0.855 976.950 1.400 ;
        RECT 978.050 0.855 979.710 1.400 ;
        RECT 980.810 0.855 982.470 1.400 ;
        RECT 983.570 0.855 985.230 1.400 ;
        RECT 986.330 0.855 987.990 1.400 ;
        RECT 989.090 0.855 990.750 1.400 ;
        RECT 991.850 0.855 993.510 1.400 ;
        RECT 994.610 0.855 996.270 1.400 ;
        RECT 997.370 0.855 999.030 1.400 ;
        RECT 1000.130 0.855 1024.790 1.400 ;
        RECT 1025.890 0.855 1050.550 1.400 ;
        RECT 1051.650 0.855 1053.310 1.400 ;
        RECT 1054.410 0.855 1056.070 1.400 ;
        RECT 1057.170 0.855 1058.830 1.400 ;
        RECT 1059.930 0.855 1061.590 1.400 ;
        RECT 1062.690 0.855 1064.350 1.400 ;
        RECT 1065.450 0.855 1067.110 1.400 ;
        RECT 1068.210 0.855 1069.870 1.400 ;
        RECT 1070.970 0.855 1072.630 1.400 ;
        RECT 1073.730 0.855 1075.390 1.400 ;
        RECT 1076.490 0.855 1078.150 1.400 ;
        RECT 1079.250 0.855 1080.910 1.400 ;
        RECT 1082.010 0.855 1083.670 1.400 ;
        RECT 1084.770 0.855 1086.430 1.400 ;
        RECT 1087.530 0.855 1089.190 1.400 ;
        RECT 1090.290 0.855 1091.950 1.400 ;
        RECT 1093.050 0.855 1094.710 1.400 ;
        RECT 1095.810 0.855 1097.470 1.400 ;
        RECT 1098.570 0.855 1100.230 1.400 ;
        RECT 1101.330 0.855 1102.990 1.400 ;
        RECT 1104.090 0.855 1105.750 1.400 ;
        RECT 1106.850 0.855 1108.510 1.400 ;
        RECT 1109.610 0.855 1111.270 1.400 ;
        RECT 1112.370 0.855 1114.030 1.400 ;
        RECT 1115.130 0.855 1116.790 1.400 ;
        RECT 1117.890 0.855 1119.550 1.400 ;
        RECT 1120.650 0.855 1122.310 1.400 ;
        RECT 1123.410 0.855 1125.070 1.400 ;
        RECT 1126.170 0.855 1127.830 1.400 ;
        RECT 1128.930 0.855 1130.590 1.400 ;
        RECT 1131.690 0.855 1133.350 1.400 ;
        RECT 1134.450 0.855 1136.110 1.400 ;
        RECT 1137.210 0.855 1138.870 1.400 ;
        RECT 1139.970 0.855 1141.630 1.400 ;
        RECT 1142.730 0.855 1144.390 1.400 ;
        RECT 1145.490 0.855 1147.150 1.400 ;
        RECT 1148.250 0.855 1149.910 1.400 ;
        RECT 1151.010 0.855 1152.670 1.400 ;
        RECT 1153.770 0.855 1155.430 1.400 ;
        RECT 1156.530 0.855 1158.190 1.400 ;
        RECT 1159.290 0.855 1160.950 1.400 ;
        RECT 1162.050 0.855 1163.710 1.400 ;
        RECT 1164.810 0.855 1166.470 1.400 ;
        RECT 1167.570 0.855 1169.230 1.400 ;
        RECT 1170.330 0.855 1194.990 1.400 ;
        RECT 1196.090 0.855 1220.750 1.400 ;
        RECT 1221.850 0.855 1223.510 1.400 ;
        RECT 1224.610 0.855 1226.270 1.400 ;
        RECT 1227.370 0.855 1229.030 1.400 ;
        RECT 1230.130 0.855 1231.790 1.400 ;
        RECT 1232.890 0.855 1234.550 1.400 ;
        RECT 1235.650 0.855 1237.310 1.400 ;
        RECT 1238.410 0.855 1240.070 1.400 ;
        RECT 1241.170 0.855 1242.830 1.400 ;
        RECT 1243.930 0.855 1245.590 1.400 ;
        RECT 1246.690 0.855 1248.350 1.400 ;
        RECT 1249.450 0.855 1251.110 1.400 ;
        RECT 1252.210 0.855 1253.870 1.400 ;
        RECT 1254.970 0.855 1256.630 1.400 ;
        RECT 1257.730 0.855 1259.390 1.400 ;
        RECT 1260.490 0.855 1262.150 1.400 ;
        RECT 1263.250 0.855 1264.910 1.400 ;
        RECT 1266.010 0.855 1267.670 1.400 ;
        RECT 1268.770 0.855 1270.430 1.400 ;
        RECT 1271.530 0.855 1273.190 1.400 ;
        RECT 1274.290 0.855 1275.950 1.400 ;
        RECT 1277.050 0.855 1278.710 1.400 ;
        RECT 1279.810 0.855 1281.470 1.400 ;
        RECT 1282.570 0.855 1284.230 1.400 ;
        RECT 1285.330 0.855 1286.990 1.400 ;
        RECT 1288.090 0.855 1289.750 1.400 ;
        RECT 1290.850 0.855 1292.510 1.400 ;
        RECT 1293.610 0.855 1295.270 1.400 ;
        RECT 1296.370 0.855 1298.030 1.400 ;
        RECT 1299.130 0.855 1300.790 1.400 ;
        RECT 1301.890 0.855 1303.550 1.400 ;
        RECT 1304.650 0.855 1306.310 1.400 ;
        RECT 1307.410 0.855 1309.070 1.400 ;
        RECT 1310.170 0.855 1311.830 1.400 ;
        RECT 1312.930 0.855 1314.590 1.400 ;
        RECT 1315.690 0.855 1317.350 1.400 ;
        RECT 1318.450 0.855 1320.110 1.400 ;
        RECT 1321.210 0.855 1322.870 1.400 ;
        RECT 1323.970 0.855 1325.630 1.400 ;
        RECT 1326.730 0.855 1328.390 1.400 ;
        RECT 1329.490 0.855 1331.150 1.400 ;
        RECT 1332.250 0.855 1333.910 1.400 ;
        RECT 1335.010 0.855 1336.670 1.400 ;
        RECT 1337.770 0.855 1339.430 1.400 ;
  END
END tt_mux
END LIBRARY

