VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_CktA_InstAmp
  CLASS BLOCK ;
  FOREIGN tt_um_CktA_InstAmp ;
  ORIGIN 0.000 0.000 ;
  SIZE 508.760 BY 225.760 ;
  PIN ui_in[0]
    ANTENNAGATEAREA 4.800000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 4.800000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ua[1]
    ANTENNAGATEAREA 10.848000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN ua[2]
    ANTENNAGATEAREA 10.848000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN ua[3]
    ANTENNADIFFAREA 66.385201 ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN uo_out[0]
    ANTENNAGATEAREA 639.591980 ;
    ANTENNADIFFAREA 1322.609009 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 639.591980 ;
    ANTENNADIFFAREA 1322.609009 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNAGATEAREA 639.591980 ;
    ANTENNADIFFAREA 1322.609009 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNAGATEAREA 639.591980 ;
    ANTENNADIFFAREA 1322.609009 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNAGATEAREA 639.591980 ;
    ANTENNADIFFAREA 1322.609009 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNAGATEAREA 639.591980 ;
    ANTENNADIFFAREA 1322.609009 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN ua[4]
    ANTENNAGATEAREA 10.848000 ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN uo_out[6]
    ANTENNAGATEAREA 639.591980 ;
    ANTENNADIFFAREA 1322.609009 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNAGATEAREA 639.591980 ;
    ANTENNADIFFAREA 1322.609009 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 639.591980 ;
    ANTENNADIFFAREA 1322.609009 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 639.591980 ;
    ANTENNADIFFAREA 1322.609009 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 639.591980 ;
    ANTENNADIFFAREA 1322.609009 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  PIN uio_out[3]
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN ua[5]
    ANTENNAGATEAREA 10.848000 ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN uio_out[4]
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uio_oe[0]
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN uio_oe[2]
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ena
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN ua[0]
    ANTENNAGATEAREA 10.848000 ;
    ANTENNADIFFAREA 66.385201 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN clk
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 74.280 186.040 147.010 209.775 ;
      LAYER pwell ;
        RECT 147.210 194.085 170.220 194.515 ;
        RECT 147.210 189.340 147.640 194.085 ;
        RECT 147.900 190.455 169.530 192.975 ;
        RECT 169.790 189.340 170.220 194.085 ;
        RECT 147.210 188.910 170.220 189.340 ;
        RECT 184.715 189.285 280.640 189.715 ;
        RECT 184.715 185.485 185.145 189.285 ;
        RECT 185.405 186.125 207.035 188.645 ;
        RECT 207.295 185.485 208.365 189.285 ;
        RECT 208.625 186.125 237.295 188.645 ;
        RECT 237.555 185.485 238.705 189.285 ;
        RECT 238.965 186.125 279.955 188.645 ;
        RECT 280.210 185.485 280.640 189.285 ;
        RECT 74.295 185.005 170.220 185.435 ;
        RECT 184.715 185.055 280.640 185.485 ;
        RECT 74.295 181.205 74.725 185.005 ;
        RECT 74.980 181.845 115.970 184.365 ;
        RECT 116.230 181.205 117.380 185.005 ;
        RECT 117.640 181.845 146.310 184.365 ;
        RECT 146.570 181.205 147.640 185.005 ;
        RECT 147.900 181.845 169.530 184.365 ;
        RECT 169.790 181.205 170.220 185.005 ;
        RECT 74.295 180.775 170.220 181.205 ;
        RECT 184.715 182.800 280.640 183.230 ;
        RECT 184.715 179.000 185.145 182.800 ;
        RECT 185.405 179.640 207.035 182.160 ;
        RECT 207.295 179.000 208.365 182.800 ;
        RECT 208.625 179.640 237.295 182.160 ;
        RECT 237.555 179.000 238.705 182.800 ;
        RECT 238.965 179.640 279.955 182.160 ;
        RECT 280.210 179.000 280.640 182.800 ;
        RECT 74.295 178.520 170.220 178.950 ;
        RECT 184.715 178.570 280.640 179.000 ;
        RECT 74.295 174.720 74.725 178.520 ;
        RECT 74.980 175.360 115.970 177.880 ;
        RECT 116.230 174.720 117.380 178.520 ;
        RECT 117.640 175.360 146.310 177.880 ;
        RECT 146.570 174.720 147.640 178.520 ;
        RECT 147.900 175.360 169.530 177.880 ;
        RECT 169.790 174.720 170.220 178.520 ;
        RECT 74.295 174.290 170.220 174.720 ;
        RECT 184.715 174.665 207.725 175.095 ;
        RECT 184.715 169.920 185.145 174.665 ;
        RECT 185.405 171.030 207.035 173.550 ;
        RECT 207.295 169.920 207.725 174.665 ;
        RECT 184.715 169.490 207.725 169.920 ;
      LAYER nwell ;
        RECT 207.925 154.230 280.655 177.965 ;
      LAYER pwell ;
        RECT 184.715 152.130 294.495 152.560 ;
        RECT 184.715 139.390 185.145 152.130 ;
        RECT 294.065 139.390 294.495 152.130 ;
        RECT 184.715 138.960 294.495 139.390 ;
        RECT 300.250 152.130 410.030 152.560 ;
        RECT 300.250 139.390 300.680 152.130 ;
        RECT 409.600 139.390 410.030 152.130 ;
        RECT 300.250 138.960 410.030 139.390 ;
        RECT 184.715 137.965 294.495 138.395 ;
        RECT 184.715 125.225 185.145 137.965 ;
        RECT 294.065 125.225 294.495 137.965 ;
        RECT 184.715 124.795 294.495 125.225 ;
        RECT 300.250 137.965 410.030 138.395 ;
        RECT 300.250 125.225 300.680 137.965 ;
        RECT 409.600 125.225 410.030 137.965 ;
        RECT 300.250 124.795 410.030 125.225 ;
        RECT 310.785 120.405 406.710 120.835 ;
        RECT 217.040 117.375 290.640 117.805 ;
      LAYER nwell ;
        RECT 184.620 112.445 213.610 115.395 ;
      LAYER pwell ;
        RECT 184.670 109.860 185.100 112.250 ;
        RECT 185.300 110.030 197.850 111.290 ;
        RECT 198.050 109.860 198.480 112.250 ;
      LAYER nwell ;
        RECT 199.700 110.055 213.610 112.445 ;
      LAYER pwell ;
        RECT 184.670 109.430 198.480 109.860 ;
        RECT 184.670 107.040 185.100 109.430 ;
        RECT 185.300 108.000 197.850 109.260 ;
        RECT 198.050 107.040 198.480 109.430 ;
      LAYER nwell ;
        RECT 184.620 99.945 198.530 106.845 ;
      LAYER pwell ;
        RECT 199.750 106.395 200.180 109.485 ;
        RECT 200.380 106.965 212.930 108.225 ;
        RECT 213.130 106.395 213.560 109.485 ;
        RECT 199.750 105.965 213.560 106.395 ;
        RECT 217.040 104.635 217.470 117.375 ;
        RECT 290.210 104.635 290.640 117.375 ;
        RECT 310.785 116.605 311.215 120.405 ;
        RECT 311.475 117.245 333.105 119.765 ;
        RECT 333.365 116.605 334.435 120.405 ;
        RECT 334.695 117.245 363.365 119.765 ;
        RECT 363.625 116.605 364.775 120.405 ;
        RECT 365.035 117.245 406.025 119.765 ;
        RECT 406.280 116.605 406.710 120.405 ;
        RECT 310.785 116.175 406.710 116.605 ;
        RECT 310.785 113.920 406.710 114.350 ;
        RECT 310.785 110.120 311.215 113.920 ;
        RECT 311.475 110.760 333.105 113.280 ;
        RECT 333.365 110.120 334.435 113.920 ;
        RECT 334.695 110.760 363.365 113.280 ;
        RECT 363.625 110.120 364.775 113.920 ;
        RECT 365.035 110.760 406.025 113.280 ;
        RECT 406.280 110.120 406.710 113.920 ;
        RECT 310.785 109.690 406.710 110.120 ;
        RECT 217.040 104.205 290.640 104.635 ;
        RECT 310.785 105.785 333.795 106.215 ;
        RECT 217.040 102.155 290.640 102.585 ;
        RECT 199.750 100.395 213.560 100.825 ;
        RECT 184.670 97.360 185.100 99.750 ;
        RECT 185.300 97.530 197.850 98.790 ;
        RECT 198.050 97.360 198.480 99.750 ;
        RECT 184.670 96.930 198.480 97.360 ;
        RECT 199.750 97.305 200.180 100.395 ;
        RECT 200.380 98.565 212.930 99.825 ;
        RECT 213.130 97.305 213.560 100.395 ;
        RECT 184.670 94.540 185.100 96.930 ;
        RECT 185.300 95.500 197.850 96.760 ;
        RECT 198.050 94.540 198.480 96.930 ;
      LAYER nwell ;
        RECT 199.700 94.345 213.610 96.735 ;
        RECT 184.620 91.395 213.610 94.345 ;
      LAYER pwell ;
        RECT 217.040 89.415 217.470 102.155 ;
        RECT 290.210 89.415 290.640 102.155 ;
        RECT 310.785 101.040 311.215 105.785 ;
        RECT 311.475 102.150 333.105 104.670 ;
        RECT 333.365 101.040 333.795 105.785 ;
        RECT 310.785 100.610 333.795 101.040 ;
        RECT 217.040 88.985 290.640 89.415 ;
      LAYER nwell ;
        RECT 333.995 85.350 406.725 109.085 ;
        RECT 443.895 108.905 505.570 119.205 ;
      LAYER pwell ;
        RECT 472.555 97.015 481.285 97.445 ;
        RECT 453.205 94.045 471.135 94.475 ;
        RECT 453.205 91.805 453.635 94.045 ;
        RECT 434.765 91.375 453.635 91.805 ;
        RECT 434.765 88.035 435.195 91.375 ;
        RECT 435.355 88.575 442.905 90.835 ;
        RECT 443.065 88.035 444.415 91.375 ;
        RECT 444.575 88.575 452.125 90.825 ;
        RECT 434.765 88.030 444.415 88.035 ;
        RECT 452.285 88.035 453.635 91.375 ;
        RECT 453.795 91.245 470.545 93.505 ;
        RECT 453.795 88.575 470.545 90.835 ;
        RECT 470.705 88.035 471.135 94.045 ;
        RECT 472.555 93.415 472.985 97.015 ;
        RECT 473.145 93.955 480.695 96.475 ;
        RECT 480.855 93.415 481.285 97.015 ;
      LAYER nwell ;
        RECT 486.930 94.610 495.840 108.905 ;
      LAYER pwell ;
        RECT 496.750 97.015 505.480 97.445 ;
        RECT 472.555 92.985 481.285 93.415 ;
        RECT 496.750 93.415 497.180 97.015 ;
        RECT 497.340 93.955 504.890 96.475 ;
        RECT 505.050 93.415 505.480 97.015 ;
        RECT 496.750 92.985 505.480 93.415 ;
        RECT 452.285 88.030 471.135 88.035 ;
        RECT 434.765 87.605 471.135 88.030 ;
        RECT 472.555 91.635 481.285 92.065 ;
        RECT 472.555 88.035 472.985 91.635 ;
        RECT 473.145 88.575 480.695 91.095 ;
        RECT 480.855 88.035 481.285 91.635 ;
        RECT 472.555 87.605 481.285 88.035 ;
        RECT 487.020 91.375 495.750 91.805 ;
        RECT 487.020 88.035 487.450 91.375 ;
        RECT 487.610 88.575 495.160 90.835 ;
        RECT 495.320 88.035 495.750 91.375 ;
        RECT 487.020 87.605 495.750 88.035 ;
        RECT 496.750 91.635 505.480 92.065 ;
        RECT 496.750 88.035 497.180 91.635 ;
        RECT 497.340 88.575 504.890 91.095 ;
        RECT 505.050 88.035 505.480 91.635 ;
        RECT 496.750 87.605 505.480 88.035 ;
        RECT 443.985 87.600 452.715 87.605 ;
        RECT 437.335 83.130 503.000 83.560 ;
        RECT 184.715 81.565 294.495 81.995 ;
        RECT 184.715 68.825 185.145 81.565 ;
        RECT 294.065 68.825 294.495 81.565 ;
        RECT 184.715 68.395 294.495 68.825 ;
        RECT 300.250 81.565 410.030 81.995 ;
        RECT 300.250 68.825 300.680 81.565 ;
        RECT 409.600 68.825 410.030 81.565 ;
        RECT 437.335 70.390 437.765 83.130 ;
        RECT 502.570 70.390 503.000 83.130 ;
        RECT 437.335 69.960 503.000 70.390 ;
        RECT 300.250 68.395 410.030 68.825 ;
        RECT 184.715 67.420 294.495 67.850 ;
        RECT 184.715 54.680 185.145 67.420 ;
        RECT 294.065 54.680 294.495 67.420 ;
        RECT 184.715 54.250 294.495 54.680 ;
        RECT 300.250 67.420 410.030 67.850 ;
        RECT 300.250 54.680 300.680 67.420 ;
        RECT 409.600 54.680 410.030 67.420 ;
        RECT 300.250 54.250 410.030 54.680 ;
        RECT 184.715 36.890 207.725 37.320 ;
        RECT 184.715 32.145 185.145 36.890 ;
        RECT 185.405 33.260 207.035 35.780 ;
        RECT 207.295 32.145 207.725 36.890 ;
        RECT 184.715 31.715 207.725 32.145 ;
      LAYER nwell ;
        RECT 207.925 28.845 280.655 52.580 ;
        RECT 330.580 28.845 403.310 52.580 ;
      LAYER pwell ;
        RECT 403.510 36.890 426.520 37.320 ;
        RECT 403.510 32.145 403.940 36.890 ;
        RECT 404.200 33.260 425.830 35.780 ;
        RECT 426.090 32.145 426.520 36.890 ;
        RECT 403.510 31.715 426.520 32.145 ;
        RECT 184.715 27.810 280.640 28.240 ;
        RECT 184.715 24.010 185.145 27.810 ;
        RECT 185.405 24.650 207.035 27.170 ;
        RECT 207.295 24.010 208.365 27.810 ;
        RECT 208.625 24.650 237.295 27.170 ;
        RECT 237.555 24.010 238.705 27.810 ;
        RECT 238.965 24.650 279.955 27.170 ;
        RECT 280.210 24.010 280.640 27.810 ;
        RECT 184.715 23.580 280.640 24.010 ;
        RECT 330.595 27.810 426.520 28.240 ;
        RECT 330.595 24.010 331.025 27.810 ;
        RECT 331.280 24.650 372.270 27.170 ;
        RECT 372.530 24.010 373.680 27.810 ;
        RECT 373.940 24.650 402.610 27.170 ;
        RECT 402.870 24.010 403.940 27.810 ;
        RECT 404.200 24.650 425.830 27.170 ;
        RECT 426.090 24.010 426.520 27.810 ;
        RECT 330.595 23.580 426.520 24.010 ;
        RECT 184.715 21.325 280.640 21.755 ;
        RECT 184.715 17.525 185.145 21.325 ;
        RECT 185.405 18.165 207.035 20.685 ;
        RECT 207.295 17.525 208.365 21.325 ;
        RECT 208.625 18.165 237.295 20.685 ;
        RECT 237.555 17.525 238.705 21.325 ;
        RECT 238.965 18.165 279.955 20.685 ;
        RECT 280.210 17.525 280.640 21.325 ;
        RECT 184.715 17.095 280.640 17.525 ;
        RECT 330.595 21.325 426.520 21.755 ;
        RECT 330.595 17.525 331.025 21.325 ;
        RECT 331.280 18.165 372.270 20.685 ;
        RECT 372.530 17.525 373.680 21.325 ;
        RECT 373.940 18.165 402.610 20.685 ;
        RECT 402.870 17.525 403.940 21.325 ;
        RECT 404.200 18.165 425.830 20.685 ;
        RECT 426.090 17.525 426.520 21.325 ;
        RECT 330.595 17.095 426.520 17.525 ;
      LAYER li1 ;
        RECT 74.400 209.365 116.550 209.655 ;
        RECT 74.400 198.815 74.690 209.365 ;
        RECT 79.010 208.775 80.260 209.105 ;
        RECT 80.770 208.775 82.020 209.105 ;
        RECT 82.530 208.775 83.780 209.105 ;
        RECT 84.290 208.775 85.540 209.105 ;
        RECT 86.050 208.775 87.300 209.105 ;
        RECT 87.810 208.775 89.060 209.105 ;
        RECT 89.570 208.775 90.820 209.105 ;
        RECT 91.330 208.775 92.580 209.105 ;
        RECT 93.090 208.775 94.340 209.105 ;
        RECT 94.850 208.775 96.100 209.105 ;
        RECT 96.610 208.775 97.860 209.105 ;
        RECT 98.370 208.775 99.620 209.105 ;
        RECT 100.130 208.775 101.380 209.105 ;
        RECT 101.890 208.775 103.140 209.105 ;
        RECT 103.650 208.775 104.900 209.105 ;
        RECT 105.410 208.775 106.660 209.105 ;
        RECT 107.170 208.775 108.420 209.105 ;
        RECT 108.930 208.775 110.180 209.105 ;
        RECT 110.690 208.775 111.940 209.105 ;
        RECT 112.450 208.775 113.700 209.105 ;
        RECT 75.150 199.575 75.320 208.605 ;
        RECT 76.030 199.575 76.200 208.605 ;
        RECT 76.910 199.575 77.080 208.605 ;
        RECT 77.790 199.575 77.960 208.605 ;
        RECT 78.670 199.575 78.840 208.605 ;
        RECT 79.550 199.575 79.720 208.605 ;
        RECT 80.430 199.575 80.600 208.605 ;
        RECT 81.310 199.575 81.480 208.605 ;
        RECT 82.190 199.575 82.360 208.605 ;
        RECT 83.070 199.575 83.240 208.605 ;
        RECT 83.950 199.575 84.120 208.605 ;
        RECT 84.830 199.575 85.000 208.605 ;
        RECT 85.710 199.575 85.880 208.605 ;
        RECT 86.590 199.575 86.760 208.605 ;
        RECT 87.470 199.575 87.640 208.605 ;
        RECT 88.350 199.575 88.520 208.605 ;
        RECT 89.230 199.575 89.400 208.605 ;
        RECT 90.110 199.575 90.280 208.605 ;
        RECT 90.990 199.575 91.160 208.605 ;
        RECT 91.870 199.575 92.040 208.605 ;
        RECT 92.750 199.575 92.920 208.605 ;
        RECT 93.630 199.575 93.800 208.605 ;
        RECT 94.510 199.575 94.680 208.605 ;
        RECT 95.390 199.575 95.560 208.605 ;
        RECT 96.270 199.575 96.440 208.605 ;
        RECT 97.150 199.575 97.320 208.605 ;
        RECT 98.030 199.575 98.200 208.605 ;
        RECT 98.910 199.575 99.080 208.605 ;
        RECT 99.790 199.575 99.960 208.605 ;
        RECT 100.670 199.575 100.840 208.605 ;
        RECT 101.550 199.575 101.720 208.605 ;
        RECT 102.430 199.575 102.600 208.605 ;
        RECT 103.310 199.575 103.480 208.605 ;
        RECT 104.190 199.575 104.360 208.605 ;
        RECT 105.070 199.575 105.240 208.605 ;
        RECT 105.950 199.575 106.120 208.605 ;
        RECT 106.830 199.575 107.000 208.605 ;
        RECT 107.710 199.575 107.880 208.605 ;
        RECT 108.590 199.575 108.760 208.605 ;
        RECT 109.470 199.575 109.640 208.605 ;
        RECT 110.350 199.575 110.520 208.605 ;
        RECT 111.230 199.575 111.400 208.605 ;
        RECT 112.110 199.575 112.280 208.605 ;
        RECT 112.990 199.575 113.160 208.605 ;
        RECT 113.870 199.575 114.040 208.605 ;
        RECT 114.750 199.575 114.920 208.605 ;
        RECT 115.630 199.575 115.800 208.605 ;
        RECT 75.490 199.075 76.740 199.405 ;
        RECT 77.250 199.075 78.500 199.405 ;
        RECT 114.210 199.075 115.460 199.405 ;
        RECT 116.260 198.815 116.550 209.365 ;
        RECT 74.400 198.525 116.550 198.815 ;
        RECT 117.060 209.365 146.890 209.655 ;
        RECT 117.060 198.815 117.350 209.365 ;
        RECT 121.670 208.775 122.920 209.105 ;
        RECT 123.430 208.775 124.680 209.105 ;
        RECT 125.190 208.775 126.440 209.105 ;
        RECT 126.950 208.775 128.200 209.105 ;
        RECT 128.710 208.775 129.960 209.105 ;
        RECT 130.470 208.775 131.720 209.105 ;
        RECT 132.230 208.775 133.480 209.105 ;
        RECT 133.990 208.775 135.240 209.105 ;
        RECT 135.750 208.775 137.000 209.105 ;
        RECT 137.510 208.775 138.760 209.105 ;
        RECT 139.270 208.775 140.520 209.105 ;
        RECT 141.030 208.775 142.280 209.105 ;
        RECT 117.810 199.575 117.980 208.605 ;
        RECT 118.690 199.575 118.860 208.605 ;
        RECT 119.570 199.575 119.740 208.605 ;
        RECT 120.450 199.575 120.620 208.605 ;
        RECT 121.330 199.575 121.500 208.605 ;
        RECT 122.210 199.575 122.380 208.605 ;
        RECT 123.090 199.575 123.260 208.605 ;
        RECT 123.970 199.575 124.140 208.605 ;
        RECT 124.850 199.575 125.020 208.605 ;
        RECT 125.730 199.575 125.900 208.605 ;
        RECT 126.610 199.575 126.780 208.605 ;
        RECT 127.490 199.575 127.660 208.605 ;
        RECT 128.370 199.575 128.540 208.605 ;
        RECT 129.250 199.575 129.420 208.605 ;
        RECT 130.130 199.575 130.300 208.605 ;
        RECT 131.010 199.575 131.180 208.605 ;
        RECT 131.890 199.575 132.060 208.605 ;
        RECT 132.770 199.575 132.940 208.605 ;
        RECT 133.650 199.575 133.820 208.605 ;
        RECT 134.530 199.575 134.700 208.605 ;
        RECT 135.410 199.575 135.580 208.605 ;
        RECT 136.290 199.575 136.460 208.605 ;
        RECT 137.170 199.575 137.340 208.605 ;
        RECT 138.050 199.575 138.220 208.605 ;
        RECT 138.930 199.575 139.100 208.605 ;
        RECT 139.810 199.575 139.980 208.605 ;
        RECT 140.690 199.575 140.860 208.605 ;
        RECT 141.570 199.575 141.740 208.605 ;
        RECT 142.450 199.575 142.620 208.605 ;
        RECT 143.330 199.575 143.500 208.605 ;
        RECT 144.210 199.575 144.380 208.605 ;
        RECT 145.090 199.575 145.260 208.605 ;
        RECT 145.970 199.575 146.140 208.605 ;
        RECT 118.150 199.075 119.400 199.405 ;
        RECT 119.910 199.075 121.160 199.405 ;
        RECT 142.790 199.075 144.040 199.405 ;
        RECT 144.550 199.075 145.800 199.405 ;
        RECT 146.600 198.815 146.890 209.365 ;
        RECT 117.060 198.525 146.890 198.815 ;
        RECT 74.400 197.000 116.550 197.290 ;
        RECT 74.400 186.450 74.690 197.000 ;
        RECT 75.490 196.410 76.740 196.740 ;
        RECT 77.250 196.410 78.500 196.740 ;
        RECT 114.210 196.410 115.460 196.740 ;
        RECT 75.150 187.210 75.320 196.240 ;
        RECT 76.030 187.210 76.200 196.240 ;
        RECT 76.910 187.210 77.080 196.240 ;
        RECT 77.790 187.210 77.960 196.240 ;
        RECT 78.670 187.210 78.840 196.240 ;
        RECT 79.550 187.210 79.720 196.240 ;
        RECT 80.430 187.210 80.600 196.240 ;
        RECT 81.310 187.210 81.480 196.240 ;
        RECT 82.190 187.210 82.360 196.240 ;
        RECT 83.070 187.210 83.240 196.240 ;
        RECT 83.950 187.210 84.120 196.240 ;
        RECT 84.830 187.210 85.000 196.240 ;
        RECT 85.710 187.210 85.880 196.240 ;
        RECT 86.590 187.210 86.760 196.240 ;
        RECT 87.470 187.210 87.640 196.240 ;
        RECT 88.350 187.210 88.520 196.240 ;
        RECT 89.230 187.210 89.400 196.240 ;
        RECT 90.110 187.210 90.280 196.240 ;
        RECT 90.990 187.210 91.160 196.240 ;
        RECT 91.870 187.210 92.040 196.240 ;
        RECT 92.750 187.210 92.920 196.240 ;
        RECT 93.630 187.210 93.800 196.240 ;
        RECT 94.510 187.210 94.680 196.240 ;
        RECT 95.390 187.210 95.560 196.240 ;
        RECT 96.270 187.210 96.440 196.240 ;
        RECT 97.150 187.210 97.320 196.240 ;
        RECT 98.030 187.210 98.200 196.240 ;
        RECT 98.910 187.210 99.080 196.240 ;
        RECT 99.790 187.210 99.960 196.240 ;
        RECT 100.670 187.210 100.840 196.240 ;
        RECT 101.550 187.210 101.720 196.240 ;
        RECT 102.430 187.210 102.600 196.240 ;
        RECT 103.310 187.210 103.480 196.240 ;
        RECT 104.190 187.210 104.360 196.240 ;
        RECT 105.070 187.210 105.240 196.240 ;
        RECT 105.950 187.210 106.120 196.240 ;
        RECT 106.830 187.210 107.000 196.240 ;
        RECT 107.710 187.210 107.880 196.240 ;
        RECT 108.590 187.210 108.760 196.240 ;
        RECT 109.470 187.210 109.640 196.240 ;
        RECT 110.350 187.210 110.520 196.240 ;
        RECT 111.230 187.210 111.400 196.240 ;
        RECT 112.110 187.210 112.280 196.240 ;
        RECT 112.990 187.210 113.160 196.240 ;
        RECT 113.870 187.210 114.040 196.240 ;
        RECT 114.750 187.210 114.920 196.240 ;
        RECT 115.630 187.210 115.800 196.240 ;
        RECT 79.010 186.710 80.260 187.040 ;
        RECT 80.770 186.710 82.020 187.040 ;
        RECT 82.530 186.710 83.780 187.040 ;
        RECT 84.290 186.710 85.540 187.040 ;
        RECT 86.050 186.710 87.300 187.040 ;
        RECT 87.810 186.710 89.060 187.040 ;
        RECT 89.570 186.710 90.820 187.040 ;
        RECT 91.330 186.710 92.580 187.040 ;
        RECT 93.090 186.710 94.340 187.040 ;
        RECT 94.850 186.710 96.100 187.040 ;
        RECT 96.610 186.710 97.860 187.040 ;
        RECT 98.370 186.710 99.620 187.040 ;
        RECT 100.130 186.710 101.380 187.040 ;
        RECT 101.890 186.710 103.140 187.040 ;
        RECT 103.650 186.710 104.900 187.040 ;
        RECT 105.410 186.710 106.660 187.040 ;
        RECT 107.170 186.710 108.420 187.040 ;
        RECT 108.930 186.710 110.180 187.040 ;
        RECT 110.690 186.710 111.940 187.040 ;
        RECT 112.450 186.710 113.700 187.040 ;
        RECT 116.260 186.450 116.550 197.000 ;
        RECT 74.400 186.160 116.550 186.450 ;
        RECT 117.060 197.000 146.890 197.290 ;
        RECT 117.060 186.450 117.350 197.000 ;
        RECT 118.150 196.410 119.400 196.740 ;
        RECT 119.910 196.410 121.160 196.740 ;
        RECT 121.670 196.410 122.920 196.740 ;
        RECT 130.470 196.410 131.720 196.740 ;
        RECT 132.230 196.410 133.480 196.740 ;
        RECT 141.030 196.410 142.280 196.740 ;
        RECT 142.790 196.410 144.040 196.740 ;
        RECT 144.550 196.410 145.800 196.740 ;
        RECT 117.810 187.210 117.980 196.240 ;
        RECT 118.690 187.210 118.860 196.240 ;
        RECT 119.570 187.210 119.740 196.240 ;
        RECT 120.450 187.210 120.620 196.240 ;
        RECT 121.330 187.210 121.500 196.240 ;
        RECT 122.210 187.210 122.380 196.240 ;
        RECT 123.090 187.210 123.260 196.240 ;
        RECT 123.970 187.210 124.140 196.240 ;
        RECT 124.850 187.210 125.020 196.240 ;
        RECT 125.730 187.210 125.900 196.240 ;
        RECT 126.610 187.210 126.780 196.240 ;
        RECT 127.490 187.210 127.660 196.240 ;
        RECT 128.370 187.210 128.540 196.240 ;
        RECT 129.250 187.210 129.420 196.240 ;
        RECT 130.130 187.210 130.300 196.240 ;
        RECT 131.010 187.210 131.180 196.240 ;
        RECT 131.890 187.210 132.060 196.240 ;
        RECT 132.770 187.210 132.940 196.240 ;
        RECT 133.650 187.210 133.820 196.240 ;
        RECT 134.530 187.210 134.700 196.240 ;
        RECT 135.410 187.210 135.580 196.240 ;
        RECT 136.290 187.210 136.460 196.240 ;
        RECT 137.170 187.210 137.340 196.240 ;
        RECT 138.050 187.210 138.220 196.240 ;
        RECT 138.930 187.210 139.100 196.240 ;
        RECT 139.810 187.210 139.980 196.240 ;
        RECT 140.690 187.210 140.860 196.240 ;
        RECT 141.570 187.210 141.740 196.240 ;
        RECT 142.450 187.210 142.620 196.240 ;
        RECT 143.330 187.210 143.500 196.240 ;
        RECT 144.210 187.210 144.380 196.240 ;
        RECT 145.090 187.210 145.260 196.240 ;
        RECT 145.970 187.210 146.140 196.240 ;
        RECT 123.430 186.710 124.680 187.040 ;
        RECT 125.190 186.710 126.440 187.040 ;
        RECT 126.950 186.710 128.200 187.040 ;
        RECT 128.710 186.710 129.960 187.040 ;
        RECT 133.990 186.710 135.240 187.040 ;
        RECT 135.750 186.710 137.000 187.040 ;
        RECT 137.510 186.710 138.760 187.040 ;
        RECT 139.270 186.710 140.520 187.040 ;
        RECT 146.600 186.450 146.890 197.000 ;
        RECT 147.340 194.215 170.090 194.385 ;
        RECT 147.340 189.210 147.510 194.215 ;
        RECT 148.410 193.015 149.660 193.345 ;
        RECT 150.170 193.015 151.420 193.345 ;
        RECT 153.690 193.015 154.940 193.345 ;
        RECT 157.210 193.015 158.460 193.345 ;
        RECT 160.730 193.015 161.980 193.345 ;
        RECT 164.250 193.015 165.500 193.345 ;
        RECT 166.010 193.015 167.260 193.345 ;
        RECT 167.770 193.015 169.020 193.345 ;
        RECT 148.070 190.585 148.240 192.845 ;
        RECT 148.950 190.585 149.120 192.845 ;
        RECT 149.830 190.585 150.000 192.845 ;
        RECT 150.710 190.585 150.880 192.845 ;
        RECT 151.590 190.585 151.760 192.845 ;
        RECT 152.470 190.585 152.640 192.845 ;
        RECT 153.350 190.585 153.520 192.845 ;
        RECT 154.230 190.585 154.400 192.845 ;
        RECT 155.110 190.585 155.280 192.845 ;
        RECT 155.990 190.585 156.160 192.845 ;
        RECT 156.870 190.585 157.040 192.845 ;
        RECT 157.750 190.585 157.920 192.845 ;
        RECT 158.630 190.585 158.800 192.845 ;
        RECT 159.510 190.585 159.680 192.845 ;
        RECT 160.390 190.585 160.560 192.845 ;
        RECT 161.270 190.585 161.440 192.845 ;
        RECT 162.150 190.585 162.320 192.845 ;
        RECT 163.030 190.585 163.200 192.845 ;
        RECT 163.910 190.585 164.080 192.845 ;
        RECT 164.790 190.585 164.960 192.845 ;
        RECT 165.670 190.585 165.840 192.845 ;
        RECT 166.550 190.585 166.720 192.845 ;
        RECT 167.430 190.585 167.600 192.845 ;
        RECT 168.310 190.585 168.480 192.845 ;
        RECT 169.190 190.585 169.360 192.845 ;
        RECT 148.410 190.085 149.660 190.415 ;
        RECT 150.170 190.085 151.420 190.415 ;
        RECT 151.930 190.085 153.180 190.415 ;
        RECT 155.450 190.085 156.700 190.415 ;
        RECT 158.970 190.085 160.220 190.415 ;
        RECT 162.490 190.085 163.740 190.415 ;
        RECT 166.010 190.085 167.260 190.415 ;
        RECT 167.770 190.085 169.020 190.415 ;
        RECT 169.920 189.210 170.090 194.215 ;
        RECT 147.340 189.040 170.090 189.210 ;
        RECT 184.845 189.415 207.595 189.585 ;
        RECT 117.060 186.160 146.890 186.450 ;
        RECT 184.845 185.355 185.015 189.415 ;
        RECT 192.955 188.685 194.205 189.015 ;
        RECT 194.715 188.685 195.965 189.015 ;
        RECT 196.475 188.685 197.725 189.015 ;
        RECT 198.235 188.685 199.485 189.015 ;
        RECT 185.575 186.255 185.745 188.515 ;
        RECT 186.455 186.255 186.625 188.515 ;
        RECT 187.335 186.255 187.505 188.515 ;
        RECT 188.215 186.255 188.385 188.515 ;
        RECT 189.095 186.255 189.265 188.515 ;
        RECT 189.975 186.255 190.145 188.515 ;
        RECT 190.855 186.255 191.025 188.515 ;
        RECT 191.735 186.255 191.905 188.515 ;
        RECT 192.615 186.255 192.785 188.515 ;
        RECT 193.495 186.255 193.665 188.515 ;
        RECT 194.375 186.255 194.545 188.515 ;
        RECT 195.255 186.255 195.425 188.515 ;
        RECT 196.135 186.255 196.305 188.515 ;
        RECT 197.015 186.255 197.185 188.515 ;
        RECT 197.895 186.255 198.065 188.515 ;
        RECT 198.775 186.255 198.945 188.515 ;
        RECT 199.655 186.255 199.825 188.515 ;
        RECT 200.535 186.255 200.705 188.515 ;
        RECT 201.415 186.255 201.585 188.515 ;
        RECT 202.295 186.255 202.465 188.515 ;
        RECT 203.175 186.255 203.345 188.515 ;
        RECT 204.055 186.255 204.225 188.515 ;
        RECT 204.935 186.255 205.105 188.515 ;
        RECT 205.815 186.255 205.985 188.515 ;
        RECT 206.695 186.255 206.865 188.515 ;
        RECT 185.915 185.755 187.165 186.085 ;
        RECT 187.675 185.755 188.925 186.085 ;
        RECT 189.435 185.755 190.685 186.085 ;
        RECT 191.195 185.755 192.445 186.085 ;
        RECT 199.995 185.755 201.245 186.085 ;
        RECT 201.755 185.755 203.005 186.085 ;
        RECT 203.515 185.755 204.765 186.085 ;
        RECT 205.275 185.755 206.525 186.085 ;
        RECT 207.425 185.355 207.595 189.415 ;
        RECT 74.425 185.135 116.530 185.305 ;
        RECT 74.425 181.075 74.595 185.135 ;
        RECT 75.490 184.405 76.740 184.735 ;
        RECT 77.250 184.405 78.500 184.735 ;
        RECT 114.210 184.405 115.460 184.735 ;
        RECT 75.150 181.975 75.320 184.235 ;
        RECT 76.030 181.975 76.200 184.235 ;
        RECT 76.910 181.975 77.080 184.235 ;
        RECT 77.790 181.975 77.960 184.235 ;
        RECT 78.670 181.975 78.840 184.235 ;
        RECT 79.550 181.975 79.720 184.235 ;
        RECT 80.430 181.975 80.600 184.235 ;
        RECT 81.310 181.975 81.480 184.235 ;
        RECT 82.190 181.975 82.360 184.235 ;
        RECT 83.070 181.975 83.240 184.235 ;
        RECT 83.950 181.975 84.120 184.235 ;
        RECT 84.830 181.975 85.000 184.235 ;
        RECT 85.710 181.975 85.880 184.235 ;
        RECT 86.590 181.975 86.760 184.235 ;
        RECT 87.470 181.975 87.640 184.235 ;
        RECT 88.350 181.975 88.520 184.235 ;
        RECT 89.230 181.975 89.400 184.235 ;
        RECT 90.110 181.975 90.280 184.235 ;
        RECT 90.990 181.975 91.160 184.235 ;
        RECT 91.870 181.975 92.040 184.235 ;
        RECT 92.750 181.975 92.920 184.235 ;
        RECT 93.630 181.975 93.800 184.235 ;
        RECT 94.510 181.975 94.680 184.235 ;
        RECT 95.390 181.975 95.560 184.235 ;
        RECT 96.270 181.975 96.440 184.235 ;
        RECT 97.150 181.975 97.320 184.235 ;
        RECT 98.030 181.975 98.200 184.235 ;
        RECT 98.910 181.975 99.080 184.235 ;
        RECT 99.790 181.975 99.960 184.235 ;
        RECT 100.670 181.975 100.840 184.235 ;
        RECT 101.550 181.975 101.720 184.235 ;
        RECT 102.430 181.975 102.600 184.235 ;
        RECT 103.310 181.975 103.480 184.235 ;
        RECT 104.190 181.975 104.360 184.235 ;
        RECT 105.070 181.975 105.240 184.235 ;
        RECT 105.950 181.975 106.120 184.235 ;
        RECT 106.830 181.975 107.000 184.235 ;
        RECT 107.710 181.975 107.880 184.235 ;
        RECT 108.590 181.975 108.760 184.235 ;
        RECT 109.470 181.975 109.640 184.235 ;
        RECT 110.350 181.975 110.520 184.235 ;
        RECT 111.230 181.975 111.400 184.235 ;
        RECT 112.110 181.975 112.280 184.235 ;
        RECT 112.990 181.975 113.160 184.235 ;
        RECT 113.870 181.975 114.040 184.235 ;
        RECT 114.750 181.975 114.920 184.235 ;
        RECT 115.630 181.975 115.800 184.235 ;
        RECT 79.010 181.475 80.260 181.805 ;
        RECT 80.770 181.475 82.020 181.805 ;
        RECT 82.530 181.475 83.780 181.805 ;
        RECT 84.290 181.475 85.540 181.805 ;
        RECT 86.050 181.475 87.300 181.805 ;
        RECT 87.810 181.475 89.060 181.805 ;
        RECT 89.570 181.475 90.820 181.805 ;
        RECT 91.330 181.475 92.580 181.805 ;
        RECT 93.090 181.475 94.340 181.805 ;
        RECT 94.850 181.475 96.100 181.805 ;
        RECT 96.610 181.475 97.860 181.805 ;
        RECT 98.370 181.475 99.620 181.805 ;
        RECT 100.130 181.475 101.380 181.805 ;
        RECT 101.890 181.475 103.140 181.805 ;
        RECT 103.650 181.475 104.900 181.805 ;
        RECT 105.410 181.475 106.660 181.805 ;
        RECT 107.170 181.475 108.420 181.805 ;
        RECT 108.930 181.475 110.180 181.805 ;
        RECT 110.690 181.475 111.940 181.805 ;
        RECT 112.450 181.475 113.700 181.805 ;
        RECT 116.360 181.075 116.530 185.135 ;
        RECT 74.425 180.905 116.530 181.075 ;
        RECT 117.080 185.135 146.870 185.305 ;
        RECT 117.080 181.075 117.250 185.135 ;
        RECT 118.150 184.405 119.400 184.735 ;
        RECT 119.910 184.405 121.160 184.735 ;
        RECT 121.670 184.405 122.920 184.735 ;
        RECT 130.470 184.405 131.720 184.735 ;
        RECT 132.230 184.405 133.480 184.735 ;
        RECT 141.030 184.405 142.280 184.735 ;
        RECT 142.790 184.405 144.040 184.735 ;
        RECT 144.550 184.405 145.800 184.735 ;
        RECT 117.810 181.975 117.980 184.235 ;
        RECT 118.690 181.975 118.860 184.235 ;
        RECT 119.570 181.975 119.740 184.235 ;
        RECT 120.450 181.975 120.620 184.235 ;
        RECT 121.330 181.975 121.500 184.235 ;
        RECT 122.210 181.975 122.380 184.235 ;
        RECT 123.090 181.975 123.260 184.235 ;
        RECT 123.970 181.975 124.140 184.235 ;
        RECT 124.850 181.975 125.020 184.235 ;
        RECT 125.730 181.975 125.900 184.235 ;
        RECT 126.610 181.975 126.780 184.235 ;
        RECT 127.490 181.975 127.660 184.235 ;
        RECT 128.370 181.975 128.540 184.235 ;
        RECT 129.250 181.975 129.420 184.235 ;
        RECT 130.130 181.975 130.300 184.235 ;
        RECT 131.010 181.975 131.180 184.235 ;
        RECT 131.890 181.975 132.060 184.235 ;
        RECT 132.770 181.975 132.940 184.235 ;
        RECT 133.650 181.975 133.820 184.235 ;
        RECT 134.530 181.975 134.700 184.235 ;
        RECT 135.410 181.975 135.580 184.235 ;
        RECT 136.290 181.975 136.460 184.235 ;
        RECT 137.170 181.975 137.340 184.235 ;
        RECT 138.050 181.975 138.220 184.235 ;
        RECT 138.930 181.975 139.100 184.235 ;
        RECT 139.810 181.975 139.980 184.235 ;
        RECT 140.690 181.975 140.860 184.235 ;
        RECT 141.570 181.975 141.740 184.235 ;
        RECT 142.450 181.975 142.620 184.235 ;
        RECT 143.330 181.975 143.500 184.235 ;
        RECT 144.210 181.975 144.380 184.235 ;
        RECT 145.090 181.975 145.260 184.235 ;
        RECT 145.970 181.975 146.140 184.235 ;
        RECT 123.430 181.475 124.680 181.805 ;
        RECT 125.190 181.475 126.440 181.805 ;
        RECT 126.950 181.475 128.200 181.805 ;
        RECT 128.710 181.475 129.960 181.805 ;
        RECT 133.990 181.475 135.240 181.805 ;
        RECT 135.750 181.475 137.000 181.805 ;
        RECT 137.510 181.475 138.760 181.805 ;
        RECT 139.270 181.475 140.520 181.805 ;
        RECT 146.700 181.075 146.870 185.135 ;
        RECT 117.080 180.905 146.870 181.075 ;
        RECT 147.340 185.135 170.090 185.305 ;
        RECT 184.845 185.185 207.595 185.355 ;
        RECT 208.065 189.415 237.855 189.585 ;
        RECT 208.065 185.355 208.235 189.415 ;
        RECT 221.455 188.685 222.705 189.015 ;
        RECT 223.215 188.685 224.465 189.015 ;
        RECT 208.795 186.255 208.965 188.515 ;
        RECT 209.675 186.255 209.845 188.515 ;
        RECT 210.555 186.255 210.725 188.515 ;
        RECT 211.435 186.255 211.605 188.515 ;
        RECT 212.315 186.255 212.485 188.515 ;
        RECT 213.195 186.255 213.365 188.515 ;
        RECT 214.075 186.255 214.245 188.515 ;
        RECT 214.955 186.255 215.125 188.515 ;
        RECT 215.835 186.255 216.005 188.515 ;
        RECT 216.715 186.255 216.885 188.515 ;
        RECT 217.595 186.255 217.765 188.515 ;
        RECT 218.475 186.255 218.645 188.515 ;
        RECT 219.355 186.255 219.525 188.515 ;
        RECT 220.235 186.255 220.405 188.515 ;
        RECT 221.115 186.255 221.285 188.515 ;
        RECT 221.995 186.255 222.165 188.515 ;
        RECT 222.875 186.255 223.045 188.515 ;
        RECT 223.755 186.255 223.925 188.515 ;
        RECT 224.635 186.255 224.805 188.515 ;
        RECT 225.515 186.255 225.685 188.515 ;
        RECT 226.395 186.255 226.565 188.515 ;
        RECT 227.275 186.255 227.445 188.515 ;
        RECT 228.155 186.255 228.325 188.515 ;
        RECT 229.035 186.255 229.205 188.515 ;
        RECT 229.915 186.255 230.085 188.515 ;
        RECT 230.795 186.255 230.965 188.515 ;
        RECT 231.675 186.255 231.845 188.515 ;
        RECT 232.555 186.255 232.725 188.515 ;
        RECT 233.435 186.255 233.605 188.515 ;
        RECT 234.315 186.255 234.485 188.515 ;
        RECT 235.195 186.255 235.365 188.515 ;
        RECT 236.075 186.255 236.245 188.515 ;
        RECT 236.955 186.255 237.125 188.515 ;
        RECT 209.135 185.755 210.385 186.085 ;
        RECT 210.895 185.755 212.145 186.085 ;
        RECT 212.655 185.755 213.905 186.085 ;
        RECT 214.415 185.755 215.665 186.085 ;
        RECT 216.175 185.755 217.425 186.085 ;
        RECT 217.935 185.755 219.185 186.085 ;
        RECT 219.695 185.755 220.945 186.085 ;
        RECT 224.975 185.755 226.225 186.085 ;
        RECT 226.735 185.755 227.985 186.085 ;
        RECT 228.495 185.755 229.745 186.085 ;
        RECT 230.255 185.755 231.505 186.085 ;
        RECT 232.015 185.755 233.265 186.085 ;
        RECT 233.775 185.755 235.025 186.085 ;
        RECT 235.535 185.755 236.785 186.085 ;
        RECT 237.685 185.355 237.855 189.415 ;
        RECT 208.065 185.185 237.855 185.355 ;
        RECT 238.405 189.415 280.510 189.585 ;
        RECT 238.405 185.355 238.575 189.415 ;
        RECT 239.135 186.255 239.305 188.515 ;
        RECT 240.015 186.255 240.185 188.515 ;
        RECT 240.895 186.255 241.065 188.515 ;
        RECT 241.775 186.255 241.945 188.515 ;
        RECT 242.655 186.255 242.825 188.515 ;
        RECT 243.535 186.255 243.705 188.515 ;
        RECT 244.415 186.255 244.585 188.515 ;
        RECT 245.295 186.255 245.465 188.515 ;
        RECT 246.175 186.255 246.345 188.515 ;
        RECT 247.055 186.255 247.225 188.515 ;
        RECT 247.935 186.255 248.105 188.515 ;
        RECT 248.815 186.255 248.985 188.515 ;
        RECT 249.695 186.255 249.865 188.515 ;
        RECT 250.575 186.255 250.745 188.515 ;
        RECT 251.455 186.255 251.625 188.515 ;
        RECT 252.335 186.255 252.505 188.515 ;
        RECT 253.215 186.255 253.385 188.515 ;
        RECT 254.095 186.255 254.265 188.515 ;
        RECT 254.975 186.255 255.145 188.515 ;
        RECT 255.855 186.255 256.025 188.515 ;
        RECT 256.735 186.255 256.905 188.515 ;
        RECT 257.615 186.255 257.785 188.515 ;
        RECT 258.495 186.255 258.665 188.515 ;
        RECT 259.375 186.255 259.545 188.515 ;
        RECT 260.255 186.255 260.425 188.515 ;
        RECT 261.135 186.255 261.305 188.515 ;
        RECT 262.015 186.255 262.185 188.515 ;
        RECT 262.895 186.255 263.065 188.515 ;
        RECT 263.775 186.255 263.945 188.515 ;
        RECT 264.655 186.255 264.825 188.515 ;
        RECT 265.535 186.255 265.705 188.515 ;
        RECT 266.415 186.255 266.585 188.515 ;
        RECT 267.295 186.255 267.465 188.515 ;
        RECT 268.175 186.255 268.345 188.515 ;
        RECT 269.055 186.255 269.225 188.515 ;
        RECT 269.935 186.255 270.105 188.515 ;
        RECT 270.815 186.255 270.985 188.515 ;
        RECT 271.695 186.255 271.865 188.515 ;
        RECT 272.575 186.255 272.745 188.515 ;
        RECT 273.455 186.255 273.625 188.515 ;
        RECT 274.335 186.255 274.505 188.515 ;
        RECT 275.215 186.255 275.385 188.515 ;
        RECT 276.095 186.255 276.265 188.515 ;
        RECT 276.975 186.255 277.145 188.515 ;
        RECT 277.855 186.255 278.025 188.515 ;
        RECT 278.735 186.255 278.905 188.515 ;
        RECT 279.615 186.255 279.785 188.515 ;
        RECT 239.475 185.755 240.725 186.085 ;
        RECT 241.235 185.755 242.485 186.085 ;
        RECT 242.995 185.755 244.245 186.085 ;
        RECT 244.755 185.755 246.005 186.085 ;
        RECT 246.515 185.755 247.765 186.085 ;
        RECT 248.275 185.755 249.525 186.085 ;
        RECT 250.035 185.755 251.285 186.085 ;
        RECT 251.795 185.755 253.045 186.085 ;
        RECT 253.555 185.755 254.805 186.085 ;
        RECT 255.315 185.755 256.565 186.085 ;
        RECT 257.075 185.755 258.325 186.085 ;
        RECT 258.835 185.755 260.085 186.085 ;
        RECT 260.595 185.755 261.845 186.085 ;
        RECT 262.355 185.755 263.605 186.085 ;
        RECT 264.115 185.755 265.365 186.085 ;
        RECT 265.875 185.755 267.125 186.085 ;
        RECT 267.635 185.755 268.885 186.085 ;
        RECT 269.395 185.755 270.645 186.085 ;
        RECT 271.155 185.755 272.405 186.085 ;
        RECT 272.915 185.755 274.165 186.085 ;
        RECT 274.675 185.755 275.925 186.085 ;
        RECT 276.435 185.755 277.685 186.085 ;
        RECT 278.195 185.755 279.445 186.085 ;
        RECT 280.340 185.355 280.510 189.415 ;
        RECT 238.405 185.185 280.510 185.355 ;
        RECT 147.340 181.075 147.510 185.135 ;
        RECT 148.410 184.405 149.660 184.735 ;
        RECT 150.170 184.405 151.420 184.735 ;
        RECT 151.930 184.405 153.180 184.735 ;
        RECT 153.690 184.405 154.940 184.735 ;
        RECT 162.490 184.405 163.740 184.735 ;
        RECT 164.250 184.405 165.500 184.735 ;
        RECT 166.010 184.405 167.260 184.735 ;
        RECT 167.770 184.405 169.020 184.735 ;
        RECT 148.070 181.975 148.240 184.235 ;
        RECT 148.950 181.975 149.120 184.235 ;
        RECT 149.830 181.975 150.000 184.235 ;
        RECT 150.710 181.975 150.880 184.235 ;
        RECT 151.590 181.975 151.760 184.235 ;
        RECT 152.470 181.975 152.640 184.235 ;
        RECT 153.350 181.975 153.520 184.235 ;
        RECT 154.230 181.975 154.400 184.235 ;
        RECT 155.110 181.975 155.280 184.235 ;
        RECT 155.990 181.975 156.160 184.235 ;
        RECT 156.870 181.975 157.040 184.235 ;
        RECT 157.750 181.975 157.920 184.235 ;
        RECT 158.630 181.975 158.800 184.235 ;
        RECT 159.510 181.975 159.680 184.235 ;
        RECT 160.390 181.975 160.560 184.235 ;
        RECT 161.270 181.975 161.440 184.235 ;
        RECT 162.150 181.975 162.320 184.235 ;
        RECT 163.030 181.975 163.200 184.235 ;
        RECT 163.910 181.975 164.080 184.235 ;
        RECT 164.790 181.975 164.960 184.235 ;
        RECT 165.670 181.975 165.840 184.235 ;
        RECT 166.550 181.975 166.720 184.235 ;
        RECT 167.430 181.975 167.600 184.235 ;
        RECT 168.310 181.975 168.480 184.235 ;
        RECT 169.190 181.975 169.360 184.235 ;
        RECT 155.450 181.475 156.700 181.805 ;
        RECT 157.210 181.475 158.460 181.805 ;
        RECT 158.970 181.475 160.220 181.805 ;
        RECT 160.730 181.475 161.980 181.805 ;
        RECT 169.920 181.075 170.090 185.135 ;
        RECT 147.340 180.905 170.090 181.075 ;
        RECT 184.845 182.930 207.595 183.100 ;
        RECT 184.845 178.870 185.015 182.930 ;
        RECT 192.955 182.200 194.205 182.530 ;
        RECT 194.715 182.200 195.965 182.530 ;
        RECT 196.475 182.200 197.725 182.530 ;
        RECT 198.235 182.200 199.485 182.530 ;
        RECT 185.575 179.770 185.745 182.030 ;
        RECT 186.455 179.770 186.625 182.030 ;
        RECT 187.335 179.770 187.505 182.030 ;
        RECT 188.215 179.770 188.385 182.030 ;
        RECT 189.095 179.770 189.265 182.030 ;
        RECT 189.975 179.770 190.145 182.030 ;
        RECT 190.855 179.770 191.025 182.030 ;
        RECT 191.735 179.770 191.905 182.030 ;
        RECT 192.615 179.770 192.785 182.030 ;
        RECT 193.495 179.770 193.665 182.030 ;
        RECT 194.375 179.770 194.545 182.030 ;
        RECT 195.255 179.770 195.425 182.030 ;
        RECT 196.135 179.770 196.305 182.030 ;
        RECT 197.015 179.770 197.185 182.030 ;
        RECT 197.895 179.770 198.065 182.030 ;
        RECT 198.775 179.770 198.945 182.030 ;
        RECT 199.655 179.770 199.825 182.030 ;
        RECT 200.535 179.770 200.705 182.030 ;
        RECT 201.415 179.770 201.585 182.030 ;
        RECT 202.295 179.770 202.465 182.030 ;
        RECT 203.175 179.770 203.345 182.030 ;
        RECT 204.055 179.770 204.225 182.030 ;
        RECT 204.935 179.770 205.105 182.030 ;
        RECT 205.815 179.770 205.985 182.030 ;
        RECT 206.695 179.770 206.865 182.030 ;
        RECT 185.915 179.270 187.165 179.600 ;
        RECT 187.675 179.270 188.925 179.600 ;
        RECT 189.435 179.270 190.685 179.600 ;
        RECT 191.195 179.270 192.445 179.600 ;
        RECT 199.995 179.270 201.245 179.600 ;
        RECT 201.755 179.270 203.005 179.600 ;
        RECT 203.515 179.270 204.765 179.600 ;
        RECT 205.275 179.270 206.525 179.600 ;
        RECT 207.425 178.870 207.595 182.930 ;
        RECT 74.425 178.650 116.530 178.820 ;
        RECT 74.425 174.590 74.595 178.650 ;
        RECT 75.490 177.920 76.740 178.250 ;
        RECT 77.250 177.920 78.500 178.250 ;
        RECT 79.010 177.920 80.260 178.250 ;
        RECT 80.770 177.920 82.020 178.250 ;
        RECT 82.530 177.920 83.780 178.250 ;
        RECT 84.290 177.920 85.540 178.250 ;
        RECT 86.050 177.920 87.300 178.250 ;
        RECT 87.810 177.920 89.060 178.250 ;
        RECT 89.570 177.920 90.820 178.250 ;
        RECT 91.330 177.920 92.580 178.250 ;
        RECT 93.090 177.920 94.340 178.250 ;
        RECT 94.850 177.920 96.100 178.250 ;
        RECT 96.610 177.920 97.860 178.250 ;
        RECT 98.370 177.920 99.620 178.250 ;
        RECT 100.130 177.920 101.380 178.250 ;
        RECT 101.890 177.920 103.140 178.250 ;
        RECT 103.650 177.920 104.900 178.250 ;
        RECT 105.410 177.920 106.660 178.250 ;
        RECT 107.170 177.920 108.420 178.250 ;
        RECT 108.930 177.920 110.180 178.250 ;
        RECT 110.690 177.920 111.940 178.250 ;
        RECT 112.450 177.920 113.700 178.250 ;
        RECT 114.210 177.920 115.460 178.250 ;
        RECT 75.150 175.490 75.320 177.750 ;
        RECT 76.030 175.490 76.200 177.750 ;
        RECT 76.910 175.490 77.080 177.750 ;
        RECT 77.790 175.490 77.960 177.750 ;
        RECT 78.670 175.490 78.840 177.750 ;
        RECT 79.550 175.490 79.720 177.750 ;
        RECT 80.430 175.490 80.600 177.750 ;
        RECT 81.310 175.490 81.480 177.750 ;
        RECT 82.190 175.490 82.360 177.750 ;
        RECT 83.070 175.490 83.240 177.750 ;
        RECT 83.950 175.490 84.120 177.750 ;
        RECT 84.830 175.490 85.000 177.750 ;
        RECT 85.710 175.490 85.880 177.750 ;
        RECT 86.590 175.490 86.760 177.750 ;
        RECT 87.470 175.490 87.640 177.750 ;
        RECT 88.350 175.490 88.520 177.750 ;
        RECT 89.230 175.490 89.400 177.750 ;
        RECT 90.110 175.490 90.280 177.750 ;
        RECT 90.990 175.490 91.160 177.750 ;
        RECT 91.870 175.490 92.040 177.750 ;
        RECT 92.750 175.490 92.920 177.750 ;
        RECT 93.630 175.490 93.800 177.750 ;
        RECT 94.510 175.490 94.680 177.750 ;
        RECT 95.390 175.490 95.560 177.750 ;
        RECT 96.270 175.490 96.440 177.750 ;
        RECT 97.150 175.490 97.320 177.750 ;
        RECT 98.030 175.490 98.200 177.750 ;
        RECT 98.910 175.490 99.080 177.750 ;
        RECT 99.790 175.490 99.960 177.750 ;
        RECT 100.670 175.490 100.840 177.750 ;
        RECT 101.550 175.490 101.720 177.750 ;
        RECT 102.430 175.490 102.600 177.750 ;
        RECT 103.310 175.490 103.480 177.750 ;
        RECT 104.190 175.490 104.360 177.750 ;
        RECT 105.070 175.490 105.240 177.750 ;
        RECT 105.950 175.490 106.120 177.750 ;
        RECT 106.830 175.490 107.000 177.750 ;
        RECT 107.710 175.490 107.880 177.750 ;
        RECT 108.590 175.490 108.760 177.750 ;
        RECT 109.470 175.490 109.640 177.750 ;
        RECT 110.350 175.490 110.520 177.750 ;
        RECT 111.230 175.490 111.400 177.750 ;
        RECT 112.110 175.490 112.280 177.750 ;
        RECT 112.990 175.490 113.160 177.750 ;
        RECT 113.870 175.490 114.040 177.750 ;
        RECT 114.750 175.490 114.920 177.750 ;
        RECT 115.630 175.490 115.800 177.750 ;
        RECT 116.360 174.590 116.530 178.650 ;
        RECT 74.425 174.420 116.530 174.590 ;
        RECT 117.080 178.650 146.870 178.820 ;
        RECT 117.080 174.590 117.250 178.650 ;
        RECT 118.150 177.920 119.400 178.250 ;
        RECT 119.910 177.920 121.160 178.250 ;
        RECT 121.670 177.920 122.920 178.250 ;
        RECT 123.430 177.920 124.680 178.250 ;
        RECT 125.190 177.920 126.440 178.250 ;
        RECT 126.950 177.920 128.200 178.250 ;
        RECT 128.710 177.920 129.960 178.250 ;
        RECT 133.990 177.920 135.240 178.250 ;
        RECT 135.750 177.920 137.000 178.250 ;
        RECT 137.510 177.920 138.760 178.250 ;
        RECT 139.270 177.920 140.520 178.250 ;
        RECT 141.030 177.920 142.280 178.250 ;
        RECT 142.790 177.920 144.040 178.250 ;
        RECT 144.550 177.920 145.800 178.250 ;
        RECT 117.810 175.490 117.980 177.750 ;
        RECT 118.690 175.490 118.860 177.750 ;
        RECT 119.570 175.490 119.740 177.750 ;
        RECT 120.450 175.490 120.620 177.750 ;
        RECT 121.330 175.490 121.500 177.750 ;
        RECT 122.210 175.490 122.380 177.750 ;
        RECT 123.090 175.490 123.260 177.750 ;
        RECT 123.970 175.490 124.140 177.750 ;
        RECT 124.850 175.490 125.020 177.750 ;
        RECT 125.730 175.490 125.900 177.750 ;
        RECT 126.610 175.490 126.780 177.750 ;
        RECT 127.490 175.490 127.660 177.750 ;
        RECT 128.370 175.490 128.540 177.750 ;
        RECT 129.250 175.490 129.420 177.750 ;
        RECT 130.130 175.490 130.300 177.750 ;
        RECT 131.010 175.490 131.180 177.750 ;
        RECT 131.890 175.490 132.060 177.750 ;
        RECT 132.770 175.490 132.940 177.750 ;
        RECT 133.650 175.490 133.820 177.750 ;
        RECT 134.530 175.490 134.700 177.750 ;
        RECT 135.410 175.490 135.580 177.750 ;
        RECT 136.290 175.490 136.460 177.750 ;
        RECT 137.170 175.490 137.340 177.750 ;
        RECT 138.050 175.490 138.220 177.750 ;
        RECT 138.930 175.490 139.100 177.750 ;
        RECT 139.810 175.490 139.980 177.750 ;
        RECT 140.690 175.490 140.860 177.750 ;
        RECT 141.570 175.490 141.740 177.750 ;
        RECT 142.450 175.490 142.620 177.750 ;
        RECT 143.330 175.490 143.500 177.750 ;
        RECT 144.210 175.490 144.380 177.750 ;
        RECT 145.090 175.490 145.260 177.750 ;
        RECT 145.970 175.490 146.140 177.750 ;
        RECT 130.470 174.990 131.720 175.320 ;
        RECT 132.230 174.990 133.480 175.320 ;
        RECT 146.700 174.590 146.870 178.650 ;
        RECT 117.080 174.420 146.870 174.590 ;
        RECT 147.340 178.650 170.090 178.820 ;
        RECT 184.845 178.700 207.595 178.870 ;
        RECT 208.065 182.930 237.855 183.100 ;
        RECT 208.065 178.870 208.235 182.930 ;
        RECT 214.415 182.200 215.665 182.530 ;
        RECT 216.175 182.200 217.425 182.530 ;
        RECT 217.935 182.200 219.185 182.530 ;
        RECT 219.695 182.200 220.945 182.530 ;
        RECT 224.975 182.200 226.225 182.530 ;
        RECT 226.735 182.200 227.985 182.530 ;
        RECT 228.495 182.200 229.745 182.530 ;
        RECT 230.255 182.200 231.505 182.530 ;
        RECT 208.795 179.770 208.965 182.030 ;
        RECT 209.675 179.770 209.845 182.030 ;
        RECT 210.555 179.770 210.725 182.030 ;
        RECT 211.435 179.770 211.605 182.030 ;
        RECT 212.315 179.770 212.485 182.030 ;
        RECT 213.195 179.770 213.365 182.030 ;
        RECT 214.075 179.770 214.245 182.030 ;
        RECT 214.955 179.770 215.125 182.030 ;
        RECT 215.835 179.770 216.005 182.030 ;
        RECT 216.715 179.770 216.885 182.030 ;
        RECT 217.595 179.770 217.765 182.030 ;
        RECT 218.475 179.770 218.645 182.030 ;
        RECT 219.355 179.770 219.525 182.030 ;
        RECT 220.235 179.770 220.405 182.030 ;
        RECT 221.115 179.770 221.285 182.030 ;
        RECT 221.995 179.770 222.165 182.030 ;
        RECT 222.875 179.770 223.045 182.030 ;
        RECT 223.755 179.770 223.925 182.030 ;
        RECT 224.635 179.770 224.805 182.030 ;
        RECT 225.515 179.770 225.685 182.030 ;
        RECT 226.395 179.770 226.565 182.030 ;
        RECT 227.275 179.770 227.445 182.030 ;
        RECT 228.155 179.770 228.325 182.030 ;
        RECT 229.035 179.770 229.205 182.030 ;
        RECT 229.915 179.770 230.085 182.030 ;
        RECT 230.795 179.770 230.965 182.030 ;
        RECT 231.675 179.770 231.845 182.030 ;
        RECT 232.555 179.770 232.725 182.030 ;
        RECT 233.435 179.770 233.605 182.030 ;
        RECT 234.315 179.770 234.485 182.030 ;
        RECT 235.195 179.770 235.365 182.030 ;
        RECT 236.075 179.770 236.245 182.030 ;
        RECT 236.955 179.770 237.125 182.030 ;
        RECT 209.135 179.270 210.385 179.600 ;
        RECT 210.895 179.270 212.145 179.600 ;
        RECT 212.655 179.270 213.905 179.600 ;
        RECT 221.455 179.270 222.705 179.600 ;
        RECT 223.215 179.270 224.465 179.600 ;
        RECT 232.015 179.270 233.265 179.600 ;
        RECT 233.775 179.270 235.025 179.600 ;
        RECT 235.535 179.270 236.785 179.600 ;
        RECT 237.685 178.870 237.855 182.930 ;
        RECT 208.065 178.700 237.855 178.870 ;
        RECT 238.405 182.930 280.510 183.100 ;
        RECT 238.405 178.870 238.575 182.930 ;
        RECT 241.235 182.200 242.485 182.530 ;
        RECT 242.995 182.200 244.245 182.530 ;
        RECT 244.755 182.200 246.005 182.530 ;
        RECT 246.515 182.200 247.765 182.530 ;
        RECT 248.275 182.200 249.525 182.530 ;
        RECT 250.035 182.200 251.285 182.530 ;
        RECT 251.795 182.200 253.045 182.530 ;
        RECT 253.555 182.200 254.805 182.530 ;
        RECT 255.315 182.200 256.565 182.530 ;
        RECT 257.075 182.200 258.325 182.530 ;
        RECT 258.835 182.200 260.085 182.530 ;
        RECT 260.595 182.200 261.845 182.530 ;
        RECT 262.355 182.200 263.605 182.530 ;
        RECT 264.115 182.200 265.365 182.530 ;
        RECT 265.875 182.200 267.125 182.530 ;
        RECT 267.635 182.200 268.885 182.530 ;
        RECT 269.395 182.200 270.645 182.530 ;
        RECT 271.155 182.200 272.405 182.530 ;
        RECT 272.915 182.200 274.165 182.530 ;
        RECT 274.675 182.200 275.925 182.530 ;
        RECT 239.135 179.770 239.305 182.030 ;
        RECT 240.015 179.770 240.185 182.030 ;
        RECT 240.895 179.770 241.065 182.030 ;
        RECT 241.775 179.770 241.945 182.030 ;
        RECT 242.655 179.770 242.825 182.030 ;
        RECT 243.535 179.770 243.705 182.030 ;
        RECT 244.415 179.770 244.585 182.030 ;
        RECT 245.295 179.770 245.465 182.030 ;
        RECT 246.175 179.770 246.345 182.030 ;
        RECT 247.055 179.770 247.225 182.030 ;
        RECT 247.935 179.770 248.105 182.030 ;
        RECT 248.815 179.770 248.985 182.030 ;
        RECT 249.695 179.770 249.865 182.030 ;
        RECT 250.575 179.770 250.745 182.030 ;
        RECT 251.455 179.770 251.625 182.030 ;
        RECT 252.335 179.770 252.505 182.030 ;
        RECT 253.215 179.770 253.385 182.030 ;
        RECT 254.095 179.770 254.265 182.030 ;
        RECT 254.975 179.770 255.145 182.030 ;
        RECT 255.855 179.770 256.025 182.030 ;
        RECT 256.735 179.770 256.905 182.030 ;
        RECT 257.615 179.770 257.785 182.030 ;
        RECT 258.495 179.770 258.665 182.030 ;
        RECT 259.375 179.770 259.545 182.030 ;
        RECT 260.255 179.770 260.425 182.030 ;
        RECT 261.135 179.770 261.305 182.030 ;
        RECT 262.015 179.770 262.185 182.030 ;
        RECT 262.895 179.770 263.065 182.030 ;
        RECT 263.775 179.770 263.945 182.030 ;
        RECT 264.655 179.770 264.825 182.030 ;
        RECT 265.535 179.770 265.705 182.030 ;
        RECT 266.415 179.770 266.585 182.030 ;
        RECT 267.295 179.770 267.465 182.030 ;
        RECT 268.175 179.770 268.345 182.030 ;
        RECT 269.055 179.770 269.225 182.030 ;
        RECT 269.935 179.770 270.105 182.030 ;
        RECT 270.815 179.770 270.985 182.030 ;
        RECT 271.695 179.770 271.865 182.030 ;
        RECT 272.575 179.770 272.745 182.030 ;
        RECT 273.455 179.770 273.625 182.030 ;
        RECT 274.335 179.770 274.505 182.030 ;
        RECT 275.215 179.770 275.385 182.030 ;
        RECT 276.095 179.770 276.265 182.030 ;
        RECT 276.975 179.770 277.145 182.030 ;
        RECT 277.855 179.770 278.025 182.030 ;
        RECT 278.735 179.770 278.905 182.030 ;
        RECT 279.615 179.770 279.785 182.030 ;
        RECT 239.475 179.270 240.725 179.600 ;
        RECT 276.435 179.270 277.685 179.600 ;
        RECT 278.195 179.270 279.445 179.600 ;
        RECT 280.340 178.870 280.510 182.930 ;
        RECT 238.405 178.700 280.510 178.870 ;
        RECT 147.340 174.590 147.510 178.650 ;
        RECT 148.410 177.920 149.660 178.250 ;
        RECT 150.170 177.920 151.420 178.250 ;
        RECT 151.930 177.920 153.180 178.250 ;
        RECT 153.690 177.920 154.940 178.250 ;
        RECT 162.490 177.920 163.740 178.250 ;
        RECT 164.250 177.920 165.500 178.250 ;
        RECT 166.010 177.920 167.260 178.250 ;
        RECT 167.770 177.920 169.020 178.250 ;
        RECT 148.070 175.490 148.240 177.750 ;
        RECT 148.950 175.490 149.120 177.750 ;
        RECT 149.830 175.490 150.000 177.750 ;
        RECT 150.710 175.490 150.880 177.750 ;
        RECT 151.590 175.490 151.760 177.750 ;
        RECT 152.470 175.490 152.640 177.750 ;
        RECT 153.350 175.490 153.520 177.750 ;
        RECT 154.230 175.490 154.400 177.750 ;
        RECT 155.110 175.490 155.280 177.750 ;
        RECT 155.990 175.490 156.160 177.750 ;
        RECT 156.870 175.490 157.040 177.750 ;
        RECT 157.750 175.490 157.920 177.750 ;
        RECT 158.630 175.490 158.800 177.750 ;
        RECT 159.510 175.490 159.680 177.750 ;
        RECT 160.390 175.490 160.560 177.750 ;
        RECT 161.270 175.490 161.440 177.750 ;
        RECT 162.150 175.490 162.320 177.750 ;
        RECT 163.030 175.490 163.200 177.750 ;
        RECT 163.910 175.490 164.080 177.750 ;
        RECT 164.790 175.490 164.960 177.750 ;
        RECT 165.670 175.490 165.840 177.750 ;
        RECT 166.550 175.490 166.720 177.750 ;
        RECT 167.430 175.490 167.600 177.750 ;
        RECT 168.310 175.490 168.480 177.750 ;
        RECT 169.190 175.490 169.360 177.750 ;
        RECT 155.450 174.990 156.700 175.320 ;
        RECT 157.210 174.990 158.460 175.320 ;
        RECT 158.970 174.990 160.220 175.320 ;
        RECT 160.730 174.990 161.980 175.320 ;
        RECT 169.920 174.590 170.090 178.650 ;
        RECT 208.045 177.555 237.875 177.845 ;
        RECT 147.340 174.420 170.090 174.590 ;
        RECT 184.845 174.795 207.595 174.965 ;
        RECT 184.845 169.790 185.015 174.795 ;
        RECT 185.915 173.590 187.165 173.920 ;
        RECT 187.675 173.590 188.925 173.920 ;
        RECT 191.195 173.590 192.445 173.920 ;
        RECT 194.715 173.590 195.965 173.920 ;
        RECT 198.235 173.590 199.485 173.920 ;
        RECT 201.755 173.590 203.005 173.920 ;
        RECT 203.515 173.590 204.765 173.920 ;
        RECT 205.275 173.590 206.525 173.920 ;
        RECT 185.575 171.160 185.745 173.420 ;
        RECT 186.455 171.160 186.625 173.420 ;
        RECT 187.335 171.160 187.505 173.420 ;
        RECT 188.215 171.160 188.385 173.420 ;
        RECT 189.095 171.160 189.265 173.420 ;
        RECT 189.975 171.160 190.145 173.420 ;
        RECT 190.855 171.160 191.025 173.420 ;
        RECT 191.735 171.160 191.905 173.420 ;
        RECT 192.615 171.160 192.785 173.420 ;
        RECT 193.495 171.160 193.665 173.420 ;
        RECT 194.375 171.160 194.545 173.420 ;
        RECT 195.255 171.160 195.425 173.420 ;
        RECT 196.135 171.160 196.305 173.420 ;
        RECT 197.015 171.160 197.185 173.420 ;
        RECT 197.895 171.160 198.065 173.420 ;
        RECT 198.775 171.160 198.945 173.420 ;
        RECT 199.655 171.160 199.825 173.420 ;
        RECT 200.535 171.160 200.705 173.420 ;
        RECT 201.415 171.160 201.585 173.420 ;
        RECT 202.295 171.160 202.465 173.420 ;
        RECT 203.175 171.160 203.345 173.420 ;
        RECT 204.055 171.160 204.225 173.420 ;
        RECT 204.935 171.160 205.105 173.420 ;
        RECT 205.815 171.160 205.985 173.420 ;
        RECT 206.695 171.160 206.865 173.420 ;
        RECT 185.915 170.660 187.165 170.990 ;
        RECT 187.675 170.660 188.925 170.990 ;
        RECT 189.435 170.660 190.685 170.990 ;
        RECT 192.955 170.660 194.205 170.990 ;
        RECT 196.475 170.660 197.725 170.990 ;
        RECT 199.995 170.660 201.245 170.990 ;
        RECT 203.515 170.660 204.765 170.990 ;
        RECT 205.275 170.660 206.525 170.990 ;
        RECT 207.425 169.790 207.595 174.795 ;
        RECT 184.845 169.620 207.595 169.790 ;
        RECT 208.045 167.005 208.335 177.555 ;
        RECT 214.415 176.965 215.665 177.295 ;
        RECT 216.175 176.965 217.425 177.295 ;
        RECT 217.935 176.965 219.185 177.295 ;
        RECT 219.695 176.965 220.945 177.295 ;
        RECT 224.975 176.965 226.225 177.295 ;
        RECT 226.735 176.965 227.985 177.295 ;
        RECT 228.495 176.965 229.745 177.295 ;
        RECT 230.255 176.965 231.505 177.295 ;
        RECT 208.795 167.765 208.965 176.795 ;
        RECT 209.675 167.765 209.845 176.795 ;
        RECT 210.555 167.765 210.725 176.795 ;
        RECT 211.435 167.765 211.605 176.795 ;
        RECT 212.315 167.765 212.485 176.795 ;
        RECT 213.195 167.765 213.365 176.795 ;
        RECT 214.075 167.765 214.245 176.795 ;
        RECT 214.955 167.765 215.125 176.795 ;
        RECT 215.835 167.765 216.005 176.795 ;
        RECT 216.715 167.765 216.885 176.795 ;
        RECT 217.595 167.765 217.765 176.795 ;
        RECT 218.475 167.765 218.645 176.795 ;
        RECT 219.355 167.765 219.525 176.795 ;
        RECT 220.235 167.765 220.405 176.795 ;
        RECT 221.115 167.765 221.285 176.795 ;
        RECT 221.995 167.765 222.165 176.795 ;
        RECT 222.875 167.765 223.045 176.795 ;
        RECT 223.755 167.765 223.925 176.795 ;
        RECT 224.635 167.765 224.805 176.795 ;
        RECT 225.515 167.765 225.685 176.795 ;
        RECT 226.395 167.765 226.565 176.795 ;
        RECT 227.275 167.765 227.445 176.795 ;
        RECT 228.155 167.765 228.325 176.795 ;
        RECT 229.035 167.765 229.205 176.795 ;
        RECT 229.915 167.765 230.085 176.795 ;
        RECT 230.795 167.765 230.965 176.795 ;
        RECT 231.675 167.765 231.845 176.795 ;
        RECT 232.555 167.765 232.725 176.795 ;
        RECT 233.435 167.765 233.605 176.795 ;
        RECT 234.315 167.765 234.485 176.795 ;
        RECT 235.195 167.765 235.365 176.795 ;
        RECT 236.075 167.765 236.245 176.795 ;
        RECT 236.955 167.765 237.125 176.795 ;
        RECT 209.135 167.265 210.385 167.595 ;
        RECT 210.895 167.265 212.145 167.595 ;
        RECT 212.655 167.265 213.905 167.595 ;
        RECT 221.455 167.265 222.705 167.595 ;
        RECT 223.215 167.265 224.465 167.595 ;
        RECT 232.015 167.265 233.265 167.595 ;
        RECT 233.775 167.265 235.025 167.595 ;
        RECT 235.535 167.265 236.785 167.595 ;
        RECT 237.585 167.005 237.875 177.555 ;
        RECT 208.045 166.715 237.875 167.005 ;
        RECT 238.385 177.555 280.535 177.845 ;
        RECT 238.385 167.005 238.675 177.555 ;
        RECT 241.235 176.965 242.485 177.295 ;
        RECT 242.995 176.965 244.245 177.295 ;
        RECT 244.755 176.965 246.005 177.295 ;
        RECT 246.515 176.965 247.765 177.295 ;
        RECT 248.275 176.965 249.525 177.295 ;
        RECT 250.035 176.965 251.285 177.295 ;
        RECT 251.795 176.965 253.045 177.295 ;
        RECT 253.555 176.965 254.805 177.295 ;
        RECT 255.315 176.965 256.565 177.295 ;
        RECT 257.075 176.965 258.325 177.295 ;
        RECT 258.835 176.965 260.085 177.295 ;
        RECT 260.595 176.965 261.845 177.295 ;
        RECT 262.355 176.965 263.605 177.295 ;
        RECT 264.115 176.965 265.365 177.295 ;
        RECT 265.875 176.965 267.125 177.295 ;
        RECT 267.635 176.965 268.885 177.295 ;
        RECT 269.395 176.965 270.645 177.295 ;
        RECT 271.155 176.965 272.405 177.295 ;
        RECT 272.915 176.965 274.165 177.295 ;
        RECT 274.675 176.965 275.925 177.295 ;
        RECT 239.135 167.765 239.305 176.795 ;
        RECT 240.015 167.765 240.185 176.795 ;
        RECT 240.895 167.765 241.065 176.795 ;
        RECT 241.775 167.765 241.945 176.795 ;
        RECT 242.655 167.765 242.825 176.795 ;
        RECT 243.535 167.765 243.705 176.795 ;
        RECT 244.415 167.765 244.585 176.795 ;
        RECT 245.295 167.765 245.465 176.795 ;
        RECT 246.175 167.765 246.345 176.795 ;
        RECT 247.055 167.765 247.225 176.795 ;
        RECT 247.935 167.765 248.105 176.795 ;
        RECT 248.815 167.765 248.985 176.795 ;
        RECT 249.695 167.765 249.865 176.795 ;
        RECT 250.575 167.765 250.745 176.795 ;
        RECT 251.455 167.765 251.625 176.795 ;
        RECT 252.335 167.765 252.505 176.795 ;
        RECT 253.215 167.765 253.385 176.795 ;
        RECT 254.095 167.765 254.265 176.795 ;
        RECT 254.975 167.765 255.145 176.795 ;
        RECT 255.855 167.765 256.025 176.795 ;
        RECT 256.735 167.765 256.905 176.795 ;
        RECT 257.615 167.765 257.785 176.795 ;
        RECT 258.495 167.765 258.665 176.795 ;
        RECT 259.375 167.765 259.545 176.795 ;
        RECT 260.255 167.765 260.425 176.795 ;
        RECT 261.135 167.765 261.305 176.795 ;
        RECT 262.015 167.765 262.185 176.795 ;
        RECT 262.895 167.765 263.065 176.795 ;
        RECT 263.775 167.765 263.945 176.795 ;
        RECT 264.655 167.765 264.825 176.795 ;
        RECT 265.535 167.765 265.705 176.795 ;
        RECT 266.415 167.765 266.585 176.795 ;
        RECT 267.295 167.765 267.465 176.795 ;
        RECT 268.175 167.765 268.345 176.795 ;
        RECT 269.055 167.765 269.225 176.795 ;
        RECT 269.935 167.765 270.105 176.795 ;
        RECT 270.815 167.765 270.985 176.795 ;
        RECT 271.695 167.765 271.865 176.795 ;
        RECT 272.575 167.765 272.745 176.795 ;
        RECT 273.455 167.765 273.625 176.795 ;
        RECT 274.335 167.765 274.505 176.795 ;
        RECT 275.215 167.765 275.385 176.795 ;
        RECT 276.095 167.765 276.265 176.795 ;
        RECT 276.975 167.765 277.145 176.795 ;
        RECT 277.855 167.765 278.025 176.795 ;
        RECT 278.735 167.765 278.905 176.795 ;
        RECT 279.615 167.765 279.785 176.795 ;
        RECT 239.475 167.265 240.725 167.595 ;
        RECT 276.435 167.265 277.685 167.595 ;
        RECT 278.195 167.265 279.445 167.595 ;
        RECT 280.245 167.005 280.535 177.555 ;
        RECT 238.385 166.715 280.535 167.005 ;
        RECT 208.045 165.190 237.875 165.480 ;
        RECT 208.045 154.640 208.335 165.190 ;
        RECT 209.135 164.600 210.385 164.930 ;
        RECT 210.895 164.600 212.145 164.930 ;
        RECT 233.775 164.600 235.025 164.930 ;
        RECT 235.535 164.600 236.785 164.930 ;
        RECT 208.795 155.400 208.965 164.430 ;
        RECT 209.675 155.400 209.845 164.430 ;
        RECT 210.555 155.400 210.725 164.430 ;
        RECT 211.435 155.400 211.605 164.430 ;
        RECT 212.315 155.400 212.485 164.430 ;
        RECT 213.195 155.400 213.365 164.430 ;
        RECT 214.075 155.400 214.245 164.430 ;
        RECT 214.955 155.400 215.125 164.430 ;
        RECT 215.835 155.400 216.005 164.430 ;
        RECT 216.715 155.400 216.885 164.430 ;
        RECT 217.595 155.400 217.765 164.430 ;
        RECT 218.475 155.400 218.645 164.430 ;
        RECT 219.355 155.400 219.525 164.430 ;
        RECT 220.235 155.400 220.405 164.430 ;
        RECT 221.115 155.400 221.285 164.430 ;
        RECT 221.995 155.400 222.165 164.430 ;
        RECT 222.875 155.400 223.045 164.430 ;
        RECT 223.755 155.400 223.925 164.430 ;
        RECT 224.635 155.400 224.805 164.430 ;
        RECT 225.515 155.400 225.685 164.430 ;
        RECT 226.395 155.400 226.565 164.430 ;
        RECT 227.275 155.400 227.445 164.430 ;
        RECT 228.155 155.400 228.325 164.430 ;
        RECT 229.035 155.400 229.205 164.430 ;
        RECT 229.915 155.400 230.085 164.430 ;
        RECT 230.795 155.400 230.965 164.430 ;
        RECT 231.675 155.400 231.845 164.430 ;
        RECT 232.555 155.400 232.725 164.430 ;
        RECT 233.435 155.400 233.605 164.430 ;
        RECT 234.315 155.400 234.485 164.430 ;
        RECT 235.195 155.400 235.365 164.430 ;
        RECT 236.075 155.400 236.245 164.430 ;
        RECT 236.955 155.400 237.125 164.430 ;
        RECT 212.655 154.900 213.905 155.230 ;
        RECT 214.415 154.900 215.665 155.230 ;
        RECT 216.175 154.900 217.425 155.230 ;
        RECT 217.935 154.900 219.185 155.230 ;
        RECT 219.695 154.900 220.945 155.230 ;
        RECT 221.455 154.900 222.705 155.230 ;
        RECT 223.215 154.900 224.465 155.230 ;
        RECT 224.975 154.900 226.225 155.230 ;
        RECT 226.735 154.900 227.985 155.230 ;
        RECT 228.495 154.900 229.745 155.230 ;
        RECT 230.255 154.900 231.505 155.230 ;
        RECT 232.015 154.900 233.265 155.230 ;
        RECT 237.585 154.640 237.875 165.190 ;
        RECT 208.045 154.350 237.875 154.640 ;
        RECT 238.385 165.190 280.535 165.480 ;
        RECT 238.385 154.640 238.675 165.190 ;
        RECT 239.475 164.600 240.725 164.930 ;
        RECT 276.435 164.600 277.685 164.930 ;
        RECT 278.195 164.600 279.445 164.930 ;
        RECT 239.135 155.400 239.305 164.430 ;
        RECT 240.015 155.400 240.185 164.430 ;
        RECT 240.895 155.400 241.065 164.430 ;
        RECT 241.775 155.400 241.945 164.430 ;
        RECT 242.655 155.400 242.825 164.430 ;
        RECT 243.535 155.400 243.705 164.430 ;
        RECT 244.415 155.400 244.585 164.430 ;
        RECT 245.295 155.400 245.465 164.430 ;
        RECT 246.175 155.400 246.345 164.430 ;
        RECT 247.055 155.400 247.225 164.430 ;
        RECT 247.935 155.400 248.105 164.430 ;
        RECT 248.815 155.400 248.985 164.430 ;
        RECT 249.695 155.400 249.865 164.430 ;
        RECT 250.575 155.400 250.745 164.430 ;
        RECT 251.455 155.400 251.625 164.430 ;
        RECT 252.335 155.400 252.505 164.430 ;
        RECT 253.215 155.400 253.385 164.430 ;
        RECT 254.095 155.400 254.265 164.430 ;
        RECT 254.975 155.400 255.145 164.430 ;
        RECT 255.855 155.400 256.025 164.430 ;
        RECT 256.735 155.400 256.905 164.430 ;
        RECT 257.615 155.400 257.785 164.430 ;
        RECT 258.495 155.400 258.665 164.430 ;
        RECT 259.375 155.400 259.545 164.430 ;
        RECT 260.255 155.400 260.425 164.430 ;
        RECT 261.135 155.400 261.305 164.430 ;
        RECT 262.015 155.400 262.185 164.430 ;
        RECT 262.895 155.400 263.065 164.430 ;
        RECT 263.775 155.400 263.945 164.430 ;
        RECT 264.655 155.400 264.825 164.430 ;
        RECT 265.535 155.400 265.705 164.430 ;
        RECT 266.415 155.400 266.585 164.430 ;
        RECT 267.295 155.400 267.465 164.430 ;
        RECT 268.175 155.400 268.345 164.430 ;
        RECT 269.055 155.400 269.225 164.430 ;
        RECT 269.935 155.400 270.105 164.430 ;
        RECT 270.815 155.400 270.985 164.430 ;
        RECT 271.695 155.400 271.865 164.430 ;
        RECT 272.575 155.400 272.745 164.430 ;
        RECT 273.455 155.400 273.625 164.430 ;
        RECT 274.335 155.400 274.505 164.430 ;
        RECT 275.215 155.400 275.385 164.430 ;
        RECT 276.095 155.400 276.265 164.430 ;
        RECT 276.975 155.400 277.145 164.430 ;
        RECT 277.855 155.400 278.025 164.430 ;
        RECT 278.735 155.400 278.905 164.430 ;
        RECT 279.615 155.400 279.785 164.430 ;
        RECT 241.235 154.900 242.485 155.230 ;
        RECT 242.995 154.900 244.245 155.230 ;
        RECT 244.755 154.900 246.005 155.230 ;
        RECT 246.515 154.900 247.765 155.230 ;
        RECT 248.275 154.900 249.525 155.230 ;
        RECT 250.035 154.900 251.285 155.230 ;
        RECT 251.795 154.900 253.045 155.230 ;
        RECT 253.555 154.900 254.805 155.230 ;
        RECT 255.315 154.900 256.565 155.230 ;
        RECT 257.075 154.900 258.325 155.230 ;
        RECT 258.835 154.900 260.085 155.230 ;
        RECT 260.595 154.900 261.845 155.230 ;
        RECT 262.355 154.900 263.605 155.230 ;
        RECT 264.115 154.900 265.365 155.230 ;
        RECT 265.875 154.900 267.125 155.230 ;
        RECT 267.635 154.900 268.885 155.230 ;
        RECT 269.395 154.900 270.645 155.230 ;
        RECT 271.155 154.900 272.405 155.230 ;
        RECT 272.915 154.900 274.165 155.230 ;
        RECT 274.675 154.900 275.925 155.230 ;
        RECT 280.245 154.640 280.535 165.190 ;
        RECT 238.385 154.350 280.535 154.640 ;
        RECT 184.845 152.260 294.365 152.430 ;
        RECT 184.845 151.060 185.015 152.260 ;
        RECT 185.635 151.060 187.045 151.640 ;
        RECT 187.645 151.060 189.055 151.640 ;
        RECT 184.845 150.060 189.055 151.060 ;
        RECT 184.845 141.465 185.015 150.060 ;
        RECT 185.635 149.480 187.045 150.060 ;
        RECT 187.645 149.480 189.055 150.060 ;
        RECT 189.655 149.480 191.065 151.640 ;
        RECT 191.665 149.480 193.075 151.640 ;
        RECT 193.675 149.480 195.085 151.640 ;
        RECT 195.685 149.480 197.095 151.640 ;
        RECT 197.695 149.480 199.105 151.640 ;
        RECT 199.705 149.480 201.115 151.640 ;
        RECT 201.715 149.480 203.125 151.640 ;
        RECT 203.725 149.480 205.135 151.640 ;
        RECT 205.735 149.480 207.145 151.640 ;
        RECT 207.745 149.480 209.155 151.640 ;
        RECT 209.755 149.480 211.165 151.640 ;
        RECT 211.765 149.480 213.175 151.640 ;
        RECT 213.775 149.480 215.185 151.640 ;
        RECT 215.785 149.480 217.195 151.640 ;
        RECT 217.795 149.480 219.205 151.640 ;
        RECT 219.805 149.480 221.215 151.640 ;
        RECT 221.815 149.480 223.225 151.640 ;
        RECT 223.825 149.480 225.235 151.640 ;
        RECT 225.835 149.480 227.245 151.640 ;
        RECT 227.845 149.480 229.255 151.640 ;
        RECT 229.855 149.480 231.265 151.640 ;
        RECT 231.865 149.480 233.275 151.640 ;
        RECT 233.875 149.480 235.285 151.640 ;
        RECT 235.885 149.480 237.295 151.640 ;
        RECT 237.895 149.480 239.305 151.640 ;
        RECT 239.905 149.480 241.315 151.640 ;
        RECT 241.915 149.480 243.325 151.640 ;
        RECT 243.925 149.480 245.335 151.640 ;
        RECT 245.935 149.480 247.345 151.640 ;
        RECT 247.945 149.480 249.355 151.640 ;
        RECT 249.955 149.480 251.365 151.640 ;
        RECT 251.965 149.480 253.375 151.640 ;
        RECT 253.975 149.480 255.385 151.640 ;
        RECT 255.985 149.480 257.395 151.640 ;
        RECT 257.995 149.480 259.405 151.640 ;
        RECT 260.005 149.480 261.415 151.640 ;
        RECT 262.015 149.480 263.425 151.640 ;
        RECT 264.025 149.480 265.435 151.640 ;
        RECT 266.035 149.480 267.445 151.640 ;
        RECT 268.045 149.480 269.455 151.640 ;
        RECT 270.055 149.480 271.465 151.640 ;
        RECT 272.065 149.480 273.475 151.640 ;
        RECT 274.075 149.480 275.485 151.640 ;
        RECT 276.085 149.480 277.495 151.640 ;
        RECT 278.095 149.480 279.505 151.640 ;
        RECT 280.105 149.480 281.515 151.640 ;
        RECT 282.115 149.480 283.525 151.640 ;
        RECT 284.125 149.480 285.535 151.640 ;
        RECT 286.135 149.480 287.545 151.640 ;
        RECT 288.145 149.480 289.555 151.640 ;
        RECT 290.155 151.060 291.565 151.640 ;
        RECT 292.165 151.060 293.575 151.640 ;
        RECT 294.195 151.060 294.365 152.260 ;
        RECT 290.155 150.060 294.365 151.060 ;
        RECT 290.155 149.480 291.565 150.060 ;
        RECT 292.165 149.480 293.575 150.060 ;
        RECT 185.635 141.465 187.045 142.040 ;
        RECT 187.645 141.465 189.055 142.040 ;
        RECT 184.845 140.465 189.055 141.465 ;
        RECT 184.845 139.260 185.015 140.465 ;
        RECT 185.635 139.880 187.045 140.465 ;
        RECT 187.645 139.880 189.055 140.465 ;
        RECT 189.655 139.880 191.065 142.040 ;
        RECT 191.665 139.880 193.075 142.040 ;
        RECT 193.675 139.880 195.085 142.040 ;
        RECT 195.685 139.880 197.095 142.040 ;
        RECT 197.695 139.880 199.105 142.040 ;
        RECT 199.705 139.880 201.115 142.040 ;
        RECT 201.715 139.880 203.125 142.040 ;
        RECT 203.725 139.880 205.135 142.040 ;
        RECT 205.735 139.880 207.145 142.040 ;
        RECT 207.745 139.880 209.155 142.040 ;
        RECT 209.755 139.880 211.165 142.040 ;
        RECT 211.765 139.880 213.175 142.040 ;
        RECT 213.775 139.880 215.185 142.040 ;
        RECT 215.785 139.880 217.195 142.040 ;
        RECT 217.795 139.880 219.205 142.040 ;
        RECT 219.805 139.880 221.215 142.040 ;
        RECT 221.815 139.880 223.225 142.040 ;
        RECT 223.825 139.880 225.235 142.040 ;
        RECT 225.835 139.880 227.245 142.040 ;
        RECT 227.845 139.880 229.255 142.040 ;
        RECT 229.855 139.880 231.265 142.040 ;
        RECT 231.865 139.880 233.275 142.040 ;
        RECT 233.875 139.880 235.285 142.040 ;
        RECT 235.885 139.880 237.295 142.040 ;
        RECT 237.895 139.880 239.305 142.040 ;
        RECT 239.905 139.880 241.315 142.040 ;
        RECT 241.915 139.880 243.325 142.040 ;
        RECT 243.925 139.880 245.335 142.040 ;
        RECT 245.935 139.880 247.345 142.040 ;
        RECT 247.945 139.880 249.355 142.040 ;
        RECT 249.955 139.880 251.365 142.040 ;
        RECT 251.965 139.880 253.375 142.040 ;
        RECT 253.975 139.880 255.385 142.040 ;
        RECT 255.985 139.880 257.395 142.040 ;
        RECT 257.995 139.880 259.405 142.040 ;
        RECT 260.005 139.880 261.415 142.040 ;
        RECT 262.015 139.880 263.425 142.040 ;
        RECT 264.025 139.880 265.435 142.040 ;
        RECT 266.035 139.880 267.445 142.040 ;
        RECT 268.045 139.880 269.455 142.040 ;
        RECT 270.055 139.880 271.465 142.040 ;
        RECT 272.065 139.880 273.475 142.040 ;
        RECT 274.075 139.880 275.485 142.040 ;
        RECT 276.085 139.880 277.495 142.040 ;
        RECT 278.095 139.880 279.505 142.040 ;
        RECT 280.105 139.880 281.515 142.040 ;
        RECT 282.115 139.880 283.525 142.040 ;
        RECT 284.125 139.880 285.535 142.040 ;
        RECT 286.135 139.880 287.545 142.040 ;
        RECT 288.145 139.880 289.555 142.040 ;
        RECT 290.155 141.465 291.565 142.040 ;
        RECT 292.165 141.465 293.575 142.040 ;
        RECT 294.195 141.465 294.365 150.060 ;
        RECT 290.155 140.465 294.365 141.465 ;
        RECT 290.155 139.880 291.565 140.465 ;
        RECT 292.165 139.880 293.575 140.465 ;
        RECT 294.195 139.260 294.365 140.465 ;
        RECT 184.845 139.090 294.365 139.260 ;
        RECT 300.380 152.260 409.900 152.430 ;
        RECT 300.380 151.060 300.550 152.260 ;
        RECT 301.170 151.060 302.580 151.640 ;
        RECT 303.180 151.060 304.590 151.640 ;
        RECT 300.380 150.060 304.590 151.060 ;
        RECT 300.380 141.465 300.550 150.060 ;
        RECT 301.170 149.480 302.580 150.060 ;
        RECT 303.180 149.480 304.590 150.060 ;
        RECT 305.190 149.480 306.600 151.640 ;
        RECT 307.200 149.480 308.610 151.640 ;
        RECT 309.210 149.480 310.620 151.640 ;
        RECT 311.220 149.480 312.630 151.640 ;
        RECT 313.230 149.480 314.640 151.640 ;
        RECT 315.240 149.480 316.650 151.640 ;
        RECT 317.250 149.480 318.660 151.640 ;
        RECT 319.260 149.480 320.670 151.640 ;
        RECT 321.270 149.480 322.680 151.640 ;
        RECT 323.280 149.480 324.690 151.640 ;
        RECT 325.290 149.480 326.700 151.640 ;
        RECT 327.300 149.480 328.710 151.640 ;
        RECT 329.310 149.480 330.720 151.640 ;
        RECT 331.320 149.480 332.730 151.640 ;
        RECT 333.330 149.480 334.740 151.640 ;
        RECT 335.340 149.480 336.750 151.640 ;
        RECT 337.350 149.480 338.760 151.640 ;
        RECT 339.360 149.480 340.770 151.640 ;
        RECT 341.370 149.480 342.780 151.640 ;
        RECT 343.380 149.480 344.790 151.640 ;
        RECT 345.390 149.480 346.800 151.640 ;
        RECT 347.400 149.480 348.810 151.640 ;
        RECT 349.410 149.480 350.820 151.640 ;
        RECT 351.420 149.480 352.830 151.640 ;
        RECT 353.430 149.480 354.840 151.640 ;
        RECT 355.440 149.480 356.850 151.640 ;
        RECT 357.450 149.480 358.860 151.640 ;
        RECT 359.460 149.480 360.870 151.640 ;
        RECT 361.470 149.480 362.880 151.640 ;
        RECT 363.480 149.480 364.890 151.640 ;
        RECT 365.490 149.480 366.900 151.640 ;
        RECT 367.500 149.480 368.910 151.640 ;
        RECT 369.510 149.480 370.920 151.640 ;
        RECT 371.520 149.480 372.930 151.640 ;
        RECT 373.530 149.480 374.940 151.640 ;
        RECT 375.540 149.480 376.950 151.640 ;
        RECT 377.550 149.480 378.960 151.640 ;
        RECT 379.560 149.480 380.970 151.640 ;
        RECT 381.570 149.480 382.980 151.640 ;
        RECT 383.580 149.480 384.990 151.640 ;
        RECT 385.590 149.480 387.000 151.640 ;
        RECT 387.600 149.480 389.010 151.640 ;
        RECT 389.610 149.480 391.020 151.640 ;
        RECT 391.620 149.480 393.030 151.640 ;
        RECT 393.630 149.480 395.040 151.640 ;
        RECT 395.640 149.480 397.050 151.640 ;
        RECT 397.650 149.480 399.060 151.640 ;
        RECT 399.660 149.480 401.070 151.640 ;
        RECT 401.670 149.480 403.080 151.640 ;
        RECT 403.680 149.480 405.090 151.640 ;
        RECT 405.690 151.060 407.100 151.640 ;
        RECT 407.700 151.060 409.110 151.640 ;
        RECT 409.730 151.060 409.900 152.260 ;
        RECT 405.690 150.060 409.900 151.060 ;
        RECT 405.690 149.480 407.100 150.060 ;
        RECT 407.700 149.480 409.110 150.060 ;
        RECT 301.170 141.465 302.580 142.040 ;
        RECT 303.180 141.465 304.590 142.040 ;
        RECT 300.380 140.465 304.590 141.465 ;
        RECT 300.380 139.260 300.550 140.465 ;
        RECT 301.170 139.880 302.580 140.465 ;
        RECT 303.180 139.880 304.590 140.465 ;
        RECT 305.190 139.880 306.600 142.040 ;
        RECT 307.200 139.880 308.610 142.040 ;
        RECT 309.210 139.880 310.620 142.040 ;
        RECT 311.220 139.880 312.630 142.040 ;
        RECT 313.230 139.880 314.640 142.040 ;
        RECT 315.240 139.880 316.650 142.040 ;
        RECT 317.250 139.880 318.660 142.040 ;
        RECT 319.260 139.880 320.670 142.040 ;
        RECT 321.270 139.880 322.680 142.040 ;
        RECT 323.280 139.880 324.690 142.040 ;
        RECT 325.290 139.880 326.700 142.040 ;
        RECT 327.300 139.880 328.710 142.040 ;
        RECT 329.310 139.880 330.720 142.040 ;
        RECT 331.320 139.880 332.730 142.040 ;
        RECT 333.330 139.880 334.740 142.040 ;
        RECT 335.340 139.880 336.750 142.040 ;
        RECT 337.350 139.880 338.760 142.040 ;
        RECT 339.360 139.880 340.770 142.040 ;
        RECT 341.370 139.880 342.780 142.040 ;
        RECT 343.380 139.880 344.790 142.040 ;
        RECT 345.390 139.880 346.800 142.040 ;
        RECT 347.400 139.880 348.810 142.040 ;
        RECT 349.410 139.880 350.820 142.040 ;
        RECT 351.420 139.880 352.830 142.040 ;
        RECT 353.430 139.880 354.840 142.040 ;
        RECT 355.440 139.880 356.850 142.040 ;
        RECT 357.450 139.880 358.860 142.040 ;
        RECT 359.460 139.880 360.870 142.040 ;
        RECT 361.470 139.880 362.880 142.040 ;
        RECT 363.480 139.880 364.890 142.040 ;
        RECT 365.490 139.880 366.900 142.040 ;
        RECT 367.500 139.880 368.910 142.040 ;
        RECT 369.510 139.880 370.920 142.040 ;
        RECT 371.520 139.880 372.930 142.040 ;
        RECT 373.530 139.880 374.940 142.040 ;
        RECT 375.540 139.880 376.950 142.040 ;
        RECT 377.550 139.880 378.960 142.040 ;
        RECT 379.560 139.880 380.970 142.040 ;
        RECT 381.570 139.880 382.980 142.040 ;
        RECT 383.580 139.880 384.990 142.040 ;
        RECT 385.590 139.880 387.000 142.040 ;
        RECT 387.600 139.880 389.010 142.040 ;
        RECT 389.610 139.880 391.020 142.040 ;
        RECT 391.620 139.880 393.030 142.040 ;
        RECT 393.630 139.880 395.040 142.040 ;
        RECT 395.640 139.880 397.050 142.040 ;
        RECT 397.650 139.880 399.060 142.040 ;
        RECT 399.660 139.880 401.070 142.040 ;
        RECT 401.670 139.880 403.080 142.040 ;
        RECT 403.680 139.880 405.090 142.040 ;
        RECT 405.690 141.465 407.100 142.040 ;
        RECT 407.700 141.465 409.110 142.040 ;
        RECT 409.730 141.465 409.900 150.060 ;
        RECT 405.690 140.465 409.900 141.465 ;
        RECT 405.690 139.880 407.100 140.465 ;
        RECT 407.700 139.880 409.110 140.465 ;
        RECT 409.730 139.260 409.900 140.465 ;
        RECT 300.380 139.090 409.900 139.260 ;
        RECT 184.845 138.095 294.365 138.265 ;
        RECT 184.845 136.895 185.015 138.095 ;
        RECT 185.635 136.895 187.045 137.475 ;
        RECT 187.645 136.895 189.055 137.475 ;
        RECT 184.845 135.895 189.055 136.895 ;
        RECT 184.845 127.300 185.015 135.895 ;
        RECT 185.635 135.315 187.045 135.895 ;
        RECT 187.645 135.315 189.055 135.895 ;
        RECT 189.655 135.315 191.065 137.475 ;
        RECT 191.665 135.315 193.075 137.475 ;
        RECT 193.675 135.315 195.085 137.475 ;
        RECT 195.685 135.315 197.095 137.475 ;
        RECT 197.695 135.315 199.105 137.475 ;
        RECT 199.705 135.315 201.115 137.475 ;
        RECT 201.715 135.315 203.125 137.475 ;
        RECT 203.725 135.315 205.135 137.475 ;
        RECT 205.735 135.315 207.145 137.475 ;
        RECT 207.745 135.315 209.155 137.475 ;
        RECT 209.755 135.315 211.165 137.475 ;
        RECT 211.765 135.315 213.175 137.475 ;
        RECT 213.775 135.315 215.185 137.475 ;
        RECT 215.785 135.315 217.195 137.475 ;
        RECT 217.795 135.315 219.205 137.475 ;
        RECT 219.805 135.315 221.215 137.475 ;
        RECT 221.815 135.315 223.225 137.475 ;
        RECT 223.825 135.315 225.235 137.475 ;
        RECT 225.835 135.315 227.245 137.475 ;
        RECT 227.845 135.315 229.255 137.475 ;
        RECT 229.855 135.315 231.265 137.475 ;
        RECT 231.865 135.315 233.275 137.475 ;
        RECT 233.875 135.315 235.285 137.475 ;
        RECT 235.885 135.315 237.295 137.475 ;
        RECT 237.895 135.315 239.305 137.475 ;
        RECT 239.905 135.315 241.315 137.475 ;
        RECT 241.915 135.315 243.325 137.475 ;
        RECT 243.925 135.315 245.335 137.475 ;
        RECT 245.935 135.315 247.345 137.475 ;
        RECT 247.945 135.315 249.355 137.475 ;
        RECT 249.955 135.315 251.365 137.475 ;
        RECT 251.965 135.315 253.375 137.475 ;
        RECT 253.975 135.315 255.385 137.475 ;
        RECT 255.985 135.315 257.395 137.475 ;
        RECT 257.995 135.315 259.405 137.475 ;
        RECT 260.005 135.315 261.415 137.475 ;
        RECT 262.015 135.315 263.425 137.475 ;
        RECT 264.025 135.315 265.435 137.475 ;
        RECT 266.035 135.315 267.445 137.475 ;
        RECT 268.045 135.315 269.455 137.475 ;
        RECT 270.055 135.315 271.465 137.475 ;
        RECT 272.065 135.315 273.475 137.475 ;
        RECT 274.075 135.315 275.485 137.475 ;
        RECT 276.085 135.315 277.495 137.475 ;
        RECT 278.095 135.315 279.505 137.475 ;
        RECT 280.105 135.315 281.515 137.475 ;
        RECT 282.115 135.315 283.525 137.475 ;
        RECT 284.125 135.315 285.535 137.475 ;
        RECT 286.135 135.315 287.545 137.475 ;
        RECT 288.145 135.315 289.555 137.475 ;
        RECT 290.155 136.895 291.565 137.475 ;
        RECT 292.165 136.895 293.575 137.475 ;
        RECT 294.195 136.895 294.365 138.095 ;
        RECT 290.155 135.895 294.365 136.895 ;
        RECT 290.155 135.315 291.565 135.895 ;
        RECT 292.165 135.315 293.575 135.895 ;
        RECT 185.635 127.300 187.045 127.875 ;
        RECT 187.645 127.300 189.055 127.875 ;
        RECT 184.845 126.300 189.055 127.300 ;
        RECT 184.845 125.095 185.015 126.300 ;
        RECT 185.635 125.715 187.045 126.300 ;
        RECT 187.645 125.715 189.055 126.300 ;
        RECT 189.655 125.715 191.065 127.875 ;
        RECT 191.665 125.715 193.075 127.875 ;
        RECT 193.675 125.715 195.085 127.875 ;
        RECT 195.685 125.715 197.095 127.875 ;
        RECT 197.695 125.715 199.105 127.875 ;
        RECT 199.705 125.715 201.115 127.875 ;
        RECT 201.715 125.715 203.125 127.875 ;
        RECT 203.725 125.715 205.135 127.875 ;
        RECT 205.735 125.715 207.145 127.875 ;
        RECT 207.745 125.715 209.155 127.875 ;
        RECT 209.755 125.715 211.165 127.875 ;
        RECT 211.765 125.715 213.175 127.875 ;
        RECT 213.775 125.715 215.185 127.875 ;
        RECT 215.785 125.715 217.195 127.875 ;
        RECT 217.795 125.715 219.205 127.875 ;
        RECT 219.805 125.715 221.215 127.875 ;
        RECT 221.815 125.715 223.225 127.875 ;
        RECT 223.825 125.715 225.235 127.875 ;
        RECT 225.835 125.715 227.245 127.875 ;
        RECT 227.845 125.715 229.255 127.875 ;
        RECT 229.855 125.715 231.265 127.875 ;
        RECT 231.865 125.715 233.275 127.875 ;
        RECT 233.875 125.715 235.285 127.875 ;
        RECT 235.885 125.715 237.295 127.875 ;
        RECT 237.895 125.715 239.305 127.875 ;
        RECT 239.905 125.715 241.315 127.875 ;
        RECT 241.915 125.715 243.325 127.875 ;
        RECT 243.925 125.715 245.335 127.875 ;
        RECT 245.935 125.715 247.345 127.875 ;
        RECT 247.945 125.715 249.355 127.875 ;
        RECT 249.955 125.715 251.365 127.875 ;
        RECT 251.965 125.715 253.375 127.875 ;
        RECT 253.975 125.715 255.385 127.875 ;
        RECT 255.985 125.715 257.395 127.875 ;
        RECT 257.995 125.715 259.405 127.875 ;
        RECT 260.005 125.715 261.415 127.875 ;
        RECT 262.015 125.715 263.425 127.875 ;
        RECT 264.025 125.715 265.435 127.875 ;
        RECT 266.035 125.715 267.445 127.875 ;
        RECT 268.045 125.715 269.455 127.875 ;
        RECT 270.055 125.715 271.465 127.875 ;
        RECT 272.065 125.715 273.475 127.875 ;
        RECT 274.075 125.715 275.485 127.875 ;
        RECT 276.085 125.715 277.495 127.875 ;
        RECT 278.095 125.715 279.505 127.875 ;
        RECT 280.105 125.715 281.515 127.875 ;
        RECT 282.115 125.715 283.525 127.875 ;
        RECT 284.125 125.715 285.535 127.875 ;
        RECT 286.135 125.715 287.545 127.875 ;
        RECT 288.145 125.715 289.555 127.875 ;
        RECT 290.155 127.300 291.565 127.875 ;
        RECT 292.165 127.300 293.575 127.875 ;
        RECT 294.195 127.300 294.365 135.895 ;
        RECT 290.155 126.300 294.365 127.300 ;
        RECT 290.155 125.715 291.565 126.300 ;
        RECT 292.165 125.715 293.575 126.300 ;
        RECT 294.195 125.095 294.365 126.300 ;
        RECT 184.845 124.925 294.365 125.095 ;
        RECT 300.380 138.095 409.900 138.265 ;
        RECT 300.380 136.895 300.550 138.095 ;
        RECT 301.170 136.895 302.580 137.475 ;
        RECT 303.180 136.895 304.590 137.475 ;
        RECT 300.380 135.895 304.590 136.895 ;
        RECT 300.380 127.300 300.550 135.895 ;
        RECT 301.170 135.315 302.580 135.895 ;
        RECT 303.180 135.315 304.590 135.895 ;
        RECT 305.190 135.315 306.600 137.475 ;
        RECT 307.200 135.315 308.610 137.475 ;
        RECT 309.210 135.315 310.620 137.475 ;
        RECT 311.220 135.315 312.630 137.475 ;
        RECT 313.230 135.315 314.640 137.475 ;
        RECT 315.240 135.315 316.650 137.475 ;
        RECT 317.250 135.315 318.660 137.475 ;
        RECT 319.260 135.315 320.670 137.475 ;
        RECT 321.270 135.315 322.680 137.475 ;
        RECT 323.280 135.315 324.690 137.475 ;
        RECT 325.290 135.315 326.700 137.475 ;
        RECT 327.300 135.315 328.710 137.475 ;
        RECT 329.310 135.315 330.720 137.475 ;
        RECT 331.320 135.315 332.730 137.475 ;
        RECT 333.330 135.315 334.740 137.475 ;
        RECT 335.340 135.315 336.750 137.475 ;
        RECT 337.350 135.315 338.760 137.475 ;
        RECT 339.360 135.315 340.770 137.475 ;
        RECT 341.370 135.315 342.780 137.475 ;
        RECT 343.380 135.315 344.790 137.475 ;
        RECT 345.390 135.315 346.800 137.475 ;
        RECT 347.400 135.315 348.810 137.475 ;
        RECT 349.410 135.315 350.820 137.475 ;
        RECT 351.420 135.315 352.830 137.475 ;
        RECT 353.430 135.315 354.840 137.475 ;
        RECT 355.440 135.315 356.850 137.475 ;
        RECT 357.450 135.315 358.860 137.475 ;
        RECT 359.460 135.315 360.870 137.475 ;
        RECT 361.470 135.315 362.880 137.475 ;
        RECT 363.480 135.315 364.890 137.475 ;
        RECT 365.490 135.315 366.900 137.475 ;
        RECT 367.500 135.315 368.910 137.475 ;
        RECT 369.510 135.315 370.920 137.475 ;
        RECT 371.520 135.315 372.930 137.475 ;
        RECT 373.530 135.315 374.940 137.475 ;
        RECT 375.540 135.315 376.950 137.475 ;
        RECT 377.550 135.315 378.960 137.475 ;
        RECT 379.560 135.315 380.970 137.475 ;
        RECT 381.570 135.315 382.980 137.475 ;
        RECT 383.580 135.315 384.990 137.475 ;
        RECT 385.590 135.315 387.000 137.475 ;
        RECT 387.600 135.315 389.010 137.475 ;
        RECT 389.610 135.315 391.020 137.475 ;
        RECT 391.620 135.315 393.030 137.475 ;
        RECT 393.630 135.315 395.040 137.475 ;
        RECT 395.640 135.315 397.050 137.475 ;
        RECT 397.650 135.315 399.060 137.475 ;
        RECT 399.660 135.315 401.070 137.475 ;
        RECT 401.670 135.315 403.080 137.475 ;
        RECT 403.680 135.315 405.090 137.475 ;
        RECT 405.690 136.895 407.100 137.475 ;
        RECT 407.700 136.895 409.110 137.475 ;
        RECT 409.730 136.895 409.900 138.095 ;
        RECT 405.690 135.895 409.900 136.895 ;
        RECT 405.690 135.315 407.100 135.895 ;
        RECT 407.700 135.315 409.110 135.895 ;
        RECT 301.170 127.300 302.580 127.875 ;
        RECT 303.180 127.300 304.590 127.875 ;
        RECT 300.380 126.300 304.590 127.300 ;
        RECT 300.380 125.095 300.550 126.300 ;
        RECT 301.170 125.715 302.580 126.300 ;
        RECT 303.180 125.715 304.590 126.300 ;
        RECT 305.190 125.715 306.600 127.875 ;
        RECT 307.200 125.715 308.610 127.875 ;
        RECT 309.210 125.715 310.620 127.875 ;
        RECT 311.220 125.715 312.630 127.875 ;
        RECT 313.230 125.715 314.640 127.875 ;
        RECT 315.240 125.715 316.650 127.875 ;
        RECT 317.250 125.715 318.660 127.875 ;
        RECT 319.260 125.715 320.670 127.875 ;
        RECT 321.270 125.715 322.680 127.875 ;
        RECT 323.280 125.715 324.690 127.875 ;
        RECT 325.290 125.715 326.700 127.875 ;
        RECT 327.300 125.715 328.710 127.875 ;
        RECT 329.310 125.715 330.720 127.875 ;
        RECT 331.320 125.715 332.730 127.875 ;
        RECT 333.330 125.715 334.740 127.875 ;
        RECT 335.340 125.715 336.750 127.875 ;
        RECT 337.350 125.715 338.760 127.875 ;
        RECT 339.360 125.715 340.770 127.875 ;
        RECT 341.370 125.715 342.780 127.875 ;
        RECT 343.380 125.715 344.790 127.875 ;
        RECT 345.390 125.715 346.800 127.875 ;
        RECT 347.400 125.715 348.810 127.875 ;
        RECT 349.410 125.715 350.820 127.875 ;
        RECT 351.420 125.715 352.830 127.875 ;
        RECT 353.430 125.715 354.840 127.875 ;
        RECT 355.440 125.715 356.850 127.875 ;
        RECT 357.450 125.715 358.860 127.875 ;
        RECT 359.460 125.715 360.870 127.875 ;
        RECT 361.470 125.715 362.880 127.875 ;
        RECT 363.480 125.715 364.890 127.875 ;
        RECT 365.490 125.715 366.900 127.875 ;
        RECT 367.500 125.715 368.910 127.875 ;
        RECT 369.510 125.715 370.920 127.875 ;
        RECT 371.520 125.715 372.930 127.875 ;
        RECT 373.530 125.715 374.940 127.875 ;
        RECT 375.540 125.715 376.950 127.875 ;
        RECT 377.550 125.715 378.960 127.875 ;
        RECT 379.560 125.715 380.970 127.875 ;
        RECT 381.570 125.715 382.980 127.875 ;
        RECT 383.580 125.715 384.990 127.875 ;
        RECT 385.590 125.715 387.000 127.875 ;
        RECT 387.600 125.715 389.010 127.875 ;
        RECT 389.610 125.715 391.020 127.875 ;
        RECT 391.620 125.715 393.030 127.875 ;
        RECT 393.630 125.715 395.040 127.875 ;
        RECT 395.640 125.715 397.050 127.875 ;
        RECT 397.650 125.715 399.060 127.875 ;
        RECT 399.660 125.715 401.070 127.875 ;
        RECT 401.670 125.715 403.080 127.875 ;
        RECT 403.680 125.715 405.090 127.875 ;
        RECT 405.690 127.300 407.100 127.875 ;
        RECT 407.700 127.300 409.110 127.875 ;
        RECT 409.730 127.300 409.900 135.895 ;
        RECT 405.690 126.300 409.900 127.300 ;
        RECT 405.690 125.715 407.100 126.300 ;
        RECT 407.700 125.715 409.110 126.300 ;
        RECT 409.730 125.095 409.900 126.300 ;
        RECT 300.380 124.925 409.900 125.095 ;
        RECT 310.915 120.535 333.665 120.705 ;
        RECT 217.170 117.505 290.510 117.675 ;
        RECT 217.170 116.305 217.340 117.505 ;
        RECT 217.960 116.305 219.370 116.885 ;
        RECT 219.970 116.305 221.380 116.885 ;
        RECT 217.170 115.305 221.380 116.305 ;
        RECT 184.800 115.045 198.350 115.215 ;
        RECT 184.800 112.625 184.970 115.045 ;
        RECT 185.470 113.585 185.640 114.585 ;
        RECT 185.900 113.585 186.070 114.585 ;
        RECT 186.330 113.585 186.500 114.585 ;
        RECT 186.760 113.585 186.930 114.585 ;
        RECT 187.190 113.585 187.360 114.585 ;
        RECT 187.620 113.585 187.790 114.585 ;
        RECT 188.050 113.585 188.220 114.585 ;
        RECT 188.480 113.585 188.650 114.585 ;
        RECT 188.910 113.585 189.080 114.585 ;
        RECT 189.340 113.585 189.510 114.585 ;
        RECT 189.770 113.585 189.940 114.585 ;
        RECT 190.200 113.585 190.370 114.585 ;
        RECT 190.630 113.585 190.800 114.585 ;
        RECT 191.060 113.585 191.230 114.585 ;
        RECT 191.490 113.585 191.660 114.585 ;
        RECT 191.920 113.585 192.090 114.585 ;
        RECT 192.350 113.585 192.520 114.585 ;
        RECT 192.780 113.585 192.950 114.585 ;
        RECT 193.210 113.585 193.380 114.585 ;
        RECT 193.640 113.585 193.810 114.585 ;
        RECT 194.070 113.585 194.240 114.585 ;
        RECT 194.500 113.585 194.670 114.585 ;
        RECT 194.930 113.585 195.100 114.585 ;
        RECT 195.360 113.585 195.530 114.585 ;
        RECT 195.790 113.585 195.960 114.585 ;
        RECT 196.220 113.585 196.390 114.585 ;
        RECT 196.650 113.585 196.820 114.585 ;
        RECT 197.080 113.585 197.250 114.585 ;
        RECT 197.510 113.585 197.680 114.585 ;
        RECT 185.695 113.145 186.275 113.375 ;
        RECT 186.555 113.145 196.595 113.375 ;
        RECT 196.875 113.145 197.455 113.375 ;
        RECT 198.180 112.625 198.350 115.045 ;
        RECT 199.880 113.185 213.430 113.355 ;
        RECT 184.800 109.730 184.970 112.120 ;
        RECT 185.695 111.370 189.715 111.600 ;
        RECT 189.995 111.370 193.155 111.600 ;
        RECT 193.435 111.370 197.455 111.600 ;
        RECT 185.470 110.160 185.640 111.160 ;
        RECT 185.900 110.160 186.070 111.160 ;
        RECT 186.330 110.160 186.500 111.160 ;
        RECT 186.760 110.160 186.930 111.160 ;
        RECT 187.190 110.160 187.360 111.160 ;
        RECT 187.620 110.160 187.790 111.160 ;
        RECT 188.050 110.160 188.220 111.160 ;
        RECT 188.480 110.160 188.650 111.160 ;
        RECT 188.910 110.160 189.080 111.160 ;
        RECT 189.340 110.160 189.510 111.160 ;
        RECT 189.770 110.160 189.940 111.160 ;
        RECT 190.200 110.160 190.370 111.160 ;
        RECT 190.630 110.160 190.800 111.160 ;
        RECT 191.060 110.160 191.230 111.160 ;
        RECT 191.490 110.160 191.660 111.160 ;
        RECT 191.920 110.160 192.090 111.160 ;
        RECT 192.350 110.160 192.520 111.160 ;
        RECT 192.780 110.160 192.950 111.160 ;
        RECT 193.210 110.160 193.380 111.160 ;
        RECT 193.640 110.160 193.810 111.160 ;
        RECT 194.070 110.160 194.240 111.160 ;
        RECT 194.500 110.160 194.670 111.160 ;
        RECT 194.930 110.160 195.100 111.160 ;
        RECT 195.360 110.160 195.530 111.160 ;
        RECT 195.790 110.160 195.960 111.160 ;
        RECT 196.220 110.160 196.390 111.160 ;
        RECT 196.650 110.160 196.820 111.160 ;
        RECT 197.080 110.160 197.250 111.160 ;
        RECT 197.510 110.160 197.680 111.160 ;
        RECT 198.180 109.730 198.350 112.120 ;
        RECT 199.880 110.235 200.050 113.185 ;
        RECT 200.800 112.365 201.330 112.695 ;
        RECT 211.980 112.365 212.510 112.695 ;
        RECT 200.550 111.195 200.720 112.195 ;
        RECT 200.980 111.195 201.150 112.195 ;
        RECT 201.410 111.195 201.580 112.195 ;
        RECT 201.840 111.195 202.010 112.195 ;
        RECT 202.270 111.195 202.440 112.195 ;
        RECT 202.700 111.195 202.870 112.195 ;
        RECT 203.130 111.195 203.300 112.195 ;
        RECT 203.560 111.195 203.730 112.195 ;
        RECT 203.990 111.195 204.160 112.195 ;
        RECT 204.420 111.195 204.590 112.195 ;
        RECT 204.850 111.195 205.020 112.195 ;
        RECT 205.280 111.195 205.450 112.195 ;
        RECT 205.710 111.195 205.880 112.195 ;
        RECT 206.140 111.195 206.310 112.195 ;
        RECT 206.570 111.195 206.740 112.195 ;
        RECT 207.000 111.195 207.170 112.195 ;
        RECT 207.430 111.195 207.600 112.195 ;
        RECT 207.860 111.195 208.030 112.195 ;
        RECT 208.290 111.195 208.460 112.195 ;
        RECT 208.720 111.195 208.890 112.195 ;
        RECT 209.150 111.195 209.320 112.195 ;
        RECT 209.580 111.195 209.750 112.195 ;
        RECT 210.010 111.195 210.180 112.195 ;
        RECT 210.440 111.195 210.610 112.195 ;
        RECT 210.870 111.195 211.040 112.195 ;
        RECT 211.300 111.195 211.470 112.195 ;
        RECT 211.730 111.195 211.900 112.195 ;
        RECT 212.160 111.195 212.330 112.195 ;
        RECT 212.590 111.195 212.760 112.195 ;
        RECT 201.635 110.755 211.675 110.985 ;
        RECT 213.260 110.235 213.430 113.185 ;
        RECT 184.800 109.560 198.350 109.730 ;
        RECT 184.800 107.170 184.970 109.560 ;
        RECT 185.470 108.130 185.640 109.130 ;
        RECT 185.900 108.130 186.070 109.130 ;
        RECT 186.330 108.130 186.500 109.130 ;
        RECT 186.760 108.130 186.930 109.130 ;
        RECT 187.190 108.130 187.360 109.130 ;
        RECT 187.620 108.130 187.790 109.130 ;
        RECT 188.050 108.130 188.220 109.130 ;
        RECT 188.480 108.130 188.650 109.130 ;
        RECT 188.910 108.130 189.080 109.130 ;
        RECT 189.340 108.130 189.510 109.130 ;
        RECT 189.770 108.130 189.940 109.130 ;
        RECT 190.200 108.130 190.370 109.130 ;
        RECT 190.630 108.130 190.800 109.130 ;
        RECT 191.060 108.130 191.230 109.130 ;
        RECT 191.490 108.130 191.660 109.130 ;
        RECT 191.920 108.130 192.090 109.130 ;
        RECT 192.350 108.130 192.520 109.130 ;
        RECT 192.780 108.130 192.950 109.130 ;
        RECT 193.210 108.130 193.380 109.130 ;
        RECT 193.640 108.130 193.810 109.130 ;
        RECT 194.070 108.130 194.240 109.130 ;
        RECT 194.500 108.130 194.670 109.130 ;
        RECT 194.930 108.130 195.100 109.130 ;
        RECT 195.360 108.130 195.530 109.130 ;
        RECT 195.790 108.130 195.960 109.130 ;
        RECT 196.220 108.130 196.390 109.130 ;
        RECT 196.650 108.130 196.820 109.130 ;
        RECT 197.080 108.130 197.250 109.130 ;
        RECT 197.510 108.130 197.680 109.130 ;
        RECT 185.695 107.690 189.715 107.920 ;
        RECT 189.995 107.690 193.155 107.920 ;
        RECT 193.435 107.690 197.455 107.920 ;
        RECT 198.180 107.170 198.350 109.560 ;
        RECT 184.800 104.245 184.970 106.665 ;
        RECT 185.695 105.915 186.275 106.145 ;
        RECT 186.555 105.915 196.595 106.145 ;
        RECT 196.875 105.915 197.455 106.145 ;
        RECT 185.470 104.705 185.640 105.705 ;
        RECT 185.900 104.705 186.070 105.705 ;
        RECT 186.330 104.705 186.500 105.705 ;
        RECT 186.760 104.705 186.930 105.705 ;
        RECT 187.190 104.705 187.360 105.705 ;
        RECT 187.620 104.705 187.790 105.705 ;
        RECT 188.050 104.705 188.220 105.705 ;
        RECT 188.480 104.705 188.650 105.705 ;
        RECT 188.910 104.705 189.080 105.705 ;
        RECT 189.340 104.705 189.510 105.705 ;
        RECT 189.770 104.705 189.940 105.705 ;
        RECT 190.200 104.705 190.370 105.705 ;
        RECT 190.630 104.705 190.800 105.705 ;
        RECT 191.060 104.705 191.230 105.705 ;
        RECT 191.490 104.705 191.660 105.705 ;
        RECT 191.920 104.705 192.090 105.705 ;
        RECT 192.350 104.705 192.520 105.705 ;
        RECT 192.780 104.705 192.950 105.705 ;
        RECT 193.210 104.705 193.380 105.705 ;
        RECT 193.640 104.705 193.810 105.705 ;
        RECT 194.070 104.705 194.240 105.705 ;
        RECT 194.500 104.705 194.670 105.705 ;
        RECT 194.930 104.705 195.100 105.705 ;
        RECT 195.360 104.705 195.530 105.705 ;
        RECT 195.790 104.705 195.960 105.705 ;
        RECT 196.220 104.705 196.390 105.705 ;
        RECT 196.650 104.705 196.820 105.705 ;
        RECT 197.080 104.705 197.250 105.705 ;
        RECT 197.510 104.705 197.680 105.705 ;
        RECT 198.180 104.245 198.350 106.665 ;
        RECT 199.880 106.265 200.050 109.355 ;
        RECT 205.075 108.305 208.235 108.535 ;
        RECT 200.550 107.095 200.720 108.095 ;
        RECT 200.980 107.095 201.150 108.095 ;
        RECT 201.410 107.095 201.580 108.095 ;
        RECT 201.840 107.095 202.010 108.095 ;
        RECT 202.270 107.095 202.440 108.095 ;
        RECT 202.700 107.095 202.870 108.095 ;
        RECT 203.130 107.095 203.300 108.095 ;
        RECT 203.560 107.095 203.730 108.095 ;
        RECT 203.990 107.095 204.160 108.095 ;
        RECT 204.420 107.095 204.590 108.095 ;
        RECT 204.850 107.095 205.020 108.095 ;
        RECT 205.280 107.095 205.450 108.095 ;
        RECT 205.710 107.095 205.880 108.095 ;
        RECT 206.140 107.095 206.310 108.095 ;
        RECT 206.570 107.095 206.740 108.095 ;
        RECT 207.000 107.095 207.170 108.095 ;
        RECT 207.430 107.095 207.600 108.095 ;
        RECT 207.860 107.095 208.030 108.095 ;
        RECT 208.290 107.095 208.460 108.095 ;
        RECT 208.720 107.095 208.890 108.095 ;
        RECT 209.150 107.095 209.320 108.095 ;
        RECT 209.580 107.095 209.750 108.095 ;
        RECT 210.010 107.095 210.180 108.095 ;
        RECT 210.440 107.095 210.610 108.095 ;
        RECT 210.870 107.095 211.040 108.095 ;
        RECT 211.300 107.095 211.470 108.095 ;
        RECT 211.730 107.095 211.900 108.095 ;
        RECT 212.160 107.095 212.330 108.095 ;
        RECT 212.590 107.095 212.760 108.095 ;
        RECT 204.635 106.885 204.805 106.925 ;
        RECT 208.505 106.885 208.675 106.925 ;
        RECT 200.775 106.655 204.835 106.885 ;
        RECT 208.475 106.655 212.535 106.885 ;
        RECT 204.635 106.595 204.805 106.655 ;
        RECT 208.505 106.595 208.675 106.655 ;
        RECT 213.260 106.265 213.430 109.355 ;
        RECT 199.880 106.095 213.430 106.265 ;
        RECT 217.170 106.705 217.340 115.305 ;
        RECT 217.960 114.725 219.370 115.305 ;
        RECT 219.970 114.725 221.380 115.305 ;
        RECT 221.980 114.725 223.390 116.885 ;
        RECT 223.990 114.725 225.400 116.885 ;
        RECT 226.000 114.725 227.410 116.885 ;
        RECT 228.010 114.725 229.420 116.885 ;
        RECT 230.020 114.725 231.430 116.885 ;
        RECT 232.030 114.725 233.440 116.885 ;
        RECT 234.040 114.725 235.450 116.885 ;
        RECT 236.050 114.725 237.460 116.885 ;
        RECT 238.060 114.725 239.470 116.885 ;
        RECT 240.070 114.725 241.480 116.885 ;
        RECT 242.080 114.725 243.490 116.885 ;
        RECT 244.090 114.725 245.500 116.885 ;
        RECT 246.100 114.725 247.510 116.885 ;
        RECT 248.110 114.725 249.520 116.885 ;
        RECT 250.120 114.725 251.530 116.885 ;
        RECT 252.130 114.725 253.540 116.885 ;
        RECT 254.140 114.725 255.550 116.885 ;
        RECT 256.150 114.725 257.560 116.885 ;
        RECT 258.160 114.725 259.570 116.885 ;
        RECT 260.170 114.725 261.580 116.885 ;
        RECT 262.180 114.725 263.590 116.885 ;
        RECT 264.190 114.725 265.600 116.885 ;
        RECT 266.200 114.725 267.610 116.885 ;
        RECT 268.210 114.725 269.620 116.885 ;
        RECT 270.220 114.725 271.630 116.885 ;
        RECT 272.230 114.725 273.640 116.885 ;
        RECT 274.240 114.725 275.650 116.885 ;
        RECT 276.250 114.725 277.660 116.885 ;
        RECT 278.260 114.725 279.670 116.885 ;
        RECT 280.270 114.725 281.680 116.885 ;
        RECT 282.280 114.725 283.690 116.885 ;
        RECT 284.290 114.725 285.700 116.885 ;
        RECT 286.300 116.305 287.710 116.885 ;
        RECT 288.310 116.305 289.720 116.885 ;
        RECT 290.340 116.305 290.510 117.505 ;
        RECT 310.915 116.475 311.085 120.535 ;
        RECT 319.025 119.805 320.275 120.135 ;
        RECT 320.785 119.805 322.035 120.135 ;
        RECT 322.545 119.805 323.795 120.135 ;
        RECT 324.305 119.805 325.555 120.135 ;
        RECT 311.645 117.375 311.815 119.635 ;
        RECT 312.525 117.375 312.695 119.635 ;
        RECT 313.405 117.375 313.575 119.635 ;
        RECT 314.285 117.375 314.455 119.635 ;
        RECT 315.165 117.375 315.335 119.635 ;
        RECT 316.045 117.375 316.215 119.635 ;
        RECT 316.925 117.375 317.095 119.635 ;
        RECT 317.805 117.375 317.975 119.635 ;
        RECT 318.685 117.375 318.855 119.635 ;
        RECT 319.565 117.375 319.735 119.635 ;
        RECT 320.445 117.375 320.615 119.635 ;
        RECT 321.325 117.375 321.495 119.635 ;
        RECT 322.205 117.375 322.375 119.635 ;
        RECT 323.085 117.375 323.255 119.635 ;
        RECT 323.965 117.375 324.135 119.635 ;
        RECT 324.845 117.375 325.015 119.635 ;
        RECT 325.725 117.375 325.895 119.635 ;
        RECT 326.605 117.375 326.775 119.635 ;
        RECT 327.485 117.375 327.655 119.635 ;
        RECT 328.365 117.375 328.535 119.635 ;
        RECT 329.245 117.375 329.415 119.635 ;
        RECT 330.125 117.375 330.295 119.635 ;
        RECT 331.005 117.375 331.175 119.635 ;
        RECT 331.885 117.375 332.055 119.635 ;
        RECT 332.765 117.375 332.935 119.635 ;
        RECT 311.985 116.875 313.235 117.205 ;
        RECT 313.745 116.875 314.995 117.205 ;
        RECT 315.505 116.875 316.755 117.205 ;
        RECT 317.265 116.875 318.515 117.205 ;
        RECT 326.065 116.875 327.315 117.205 ;
        RECT 327.825 116.875 329.075 117.205 ;
        RECT 329.585 116.875 330.835 117.205 ;
        RECT 331.345 116.875 332.595 117.205 ;
        RECT 333.495 116.475 333.665 120.535 ;
        RECT 310.915 116.305 333.665 116.475 ;
        RECT 334.135 120.535 363.925 120.705 ;
        RECT 334.135 116.475 334.305 120.535 ;
        RECT 347.525 119.805 348.775 120.135 ;
        RECT 349.285 119.805 350.535 120.135 ;
        RECT 334.865 117.375 335.035 119.635 ;
        RECT 335.745 117.375 335.915 119.635 ;
        RECT 336.625 117.375 336.795 119.635 ;
        RECT 337.505 117.375 337.675 119.635 ;
        RECT 338.385 117.375 338.555 119.635 ;
        RECT 339.265 117.375 339.435 119.635 ;
        RECT 340.145 117.375 340.315 119.635 ;
        RECT 341.025 117.375 341.195 119.635 ;
        RECT 341.905 117.375 342.075 119.635 ;
        RECT 342.785 117.375 342.955 119.635 ;
        RECT 343.665 117.375 343.835 119.635 ;
        RECT 344.545 117.375 344.715 119.635 ;
        RECT 345.425 117.375 345.595 119.635 ;
        RECT 346.305 117.375 346.475 119.635 ;
        RECT 347.185 117.375 347.355 119.635 ;
        RECT 348.065 117.375 348.235 119.635 ;
        RECT 348.945 117.375 349.115 119.635 ;
        RECT 349.825 117.375 349.995 119.635 ;
        RECT 350.705 117.375 350.875 119.635 ;
        RECT 351.585 117.375 351.755 119.635 ;
        RECT 352.465 117.375 352.635 119.635 ;
        RECT 353.345 117.375 353.515 119.635 ;
        RECT 354.225 117.375 354.395 119.635 ;
        RECT 355.105 117.375 355.275 119.635 ;
        RECT 355.985 117.375 356.155 119.635 ;
        RECT 356.865 117.375 357.035 119.635 ;
        RECT 357.745 117.375 357.915 119.635 ;
        RECT 358.625 117.375 358.795 119.635 ;
        RECT 359.505 117.375 359.675 119.635 ;
        RECT 360.385 117.375 360.555 119.635 ;
        RECT 361.265 117.375 361.435 119.635 ;
        RECT 362.145 117.375 362.315 119.635 ;
        RECT 363.025 117.375 363.195 119.635 ;
        RECT 335.205 116.875 336.455 117.205 ;
        RECT 336.965 116.875 338.215 117.205 ;
        RECT 338.725 116.875 339.975 117.205 ;
        RECT 340.485 116.875 341.735 117.205 ;
        RECT 342.245 116.875 343.495 117.205 ;
        RECT 344.005 116.875 345.255 117.205 ;
        RECT 345.765 116.875 347.015 117.205 ;
        RECT 351.045 116.875 352.295 117.205 ;
        RECT 352.805 116.875 354.055 117.205 ;
        RECT 354.565 116.875 355.815 117.205 ;
        RECT 356.325 116.875 357.575 117.205 ;
        RECT 358.085 116.875 359.335 117.205 ;
        RECT 359.845 116.875 361.095 117.205 ;
        RECT 361.605 116.875 362.855 117.205 ;
        RECT 363.755 116.475 363.925 120.535 ;
        RECT 334.135 116.305 363.925 116.475 ;
        RECT 364.475 120.535 406.580 120.705 ;
        RECT 364.475 116.475 364.645 120.535 ;
        RECT 365.205 117.375 365.375 119.635 ;
        RECT 366.085 117.375 366.255 119.635 ;
        RECT 366.965 117.375 367.135 119.635 ;
        RECT 367.845 117.375 368.015 119.635 ;
        RECT 368.725 117.375 368.895 119.635 ;
        RECT 369.605 117.375 369.775 119.635 ;
        RECT 370.485 117.375 370.655 119.635 ;
        RECT 371.365 117.375 371.535 119.635 ;
        RECT 372.245 117.375 372.415 119.635 ;
        RECT 373.125 117.375 373.295 119.635 ;
        RECT 374.005 117.375 374.175 119.635 ;
        RECT 374.885 117.375 375.055 119.635 ;
        RECT 375.765 117.375 375.935 119.635 ;
        RECT 376.645 117.375 376.815 119.635 ;
        RECT 377.525 117.375 377.695 119.635 ;
        RECT 378.405 117.375 378.575 119.635 ;
        RECT 379.285 117.375 379.455 119.635 ;
        RECT 380.165 117.375 380.335 119.635 ;
        RECT 381.045 117.375 381.215 119.635 ;
        RECT 381.925 117.375 382.095 119.635 ;
        RECT 382.805 117.375 382.975 119.635 ;
        RECT 383.685 117.375 383.855 119.635 ;
        RECT 384.565 117.375 384.735 119.635 ;
        RECT 385.445 117.375 385.615 119.635 ;
        RECT 386.325 117.375 386.495 119.635 ;
        RECT 387.205 117.375 387.375 119.635 ;
        RECT 388.085 117.375 388.255 119.635 ;
        RECT 388.965 117.375 389.135 119.635 ;
        RECT 389.845 117.375 390.015 119.635 ;
        RECT 390.725 117.375 390.895 119.635 ;
        RECT 391.605 117.375 391.775 119.635 ;
        RECT 392.485 117.375 392.655 119.635 ;
        RECT 393.365 117.375 393.535 119.635 ;
        RECT 394.245 117.375 394.415 119.635 ;
        RECT 395.125 117.375 395.295 119.635 ;
        RECT 396.005 117.375 396.175 119.635 ;
        RECT 396.885 117.375 397.055 119.635 ;
        RECT 397.765 117.375 397.935 119.635 ;
        RECT 398.645 117.375 398.815 119.635 ;
        RECT 399.525 117.375 399.695 119.635 ;
        RECT 400.405 117.375 400.575 119.635 ;
        RECT 401.285 117.375 401.455 119.635 ;
        RECT 402.165 117.375 402.335 119.635 ;
        RECT 403.045 117.375 403.215 119.635 ;
        RECT 403.925 117.375 404.095 119.635 ;
        RECT 404.805 117.375 404.975 119.635 ;
        RECT 405.685 117.375 405.855 119.635 ;
        RECT 365.545 116.875 366.795 117.205 ;
        RECT 367.305 116.875 368.555 117.205 ;
        RECT 369.065 116.875 370.315 117.205 ;
        RECT 370.825 116.875 372.075 117.205 ;
        RECT 372.585 116.875 373.835 117.205 ;
        RECT 374.345 116.875 375.595 117.205 ;
        RECT 376.105 116.875 377.355 117.205 ;
        RECT 377.865 116.875 379.115 117.205 ;
        RECT 379.625 116.875 380.875 117.205 ;
        RECT 381.385 116.875 382.635 117.205 ;
        RECT 383.145 116.875 384.395 117.205 ;
        RECT 384.905 116.875 386.155 117.205 ;
        RECT 386.665 116.875 387.915 117.205 ;
        RECT 388.425 116.875 389.675 117.205 ;
        RECT 390.185 116.875 391.435 117.205 ;
        RECT 391.945 116.875 393.195 117.205 ;
        RECT 393.705 116.875 394.955 117.205 ;
        RECT 395.465 116.875 396.715 117.205 ;
        RECT 397.225 116.875 398.475 117.205 ;
        RECT 398.985 116.875 400.235 117.205 ;
        RECT 400.745 116.875 401.995 117.205 ;
        RECT 402.505 116.875 403.755 117.205 ;
        RECT 404.265 116.875 405.515 117.205 ;
        RECT 406.410 116.475 406.580 120.535 ;
        RECT 364.475 116.305 406.580 116.475 ;
        RECT 444.015 118.795 452.685 119.085 ;
        RECT 286.300 115.305 290.510 116.305 ;
        RECT 286.300 114.725 287.710 115.305 ;
        RECT 288.310 114.725 289.720 115.305 ;
        RECT 217.960 106.705 219.370 107.285 ;
        RECT 219.970 106.705 221.380 107.285 ;
        RECT 217.170 105.705 221.380 106.705 ;
        RECT 217.170 104.505 217.340 105.705 ;
        RECT 217.960 105.125 219.370 105.705 ;
        RECT 219.970 105.125 221.380 105.705 ;
        RECT 221.980 105.125 223.390 107.285 ;
        RECT 223.990 105.125 225.400 107.285 ;
        RECT 226.000 105.125 227.410 107.285 ;
        RECT 228.010 105.125 229.420 107.285 ;
        RECT 230.020 105.125 231.430 107.285 ;
        RECT 232.030 105.125 233.440 107.285 ;
        RECT 234.040 105.125 235.450 107.285 ;
        RECT 236.050 105.125 237.460 107.285 ;
        RECT 238.060 105.125 239.470 107.285 ;
        RECT 240.070 105.125 241.480 107.285 ;
        RECT 242.080 105.125 243.490 107.285 ;
        RECT 244.090 105.125 245.500 107.285 ;
        RECT 246.100 105.125 247.510 107.285 ;
        RECT 248.110 105.125 249.520 107.285 ;
        RECT 250.120 105.125 251.530 107.285 ;
        RECT 252.130 105.125 253.540 107.285 ;
        RECT 254.140 105.125 255.550 107.285 ;
        RECT 256.150 105.125 257.560 107.285 ;
        RECT 258.160 105.125 259.570 107.285 ;
        RECT 260.170 105.125 261.580 107.285 ;
        RECT 262.180 105.125 263.590 107.285 ;
        RECT 264.190 105.125 265.600 107.285 ;
        RECT 266.200 105.125 267.610 107.285 ;
        RECT 268.210 105.125 269.620 107.285 ;
        RECT 270.220 105.125 271.630 107.285 ;
        RECT 272.230 105.125 273.640 107.285 ;
        RECT 274.240 105.125 275.650 107.285 ;
        RECT 276.250 105.125 277.660 107.285 ;
        RECT 278.260 105.125 279.670 107.285 ;
        RECT 280.270 105.125 281.680 107.285 ;
        RECT 282.280 105.125 283.690 107.285 ;
        RECT 284.290 105.125 285.700 107.285 ;
        RECT 286.300 106.705 287.710 107.285 ;
        RECT 288.310 106.705 289.720 107.285 ;
        RECT 290.340 106.705 290.510 115.305 ;
        RECT 310.915 114.050 333.665 114.220 ;
        RECT 310.915 109.990 311.085 114.050 ;
        RECT 319.025 113.320 320.275 113.650 ;
        RECT 320.785 113.320 322.035 113.650 ;
        RECT 322.545 113.320 323.795 113.650 ;
        RECT 324.305 113.320 325.555 113.650 ;
        RECT 311.645 110.890 311.815 113.150 ;
        RECT 312.525 110.890 312.695 113.150 ;
        RECT 313.405 110.890 313.575 113.150 ;
        RECT 314.285 110.890 314.455 113.150 ;
        RECT 315.165 110.890 315.335 113.150 ;
        RECT 316.045 110.890 316.215 113.150 ;
        RECT 316.925 110.890 317.095 113.150 ;
        RECT 317.805 110.890 317.975 113.150 ;
        RECT 318.685 110.890 318.855 113.150 ;
        RECT 319.565 110.890 319.735 113.150 ;
        RECT 320.445 110.890 320.615 113.150 ;
        RECT 321.325 110.890 321.495 113.150 ;
        RECT 322.205 110.890 322.375 113.150 ;
        RECT 323.085 110.890 323.255 113.150 ;
        RECT 323.965 110.890 324.135 113.150 ;
        RECT 324.845 110.890 325.015 113.150 ;
        RECT 325.725 110.890 325.895 113.150 ;
        RECT 326.605 110.890 326.775 113.150 ;
        RECT 327.485 110.890 327.655 113.150 ;
        RECT 328.365 110.890 328.535 113.150 ;
        RECT 329.245 110.890 329.415 113.150 ;
        RECT 330.125 110.890 330.295 113.150 ;
        RECT 331.005 110.890 331.175 113.150 ;
        RECT 331.885 110.890 332.055 113.150 ;
        RECT 332.765 110.890 332.935 113.150 ;
        RECT 311.985 110.390 313.235 110.720 ;
        RECT 313.745 110.390 314.995 110.720 ;
        RECT 315.505 110.390 316.755 110.720 ;
        RECT 317.265 110.390 318.515 110.720 ;
        RECT 326.065 110.390 327.315 110.720 ;
        RECT 327.825 110.390 329.075 110.720 ;
        RECT 329.585 110.390 330.835 110.720 ;
        RECT 331.345 110.390 332.595 110.720 ;
        RECT 333.495 109.990 333.665 114.050 ;
        RECT 310.915 109.820 333.665 109.990 ;
        RECT 334.135 114.050 363.925 114.220 ;
        RECT 334.135 109.990 334.305 114.050 ;
        RECT 340.485 113.320 341.735 113.650 ;
        RECT 342.245 113.320 343.495 113.650 ;
        RECT 344.005 113.320 345.255 113.650 ;
        RECT 345.765 113.320 347.015 113.650 ;
        RECT 351.045 113.320 352.295 113.650 ;
        RECT 352.805 113.320 354.055 113.650 ;
        RECT 354.565 113.320 355.815 113.650 ;
        RECT 356.325 113.320 357.575 113.650 ;
        RECT 334.865 110.890 335.035 113.150 ;
        RECT 335.745 110.890 335.915 113.150 ;
        RECT 336.625 110.890 336.795 113.150 ;
        RECT 337.505 110.890 337.675 113.150 ;
        RECT 338.385 110.890 338.555 113.150 ;
        RECT 339.265 110.890 339.435 113.150 ;
        RECT 340.145 110.890 340.315 113.150 ;
        RECT 341.025 110.890 341.195 113.150 ;
        RECT 341.905 110.890 342.075 113.150 ;
        RECT 342.785 110.890 342.955 113.150 ;
        RECT 343.665 110.890 343.835 113.150 ;
        RECT 344.545 110.890 344.715 113.150 ;
        RECT 345.425 110.890 345.595 113.150 ;
        RECT 346.305 110.890 346.475 113.150 ;
        RECT 347.185 110.890 347.355 113.150 ;
        RECT 348.065 110.890 348.235 113.150 ;
        RECT 348.945 110.890 349.115 113.150 ;
        RECT 349.825 110.890 349.995 113.150 ;
        RECT 350.705 110.890 350.875 113.150 ;
        RECT 351.585 110.890 351.755 113.150 ;
        RECT 352.465 110.890 352.635 113.150 ;
        RECT 353.345 110.890 353.515 113.150 ;
        RECT 354.225 110.890 354.395 113.150 ;
        RECT 355.105 110.890 355.275 113.150 ;
        RECT 355.985 110.890 356.155 113.150 ;
        RECT 356.865 110.890 357.035 113.150 ;
        RECT 357.745 110.890 357.915 113.150 ;
        RECT 358.625 110.890 358.795 113.150 ;
        RECT 359.505 110.890 359.675 113.150 ;
        RECT 360.385 110.890 360.555 113.150 ;
        RECT 361.265 110.890 361.435 113.150 ;
        RECT 362.145 110.890 362.315 113.150 ;
        RECT 363.025 110.890 363.195 113.150 ;
        RECT 335.205 110.390 336.455 110.720 ;
        RECT 336.965 110.390 338.215 110.720 ;
        RECT 338.725 110.390 339.975 110.720 ;
        RECT 347.525 110.390 348.775 110.720 ;
        RECT 349.285 110.390 350.535 110.720 ;
        RECT 358.085 110.390 359.335 110.720 ;
        RECT 359.845 110.390 361.095 110.720 ;
        RECT 361.605 110.390 362.855 110.720 ;
        RECT 363.755 109.990 363.925 114.050 ;
        RECT 334.135 109.820 363.925 109.990 ;
        RECT 364.475 114.050 406.580 114.220 ;
        RECT 364.475 109.990 364.645 114.050 ;
        RECT 367.305 113.320 368.555 113.650 ;
        RECT 369.065 113.320 370.315 113.650 ;
        RECT 370.825 113.320 372.075 113.650 ;
        RECT 372.585 113.320 373.835 113.650 ;
        RECT 374.345 113.320 375.595 113.650 ;
        RECT 376.105 113.320 377.355 113.650 ;
        RECT 377.865 113.320 379.115 113.650 ;
        RECT 379.625 113.320 380.875 113.650 ;
        RECT 381.385 113.320 382.635 113.650 ;
        RECT 383.145 113.320 384.395 113.650 ;
        RECT 384.905 113.320 386.155 113.650 ;
        RECT 386.665 113.320 387.915 113.650 ;
        RECT 388.425 113.320 389.675 113.650 ;
        RECT 390.185 113.320 391.435 113.650 ;
        RECT 391.945 113.320 393.195 113.650 ;
        RECT 393.705 113.320 394.955 113.650 ;
        RECT 395.465 113.320 396.715 113.650 ;
        RECT 397.225 113.320 398.475 113.650 ;
        RECT 398.985 113.320 400.235 113.650 ;
        RECT 400.745 113.320 401.995 113.650 ;
        RECT 365.205 110.890 365.375 113.150 ;
        RECT 366.085 110.890 366.255 113.150 ;
        RECT 366.965 110.890 367.135 113.150 ;
        RECT 367.845 110.890 368.015 113.150 ;
        RECT 368.725 110.890 368.895 113.150 ;
        RECT 369.605 110.890 369.775 113.150 ;
        RECT 370.485 110.890 370.655 113.150 ;
        RECT 371.365 110.890 371.535 113.150 ;
        RECT 372.245 110.890 372.415 113.150 ;
        RECT 373.125 110.890 373.295 113.150 ;
        RECT 374.005 110.890 374.175 113.150 ;
        RECT 374.885 110.890 375.055 113.150 ;
        RECT 375.765 110.890 375.935 113.150 ;
        RECT 376.645 110.890 376.815 113.150 ;
        RECT 377.525 110.890 377.695 113.150 ;
        RECT 378.405 110.890 378.575 113.150 ;
        RECT 379.285 110.890 379.455 113.150 ;
        RECT 380.165 110.890 380.335 113.150 ;
        RECT 381.045 110.890 381.215 113.150 ;
        RECT 381.925 110.890 382.095 113.150 ;
        RECT 382.805 110.890 382.975 113.150 ;
        RECT 383.685 110.890 383.855 113.150 ;
        RECT 384.565 110.890 384.735 113.150 ;
        RECT 385.445 110.890 385.615 113.150 ;
        RECT 386.325 110.890 386.495 113.150 ;
        RECT 387.205 110.890 387.375 113.150 ;
        RECT 388.085 110.890 388.255 113.150 ;
        RECT 388.965 110.890 389.135 113.150 ;
        RECT 389.845 110.890 390.015 113.150 ;
        RECT 390.725 110.890 390.895 113.150 ;
        RECT 391.605 110.890 391.775 113.150 ;
        RECT 392.485 110.890 392.655 113.150 ;
        RECT 393.365 110.890 393.535 113.150 ;
        RECT 394.245 110.890 394.415 113.150 ;
        RECT 395.125 110.890 395.295 113.150 ;
        RECT 396.005 110.890 396.175 113.150 ;
        RECT 396.885 110.890 397.055 113.150 ;
        RECT 397.765 110.890 397.935 113.150 ;
        RECT 398.645 110.890 398.815 113.150 ;
        RECT 399.525 110.890 399.695 113.150 ;
        RECT 400.405 110.890 400.575 113.150 ;
        RECT 401.285 110.890 401.455 113.150 ;
        RECT 402.165 110.890 402.335 113.150 ;
        RECT 403.045 110.890 403.215 113.150 ;
        RECT 403.925 110.890 404.095 113.150 ;
        RECT 404.805 110.890 404.975 113.150 ;
        RECT 405.685 110.890 405.855 113.150 ;
        RECT 365.545 110.390 366.795 110.720 ;
        RECT 402.505 110.390 403.755 110.720 ;
        RECT 404.265 110.390 405.515 110.720 ;
        RECT 406.410 109.990 406.580 114.050 ;
        RECT 364.475 109.820 406.580 109.990 ;
        RECT 444.015 109.315 444.305 118.795 ;
        RECT 446.845 118.225 448.095 118.555 ;
        RECT 448.605 118.225 449.855 118.555 ;
        RECT 444.745 110.055 444.915 118.055 ;
        RECT 445.625 110.055 445.795 118.055 ;
        RECT 446.505 110.055 446.675 118.055 ;
        RECT 447.385 110.055 447.555 118.055 ;
        RECT 448.265 110.055 448.435 118.055 ;
        RECT 449.145 110.055 449.315 118.055 ;
        RECT 450.025 110.055 450.195 118.055 ;
        RECT 450.905 110.055 451.075 118.055 ;
        RECT 451.785 110.055 451.955 118.055 ;
        RECT 445.085 109.555 446.335 109.885 ;
        RECT 450.365 109.555 451.615 109.885 ;
        RECT 452.395 109.315 452.685 118.795 ;
        RECT 444.015 109.025 452.685 109.315 ;
        RECT 457.835 118.795 466.505 119.085 ;
        RECT 457.835 109.315 458.125 118.795 ;
        RECT 460.665 118.225 461.915 118.555 ;
        RECT 462.425 118.225 463.675 118.555 ;
        RECT 458.565 110.055 458.735 118.055 ;
        RECT 459.445 110.055 459.615 118.055 ;
        RECT 460.325 110.055 460.495 118.055 ;
        RECT 461.205 110.055 461.375 118.055 ;
        RECT 462.085 110.055 462.255 118.055 ;
        RECT 462.965 110.055 463.135 118.055 ;
        RECT 463.845 110.055 464.015 118.055 ;
        RECT 464.725 110.055 464.895 118.055 ;
        RECT 465.605 110.055 465.775 118.055 ;
        RECT 458.905 109.555 460.155 109.885 ;
        RECT 464.185 109.555 465.435 109.885 ;
        RECT 466.215 109.315 466.505 118.795 ;
        RECT 457.835 109.025 466.505 109.315 ;
        RECT 467.575 118.795 486.265 119.085 ;
        RECT 467.575 109.315 467.865 118.795 ;
        RECT 468.305 110.055 468.475 118.055 ;
        RECT 469.585 110.055 469.755 118.055 ;
        RECT 470.865 110.055 471.035 118.055 ;
        RECT 473.850 110.055 474.020 118.055 ;
        RECT 476.835 110.055 477.005 118.055 ;
        RECT 479.820 110.055 479.990 118.055 ;
        RECT 482.805 110.055 482.975 118.055 ;
        RECT 484.085 110.055 484.255 118.055 ;
        RECT 485.365 110.055 485.535 118.055 ;
        RECT 468.765 109.555 469.295 109.885 ;
        RECT 470.045 109.555 470.575 109.885 ;
        RECT 471.150 109.555 476.720 109.885 ;
        RECT 477.120 109.555 482.690 109.885 ;
        RECT 483.265 109.555 483.795 109.885 ;
        RECT 484.545 109.555 485.075 109.885 ;
        RECT 485.975 109.315 486.265 118.795 ;
        RECT 467.575 109.025 486.265 109.315 ;
        RECT 487.050 118.795 495.720 119.085 ;
        RECT 286.300 105.705 290.510 106.705 ;
        RECT 334.115 108.675 363.945 108.965 ;
        RECT 286.300 105.125 287.710 105.705 ;
        RECT 288.310 105.125 289.720 105.705 ;
        RECT 290.340 104.505 290.510 105.705 ;
        RECT 217.170 104.335 290.510 104.505 ;
        RECT 310.915 105.915 333.665 106.085 ;
        RECT 184.800 104.075 198.350 104.245 ;
        RECT 184.800 102.545 198.350 102.715 ;
        RECT 184.800 100.125 184.970 102.545 ;
        RECT 185.470 101.085 185.640 102.085 ;
        RECT 185.900 101.085 186.070 102.085 ;
        RECT 186.330 101.085 186.500 102.085 ;
        RECT 186.760 101.085 186.930 102.085 ;
        RECT 187.190 101.085 187.360 102.085 ;
        RECT 187.620 101.085 187.790 102.085 ;
        RECT 188.050 101.085 188.220 102.085 ;
        RECT 188.480 101.085 188.650 102.085 ;
        RECT 188.910 101.085 189.080 102.085 ;
        RECT 189.340 101.085 189.510 102.085 ;
        RECT 189.770 101.085 189.940 102.085 ;
        RECT 190.200 101.085 190.370 102.085 ;
        RECT 190.630 101.085 190.800 102.085 ;
        RECT 191.060 101.085 191.230 102.085 ;
        RECT 191.490 101.085 191.660 102.085 ;
        RECT 191.920 101.085 192.090 102.085 ;
        RECT 192.350 101.085 192.520 102.085 ;
        RECT 192.780 101.085 192.950 102.085 ;
        RECT 193.210 101.085 193.380 102.085 ;
        RECT 193.640 101.085 193.810 102.085 ;
        RECT 194.070 101.085 194.240 102.085 ;
        RECT 194.500 101.085 194.670 102.085 ;
        RECT 194.930 101.085 195.100 102.085 ;
        RECT 195.360 101.085 195.530 102.085 ;
        RECT 195.790 101.085 195.960 102.085 ;
        RECT 196.220 101.085 196.390 102.085 ;
        RECT 196.650 101.085 196.820 102.085 ;
        RECT 197.080 101.085 197.250 102.085 ;
        RECT 197.510 101.085 197.680 102.085 ;
        RECT 185.695 100.645 186.275 100.875 ;
        RECT 186.555 100.645 196.595 100.875 ;
        RECT 196.875 100.645 197.455 100.875 ;
        RECT 198.180 100.125 198.350 102.545 ;
        RECT 217.170 102.285 290.510 102.455 ;
        RECT 217.170 101.085 217.340 102.285 ;
        RECT 217.960 101.085 219.370 101.665 ;
        RECT 219.970 101.085 221.380 101.665 ;
        RECT 199.880 100.525 213.430 100.695 ;
        RECT 184.800 97.230 184.970 99.620 ;
        RECT 185.695 98.870 189.715 99.100 ;
        RECT 189.995 98.870 193.155 99.100 ;
        RECT 193.435 98.870 197.455 99.100 ;
        RECT 185.470 97.660 185.640 98.660 ;
        RECT 185.900 97.660 186.070 98.660 ;
        RECT 186.330 97.660 186.500 98.660 ;
        RECT 186.760 97.660 186.930 98.660 ;
        RECT 187.190 97.660 187.360 98.660 ;
        RECT 187.620 97.660 187.790 98.660 ;
        RECT 188.050 97.660 188.220 98.660 ;
        RECT 188.480 97.660 188.650 98.660 ;
        RECT 188.910 97.660 189.080 98.660 ;
        RECT 189.340 97.660 189.510 98.660 ;
        RECT 189.770 97.660 189.940 98.660 ;
        RECT 190.200 97.660 190.370 98.660 ;
        RECT 190.630 97.660 190.800 98.660 ;
        RECT 191.060 97.660 191.230 98.660 ;
        RECT 191.490 97.660 191.660 98.660 ;
        RECT 191.920 97.660 192.090 98.660 ;
        RECT 192.350 97.660 192.520 98.660 ;
        RECT 192.780 97.660 192.950 98.660 ;
        RECT 193.210 97.660 193.380 98.660 ;
        RECT 193.640 97.660 193.810 98.660 ;
        RECT 194.070 97.660 194.240 98.660 ;
        RECT 194.500 97.660 194.670 98.660 ;
        RECT 194.930 97.660 195.100 98.660 ;
        RECT 195.360 97.660 195.530 98.660 ;
        RECT 195.790 97.660 195.960 98.660 ;
        RECT 196.220 97.660 196.390 98.660 ;
        RECT 196.650 97.660 196.820 98.660 ;
        RECT 197.080 97.660 197.250 98.660 ;
        RECT 197.510 97.660 197.680 98.660 ;
        RECT 198.180 97.230 198.350 99.620 ;
        RECT 199.880 97.435 200.050 100.525 ;
        RECT 204.635 100.135 204.805 100.195 ;
        RECT 208.505 100.135 208.675 100.195 ;
        RECT 200.775 99.905 204.835 100.135 ;
        RECT 208.475 99.905 212.535 100.135 ;
        RECT 204.635 99.865 204.805 99.905 ;
        RECT 208.505 99.865 208.675 99.905 ;
        RECT 200.550 98.695 200.720 99.695 ;
        RECT 200.980 98.695 201.150 99.695 ;
        RECT 201.410 98.695 201.580 99.695 ;
        RECT 201.840 98.695 202.010 99.695 ;
        RECT 202.270 98.695 202.440 99.695 ;
        RECT 202.700 98.695 202.870 99.695 ;
        RECT 203.130 98.695 203.300 99.695 ;
        RECT 203.560 98.695 203.730 99.695 ;
        RECT 203.990 98.695 204.160 99.695 ;
        RECT 204.420 98.695 204.590 99.695 ;
        RECT 204.850 98.695 205.020 99.695 ;
        RECT 205.280 98.695 205.450 99.695 ;
        RECT 205.710 98.695 205.880 99.695 ;
        RECT 206.140 98.695 206.310 99.695 ;
        RECT 206.570 98.695 206.740 99.695 ;
        RECT 207.000 98.695 207.170 99.695 ;
        RECT 207.430 98.695 207.600 99.695 ;
        RECT 207.860 98.695 208.030 99.695 ;
        RECT 208.290 98.695 208.460 99.695 ;
        RECT 208.720 98.695 208.890 99.695 ;
        RECT 209.150 98.695 209.320 99.695 ;
        RECT 209.580 98.695 209.750 99.695 ;
        RECT 210.010 98.695 210.180 99.695 ;
        RECT 210.440 98.695 210.610 99.695 ;
        RECT 210.870 98.695 211.040 99.695 ;
        RECT 211.300 98.695 211.470 99.695 ;
        RECT 211.730 98.695 211.900 99.695 ;
        RECT 212.160 98.695 212.330 99.695 ;
        RECT 212.590 98.695 212.760 99.695 ;
        RECT 205.075 98.255 208.235 98.485 ;
        RECT 213.260 97.435 213.430 100.525 ;
        RECT 217.170 100.085 221.380 101.085 ;
        RECT 184.800 97.060 198.350 97.230 ;
        RECT 184.800 94.670 184.970 97.060 ;
        RECT 185.470 95.630 185.640 96.630 ;
        RECT 185.900 95.630 186.070 96.630 ;
        RECT 186.330 95.630 186.500 96.630 ;
        RECT 186.760 95.630 186.930 96.630 ;
        RECT 187.190 95.630 187.360 96.630 ;
        RECT 187.620 95.630 187.790 96.630 ;
        RECT 188.050 95.630 188.220 96.630 ;
        RECT 188.480 95.630 188.650 96.630 ;
        RECT 188.910 95.630 189.080 96.630 ;
        RECT 189.340 95.630 189.510 96.630 ;
        RECT 189.770 95.630 189.940 96.630 ;
        RECT 190.200 95.630 190.370 96.630 ;
        RECT 190.630 95.630 190.800 96.630 ;
        RECT 191.060 95.630 191.230 96.630 ;
        RECT 191.490 95.630 191.660 96.630 ;
        RECT 191.920 95.630 192.090 96.630 ;
        RECT 192.350 95.630 192.520 96.630 ;
        RECT 192.780 95.630 192.950 96.630 ;
        RECT 193.210 95.630 193.380 96.630 ;
        RECT 193.640 95.630 193.810 96.630 ;
        RECT 194.070 95.630 194.240 96.630 ;
        RECT 194.500 95.630 194.670 96.630 ;
        RECT 194.930 95.630 195.100 96.630 ;
        RECT 195.360 95.630 195.530 96.630 ;
        RECT 195.790 95.630 195.960 96.630 ;
        RECT 196.220 95.630 196.390 96.630 ;
        RECT 196.650 95.630 196.820 96.630 ;
        RECT 197.080 95.630 197.250 96.630 ;
        RECT 197.510 95.630 197.680 96.630 ;
        RECT 185.695 95.190 189.715 95.420 ;
        RECT 189.995 95.190 193.155 95.420 ;
        RECT 193.435 95.190 197.455 95.420 ;
        RECT 198.180 94.670 198.350 97.060 ;
        RECT 184.800 91.745 184.970 94.165 ;
        RECT 185.695 93.415 186.275 93.645 ;
        RECT 186.555 93.415 196.595 93.645 ;
        RECT 196.875 93.415 197.455 93.645 ;
        RECT 185.470 92.205 185.640 93.205 ;
        RECT 185.900 92.205 186.070 93.205 ;
        RECT 186.330 92.205 186.500 93.205 ;
        RECT 186.760 92.205 186.930 93.205 ;
        RECT 187.190 92.205 187.360 93.205 ;
        RECT 187.620 92.205 187.790 93.205 ;
        RECT 188.050 92.205 188.220 93.205 ;
        RECT 188.480 92.205 188.650 93.205 ;
        RECT 188.910 92.205 189.080 93.205 ;
        RECT 189.340 92.205 189.510 93.205 ;
        RECT 189.770 92.205 189.940 93.205 ;
        RECT 190.200 92.205 190.370 93.205 ;
        RECT 190.630 92.205 190.800 93.205 ;
        RECT 191.060 92.205 191.230 93.205 ;
        RECT 191.490 92.205 191.660 93.205 ;
        RECT 191.920 92.205 192.090 93.205 ;
        RECT 192.350 92.205 192.520 93.205 ;
        RECT 192.780 92.205 192.950 93.205 ;
        RECT 193.210 92.205 193.380 93.205 ;
        RECT 193.640 92.205 193.810 93.205 ;
        RECT 194.070 92.205 194.240 93.205 ;
        RECT 194.500 92.205 194.670 93.205 ;
        RECT 194.930 92.205 195.100 93.205 ;
        RECT 195.360 92.205 195.530 93.205 ;
        RECT 195.790 92.205 195.960 93.205 ;
        RECT 196.220 92.205 196.390 93.205 ;
        RECT 196.650 92.205 196.820 93.205 ;
        RECT 197.080 92.205 197.250 93.205 ;
        RECT 197.510 92.205 197.680 93.205 ;
        RECT 198.180 91.745 198.350 94.165 ;
        RECT 199.880 93.605 200.050 96.555 ;
        RECT 201.635 95.805 211.675 96.035 ;
        RECT 200.550 94.595 200.720 95.595 ;
        RECT 200.980 94.595 201.150 95.595 ;
        RECT 201.410 94.595 201.580 95.595 ;
        RECT 201.840 94.595 202.010 95.595 ;
        RECT 202.270 94.595 202.440 95.595 ;
        RECT 202.700 94.595 202.870 95.595 ;
        RECT 203.130 94.595 203.300 95.595 ;
        RECT 203.560 94.595 203.730 95.595 ;
        RECT 203.990 94.595 204.160 95.595 ;
        RECT 204.420 94.595 204.590 95.595 ;
        RECT 204.850 94.595 205.020 95.595 ;
        RECT 205.280 94.595 205.450 95.595 ;
        RECT 205.710 94.595 205.880 95.595 ;
        RECT 206.140 94.595 206.310 95.595 ;
        RECT 206.570 94.595 206.740 95.595 ;
        RECT 207.000 94.595 207.170 95.595 ;
        RECT 207.430 94.595 207.600 95.595 ;
        RECT 207.860 94.595 208.030 95.595 ;
        RECT 208.290 94.595 208.460 95.595 ;
        RECT 208.720 94.595 208.890 95.595 ;
        RECT 209.150 94.595 209.320 95.595 ;
        RECT 209.580 94.595 209.750 95.595 ;
        RECT 210.010 94.595 210.180 95.595 ;
        RECT 210.440 94.595 210.610 95.595 ;
        RECT 210.870 94.595 211.040 95.595 ;
        RECT 211.300 94.595 211.470 95.595 ;
        RECT 211.730 94.595 211.900 95.595 ;
        RECT 212.160 94.595 212.330 95.595 ;
        RECT 212.590 94.595 212.760 95.595 ;
        RECT 200.800 94.095 201.330 94.425 ;
        RECT 211.980 94.095 212.510 94.425 ;
        RECT 213.260 93.605 213.430 96.555 ;
        RECT 199.880 93.435 213.430 93.605 ;
        RECT 184.800 91.575 198.350 91.745 ;
        RECT 217.170 91.485 217.340 100.085 ;
        RECT 217.960 99.505 219.370 100.085 ;
        RECT 219.970 99.505 221.380 100.085 ;
        RECT 221.980 99.505 223.390 101.665 ;
        RECT 223.990 99.505 225.400 101.665 ;
        RECT 226.000 99.505 227.410 101.665 ;
        RECT 228.010 99.505 229.420 101.665 ;
        RECT 230.020 99.505 231.430 101.665 ;
        RECT 232.030 99.505 233.440 101.665 ;
        RECT 234.040 99.505 235.450 101.665 ;
        RECT 236.050 99.505 237.460 101.665 ;
        RECT 238.060 99.505 239.470 101.665 ;
        RECT 240.070 99.505 241.480 101.665 ;
        RECT 242.080 99.505 243.490 101.665 ;
        RECT 244.090 99.505 245.500 101.665 ;
        RECT 246.100 99.505 247.510 101.665 ;
        RECT 248.110 99.505 249.520 101.665 ;
        RECT 250.120 99.505 251.530 101.665 ;
        RECT 252.130 99.505 253.540 101.665 ;
        RECT 254.140 99.505 255.550 101.665 ;
        RECT 256.150 99.505 257.560 101.665 ;
        RECT 258.160 99.505 259.570 101.665 ;
        RECT 260.170 99.505 261.580 101.665 ;
        RECT 262.180 99.505 263.590 101.665 ;
        RECT 264.190 99.505 265.600 101.665 ;
        RECT 266.200 99.505 267.610 101.665 ;
        RECT 268.210 99.505 269.620 101.665 ;
        RECT 270.220 99.505 271.630 101.665 ;
        RECT 272.230 99.505 273.640 101.665 ;
        RECT 274.240 99.505 275.650 101.665 ;
        RECT 276.250 99.505 277.660 101.665 ;
        RECT 278.260 99.505 279.670 101.665 ;
        RECT 280.270 99.505 281.680 101.665 ;
        RECT 282.280 99.505 283.690 101.665 ;
        RECT 284.290 99.505 285.700 101.665 ;
        RECT 286.300 101.085 287.710 101.665 ;
        RECT 288.310 101.085 289.720 101.665 ;
        RECT 290.340 101.085 290.510 102.285 ;
        RECT 286.300 100.085 290.510 101.085 ;
        RECT 310.915 100.910 311.085 105.915 ;
        RECT 311.985 104.710 313.235 105.040 ;
        RECT 313.745 104.710 314.995 105.040 ;
        RECT 317.265 104.710 318.515 105.040 ;
        RECT 320.785 104.710 322.035 105.040 ;
        RECT 324.305 104.710 325.555 105.040 ;
        RECT 327.825 104.710 329.075 105.040 ;
        RECT 329.585 104.710 330.835 105.040 ;
        RECT 331.345 104.710 332.595 105.040 ;
        RECT 311.645 102.280 311.815 104.540 ;
        RECT 312.525 102.280 312.695 104.540 ;
        RECT 313.405 102.280 313.575 104.540 ;
        RECT 314.285 102.280 314.455 104.540 ;
        RECT 315.165 102.280 315.335 104.540 ;
        RECT 316.045 102.280 316.215 104.540 ;
        RECT 316.925 102.280 317.095 104.540 ;
        RECT 317.805 102.280 317.975 104.540 ;
        RECT 318.685 102.280 318.855 104.540 ;
        RECT 319.565 102.280 319.735 104.540 ;
        RECT 320.445 102.280 320.615 104.540 ;
        RECT 321.325 102.280 321.495 104.540 ;
        RECT 322.205 102.280 322.375 104.540 ;
        RECT 323.085 102.280 323.255 104.540 ;
        RECT 323.965 102.280 324.135 104.540 ;
        RECT 324.845 102.280 325.015 104.540 ;
        RECT 325.725 102.280 325.895 104.540 ;
        RECT 326.605 102.280 326.775 104.540 ;
        RECT 327.485 102.280 327.655 104.540 ;
        RECT 328.365 102.280 328.535 104.540 ;
        RECT 329.245 102.280 329.415 104.540 ;
        RECT 330.125 102.280 330.295 104.540 ;
        RECT 331.005 102.280 331.175 104.540 ;
        RECT 331.885 102.280 332.055 104.540 ;
        RECT 332.765 102.280 332.935 104.540 ;
        RECT 311.985 101.780 313.235 102.110 ;
        RECT 313.745 101.780 314.995 102.110 ;
        RECT 315.505 101.780 316.755 102.110 ;
        RECT 319.025 101.780 320.275 102.110 ;
        RECT 322.545 101.780 323.795 102.110 ;
        RECT 326.065 101.780 327.315 102.110 ;
        RECT 329.585 101.780 330.835 102.110 ;
        RECT 331.345 101.780 332.595 102.110 ;
        RECT 333.495 100.910 333.665 105.915 ;
        RECT 310.915 100.740 333.665 100.910 ;
        RECT 286.300 99.505 287.710 100.085 ;
        RECT 288.310 99.505 289.720 100.085 ;
        RECT 217.960 91.485 219.370 92.065 ;
        RECT 219.970 91.485 221.380 92.065 ;
        RECT 217.170 90.485 221.380 91.485 ;
        RECT 217.170 89.285 217.340 90.485 ;
        RECT 217.960 89.905 219.370 90.485 ;
        RECT 219.970 89.905 221.380 90.485 ;
        RECT 221.980 89.905 223.390 92.065 ;
        RECT 223.990 89.905 225.400 92.065 ;
        RECT 226.000 89.905 227.410 92.065 ;
        RECT 228.010 89.905 229.420 92.065 ;
        RECT 230.020 89.905 231.430 92.065 ;
        RECT 232.030 89.905 233.440 92.065 ;
        RECT 234.040 89.905 235.450 92.065 ;
        RECT 236.050 89.905 237.460 92.065 ;
        RECT 238.060 89.905 239.470 92.065 ;
        RECT 240.070 89.905 241.480 92.065 ;
        RECT 242.080 89.905 243.490 92.065 ;
        RECT 244.090 89.905 245.500 92.065 ;
        RECT 246.100 89.905 247.510 92.065 ;
        RECT 248.110 89.905 249.520 92.065 ;
        RECT 250.120 89.905 251.530 92.065 ;
        RECT 252.130 89.905 253.540 92.065 ;
        RECT 254.140 89.905 255.550 92.065 ;
        RECT 256.150 89.905 257.560 92.065 ;
        RECT 258.160 89.905 259.570 92.065 ;
        RECT 260.170 89.905 261.580 92.065 ;
        RECT 262.180 89.905 263.590 92.065 ;
        RECT 264.190 89.905 265.600 92.065 ;
        RECT 266.200 89.905 267.610 92.065 ;
        RECT 268.210 89.905 269.620 92.065 ;
        RECT 270.220 89.905 271.630 92.065 ;
        RECT 272.230 89.905 273.640 92.065 ;
        RECT 274.240 89.905 275.650 92.065 ;
        RECT 276.250 89.905 277.660 92.065 ;
        RECT 278.260 89.905 279.670 92.065 ;
        RECT 280.270 89.905 281.680 92.065 ;
        RECT 282.280 89.905 283.690 92.065 ;
        RECT 284.290 89.905 285.700 92.065 ;
        RECT 286.300 91.485 287.710 92.065 ;
        RECT 288.310 91.485 289.720 92.065 ;
        RECT 290.340 91.485 290.510 100.085 ;
        RECT 334.115 98.125 334.405 108.675 ;
        RECT 340.485 108.085 341.735 108.415 ;
        RECT 342.245 108.085 343.495 108.415 ;
        RECT 344.005 108.085 345.255 108.415 ;
        RECT 345.765 108.085 347.015 108.415 ;
        RECT 351.045 108.085 352.295 108.415 ;
        RECT 352.805 108.085 354.055 108.415 ;
        RECT 354.565 108.085 355.815 108.415 ;
        RECT 356.325 108.085 357.575 108.415 ;
        RECT 334.865 98.885 335.035 107.915 ;
        RECT 335.745 98.885 335.915 107.915 ;
        RECT 336.625 98.885 336.795 107.915 ;
        RECT 337.505 98.885 337.675 107.915 ;
        RECT 338.385 98.885 338.555 107.915 ;
        RECT 339.265 98.885 339.435 107.915 ;
        RECT 340.145 98.885 340.315 107.915 ;
        RECT 341.025 98.885 341.195 107.915 ;
        RECT 341.905 98.885 342.075 107.915 ;
        RECT 342.785 98.885 342.955 107.915 ;
        RECT 343.665 98.885 343.835 107.915 ;
        RECT 344.545 98.885 344.715 107.915 ;
        RECT 345.425 98.885 345.595 107.915 ;
        RECT 346.305 98.885 346.475 107.915 ;
        RECT 347.185 98.885 347.355 107.915 ;
        RECT 348.065 98.885 348.235 107.915 ;
        RECT 348.945 98.885 349.115 107.915 ;
        RECT 349.825 98.885 349.995 107.915 ;
        RECT 350.705 98.885 350.875 107.915 ;
        RECT 351.585 98.885 351.755 107.915 ;
        RECT 352.465 98.885 352.635 107.915 ;
        RECT 353.345 98.885 353.515 107.915 ;
        RECT 354.225 98.885 354.395 107.915 ;
        RECT 355.105 98.885 355.275 107.915 ;
        RECT 355.985 98.885 356.155 107.915 ;
        RECT 356.865 98.885 357.035 107.915 ;
        RECT 357.745 98.885 357.915 107.915 ;
        RECT 358.625 98.885 358.795 107.915 ;
        RECT 359.505 98.885 359.675 107.915 ;
        RECT 360.385 98.885 360.555 107.915 ;
        RECT 361.265 98.885 361.435 107.915 ;
        RECT 362.145 98.885 362.315 107.915 ;
        RECT 363.025 98.885 363.195 107.915 ;
        RECT 335.205 98.385 336.455 98.715 ;
        RECT 336.965 98.385 338.215 98.715 ;
        RECT 338.725 98.385 339.975 98.715 ;
        RECT 347.525 98.385 348.775 98.715 ;
        RECT 349.285 98.385 350.535 98.715 ;
        RECT 358.085 98.385 359.335 98.715 ;
        RECT 359.845 98.385 361.095 98.715 ;
        RECT 361.605 98.385 362.855 98.715 ;
        RECT 363.655 98.125 363.945 108.675 ;
        RECT 334.115 97.835 363.945 98.125 ;
        RECT 364.455 108.675 406.605 108.965 ;
        RECT 364.455 98.125 364.745 108.675 ;
        RECT 367.305 108.085 368.555 108.415 ;
        RECT 369.065 108.085 370.315 108.415 ;
        RECT 370.825 108.085 372.075 108.415 ;
        RECT 372.585 108.085 373.835 108.415 ;
        RECT 374.345 108.085 375.595 108.415 ;
        RECT 376.105 108.085 377.355 108.415 ;
        RECT 377.865 108.085 379.115 108.415 ;
        RECT 379.625 108.085 380.875 108.415 ;
        RECT 381.385 108.085 382.635 108.415 ;
        RECT 383.145 108.085 384.395 108.415 ;
        RECT 384.905 108.085 386.155 108.415 ;
        RECT 386.665 108.085 387.915 108.415 ;
        RECT 388.425 108.085 389.675 108.415 ;
        RECT 390.185 108.085 391.435 108.415 ;
        RECT 391.945 108.085 393.195 108.415 ;
        RECT 393.705 108.085 394.955 108.415 ;
        RECT 395.465 108.085 396.715 108.415 ;
        RECT 397.225 108.085 398.475 108.415 ;
        RECT 398.985 108.085 400.235 108.415 ;
        RECT 400.745 108.085 401.995 108.415 ;
        RECT 365.205 98.885 365.375 107.915 ;
        RECT 366.085 98.885 366.255 107.915 ;
        RECT 366.965 98.885 367.135 107.915 ;
        RECT 367.845 98.885 368.015 107.915 ;
        RECT 368.725 98.885 368.895 107.915 ;
        RECT 369.605 98.885 369.775 107.915 ;
        RECT 370.485 98.885 370.655 107.915 ;
        RECT 371.365 98.885 371.535 107.915 ;
        RECT 372.245 98.885 372.415 107.915 ;
        RECT 373.125 98.885 373.295 107.915 ;
        RECT 374.005 98.885 374.175 107.915 ;
        RECT 374.885 98.885 375.055 107.915 ;
        RECT 375.765 98.885 375.935 107.915 ;
        RECT 376.645 98.885 376.815 107.915 ;
        RECT 377.525 98.885 377.695 107.915 ;
        RECT 378.405 98.885 378.575 107.915 ;
        RECT 379.285 98.885 379.455 107.915 ;
        RECT 380.165 98.885 380.335 107.915 ;
        RECT 381.045 98.885 381.215 107.915 ;
        RECT 381.925 98.885 382.095 107.915 ;
        RECT 382.805 98.885 382.975 107.915 ;
        RECT 383.685 98.885 383.855 107.915 ;
        RECT 384.565 98.885 384.735 107.915 ;
        RECT 385.445 98.885 385.615 107.915 ;
        RECT 386.325 98.885 386.495 107.915 ;
        RECT 387.205 98.885 387.375 107.915 ;
        RECT 388.085 98.885 388.255 107.915 ;
        RECT 388.965 98.885 389.135 107.915 ;
        RECT 389.845 98.885 390.015 107.915 ;
        RECT 390.725 98.885 390.895 107.915 ;
        RECT 391.605 98.885 391.775 107.915 ;
        RECT 392.485 98.885 392.655 107.915 ;
        RECT 393.365 98.885 393.535 107.915 ;
        RECT 394.245 98.885 394.415 107.915 ;
        RECT 395.125 98.885 395.295 107.915 ;
        RECT 396.005 98.885 396.175 107.915 ;
        RECT 396.885 98.885 397.055 107.915 ;
        RECT 397.765 98.885 397.935 107.915 ;
        RECT 398.645 98.885 398.815 107.915 ;
        RECT 399.525 98.885 399.695 107.915 ;
        RECT 400.405 98.885 400.575 107.915 ;
        RECT 401.285 98.885 401.455 107.915 ;
        RECT 402.165 98.885 402.335 107.915 ;
        RECT 403.045 98.885 403.215 107.915 ;
        RECT 403.925 98.885 404.095 107.915 ;
        RECT 404.805 98.885 404.975 107.915 ;
        RECT 405.685 98.885 405.855 107.915 ;
        RECT 365.545 98.385 366.795 98.715 ;
        RECT 402.505 98.385 403.755 98.715 ;
        RECT 404.265 98.385 405.515 98.715 ;
        RECT 406.315 98.125 406.605 108.675 ;
        RECT 487.050 108.285 487.340 118.795 ;
        RECT 489.880 118.225 491.130 118.555 ;
        RECT 491.640 118.225 492.890 118.555 ;
        RECT 487.780 109.025 487.950 118.055 ;
        RECT 488.660 109.025 488.830 118.055 ;
        RECT 489.540 109.025 489.710 118.055 ;
        RECT 490.420 109.025 490.590 118.055 ;
        RECT 491.300 109.025 491.470 118.055 ;
        RECT 492.180 109.025 492.350 118.055 ;
        RECT 493.060 109.025 493.230 118.055 ;
        RECT 493.940 109.025 494.110 118.055 ;
        RECT 494.820 109.025 494.990 118.055 ;
        RECT 488.120 108.525 489.370 108.855 ;
        RECT 493.400 108.525 494.650 108.855 ;
        RECT 495.430 108.285 495.720 118.795 ;
        RECT 496.780 118.795 505.450 119.085 ;
        RECT 496.780 109.315 497.070 118.795 ;
        RECT 497.510 110.055 497.680 118.055 ;
        RECT 498.390 110.055 498.560 118.055 ;
        RECT 499.270 110.055 499.440 118.055 ;
        RECT 500.150 110.055 500.320 118.055 ;
        RECT 501.030 110.055 501.200 118.055 ;
        RECT 501.910 110.055 502.080 118.055 ;
        RECT 502.790 110.055 502.960 118.055 ;
        RECT 503.670 110.055 503.840 118.055 ;
        RECT 504.550 110.055 504.720 118.055 ;
        RECT 497.850 109.555 499.100 109.885 ;
        RECT 499.610 109.555 500.860 109.885 ;
        RECT 501.370 109.555 502.620 109.885 ;
        RECT 503.130 109.555 504.380 109.885 ;
        RECT 505.160 109.315 505.450 118.795 ;
        RECT 496.780 109.025 505.450 109.315 ;
        RECT 487.050 107.995 495.720 108.285 ;
        RECT 364.455 97.835 406.605 98.125 ;
        RECT 487.050 105.530 495.720 105.820 ;
        RECT 472.625 97.085 481.215 97.375 ;
        RECT 286.300 90.485 290.510 91.485 ;
        RECT 286.300 89.905 287.710 90.485 ;
        RECT 288.310 89.905 289.720 90.485 ;
        RECT 290.340 89.285 290.510 90.485 ;
        RECT 217.170 89.115 290.510 89.285 ;
        RECT 334.115 96.310 363.945 96.600 ;
        RECT 334.115 85.760 334.405 96.310 ;
        RECT 335.205 95.720 336.455 96.050 ;
        RECT 336.965 95.720 338.215 96.050 ;
        RECT 359.845 95.720 361.095 96.050 ;
        RECT 361.605 95.720 362.855 96.050 ;
        RECT 334.865 86.520 335.035 95.550 ;
        RECT 335.745 86.520 335.915 95.550 ;
        RECT 336.625 86.520 336.795 95.550 ;
        RECT 337.505 86.520 337.675 95.550 ;
        RECT 338.385 86.520 338.555 95.550 ;
        RECT 339.265 86.520 339.435 95.550 ;
        RECT 340.145 86.520 340.315 95.550 ;
        RECT 341.025 86.520 341.195 95.550 ;
        RECT 341.905 86.520 342.075 95.550 ;
        RECT 342.785 86.520 342.955 95.550 ;
        RECT 343.665 86.520 343.835 95.550 ;
        RECT 344.545 86.520 344.715 95.550 ;
        RECT 345.425 86.520 345.595 95.550 ;
        RECT 346.305 86.520 346.475 95.550 ;
        RECT 347.185 86.520 347.355 95.550 ;
        RECT 348.065 86.520 348.235 95.550 ;
        RECT 348.945 86.520 349.115 95.550 ;
        RECT 349.825 86.520 349.995 95.550 ;
        RECT 350.705 86.520 350.875 95.550 ;
        RECT 351.585 86.520 351.755 95.550 ;
        RECT 352.465 86.520 352.635 95.550 ;
        RECT 353.345 86.520 353.515 95.550 ;
        RECT 354.225 86.520 354.395 95.550 ;
        RECT 355.105 86.520 355.275 95.550 ;
        RECT 355.985 86.520 356.155 95.550 ;
        RECT 356.865 86.520 357.035 95.550 ;
        RECT 357.745 86.520 357.915 95.550 ;
        RECT 358.625 86.520 358.795 95.550 ;
        RECT 359.505 86.520 359.675 95.550 ;
        RECT 360.385 86.520 360.555 95.550 ;
        RECT 361.265 86.520 361.435 95.550 ;
        RECT 362.145 86.520 362.315 95.550 ;
        RECT 363.025 86.520 363.195 95.550 ;
        RECT 338.725 86.020 339.975 86.350 ;
        RECT 340.485 86.020 341.735 86.350 ;
        RECT 342.245 86.020 343.495 86.350 ;
        RECT 344.005 86.020 345.255 86.350 ;
        RECT 345.765 86.020 347.015 86.350 ;
        RECT 347.525 86.020 348.775 86.350 ;
        RECT 349.285 86.020 350.535 86.350 ;
        RECT 351.045 86.020 352.295 86.350 ;
        RECT 352.805 86.020 354.055 86.350 ;
        RECT 354.565 86.020 355.815 86.350 ;
        RECT 356.325 86.020 357.575 86.350 ;
        RECT 358.085 86.020 359.335 86.350 ;
        RECT 363.655 85.760 363.945 96.310 ;
        RECT 334.115 85.470 363.945 85.760 ;
        RECT 364.455 96.310 406.605 96.600 ;
        RECT 364.455 85.760 364.745 96.310 ;
        RECT 365.545 95.720 366.795 96.050 ;
        RECT 402.505 95.720 403.755 96.050 ;
        RECT 404.265 95.720 405.515 96.050 ;
        RECT 365.205 86.520 365.375 95.550 ;
        RECT 366.085 86.520 366.255 95.550 ;
        RECT 366.965 86.520 367.135 95.550 ;
        RECT 367.845 86.520 368.015 95.550 ;
        RECT 368.725 86.520 368.895 95.550 ;
        RECT 369.605 86.520 369.775 95.550 ;
        RECT 370.485 86.520 370.655 95.550 ;
        RECT 371.365 86.520 371.535 95.550 ;
        RECT 372.245 86.520 372.415 95.550 ;
        RECT 373.125 86.520 373.295 95.550 ;
        RECT 374.005 86.520 374.175 95.550 ;
        RECT 374.885 86.520 375.055 95.550 ;
        RECT 375.765 86.520 375.935 95.550 ;
        RECT 376.645 86.520 376.815 95.550 ;
        RECT 377.525 86.520 377.695 95.550 ;
        RECT 378.405 86.520 378.575 95.550 ;
        RECT 379.285 86.520 379.455 95.550 ;
        RECT 380.165 86.520 380.335 95.550 ;
        RECT 381.045 86.520 381.215 95.550 ;
        RECT 381.925 86.520 382.095 95.550 ;
        RECT 382.805 86.520 382.975 95.550 ;
        RECT 383.685 86.520 383.855 95.550 ;
        RECT 384.565 86.520 384.735 95.550 ;
        RECT 385.445 86.520 385.615 95.550 ;
        RECT 386.325 86.520 386.495 95.550 ;
        RECT 387.205 86.520 387.375 95.550 ;
        RECT 388.085 86.520 388.255 95.550 ;
        RECT 388.965 86.520 389.135 95.550 ;
        RECT 389.845 86.520 390.015 95.550 ;
        RECT 390.725 86.520 390.895 95.550 ;
        RECT 391.605 86.520 391.775 95.550 ;
        RECT 392.485 86.520 392.655 95.550 ;
        RECT 393.365 86.520 393.535 95.550 ;
        RECT 394.245 86.520 394.415 95.550 ;
        RECT 395.125 86.520 395.295 95.550 ;
        RECT 396.005 86.520 396.175 95.550 ;
        RECT 396.885 86.520 397.055 95.550 ;
        RECT 397.765 86.520 397.935 95.550 ;
        RECT 398.645 86.520 398.815 95.550 ;
        RECT 399.525 86.520 399.695 95.550 ;
        RECT 400.405 86.520 400.575 95.550 ;
        RECT 401.285 86.520 401.455 95.550 ;
        RECT 402.165 86.520 402.335 95.550 ;
        RECT 403.045 86.520 403.215 95.550 ;
        RECT 403.925 86.520 404.095 95.550 ;
        RECT 404.805 86.520 404.975 95.550 ;
        RECT 405.685 86.520 405.855 95.550 ;
        RECT 367.305 86.020 368.555 86.350 ;
        RECT 369.065 86.020 370.315 86.350 ;
        RECT 370.825 86.020 372.075 86.350 ;
        RECT 372.585 86.020 373.835 86.350 ;
        RECT 374.345 86.020 375.595 86.350 ;
        RECT 376.105 86.020 377.355 86.350 ;
        RECT 377.865 86.020 379.115 86.350 ;
        RECT 379.625 86.020 380.875 86.350 ;
        RECT 381.385 86.020 382.635 86.350 ;
        RECT 383.145 86.020 384.395 86.350 ;
        RECT 384.905 86.020 386.155 86.350 ;
        RECT 386.665 86.020 387.915 86.350 ;
        RECT 388.425 86.020 389.675 86.350 ;
        RECT 390.185 86.020 391.435 86.350 ;
        RECT 391.945 86.020 393.195 86.350 ;
        RECT 393.705 86.020 394.955 86.350 ;
        RECT 395.465 86.020 396.715 86.350 ;
        RECT 397.225 86.020 398.475 86.350 ;
        RECT 398.985 86.020 400.235 86.350 ;
        RECT 400.745 86.020 401.995 86.350 ;
        RECT 406.315 85.760 406.605 96.310 ;
        RECT 453.275 94.115 471.065 94.405 ;
        RECT 434.835 91.445 443.425 91.735 ;
        RECT 434.835 87.965 435.125 91.445 ;
        RECT 435.865 90.875 437.115 91.205 ;
        RECT 441.145 90.875 442.395 91.205 ;
        RECT 435.525 88.705 435.695 90.705 ;
        RECT 436.405 88.705 436.575 90.705 ;
        RECT 437.285 88.705 437.455 90.705 ;
        RECT 438.165 88.705 438.335 90.705 ;
        RECT 439.045 88.705 439.215 90.705 ;
        RECT 439.925 88.705 440.095 90.705 ;
        RECT 440.805 88.705 440.975 90.705 ;
        RECT 441.685 88.705 441.855 90.705 ;
        RECT 442.565 88.705 442.735 90.705 ;
        RECT 437.625 88.205 438.875 88.535 ;
        RECT 439.385 88.205 440.635 88.535 ;
        RECT 443.135 87.965 443.425 91.445 ;
        RECT 434.835 87.675 443.425 87.965 ;
        RECT 444.055 91.445 452.645 91.735 ;
        RECT 444.055 87.960 444.345 91.445 ;
        RECT 445.085 90.865 446.335 91.195 ;
        RECT 450.365 90.865 451.615 91.195 ;
        RECT 444.745 88.705 444.915 90.695 ;
        RECT 445.625 88.705 445.795 90.695 ;
        RECT 446.505 88.705 446.675 90.695 ;
        RECT 447.385 88.705 447.555 90.695 ;
        RECT 448.265 88.705 448.435 90.695 ;
        RECT 449.145 88.705 449.315 90.695 ;
        RECT 450.025 88.705 450.195 90.695 ;
        RECT 450.905 88.705 451.075 90.695 ;
        RECT 451.785 88.705 451.955 90.695 ;
        RECT 446.845 88.205 448.095 88.535 ;
        RECT 448.605 88.205 449.855 88.535 ;
        RECT 452.355 87.960 452.645 91.445 ;
        RECT 444.055 87.670 452.645 87.960 ;
        RECT 453.275 87.965 453.565 94.115 ;
        RECT 454.245 93.545 455.135 93.875 ;
        RECT 455.525 93.545 456.415 93.875 ;
        RECT 456.965 93.545 461.815 93.875 ;
        RECT 462.525 93.545 467.375 93.875 ;
        RECT 467.925 93.545 468.815 93.875 ;
        RECT 469.205 93.545 470.095 93.875 ;
        RECT 453.965 91.375 454.135 93.375 ;
        RECT 455.245 91.375 455.415 93.375 ;
        RECT 456.525 91.375 456.695 93.375 ;
        RECT 462.085 91.375 462.255 93.375 ;
        RECT 467.645 91.375 467.815 93.375 ;
        RECT 468.925 91.375 469.095 93.375 ;
        RECT 470.205 91.375 470.375 93.375 ;
        RECT 454.245 90.875 455.135 91.205 ;
        RECT 455.525 90.875 456.415 91.205 ;
        RECT 456.965 90.875 461.815 91.205 ;
        RECT 462.525 90.875 467.375 91.205 ;
        RECT 467.925 90.875 468.815 91.205 ;
        RECT 469.205 90.875 470.095 91.205 ;
        RECT 453.965 88.705 454.135 90.705 ;
        RECT 455.245 88.705 455.415 90.705 ;
        RECT 456.525 88.705 456.695 90.705 ;
        RECT 462.085 88.705 462.255 90.705 ;
        RECT 467.645 88.705 467.815 90.705 ;
        RECT 468.925 88.705 469.095 90.705 ;
        RECT 470.205 88.705 470.375 90.705 ;
        RECT 456.965 88.205 461.815 88.535 ;
        RECT 462.525 88.205 467.375 88.535 ;
        RECT 470.775 87.965 471.065 94.115 ;
        RECT 472.625 93.345 472.915 97.085 ;
        RECT 473.655 96.515 474.905 96.845 ;
        RECT 478.935 96.515 480.185 96.845 ;
        RECT 473.315 94.085 473.485 96.345 ;
        RECT 474.195 94.085 474.365 96.345 ;
        RECT 475.075 94.085 475.245 96.345 ;
        RECT 475.955 94.085 476.125 96.345 ;
        RECT 476.835 94.085 477.005 96.345 ;
        RECT 477.715 94.085 477.885 96.345 ;
        RECT 478.595 94.085 478.765 96.345 ;
        RECT 479.475 94.085 479.645 96.345 ;
        RECT 480.355 94.085 480.525 96.345 ;
        RECT 475.415 93.585 476.665 93.915 ;
        RECT 477.175 93.585 478.425 93.915 ;
        RECT 480.925 93.345 481.215 97.085 ;
        RECT 487.050 95.020 487.340 105.530 ;
        RECT 489.880 104.960 491.130 105.290 ;
        RECT 491.640 104.960 492.890 105.290 ;
        RECT 487.780 95.760 487.950 104.790 ;
        RECT 488.660 95.760 488.830 104.790 ;
        RECT 489.540 95.760 489.710 104.790 ;
        RECT 490.420 95.760 490.590 104.790 ;
        RECT 491.300 95.760 491.470 104.790 ;
        RECT 492.180 95.760 492.350 104.790 ;
        RECT 493.060 95.760 493.230 104.790 ;
        RECT 493.940 95.760 494.110 104.790 ;
        RECT 494.820 95.760 494.990 104.790 ;
        RECT 488.120 95.260 489.370 95.590 ;
        RECT 493.400 95.260 494.650 95.590 ;
        RECT 495.430 95.020 495.720 105.530 ;
        RECT 487.050 94.730 495.720 95.020 ;
        RECT 496.820 97.085 505.410 97.375 ;
        RECT 472.625 93.055 481.215 93.345 ;
        RECT 496.820 93.345 497.110 97.085 ;
        RECT 497.850 96.515 499.100 96.845 ;
        RECT 503.130 96.515 504.380 96.845 ;
        RECT 497.510 94.085 497.680 96.345 ;
        RECT 498.390 94.085 498.560 96.345 ;
        RECT 499.270 94.085 499.440 96.345 ;
        RECT 500.150 94.085 500.320 96.345 ;
        RECT 501.030 94.085 501.200 96.345 ;
        RECT 501.910 94.085 502.080 96.345 ;
        RECT 502.790 94.085 502.960 96.345 ;
        RECT 503.670 94.085 503.840 96.345 ;
        RECT 504.550 94.085 504.720 96.345 ;
        RECT 499.610 93.585 500.860 93.915 ;
        RECT 501.370 93.585 502.620 93.915 ;
        RECT 505.120 93.345 505.410 97.085 ;
        RECT 496.820 93.055 505.410 93.345 ;
        RECT 453.275 87.675 471.065 87.965 ;
        RECT 472.625 91.705 481.215 91.995 ;
        RECT 472.625 87.965 472.915 91.705 ;
        RECT 473.655 91.135 474.905 91.465 ;
        RECT 478.935 91.135 480.185 91.465 ;
        RECT 473.315 88.705 473.485 90.965 ;
        RECT 474.195 88.705 474.365 90.965 ;
        RECT 475.075 88.705 475.245 90.965 ;
        RECT 475.955 88.705 476.125 90.965 ;
        RECT 476.835 88.705 477.005 90.965 ;
        RECT 477.715 88.705 477.885 90.965 ;
        RECT 478.595 88.705 478.765 90.965 ;
        RECT 479.475 88.705 479.645 90.965 ;
        RECT 480.355 88.705 480.525 90.965 ;
        RECT 475.415 88.205 476.665 88.535 ;
        RECT 477.175 88.205 478.425 88.535 ;
        RECT 480.925 87.965 481.215 91.705 ;
        RECT 472.625 87.675 481.215 87.965 ;
        RECT 487.090 91.445 495.680 91.735 ;
        RECT 487.090 87.965 487.380 91.445 ;
        RECT 489.880 90.875 491.130 91.205 ;
        RECT 491.640 90.875 492.890 91.205 ;
        RECT 487.780 88.705 487.950 90.705 ;
        RECT 488.660 88.705 488.830 90.705 ;
        RECT 489.540 88.705 489.710 90.705 ;
        RECT 490.420 88.705 490.590 90.705 ;
        RECT 491.300 88.705 491.470 90.705 ;
        RECT 492.180 88.705 492.350 90.705 ;
        RECT 493.060 88.705 493.230 90.705 ;
        RECT 493.940 88.705 494.110 90.705 ;
        RECT 494.820 88.705 494.990 90.705 ;
        RECT 488.120 88.205 489.370 88.535 ;
        RECT 493.400 88.205 494.650 88.535 ;
        RECT 495.390 87.965 495.680 91.445 ;
        RECT 487.090 87.675 495.680 87.965 ;
        RECT 496.820 91.705 505.410 91.995 ;
        RECT 496.820 87.965 497.110 91.705 ;
        RECT 497.850 91.135 499.100 91.465 ;
        RECT 503.130 91.135 504.380 91.465 ;
        RECT 497.510 88.705 497.680 90.965 ;
        RECT 498.390 88.705 498.560 90.965 ;
        RECT 499.270 88.705 499.440 90.965 ;
        RECT 500.150 88.705 500.320 90.965 ;
        RECT 501.030 88.705 501.200 90.965 ;
        RECT 501.910 88.705 502.080 90.965 ;
        RECT 502.790 88.705 502.960 90.965 ;
        RECT 503.670 88.705 503.840 90.965 ;
        RECT 504.550 88.705 504.720 90.965 ;
        RECT 499.610 88.205 500.860 88.535 ;
        RECT 501.370 88.205 502.620 88.535 ;
        RECT 505.120 87.965 505.410 91.705 ;
        RECT 496.820 87.675 505.410 87.965 ;
        RECT 364.455 85.470 406.605 85.760 ;
        RECT 437.465 83.260 502.870 83.430 ;
        RECT 437.465 82.060 437.635 83.260 ;
        RECT 438.360 82.060 439.770 82.640 ;
        RECT 440.370 82.060 441.780 82.640 ;
        RECT 184.845 81.695 294.365 81.865 ;
        RECT 184.845 80.490 185.015 81.695 ;
        RECT 185.635 80.490 187.045 81.075 ;
        RECT 187.645 80.490 189.055 81.075 ;
        RECT 184.845 79.490 189.055 80.490 ;
        RECT 184.845 70.895 185.015 79.490 ;
        RECT 185.635 78.915 187.045 79.490 ;
        RECT 187.645 78.915 189.055 79.490 ;
        RECT 189.655 78.915 191.065 81.075 ;
        RECT 191.665 78.915 193.075 81.075 ;
        RECT 193.675 78.915 195.085 81.075 ;
        RECT 195.685 78.915 197.095 81.075 ;
        RECT 197.695 78.915 199.105 81.075 ;
        RECT 199.705 78.915 201.115 81.075 ;
        RECT 201.715 78.915 203.125 81.075 ;
        RECT 203.725 78.915 205.135 81.075 ;
        RECT 205.735 78.915 207.145 81.075 ;
        RECT 207.745 78.915 209.155 81.075 ;
        RECT 209.755 78.915 211.165 81.075 ;
        RECT 211.765 78.915 213.175 81.075 ;
        RECT 213.775 78.915 215.185 81.075 ;
        RECT 215.785 78.915 217.195 81.075 ;
        RECT 217.795 78.915 219.205 81.075 ;
        RECT 219.805 78.915 221.215 81.075 ;
        RECT 221.815 78.915 223.225 81.075 ;
        RECT 223.825 78.915 225.235 81.075 ;
        RECT 225.835 78.915 227.245 81.075 ;
        RECT 227.845 78.915 229.255 81.075 ;
        RECT 229.855 78.915 231.265 81.075 ;
        RECT 231.865 78.915 233.275 81.075 ;
        RECT 233.875 78.915 235.285 81.075 ;
        RECT 235.885 78.915 237.295 81.075 ;
        RECT 237.895 78.915 239.305 81.075 ;
        RECT 239.905 78.915 241.315 81.075 ;
        RECT 241.915 78.915 243.325 81.075 ;
        RECT 243.925 78.915 245.335 81.075 ;
        RECT 245.935 78.915 247.345 81.075 ;
        RECT 247.945 78.915 249.355 81.075 ;
        RECT 249.955 78.915 251.365 81.075 ;
        RECT 251.965 78.915 253.375 81.075 ;
        RECT 253.975 78.915 255.385 81.075 ;
        RECT 255.985 78.915 257.395 81.075 ;
        RECT 257.995 78.915 259.405 81.075 ;
        RECT 260.005 78.915 261.415 81.075 ;
        RECT 262.015 78.915 263.425 81.075 ;
        RECT 264.025 78.915 265.435 81.075 ;
        RECT 266.035 78.915 267.445 81.075 ;
        RECT 268.045 78.915 269.455 81.075 ;
        RECT 270.055 78.915 271.465 81.075 ;
        RECT 272.065 78.915 273.475 81.075 ;
        RECT 274.075 78.915 275.485 81.075 ;
        RECT 276.085 78.915 277.495 81.075 ;
        RECT 278.095 78.915 279.505 81.075 ;
        RECT 280.105 78.915 281.515 81.075 ;
        RECT 282.115 78.915 283.525 81.075 ;
        RECT 284.125 78.915 285.535 81.075 ;
        RECT 286.135 78.915 287.545 81.075 ;
        RECT 288.145 78.915 289.555 81.075 ;
        RECT 290.155 80.490 291.565 81.075 ;
        RECT 292.165 80.490 293.575 81.075 ;
        RECT 294.195 80.490 294.365 81.695 ;
        RECT 290.155 79.490 294.365 80.490 ;
        RECT 290.155 78.915 291.565 79.490 ;
        RECT 292.165 78.915 293.575 79.490 ;
        RECT 185.635 70.895 187.045 71.475 ;
        RECT 187.645 70.895 189.055 71.475 ;
        RECT 184.845 69.895 189.055 70.895 ;
        RECT 184.845 68.695 185.015 69.895 ;
        RECT 185.635 69.315 187.045 69.895 ;
        RECT 187.645 69.315 189.055 69.895 ;
        RECT 189.655 69.315 191.065 71.475 ;
        RECT 191.665 69.315 193.075 71.475 ;
        RECT 193.675 69.315 195.085 71.475 ;
        RECT 195.685 69.315 197.095 71.475 ;
        RECT 197.695 69.315 199.105 71.475 ;
        RECT 199.705 69.315 201.115 71.475 ;
        RECT 201.715 69.315 203.125 71.475 ;
        RECT 203.725 69.315 205.135 71.475 ;
        RECT 205.735 69.315 207.145 71.475 ;
        RECT 207.745 69.315 209.155 71.475 ;
        RECT 209.755 69.315 211.165 71.475 ;
        RECT 211.765 69.315 213.175 71.475 ;
        RECT 213.775 69.315 215.185 71.475 ;
        RECT 215.785 69.315 217.195 71.475 ;
        RECT 217.795 69.315 219.205 71.475 ;
        RECT 219.805 69.315 221.215 71.475 ;
        RECT 221.815 69.315 223.225 71.475 ;
        RECT 223.825 69.315 225.235 71.475 ;
        RECT 225.835 69.315 227.245 71.475 ;
        RECT 227.845 69.315 229.255 71.475 ;
        RECT 229.855 69.315 231.265 71.475 ;
        RECT 231.865 69.315 233.275 71.475 ;
        RECT 233.875 69.315 235.285 71.475 ;
        RECT 235.885 69.315 237.295 71.475 ;
        RECT 237.895 69.315 239.305 71.475 ;
        RECT 239.905 69.315 241.315 71.475 ;
        RECT 241.915 69.315 243.325 71.475 ;
        RECT 243.925 69.315 245.335 71.475 ;
        RECT 245.935 69.315 247.345 71.475 ;
        RECT 247.945 69.315 249.355 71.475 ;
        RECT 249.955 69.315 251.365 71.475 ;
        RECT 251.965 69.315 253.375 71.475 ;
        RECT 253.975 69.315 255.385 71.475 ;
        RECT 255.985 69.315 257.395 71.475 ;
        RECT 257.995 69.315 259.405 71.475 ;
        RECT 260.005 69.315 261.415 71.475 ;
        RECT 262.015 69.315 263.425 71.475 ;
        RECT 264.025 69.315 265.435 71.475 ;
        RECT 266.035 69.315 267.445 71.475 ;
        RECT 268.045 69.315 269.455 71.475 ;
        RECT 270.055 69.315 271.465 71.475 ;
        RECT 272.065 69.315 273.475 71.475 ;
        RECT 274.075 69.315 275.485 71.475 ;
        RECT 276.085 69.315 277.495 71.475 ;
        RECT 278.095 69.315 279.505 71.475 ;
        RECT 280.105 69.315 281.515 71.475 ;
        RECT 282.115 69.315 283.525 71.475 ;
        RECT 284.125 69.315 285.535 71.475 ;
        RECT 286.135 69.315 287.545 71.475 ;
        RECT 288.145 69.315 289.555 71.475 ;
        RECT 290.155 70.895 291.565 71.475 ;
        RECT 292.165 70.895 293.575 71.475 ;
        RECT 294.195 70.895 294.365 79.490 ;
        RECT 290.155 69.895 294.365 70.895 ;
        RECT 290.155 69.315 291.565 69.895 ;
        RECT 292.165 69.315 293.575 69.895 ;
        RECT 294.195 68.695 294.365 69.895 ;
        RECT 184.845 68.525 294.365 68.695 ;
        RECT 300.380 81.695 409.900 81.865 ;
        RECT 300.380 80.490 300.550 81.695 ;
        RECT 301.170 80.490 302.580 81.075 ;
        RECT 303.180 80.490 304.590 81.075 ;
        RECT 300.380 79.490 304.590 80.490 ;
        RECT 300.380 70.895 300.550 79.490 ;
        RECT 301.170 78.915 302.580 79.490 ;
        RECT 303.180 78.915 304.590 79.490 ;
        RECT 305.190 78.915 306.600 81.075 ;
        RECT 307.200 78.915 308.610 81.075 ;
        RECT 309.210 78.915 310.620 81.075 ;
        RECT 311.220 78.915 312.630 81.075 ;
        RECT 313.230 78.915 314.640 81.075 ;
        RECT 315.240 78.915 316.650 81.075 ;
        RECT 317.250 78.915 318.660 81.075 ;
        RECT 319.260 78.915 320.670 81.075 ;
        RECT 321.270 78.915 322.680 81.075 ;
        RECT 323.280 78.915 324.690 81.075 ;
        RECT 325.290 78.915 326.700 81.075 ;
        RECT 327.300 78.915 328.710 81.075 ;
        RECT 329.310 78.915 330.720 81.075 ;
        RECT 331.320 78.915 332.730 81.075 ;
        RECT 333.330 78.915 334.740 81.075 ;
        RECT 335.340 78.915 336.750 81.075 ;
        RECT 337.350 78.915 338.760 81.075 ;
        RECT 339.360 78.915 340.770 81.075 ;
        RECT 341.370 78.915 342.780 81.075 ;
        RECT 343.380 78.915 344.790 81.075 ;
        RECT 345.390 78.915 346.800 81.075 ;
        RECT 347.400 78.915 348.810 81.075 ;
        RECT 349.410 78.915 350.820 81.075 ;
        RECT 351.420 78.915 352.830 81.075 ;
        RECT 353.430 78.915 354.840 81.075 ;
        RECT 355.440 78.915 356.850 81.075 ;
        RECT 357.450 78.915 358.860 81.075 ;
        RECT 359.460 78.915 360.870 81.075 ;
        RECT 361.470 78.915 362.880 81.075 ;
        RECT 363.480 78.915 364.890 81.075 ;
        RECT 365.490 78.915 366.900 81.075 ;
        RECT 367.500 78.915 368.910 81.075 ;
        RECT 369.510 78.915 370.920 81.075 ;
        RECT 371.520 78.915 372.930 81.075 ;
        RECT 373.530 78.915 374.940 81.075 ;
        RECT 375.540 78.915 376.950 81.075 ;
        RECT 377.550 78.915 378.960 81.075 ;
        RECT 379.560 78.915 380.970 81.075 ;
        RECT 381.570 78.915 382.980 81.075 ;
        RECT 383.580 78.915 384.990 81.075 ;
        RECT 385.590 78.915 387.000 81.075 ;
        RECT 387.600 78.915 389.010 81.075 ;
        RECT 389.610 78.915 391.020 81.075 ;
        RECT 391.620 78.915 393.030 81.075 ;
        RECT 393.630 78.915 395.040 81.075 ;
        RECT 395.640 78.915 397.050 81.075 ;
        RECT 397.650 78.915 399.060 81.075 ;
        RECT 399.660 78.915 401.070 81.075 ;
        RECT 401.670 78.915 403.080 81.075 ;
        RECT 403.680 78.915 405.090 81.075 ;
        RECT 405.690 80.490 407.100 81.075 ;
        RECT 407.700 80.490 409.110 81.075 ;
        RECT 409.730 80.490 409.900 81.695 ;
        RECT 405.690 79.490 409.900 80.490 ;
        RECT 405.690 78.915 407.100 79.490 ;
        RECT 407.700 78.915 409.110 79.490 ;
        RECT 301.170 70.895 302.580 71.475 ;
        RECT 303.180 70.895 304.590 71.475 ;
        RECT 300.380 69.895 304.590 70.895 ;
        RECT 300.380 68.695 300.550 69.895 ;
        RECT 301.170 69.315 302.580 69.895 ;
        RECT 303.180 69.315 304.590 69.895 ;
        RECT 305.190 69.315 306.600 71.475 ;
        RECT 307.200 69.315 308.610 71.475 ;
        RECT 309.210 69.315 310.620 71.475 ;
        RECT 311.220 69.315 312.630 71.475 ;
        RECT 313.230 69.315 314.640 71.475 ;
        RECT 315.240 69.315 316.650 71.475 ;
        RECT 317.250 69.315 318.660 71.475 ;
        RECT 319.260 69.315 320.670 71.475 ;
        RECT 321.270 69.315 322.680 71.475 ;
        RECT 323.280 69.315 324.690 71.475 ;
        RECT 325.290 69.315 326.700 71.475 ;
        RECT 327.300 69.315 328.710 71.475 ;
        RECT 329.310 69.315 330.720 71.475 ;
        RECT 331.320 69.315 332.730 71.475 ;
        RECT 333.330 69.315 334.740 71.475 ;
        RECT 335.340 69.315 336.750 71.475 ;
        RECT 337.350 69.315 338.760 71.475 ;
        RECT 339.360 69.315 340.770 71.475 ;
        RECT 341.370 69.315 342.780 71.475 ;
        RECT 343.380 69.315 344.790 71.475 ;
        RECT 345.390 69.315 346.800 71.475 ;
        RECT 347.400 69.315 348.810 71.475 ;
        RECT 349.410 69.315 350.820 71.475 ;
        RECT 351.420 69.315 352.830 71.475 ;
        RECT 353.430 69.315 354.840 71.475 ;
        RECT 355.440 69.315 356.850 71.475 ;
        RECT 357.450 69.315 358.860 71.475 ;
        RECT 359.460 69.315 360.870 71.475 ;
        RECT 361.470 69.315 362.880 71.475 ;
        RECT 363.480 69.315 364.890 71.475 ;
        RECT 365.490 69.315 366.900 71.475 ;
        RECT 367.500 69.315 368.910 71.475 ;
        RECT 369.510 69.315 370.920 71.475 ;
        RECT 371.520 69.315 372.930 71.475 ;
        RECT 373.530 69.315 374.940 71.475 ;
        RECT 375.540 69.315 376.950 71.475 ;
        RECT 377.550 69.315 378.960 71.475 ;
        RECT 379.560 69.315 380.970 71.475 ;
        RECT 381.570 69.315 382.980 71.475 ;
        RECT 383.580 69.315 384.990 71.475 ;
        RECT 385.590 69.315 387.000 71.475 ;
        RECT 387.600 69.315 389.010 71.475 ;
        RECT 389.610 69.315 391.020 71.475 ;
        RECT 391.620 69.315 393.030 71.475 ;
        RECT 393.630 69.315 395.040 71.475 ;
        RECT 395.640 69.315 397.050 71.475 ;
        RECT 397.650 69.315 399.060 71.475 ;
        RECT 399.660 69.315 401.070 71.475 ;
        RECT 401.670 69.315 403.080 71.475 ;
        RECT 403.680 69.315 405.090 71.475 ;
        RECT 405.690 70.895 407.100 71.475 ;
        RECT 407.700 70.895 409.110 71.475 ;
        RECT 409.730 70.895 409.900 79.490 ;
        RECT 405.690 69.895 409.900 70.895 ;
        RECT 437.465 81.060 441.780 82.060 ;
        RECT 437.465 75.900 437.635 81.060 ;
        RECT 438.360 80.480 439.770 81.060 ;
        RECT 440.370 80.480 441.780 81.060 ;
        RECT 442.380 80.480 443.790 82.640 ;
        RECT 444.390 80.480 445.800 82.640 ;
        RECT 446.400 80.480 447.810 82.640 ;
        RECT 448.410 80.480 449.820 82.640 ;
        RECT 450.420 80.480 451.830 82.640 ;
        RECT 452.430 80.480 453.840 82.640 ;
        RECT 454.440 80.480 455.850 82.640 ;
        RECT 456.450 80.480 457.860 82.640 ;
        RECT 458.460 80.480 459.870 82.640 ;
        RECT 460.470 80.480 461.880 82.640 ;
        RECT 462.480 80.480 463.890 82.640 ;
        RECT 464.490 80.480 465.900 82.640 ;
        RECT 466.500 80.480 467.910 82.640 ;
        RECT 468.510 80.480 469.920 82.640 ;
        RECT 470.520 80.480 471.930 82.640 ;
        RECT 472.530 80.480 473.940 82.640 ;
        RECT 474.540 80.480 475.950 82.640 ;
        RECT 476.550 80.480 477.960 82.640 ;
        RECT 478.560 80.480 479.970 82.640 ;
        RECT 480.570 80.480 481.980 82.640 ;
        RECT 482.580 80.480 483.990 82.640 ;
        RECT 484.590 80.480 486.000 82.640 ;
        RECT 486.600 80.480 488.010 82.640 ;
        RECT 488.610 80.480 490.020 82.640 ;
        RECT 490.620 80.480 492.030 82.640 ;
        RECT 492.630 80.480 494.040 82.640 ;
        RECT 494.640 80.480 496.050 82.640 ;
        RECT 496.650 80.480 498.060 82.640 ;
        RECT 498.660 82.060 500.070 82.640 ;
        RECT 500.670 82.060 502.080 82.640 ;
        RECT 502.700 82.060 502.870 83.260 ;
        RECT 498.660 81.060 502.870 82.060 ;
        RECT 498.660 80.480 500.070 81.060 ;
        RECT 500.670 80.480 502.080 81.060 ;
        RECT 437.465 73.900 437.740 75.900 ;
        RECT 437.465 72.460 437.635 73.900 ;
        RECT 438.360 72.460 439.770 73.040 ;
        RECT 440.370 72.460 441.780 73.040 ;
        RECT 437.465 71.460 441.780 72.460 ;
        RECT 437.465 70.260 437.635 71.460 ;
        RECT 438.360 70.880 439.770 71.460 ;
        RECT 440.370 70.880 441.780 71.460 ;
        RECT 442.380 70.880 443.790 73.040 ;
        RECT 444.390 70.880 445.800 73.040 ;
        RECT 446.400 70.880 447.810 73.040 ;
        RECT 448.410 70.880 449.820 73.040 ;
        RECT 450.420 70.880 451.830 73.040 ;
        RECT 452.430 70.880 453.840 73.040 ;
        RECT 454.440 70.880 455.850 73.040 ;
        RECT 456.450 70.880 457.860 73.040 ;
        RECT 458.460 70.880 459.870 73.040 ;
        RECT 460.470 70.880 461.880 73.040 ;
        RECT 462.480 70.880 463.890 73.040 ;
        RECT 464.490 70.880 465.900 73.040 ;
        RECT 466.500 70.880 467.910 73.040 ;
        RECT 468.510 70.880 469.920 73.040 ;
        RECT 470.520 70.880 471.930 73.040 ;
        RECT 472.530 70.880 473.940 73.040 ;
        RECT 474.540 70.880 475.950 73.040 ;
        RECT 476.550 70.880 477.960 73.040 ;
        RECT 478.560 70.880 479.970 73.040 ;
        RECT 480.570 70.880 481.980 73.040 ;
        RECT 482.580 70.880 483.990 73.040 ;
        RECT 484.590 70.880 486.000 73.040 ;
        RECT 486.600 70.880 488.010 73.040 ;
        RECT 488.610 70.880 490.020 73.040 ;
        RECT 490.620 70.880 492.030 73.040 ;
        RECT 492.630 70.880 494.040 73.040 ;
        RECT 494.640 70.880 496.050 73.040 ;
        RECT 496.650 70.880 498.060 73.040 ;
        RECT 498.660 72.460 500.070 73.040 ;
        RECT 500.670 72.460 502.080 73.040 ;
        RECT 502.700 72.460 502.870 81.060 ;
        RECT 498.660 71.460 502.870 72.460 ;
        RECT 498.660 70.880 500.070 71.460 ;
        RECT 500.670 70.880 502.080 71.460 ;
        RECT 502.700 70.260 502.870 71.460 ;
        RECT 437.465 70.090 502.870 70.260 ;
        RECT 405.690 69.315 407.100 69.895 ;
        RECT 407.700 69.315 409.110 69.895 ;
        RECT 409.730 68.695 409.900 69.895 ;
        RECT 300.380 68.525 409.900 68.695 ;
        RECT 184.845 67.550 294.365 67.720 ;
        RECT 184.845 66.345 185.015 67.550 ;
        RECT 185.635 66.345 187.045 66.930 ;
        RECT 187.645 66.345 189.055 66.930 ;
        RECT 184.845 65.345 189.055 66.345 ;
        RECT 184.845 56.750 185.015 65.345 ;
        RECT 185.635 64.770 187.045 65.345 ;
        RECT 187.645 64.770 189.055 65.345 ;
        RECT 189.655 64.770 191.065 66.930 ;
        RECT 191.665 64.770 193.075 66.930 ;
        RECT 193.675 64.770 195.085 66.930 ;
        RECT 195.685 64.770 197.095 66.930 ;
        RECT 197.695 64.770 199.105 66.930 ;
        RECT 199.705 64.770 201.115 66.930 ;
        RECT 201.715 64.770 203.125 66.930 ;
        RECT 203.725 64.770 205.135 66.930 ;
        RECT 205.735 64.770 207.145 66.930 ;
        RECT 207.745 64.770 209.155 66.930 ;
        RECT 209.755 64.770 211.165 66.930 ;
        RECT 211.765 64.770 213.175 66.930 ;
        RECT 213.775 64.770 215.185 66.930 ;
        RECT 215.785 64.770 217.195 66.930 ;
        RECT 217.795 64.770 219.205 66.930 ;
        RECT 219.805 64.770 221.215 66.930 ;
        RECT 221.815 64.770 223.225 66.930 ;
        RECT 223.825 64.770 225.235 66.930 ;
        RECT 225.835 64.770 227.245 66.930 ;
        RECT 227.845 64.770 229.255 66.930 ;
        RECT 229.855 64.770 231.265 66.930 ;
        RECT 231.865 64.770 233.275 66.930 ;
        RECT 233.875 64.770 235.285 66.930 ;
        RECT 235.885 64.770 237.295 66.930 ;
        RECT 237.895 64.770 239.305 66.930 ;
        RECT 239.905 64.770 241.315 66.930 ;
        RECT 241.915 64.770 243.325 66.930 ;
        RECT 243.925 64.770 245.335 66.930 ;
        RECT 245.935 64.770 247.345 66.930 ;
        RECT 247.945 64.770 249.355 66.930 ;
        RECT 249.955 64.770 251.365 66.930 ;
        RECT 251.965 64.770 253.375 66.930 ;
        RECT 253.975 64.770 255.385 66.930 ;
        RECT 255.985 64.770 257.395 66.930 ;
        RECT 257.995 64.770 259.405 66.930 ;
        RECT 260.005 64.770 261.415 66.930 ;
        RECT 262.015 64.770 263.425 66.930 ;
        RECT 264.025 64.770 265.435 66.930 ;
        RECT 266.035 64.770 267.445 66.930 ;
        RECT 268.045 64.770 269.455 66.930 ;
        RECT 270.055 64.770 271.465 66.930 ;
        RECT 272.065 64.770 273.475 66.930 ;
        RECT 274.075 64.770 275.485 66.930 ;
        RECT 276.085 64.770 277.495 66.930 ;
        RECT 278.095 64.770 279.505 66.930 ;
        RECT 280.105 64.770 281.515 66.930 ;
        RECT 282.115 64.770 283.525 66.930 ;
        RECT 284.125 64.770 285.535 66.930 ;
        RECT 286.135 64.770 287.545 66.930 ;
        RECT 288.145 64.770 289.555 66.930 ;
        RECT 290.155 66.345 291.565 66.930 ;
        RECT 292.165 66.345 293.575 66.930 ;
        RECT 294.195 66.345 294.365 67.550 ;
        RECT 290.155 65.345 294.365 66.345 ;
        RECT 290.155 64.770 291.565 65.345 ;
        RECT 292.165 64.770 293.575 65.345 ;
        RECT 185.635 56.750 187.045 57.330 ;
        RECT 187.645 56.750 189.055 57.330 ;
        RECT 184.845 55.750 189.055 56.750 ;
        RECT 184.845 54.550 185.015 55.750 ;
        RECT 185.635 55.170 187.045 55.750 ;
        RECT 187.645 55.170 189.055 55.750 ;
        RECT 189.655 55.170 191.065 57.330 ;
        RECT 191.665 55.170 193.075 57.330 ;
        RECT 193.675 55.170 195.085 57.330 ;
        RECT 195.685 55.170 197.095 57.330 ;
        RECT 197.695 55.170 199.105 57.330 ;
        RECT 199.705 55.170 201.115 57.330 ;
        RECT 201.715 55.170 203.125 57.330 ;
        RECT 203.725 55.170 205.135 57.330 ;
        RECT 205.735 55.170 207.145 57.330 ;
        RECT 207.745 55.170 209.155 57.330 ;
        RECT 209.755 55.170 211.165 57.330 ;
        RECT 211.765 55.170 213.175 57.330 ;
        RECT 213.775 55.170 215.185 57.330 ;
        RECT 215.785 55.170 217.195 57.330 ;
        RECT 217.795 55.170 219.205 57.330 ;
        RECT 219.805 55.170 221.215 57.330 ;
        RECT 221.815 55.170 223.225 57.330 ;
        RECT 223.825 55.170 225.235 57.330 ;
        RECT 225.835 55.170 227.245 57.330 ;
        RECT 227.845 55.170 229.255 57.330 ;
        RECT 229.855 55.170 231.265 57.330 ;
        RECT 231.865 55.170 233.275 57.330 ;
        RECT 233.875 55.170 235.285 57.330 ;
        RECT 235.885 55.170 237.295 57.330 ;
        RECT 237.895 55.170 239.305 57.330 ;
        RECT 239.905 55.170 241.315 57.330 ;
        RECT 241.915 55.170 243.325 57.330 ;
        RECT 243.925 55.170 245.335 57.330 ;
        RECT 245.935 55.170 247.345 57.330 ;
        RECT 247.945 55.170 249.355 57.330 ;
        RECT 249.955 55.170 251.365 57.330 ;
        RECT 251.965 55.170 253.375 57.330 ;
        RECT 253.975 55.170 255.385 57.330 ;
        RECT 255.985 55.170 257.395 57.330 ;
        RECT 257.995 55.170 259.405 57.330 ;
        RECT 260.005 55.170 261.415 57.330 ;
        RECT 262.015 55.170 263.425 57.330 ;
        RECT 264.025 55.170 265.435 57.330 ;
        RECT 266.035 55.170 267.445 57.330 ;
        RECT 268.045 55.170 269.455 57.330 ;
        RECT 270.055 55.170 271.465 57.330 ;
        RECT 272.065 55.170 273.475 57.330 ;
        RECT 274.075 55.170 275.485 57.330 ;
        RECT 276.085 55.170 277.495 57.330 ;
        RECT 278.095 55.170 279.505 57.330 ;
        RECT 280.105 55.170 281.515 57.330 ;
        RECT 282.115 55.170 283.525 57.330 ;
        RECT 284.125 55.170 285.535 57.330 ;
        RECT 286.135 55.170 287.545 57.330 ;
        RECT 288.145 55.170 289.555 57.330 ;
        RECT 290.155 56.750 291.565 57.330 ;
        RECT 292.165 56.750 293.575 57.330 ;
        RECT 294.195 56.750 294.365 65.345 ;
        RECT 290.155 55.750 294.365 56.750 ;
        RECT 290.155 55.170 291.565 55.750 ;
        RECT 292.165 55.170 293.575 55.750 ;
        RECT 294.195 54.550 294.365 55.750 ;
        RECT 184.845 54.380 294.365 54.550 ;
        RECT 300.380 67.550 409.900 67.720 ;
        RECT 300.380 66.345 300.550 67.550 ;
        RECT 301.170 66.345 302.580 66.930 ;
        RECT 303.180 66.345 304.590 66.930 ;
        RECT 300.380 65.345 304.590 66.345 ;
        RECT 300.380 56.750 300.550 65.345 ;
        RECT 301.170 64.770 302.580 65.345 ;
        RECT 303.180 64.770 304.590 65.345 ;
        RECT 305.190 64.770 306.600 66.930 ;
        RECT 307.200 64.770 308.610 66.930 ;
        RECT 309.210 64.770 310.620 66.930 ;
        RECT 311.220 64.770 312.630 66.930 ;
        RECT 313.230 64.770 314.640 66.930 ;
        RECT 315.240 64.770 316.650 66.930 ;
        RECT 317.250 64.770 318.660 66.930 ;
        RECT 319.260 64.770 320.670 66.930 ;
        RECT 321.270 64.770 322.680 66.930 ;
        RECT 323.280 64.770 324.690 66.930 ;
        RECT 325.290 64.770 326.700 66.930 ;
        RECT 327.300 64.770 328.710 66.930 ;
        RECT 329.310 64.770 330.720 66.930 ;
        RECT 331.320 64.770 332.730 66.930 ;
        RECT 333.330 64.770 334.740 66.930 ;
        RECT 335.340 64.770 336.750 66.930 ;
        RECT 337.350 64.770 338.760 66.930 ;
        RECT 339.360 64.770 340.770 66.930 ;
        RECT 341.370 64.770 342.780 66.930 ;
        RECT 343.380 64.770 344.790 66.930 ;
        RECT 345.390 64.770 346.800 66.930 ;
        RECT 347.400 64.770 348.810 66.930 ;
        RECT 349.410 64.770 350.820 66.930 ;
        RECT 351.420 64.770 352.830 66.930 ;
        RECT 353.430 64.770 354.840 66.930 ;
        RECT 355.440 64.770 356.850 66.930 ;
        RECT 357.450 64.770 358.860 66.930 ;
        RECT 359.460 64.770 360.870 66.930 ;
        RECT 361.470 64.770 362.880 66.930 ;
        RECT 363.480 64.770 364.890 66.930 ;
        RECT 365.490 64.770 366.900 66.930 ;
        RECT 367.500 64.770 368.910 66.930 ;
        RECT 369.510 64.770 370.920 66.930 ;
        RECT 371.520 64.770 372.930 66.930 ;
        RECT 373.530 64.770 374.940 66.930 ;
        RECT 375.540 64.770 376.950 66.930 ;
        RECT 377.550 64.770 378.960 66.930 ;
        RECT 379.560 64.770 380.970 66.930 ;
        RECT 381.570 64.770 382.980 66.930 ;
        RECT 383.580 64.770 384.990 66.930 ;
        RECT 385.590 64.770 387.000 66.930 ;
        RECT 387.600 64.770 389.010 66.930 ;
        RECT 389.610 64.770 391.020 66.930 ;
        RECT 391.620 64.770 393.030 66.930 ;
        RECT 393.630 64.770 395.040 66.930 ;
        RECT 395.640 64.770 397.050 66.930 ;
        RECT 397.650 64.770 399.060 66.930 ;
        RECT 399.660 64.770 401.070 66.930 ;
        RECT 401.670 64.770 403.080 66.930 ;
        RECT 403.680 64.770 405.090 66.930 ;
        RECT 405.690 66.345 407.100 66.930 ;
        RECT 407.700 66.345 409.110 66.930 ;
        RECT 409.730 66.345 409.900 67.550 ;
        RECT 405.690 65.345 409.900 66.345 ;
        RECT 405.690 64.770 407.100 65.345 ;
        RECT 407.700 64.770 409.110 65.345 ;
        RECT 301.170 56.750 302.580 57.330 ;
        RECT 303.180 56.750 304.590 57.330 ;
        RECT 300.380 55.750 304.590 56.750 ;
        RECT 300.380 54.550 300.550 55.750 ;
        RECT 301.170 55.170 302.580 55.750 ;
        RECT 303.180 55.170 304.590 55.750 ;
        RECT 305.190 55.170 306.600 57.330 ;
        RECT 307.200 55.170 308.610 57.330 ;
        RECT 309.210 55.170 310.620 57.330 ;
        RECT 311.220 55.170 312.630 57.330 ;
        RECT 313.230 55.170 314.640 57.330 ;
        RECT 315.240 55.170 316.650 57.330 ;
        RECT 317.250 55.170 318.660 57.330 ;
        RECT 319.260 55.170 320.670 57.330 ;
        RECT 321.270 55.170 322.680 57.330 ;
        RECT 323.280 55.170 324.690 57.330 ;
        RECT 325.290 55.170 326.700 57.330 ;
        RECT 327.300 55.170 328.710 57.330 ;
        RECT 329.310 55.170 330.720 57.330 ;
        RECT 331.320 55.170 332.730 57.330 ;
        RECT 333.330 55.170 334.740 57.330 ;
        RECT 335.340 55.170 336.750 57.330 ;
        RECT 337.350 55.170 338.760 57.330 ;
        RECT 339.360 55.170 340.770 57.330 ;
        RECT 341.370 55.170 342.780 57.330 ;
        RECT 343.380 55.170 344.790 57.330 ;
        RECT 345.390 55.170 346.800 57.330 ;
        RECT 347.400 55.170 348.810 57.330 ;
        RECT 349.410 55.170 350.820 57.330 ;
        RECT 351.420 55.170 352.830 57.330 ;
        RECT 353.430 55.170 354.840 57.330 ;
        RECT 355.440 55.170 356.850 57.330 ;
        RECT 357.450 55.170 358.860 57.330 ;
        RECT 359.460 55.170 360.870 57.330 ;
        RECT 361.470 55.170 362.880 57.330 ;
        RECT 363.480 55.170 364.890 57.330 ;
        RECT 365.490 55.170 366.900 57.330 ;
        RECT 367.500 55.170 368.910 57.330 ;
        RECT 369.510 55.170 370.920 57.330 ;
        RECT 371.520 55.170 372.930 57.330 ;
        RECT 373.530 55.170 374.940 57.330 ;
        RECT 375.540 55.170 376.950 57.330 ;
        RECT 377.550 55.170 378.960 57.330 ;
        RECT 379.560 55.170 380.970 57.330 ;
        RECT 381.570 55.170 382.980 57.330 ;
        RECT 383.580 55.170 384.990 57.330 ;
        RECT 385.590 55.170 387.000 57.330 ;
        RECT 387.600 55.170 389.010 57.330 ;
        RECT 389.610 55.170 391.020 57.330 ;
        RECT 391.620 55.170 393.030 57.330 ;
        RECT 393.630 55.170 395.040 57.330 ;
        RECT 395.640 55.170 397.050 57.330 ;
        RECT 397.650 55.170 399.060 57.330 ;
        RECT 399.660 55.170 401.070 57.330 ;
        RECT 401.670 55.170 403.080 57.330 ;
        RECT 403.680 55.170 405.090 57.330 ;
        RECT 405.690 56.750 407.100 57.330 ;
        RECT 407.700 56.750 409.110 57.330 ;
        RECT 409.730 56.750 409.900 65.345 ;
        RECT 405.690 55.750 409.900 56.750 ;
        RECT 405.690 55.170 407.100 55.750 ;
        RECT 407.700 55.170 409.110 55.750 ;
        RECT 409.730 54.550 409.900 55.750 ;
        RECT 300.380 54.380 409.900 54.550 ;
        RECT 208.045 52.170 237.875 52.460 ;
        RECT 208.045 41.620 208.335 52.170 ;
        RECT 212.655 51.580 213.905 51.910 ;
        RECT 214.415 51.580 215.665 51.910 ;
        RECT 216.175 51.580 217.425 51.910 ;
        RECT 217.935 51.580 219.185 51.910 ;
        RECT 219.695 51.580 220.945 51.910 ;
        RECT 221.455 51.580 222.705 51.910 ;
        RECT 223.215 51.580 224.465 51.910 ;
        RECT 224.975 51.580 226.225 51.910 ;
        RECT 226.735 51.580 227.985 51.910 ;
        RECT 228.495 51.580 229.745 51.910 ;
        RECT 230.255 51.580 231.505 51.910 ;
        RECT 232.015 51.580 233.265 51.910 ;
        RECT 208.795 42.380 208.965 51.410 ;
        RECT 209.675 42.380 209.845 51.410 ;
        RECT 210.555 42.380 210.725 51.410 ;
        RECT 211.435 42.380 211.605 51.410 ;
        RECT 212.315 42.380 212.485 51.410 ;
        RECT 213.195 42.380 213.365 51.410 ;
        RECT 214.075 42.380 214.245 51.410 ;
        RECT 214.955 42.380 215.125 51.410 ;
        RECT 215.835 42.380 216.005 51.410 ;
        RECT 216.715 42.380 216.885 51.410 ;
        RECT 217.595 42.380 217.765 51.410 ;
        RECT 218.475 42.380 218.645 51.410 ;
        RECT 219.355 42.380 219.525 51.410 ;
        RECT 220.235 42.380 220.405 51.410 ;
        RECT 221.115 42.380 221.285 51.410 ;
        RECT 221.995 42.380 222.165 51.410 ;
        RECT 222.875 42.380 223.045 51.410 ;
        RECT 223.755 42.380 223.925 51.410 ;
        RECT 224.635 42.380 224.805 51.410 ;
        RECT 225.515 42.380 225.685 51.410 ;
        RECT 226.395 42.380 226.565 51.410 ;
        RECT 227.275 42.380 227.445 51.410 ;
        RECT 228.155 42.380 228.325 51.410 ;
        RECT 229.035 42.380 229.205 51.410 ;
        RECT 229.915 42.380 230.085 51.410 ;
        RECT 230.795 42.380 230.965 51.410 ;
        RECT 231.675 42.380 231.845 51.410 ;
        RECT 232.555 42.380 232.725 51.410 ;
        RECT 233.435 42.380 233.605 51.410 ;
        RECT 234.315 42.380 234.485 51.410 ;
        RECT 235.195 42.380 235.365 51.410 ;
        RECT 236.075 42.380 236.245 51.410 ;
        RECT 236.955 42.380 237.125 51.410 ;
        RECT 209.135 41.880 210.385 42.210 ;
        RECT 210.895 41.880 212.145 42.210 ;
        RECT 233.775 41.880 235.025 42.210 ;
        RECT 235.535 41.880 236.785 42.210 ;
        RECT 237.585 41.620 237.875 52.170 ;
        RECT 208.045 41.330 237.875 41.620 ;
        RECT 238.385 52.170 280.535 52.460 ;
        RECT 238.385 41.620 238.675 52.170 ;
        RECT 241.235 51.580 242.485 51.910 ;
        RECT 242.995 51.580 244.245 51.910 ;
        RECT 244.755 51.580 246.005 51.910 ;
        RECT 246.515 51.580 247.765 51.910 ;
        RECT 248.275 51.580 249.525 51.910 ;
        RECT 250.035 51.580 251.285 51.910 ;
        RECT 251.795 51.580 253.045 51.910 ;
        RECT 253.555 51.580 254.805 51.910 ;
        RECT 255.315 51.580 256.565 51.910 ;
        RECT 257.075 51.580 258.325 51.910 ;
        RECT 258.835 51.580 260.085 51.910 ;
        RECT 260.595 51.580 261.845 51.910 ;
        RECT 262.355 51.580 263.605 51.910 ;
        RECT 264.115 51.580 265.365 51.910 ;
        RECT 265.875 51.580 267.125 51.910 ;
        RECT 267.635 51.580 268.885 51.910 ;
        RECT 269.395 51.580 270.645 51.910 ;
        RECT 271.155 51.580 272.405 51.910 ;
        RECT 272.915 51.580 274.165 51.910 ;
        RECT 274.675 51.580 275.925 51.910 ;
        RECT 239.135 42.380 239.305 51.410 ;
        RECT 240.015 42.380 240.185 51.410 ;
        RECT 240.895 42.380 241.065 51.410 ;
        RECT 241.775 42.380 241.945 51.410 ;
        RECT 242.655 42.380 242.825 51.410 ;
        RECT 243.535 42.380 243.705 51.410 ;
        RECT 244.415 42.380 244.585 51.410 ;
        RECT 245.295 42.380 245.465 51.410 ;
        RECT 246.175 42.380 246.345 51.410 ;
        RECT 247.055 42.380 247.225 51.410 ;
        RECT 247.935 42.380 248.105 51.410 ;
        RECT 248.815 42.380 248.985 51.410 ;
        RECT 249.695 42.380 249.865 51.410 ;
        RECT 250.575 42.380 250.745 51.410 ;
        RECT 251.455 42.380 251.625 51.410 ;
        RECT 252.335 42.380 252.505 51.410 ;
        RECT 253.215 42.380 253.385 51.410 ;
        RECT 254.095 42.380 254.265 51.410 ;
        RECT 254.975 42.380 255.145 51.410 ;
        RECT 255.855 42.380 256.025 51.410 ;
        RECT 256.735 42.380 256.905 51.410 ;
        RECT 257.615 42.380 257.785 51.410 ;
        RECT 258.495 42.380 258.665 51.410 ;
        RECT 259.375 42.380 259.545 51.410 ;
        RECT 260.255 42.380 260.425 51.410 ;
        RECT 261.135 42.380 261.305 51.410 ;
        RECT 262.015 42.380 262.185 51.410 ;
        RECT 262.895 42.380 263.065 51.410 ;
        RECT 263.775 42.380 263.945 51.410 ;
        RECT 264.655 42.380 264.825 51.410 ;
        RECT 265.535 42.380 265.705 51.410 ;
        RECT 266.415 42.380 266.585 51.410 ;
        RECT 267.295 42.380 267.465 51.410 ;
        RECT 268.175 42.380 268.345 51.410 ;
        RECT 269.055 42.380 269.225 51.410 ;
        RECT 269.935 42.380 270.105 51.410 ;
        RECT 270.815 42.380 270.985 51.410 ;
        RECT 271.695 42.380 271.865 51.410 ;
        RECT 272.575 42.380 272.745 51.410 ;
        RECT 273.455 42.380 273.625 51.410 ;
        RECT 274.335 42.380 274.505 51.410 ;
        RECT 275.215 42.380 275.385 51.410 ;
        RECT 276.095 42.380 276.265 51.410 ;
        RECT 276.975 42.380 277.145 51.410 ;
        RECT 277.855 42.380 278.025 51.410 ;
        RECT 278.735 42.380 278.905 51.410 ;
        RECT 279.615 42.380 279.785 51.410 ;
        RECT 239.475 41.880 240.725 42.210 ;
        RECT 276.435 41.880 277.685 42.210 ;
        RECT 278.195 41.880 279.445 42.210 ;
        RECT 280.245 41.620 280.535 52.170 ;
        RECT 238.385 41.330 280.535 41.620 ;
        RECT 330.700 52.170 372.850 52.460 ;
        RECT 330.700 41.620 330.990 52.170 ;
        RECT 335.310 51.580 336.560 51.910 ;
        RECT 337.070 51.580 338.320 51.910 ;
        RECT 338.830 51.580 340.080 51.910 ;
        RECT 340.590 51.580 341.840 51.910 ;
        RECT 342.350 51.580 343.600 51.910 ;
        RECT 344.110 51.580 345.360 51.910 ;
        RECT 345.870 51.580 347.120 51.910 ;
        RECT 347.630 51.580 348.880 51.910 ;
        RECT 349.390 51.580 350.640 51.910 ;
        RECT 351.150 51.580 352.400 51.910 ;
        RECT 352.910 51.580 354.160 51.910 ;
        RECT 354.670 51.580 355.920 51.910 ;
        RECT 356.430 51.580 357.680 51.910 ;
        RECT 358.190 51.580 359.440 51.910 ;
        RECT 359.950 51.580 361.200 51.910 ;
        RECT 361.710 51.580 362.960 51.910 ;
        RECT 363.470 51.580 364.720 51.910 ;
        RECT 365.230 51.580 366.480 51.910 ;
        RECT 366.990 51.580 368.240 51.910 ;
        RECT 368.750 51.580 370.000 51.910 ;
        RECT 331.450 42.380 331.620 51.410 ;
        RECT 332.330 42.380 332.500 51.410 ;
        RECT 333.210 42.380 333.380 51.410 ;
        RECT 334.090 42.380 334.260 51.410 ;
        RECT 334.970 42.380 335.140 51.410 ;
        RECT 335.850 42.380 336.020 51.410 ;
        RECT 336.730 42.380 336.900 51.410 ;
        RECT 337.610 42.380 337.780 51.410 ;
        RECT 338.490 42.380 338.660 51.410 ;
        RECT 339.370 42.380 339.540 51.410 ;
        RECT 340.250 42.380 340.420 51.410 ;
        RECT 341.130 42.380 341.300 51.410 ;
        RECT 342.010 42.380 342.180 51.410 ;
        RECT 342.890 42.380 343.060 51.410 ;
        RECT 343.770 42.380 343.940 51.410 ;
        RECT 344.650 42.380 344.820 51.410 ;
        RECT 345.530 42.380 345.700 51.410 ;
        RECT 346.410 42.380 346.580 51.410 ;
        RECT 347.290 42.380 347.460 51.410 ;
        RECT 348.170 42.380 348.340 51.410 ;
        RECT 349.050 42.380 349.220 51.410 ;
        RECT 349.930 42.380 350.100 51.410 ;
        RECT 350.810 42.380 350.980 51.410 ;
        RECT 351.690 42.380 351.860 51.410 ;
        RECT 352.570 42.380 352.740 51.410 ;
        RECT 353.450 42.380 353.620 51.410 ;
        RECT 354.330 42.380 354.500 51.410 ;
        RECT 355.210 42.380 355.380 51.410 ;
        RECT 356.090 42.380 356.260 51.410 ;
        RECT 356.970 42.380 357.140 51.410 ;
        RECT 357.850 42.380 358.020 51.410 ;
        RECT 358.730 42.380 358.900 51.410 ;
        RECT 359.610 42.380 359.780 51.410 ;
        RECT 360.490 42.380 360.660 51.410 ;
        RECT 361.370 42.380 361.540 51.410 ;
        RECT 362.250 42.380 362.420 51.410 ;
        RECT 363.130 42.380 363.300 51.410 ;
        RECT 364.010 42.380 364.180 51.410 ;
        RECT 364.890 42.380 365.060 51.410 ;
        RECT 365.770 42.380 365.940 51.410 ;
        RECT 366.650 42.380 366.820 51.410 ;
        RECT 367.530 42.380 367.700 51.410 ;
        RECT 368.410 42.380 368.580 51.410 ;
        RECT 369.290 42.380 369.460 51.410 ;
        RECT 370.170 42.380 370.340 51.410 ;
        RECT 371.050 42.380 371.220 51.410 ;
        RECT 371.930 42.380 372.100 51.410 ;
        RECT 331.790 41.880 333.040 42.210 ;
        RECT 333.550 41.880 334.800 42.210 ;
        RECT 370.510 41.880 371.760 42.210 ;
        RECT 372.560 41.620 372.850 52.170 ;
        RECT 330.700 41.330 372.850 41.620 ;
        RECT 373.360 52.170 403.190 52.460 ;
        RECT 373.360 41.620 373.650 52.170 ;
        RECT 377.970 51.580 379.220 51.910 ;
        RECT 379.730 51.580 380.980 51.910 ;
        RECT 381.490 51.580 382.740 51.910 ;
        RECT 383.250 51.580 384.500 51.910 ;
        RECT 385.010 51.580 386.260 51.910 ;
        RECT 386.770 51.580 388.020 51.910 ;
        RECT 388.530 51.580 389.780 51.910 ;
        RECT 390.290 51.580 391.540 51.910 ;
        RECT 392.050 51.580 393.300 51.910 ;
        RECT 393.810 51.580 395.060 51.910 ;
        RECT 395.570 51.580 396.820 51.910 ;
        RECT 397.330 51.580 398.580 51.910 ;
        RECT 374.110 42.380 374.280 51.410 ;
        RECT 374.990 42.380 375.160 51.410 ;
        RECT 375.870 42.380 376.040 51.410 ;
        RECT 376.750 42.380 376.920 51.410 ;
        RECT 377.630 42.380 377.800 51.410 ;
        RECT 378.510 42.380 378.680 51.410 ;
        RECT 379.390 42.380 379.560 51.410 ;
        RECT 380.270 42.380 380.440 51.410 ;
        RECT 381.150 42.380 381.320 51.410 ;
        RECT 382.030 42.380 382.200 51.410 ;
        RECT 382.910 42.380 383.080 51.410 ;
        RECT 383.790 42.380 383.960 51.410 ;
        RECT 384.670 42.380 384.840 51.410 ;
        RECT 385.550 42.380 385.720 51.410 ;
        RECT 386.430 42.380 386.600 51.410 ;
        RECT 387.310 42.380 387.480 51.410 ;
        RECT 388.190 42.380 388.360 51.410 ;
        RECT 389.070 42.380 389.240 51.410 ;
        RECT 389.950 42.380 390.120 51.410 ;
        RECT 390.830 42.380 391.000 51.410 ;
        RECT 391.710 42.380 391.880 51.410 ;
        RECT 392.590 42.380 392.760 51.410 ;
        RECT 393.470 42.380 393.640 51.410 ;
        RECT 394.350 42.380 394.520 51.410 ;
        RECT 395.230 42.380 395.400 51.410 ;
        RECT 396.110 42.380 396.280 51.410 ;
        RECT 396.990 42.380 397.160 51.410 ;
        RECT 397.870 42.380 398.040 51.410 ;
        RECT 398.750 42.380 398.920 51.410 ;
        RECT 399.630 42.380 399.800 51.410 ;
        RECT 400.510 42.380 400.680 51.410 ;
        RECT 401.390 42.380 401.560 51.410 ;
        RECT 402.270 42.380 402.440 51.410 ;
        RECT 374.450 41.880 375.700 42.210 ;
        RECT 376.210 41.880 377.460 42.210 ;
        RECT 399.090 41.880 400.340 42.210 ;
        RECT 400.850 41.880 402.100 42.210 ;
        RECT 402.900 41.620 403.190 52.170 ;
        RECT 373.360 41.330 403.190 41.620 ;
        RECT 208.045 39.805 237.875 40.095 ;
        RECT 184.845 37.020 207.595 37.190 ;
        RECT 184.845 32.015 185.015 37.020 ;
        RECT 185.915 35.820 187.165 36.150 ;
        RECT 187.675 35.820 188.925 36.150 ;
        RECT 189.435 35.820 190.685 36.150 ;
        RECT 192.955 35.820 194.205 36.150 ;
        RECT 196.475 35.820 197.725 36.150 ;
        RECT 199.995 35.820 201.245 36.150 ;
        RECT 203.515 35.820 204.765 36.150 ;
        RECT 205.275 35.820 206.525 36.150 ;
        RECT 185.575 33.390 185.745 35.650 ;
        RECT 186.455 33.390 186.625 35.650 ;
        RECT 187.335 33.390 187.505 35.650 ;
        RECT 188.215 33.390 188.385 35.650 ;
        RECT 189.095 33.390 189.265 35.650 ;
        RECT 189.975 33.390 190.145 35.650 ;
        RECT 190.855 33.390 191.025 35.650 ;
        RECT 191.735 33.390 191.905 35.650 ;
        RECT 192.615 33.390 192.785 35.650 ;
        RECT 193.495 33.390 193.665 35.650 ;
        RECT 194.375 33.390 194.545 35.650 ;
        RECT 195.255 33.390 195.425 35.650 ;
        RECT 196.135 33.390 196.305 35.650 ;
        RECT 197.015 33.390 197.185 35.650 ;
        RECT 197.895 33.390 198.065 35.650 ;
        RECT 198.775 33.390 198.945 35.650 ;
        RECT 199.655 33.390 199.825 35.650 ;
        RECT 200.535 33.390 200.705 35.650 ;
        RECT 201.415 33.390 201.585 35.650 ;
        RECT 202.295 33.390 202.465 35.650 ;
        RECT 203.175 33.390 203.345 35.650 ;
        RECT 204.055 33.390 204.225 35.650 ;
        RECT 204.935 33.390 205.105 35.650 ;
        RECT 205.815 33.390 205.985 35.650 ;
        RECT 206.695 33.390 206.865 35.650 ;
        RECT 185.915 32.890 187.165 33.220 ;
        RECT 187.675 32.890 188.925 33.220 ;
        RECT 191.195 32.890 192.445 33.220 ;
        RECT 194.715 32.890 195.965 33.220 ;
        RECT 198.235 32.890 199.485 33.220 ;
        RECT 201.755 32.890 203.005 33.220 ;
        RECT 203.515 32.890 204.765 33.220 ;
        RECT 205.275 32.890 206.525 33.220 ;
        RECT 207.425 32.015 207.595 37.020 ;
        RECT 184.845 31.845 207.595 32.015 ;
        RECT 208.045 29.255 208.335 39.805 ;
        RECT 209.135 39.215 210.385 39.545 ;
        RECT 210.895 39.215 212.145 39.545 ;
        RECT 212.655 39.215 213.905 39.545 ;
        RECT 221.455 39.215 222.705 39.545 ;
        RECT 223.215 39.215 224.465 39.545 ;
        RECT 232.015 39.215 233.265 39.545 ;
        RECT 233.775 39.215 235.025 39.545 ;
        RECT 235.535 39.215 236.785 39.545 ;
        RECT 208.795 30.015 208.965 39.045 ;
        RECT 209.675 30.015 209.845 39.045 ;
        RECT 210.555 30.015 210.725 39.045 ;
        RECT 211.435 30.015 211.605 39.045 ;
        RECT 212.315 30.015 212.485 39.045 ;
        RECT 213.195 30.015 213.365 39.045 ;
        RECT 214.075 30.015 214.245 39.045 ;
        RECT 214.955 30.015 215.125 39.045 ;
        RECT 215.835 30.015 216.005 39.045 ;
        RECT 216.715 30.015 216.885 39.045 ;
        RECT 217.595 30.015 217.765 39.045 ;
        RECT 218.475 30.015 218.645 39.045 ;
        RECT 219.355 30.015 219.525 39.045 ;
        RECT 220.235 30.015 220.405 39.045 ;
        RECT 221.115 30.015 221.285 39.045 ;
        RECT 221.995 30.015 222.165 39.045 ;
        RECT 222.875 30.015 223.045 39.045 ;
        RECT 223.755 30.015 223.925 39.045 ;
        RECT 224.635 30.015 224.805 39.045 ;
        RECT 225.515 30.015 225.685 39.045 ;
        RECT 226.395 30.015 226.565 39.045 ;
        RECT 227.275 30.015 227.445 39.045 ;
        RECT 228.155 30.015 228.325 39.045 ;
        RECT 229.035 30.015 229.205 39.045 ;
        RECT 229.915 30.015 230.085 39.045 ;
        RECT 230.795 30.015 230.965 39.045 ;
        RECT 231.675 30.015 231.845 39.045 ;
        RECT 232.555 30.015 232.725 39.045 ;
        RECT 233.435 30.015 233.605 39.045 ;
        RECT 234.315 30.015 234.485 39.045 ;
        RECT 235.195 30.015 235.365 39.045 ;
        RECT 236.075 30.015 236.245 39.045 ;
        RECT 236.955 30.015 237.125 39.045 ;
        RECT 214.415 29.515 215.665 29.845 ;
        RECT 216.175 29.515 217.425 29.845 ;
        RECT 217.935 29.515 219.185 29.845 ;
        RECT 219.695 29.515 220.945 29.845 ;
        RECT 224.975 29.515 226.225 29.845 ;
        RECT 226.735 29.515 227.985 29.845 ;
        RECT 228.495 29.515 229.745 29.845 ;
        RECT 230.255 29.515 231.505 29.845 ;
        RECT 237.585 29.255 237.875 39.805 ;
        RECT 208.045 28.965 237.875 29.255 ;
        RECT 238.385 39.805 280.535 40.095 ;
        RECT 238.385 29.255 238.675 39.805 ;
        RECT 239.475 39.215 240.725 39.545 ;
        RECT 276.435 39.215 277.685 39.545 ;
        RECT 278.195 39.215 279.445 39.545 ;
        RECT 239.135 30.015 239.305 39.045 ;
        RECT 240.015 30.015 240.185 39.045 ;
        RECT 240.895 30.015 241.065 39.045 ;
        RECT 241.775 30.015 241.945 39.045 ;
        RECT 242.655 30.015 242.825 39.045 ;
        RECT 243.535 30.015 243.705 39.045 ;
        RECT 244.415 30.015 244.585 39.045 ;
        RECT 245.295 30.015 245.465 39.045 ;
        RECT 246.175 30.015 246.345 39.045 ;
        RECT 247.055 30.015 247.225 39.045 ;
        RECT 247.935 30.015 248.105 39.045 ;
        RECT 248.815 30.015 248.985 39.045 ;
        RECT 249.695 30.015 249.865 39.045 ;
        RECT 250.575 30.015 250.745 39.045 ;
        RECT 251.455 30.015 251.625 39.045 ;
        RECT 252.335 30.015 252.505 39.045 ;
        RECT 253.215 30.015 253.385 39.045 ;
        RECT 254.095 30.015 254.265 39.045 ;
        RECT 254.975 30.015 255.145 39.045 ;
        RECT 255.855 30.015 256.025 39.045 ;
        RECT 256.735 30.015 256.905 39.045 ;
        RECT 257.615 30.015 257.785 39.045 ;
        RECT 258.495 30.015 258.665 39.045 ;
        RECT 259.375 30.015 259.545 39.045 ;
        RECT 260.255 30.015 260.425 39.045 ;
        RECT 261.135 30.015 261.305 39.045 ;
        RECT 262.015 30.015 262.185 39.045 ;
        RECT 262.895 30.015 263.065 39.045 ;
        RECT 263.775 30.015 263.945 39.045 ;
        RECT 264.655 30.015 264.825 39.045 ;
        RECT 265.535 30.015 265.705 39.045 ;
        RECT 266.415 30.015 266.585 39.045 ;
        RECT 267.295 30.015 267.465 39.045 ;
        RECT 268.175 30.015 268.345 39.045 ;
        RECT 269.055 30.015 269.225 39.045 ;
        RECT 269.935 30.015 270.105 39.045 ;
        RECT 270.815 30.015 270.985 39.045 ;
        RECT 271.695 30.015 271.865 39.045 ;
        RECT 272.575 30.015 272.745 39.045 ;
        RECT 273.455 30.015 273.625 39.045 ;
        RECT 274.335 30.015 274.505 39.045 ;
        RECT 275.215 30.015 275.385 39.045 ;
        RECT 276.095 30.015 276.265 39.045 ;
        RECT 276.975 30.015 277.145 39.045 ;
        RECT 277.855 30.015 278.025 39.045 ;
        RECT 278.735 30.015 278.905 39.045 ;
        RECT 279.615 30.015 279.785 39.045 ;
        RECT 241.235 29.515 242.485 29.845 ;
        RECT 242.995 29.515 244.245 29.845 ;
        RECT 244.755 29.515 246.005 29.845 ;
        RECT 246.515 29.515 247.765 29.845 ;
        RECT 248.275 29.515 249.525 29.845 ;
        RECT 250.035 29.515 251.285 29.845 ;
        RECT 251.795 29.515 253.045 29.845 ;
        RECT 253.555 29.515 254.805 29.845 ;
        RECT 255.315 29.515 256.565 29.845 ;
        RECT 257.075 29.515 258.325 29.845 ;
        RECT 258.835 29.515 260.085 29.845 ;
        RECT 260.595 29.515 261.845 29.845 ;
        RECT 262.355 29.515 263.605 29.845 ;
        RECT 264.115 29.515 265.365 29.845 ;
        RECT 265.875 29.515 267.125 29.845 ;
        RECT 267.635 29.515 268.885 29.845 ;
        RECT 269.395 29.515 270.645 29.845 ;
        RECT 271.155 29.515 272.405 29.845 ;
        RECT 272.915 29.515 274.165 29.845 ;
        RECT 274.675 29.515 275.925 29.845 ;
        RECT 280.245 29.255 280.535 39.805 ;
        RECT 238.385 28.965 280.535 29.255 ;
        RECT 330.700 39.805 372.850 40.095 ;
        RECT 330.700 29.255 330.990 39.805 ;
        RECT 331.790 39.215 333.040 39.545 ;
        RECT 333.550 39.215 334.800 39.545 ;
        RECT 370.510 39.215 371.760 39.545 ;
        RECT 331.450 30.015 331.620 39.045 ;
        RECT 332.330 30.015 332.500 39.045 ;
        RECT 333.210 30.015 333.380 39.045 ;
        RECT 334.090 30.015 334.260 39.045 ;
        RECT 334.970 30.015 335.140 39.045 ;
        RECT 335.850 30.015 336.020 39.045 ;
        RECT 336.730 30.015 336.900 39.045 ;
        RECT 337.610 30.015 337.780 39.045 ;
        RECT 338.490 30.015 338.660 39.045 ;
        RECT 339.370 30.015 339.540 39.045 ;
        RECT 340.250 30.015 340.420 39.045 ;
        RECT 341.130 30.015 341.300 39.045 ;
        RECT 342.010 30.015 342.180 39.045 ;
        RECT 342.890 30.015 343.060 39.045 ;
        RECT 343.770 30.015 343.940 39.045 ;
        RECT 344.650 30.015 344.820 39.045 ;
        RECT 345.530 30.015 345.700 39.045 ;
        RECT 346.410 30.015 346.580 39.045 ;
        RECT 347.290 30.015 347.460 39.045 ;
        RECT 348.170 30.015 348.340 39.045 ;
        RECT 349.050 30.015 349.220 39.045 ;
        RECT 349.930 30.015 350.100 39.045 ;
        RECT 350.810 30.015 350.980 39.045 ;
        RECT 351.690 30.015 351.860 39.045 ;
        RECT 352.570 30.015 352.740 39.045 ;
        RECT 353.450 30.015 353.620 39.045 ;
        RECT 354.330 30.015 354.500 39.045 ;
        RECT 355.210 30.015 355.380 39.045 ;
        RECT 356.090 30.015 356.260 39.045 ;
        RECT 356.970 30.015 357.140 39.045 ;
        RECT 357.850 30.015 358.020 39.045 ;
        RECT 358.730 30.015 358.900 39.045 ;
        RECT 359.610 30.015 359.780 39.045 ;
        RECT 360.490 30.015 360.660 39.045 ;
        RECT 361.370 30.015 361.540 39.045 ;
        RECT 362.250 30.015 362.420 39.045 ;
        RECT 363.130 30.015 363.300 39.045 ;
        RECT 364.010 30.015 364.180 39.045 ;
        RECT 364.890 30.015 365.060 39.045 ;
        RECT 365.770 30.015 365.940 39.045 ;
        RECT 366.650 30.015 366.820 39.045 ;
        RECT 367.530 30.015 367.700 39.045 ;
        RECT 368.410 30.015 368.580 39.045 ;
        RECT 369.290 30.015 369.460 39.045 ;
        RECT 370.170 30.015 370.340 39.045 ;
        RECT 371.050 30.015 371.220 39.045 ;
        RECT 371.930 30.015 372.100 39.045 ;
        RECT 335.310 29.515 336.560 29.845 ;
        RECT 337.070 29.515 338.320 29.845 ;
        RECT 338.830 29.515 340.080 29.845 ;
        RECT 340.590 29.515 341.840 29.845 ;
        RECT 342.350 29.515 343.600 29.845 ;
        RECT 344.110 29.515 345.360 29.845 ;
        RECT 345.870 29.515 347.120 29.845 ;
        RECT 347.630 29.515 348.880 29.845 ;
        RECT 349.390 29.515 350.640 29.845 ;
        RECT 351.150 29.515 352.400 29.845 ;
        RECT 352.910 29.515 354.160 29.845 ;
        RECT 354.670 29.515 355.920 29.845 ;
        RECT 356.430 29.515 357.680 29.845 ;
        RECT 358.190 29.515 359.440 29.845 ;
        RECT 359.950 29.515 361.200 29.845 ;
        RECT 361.710 29.515 362.960 29.845 ;
        RECT 363.470 29.515 364.720 29.845 ;
        RECT 365.230 29.515 366.480 29.845 ;
        RECT 366.990 29.515 368.240 29.845 ;
        RECT 368.750 29.515 370.000 29.845 ;
        RECT 372.560 29.255 372.850 39.805 ;
        RECT 330.700 28.965 372.850 29.255 ;
        RECT 373.360 39.805 403.190 40.095 ;
        RECT 373.360 29.255 373.650 39.805 ;
        RECT 374.450 39.215 375.700 39.545 ;
        RECT 376.210 39.215 377.460 39.545 ;
        RECT 377.970 39.215 379.220 39.545 ;
        RECT 386.770 39.215 388.020 39.545 ;
        RECT 388.530 39.215 389.780 39.545 ;
        RECT 397.330 39.215 398.580 39.545 ;
        RECT 399.090 39.215 400.340 39.545 ;
        RECT 400.850 39.215 402.100 39.545 ;
        RECT 374.110 30.015 374.280 39.045 ;
        RECT 374.990 30.015 375.160 39.045 ;
        RECT 375.870 30.015 376.040 39.045 ;
        RECT 376.750 30.015 376.920 39.045 ;
        RECT 377.630 30.015 377.800 39.045 ;
        RECT 378.510 30.015 378.680 39.045 ;
        RECT 379.390 30.015 379.560 39.045 ;
        RECT 380.270 30.015 380.440 39.045 ;
        RECT 381.150 30.015 381.320 39.045 ;
        RECT 382.030 30.015 382.200 39.045 ;
        RECT 382.910 30.015 383.080 39.045 ;
        RECT 383.790 30.015 383.960 39.045 ;
        RECT 384.670 30.015 384.840 39.045 ;
        RECT 385.550 30.015 385.720 39.045 ;
        RECT 386.430 30.015 386.600 39.045 ;
        RECT 387.310 30.015 387.480 39.045 ;
        RECT 388.190 30.015 388.360 39.045 ;
        RECT 389.070 30.015 389.240 39.045 ;
        RECT 389.950 30.015 390.120 39.045 ;
        RECT 390.830 30.015 391.000 39.045 ;
        RECT 391.710 30.015 391.880 39.045 ;
        RECT 392.590 30.015 392.760 39.045 ;
        RECT 393.470 30.015 393.640 39.045 ;
        RECT 394.350 30.015 394.520 39.045 ;
        RECT 395.230 30.015 395.400 39.045 ;
        RECT 396.110 30.015 396.280 39.045 ;
        RECT 396.990 30.015 397.160 39.045 ;
        RECT 397.870 30.015 398.040 39.045 ;
        RECT 398.750 30.015 398.920 39.045 ;
        RECT 399.630 30.015 399.800 39.045 ;
        RECT 400.510 30.015 400.680 39.045 ;
        RECT 401.390 30.015 401.560 39.045 ;
        RECT 402.270 30.015 402.440 39.045 ;
        RECT 379.730 29.515 380.980 29.845 ;
        RECT 381.490 29.515 382.740 29.845 ;
        RECT 383.250 29.515 384.500 29.845 ;
        RECT 385.010 29.515 386.260 29.845 ;
        RECT 390.290 29.515 391.540 29.845 ;
        RECT 392.050 29.515 393.300 29.845 ;
        RECT 393.810 29.515 395.060 29.845 ;
        RECT 395.570 29.515 396.820 29.845 ;
        RECT 402.900 29.255 403.190 39.805 ;
        RECT 403.640 37.020 426.390 37.190 ;
        RECT 403.640 32.015 403.810 37.020 ;
        RECT 404.710 35.820 405.960 36.150 ;
        RECT 406.470 35.820 407.720 36.150 ;
        RECT 409.990 35.820 411.240 36.150 ;
        RECT 413.510 35.820 414.760 36.150 ;
        RECT 417.030 35.820 418.280 36.150 ;
        RECT 420.550 35.820 421.800 36.150 ;
        RECT 422.310 35.820 423.560 36.150 ;
        RECT 424.070 35.820 425.320 36.150 ;
        RECT 404.370 33.390 404.540 35.650 ;
        RECT 405.250 33.390 405.420 35.650 ;
        RECT 406.130 33.390 406.300 35.650 ;
        RECT 407.010 33.390 407.180 35.650 ;
        RECT 407.890 33.390 408.060 35.650 ;
        RECT 408.770 33.390 408.940 35.650 ;
        RECT 409.650 33.390 409.820 35.650 ;
        RECT 410.530 33.390 410.700 35.650 ;
        RECT 411.410 33.390 411.580 35.650 ;
        RECT 412.290 33.390 412.460 35.650 ;
        RECT 413.170 33.390 413.340 35.650 ;
        RECT 414.050 33.390 414.220 35.650 ;
        RECT 414.930 33.390 415.100 35.650 ;
        RECT 415.810 33.390 415.980 35.650 ;
        RECT 416.690 33.390 416.860 35.650 ;
        RECT 417.570 33.390 417.740 35.650 ;
        RECT 418.450 33.390 418.620 35.650 ;
        RECT 419.330 33.390 419.500 35.650 ;
        RECT 420.210 33.390 420.380 35.650 ;
        RECT 421.090 33.390 421.260 35.650 ;
        RECT 421.970 33.390 422.140 35.650 ;
        RECT 422.850 33.390 423.020 35.650 ;
        RECT 423.730 33.390 423.900 35.650 ;
        RECT 424.610 33.390 424.780 35.650 ;
        RECT 425.490 33.390 425.660 35.650 ;
        RECT 404.710 32.890 405.960 33.220 ;
        RECT 406.470 32.890 407.720 33.220 ;
        RECT 408.230 32.890 409.480 33.220 ;
        RECT 411.750 32.890 413.000 33.220 ;
        RECT 415.270 32.890 416.520 33.220 ;
        RECT 418.790 32.890 420.040 33.220 ;
        RECT 422.310 32.890 423.560 33.220 ;
        RECT 424.070 32.890 425.320 33.220 ;
        RECT 426.220 32.015 426.390 37.020 ;
        RECT 403.640 31.845 426.390 32.015 ;
        RECT 373.360 28.965 403.190 29.255 ;
        RECT 184.845 27.940 207.595 28.110 ;
        RECT 184.845 23.880 185.015 27.940 ;
        RECT 185.915 27.210 187.165 27.540 ;
        RECT 187.675 27.210 188.925 27.540 ;
        RECT 189.435 27.210 190.685 27.540 ;
        RECT 191.195 27.210 192.445 27.540 ;
        RECT 199.995 27.210 201.245 27.540 ;
        RECT 201.755 27.210 203.005 27.540 ;
        RECT 203.515 27.210 204.765 27.540 ;
        RECT 205.275 27.210 206.525 27.540 ;
        RECT 185.575 24.780 185.745 27.040 ;
        RECT 186.455 24.780 186.625 27.040 ;
        RECT 187.335 24.780 187.505 27.040 ;
        RECT 188.215 24.780 188.385 27.040 ;
        RECT 189.095 24.780 189.265 27.040 ;
        RECT 189.975 24.780 190.145 27.040 ;
        RECT 190.855 24.780 191.025 27.040 ;
        RECT 191.735 24.780 191.905 27.040 ;
        RECT 192.615 24.780 192.785 27.040 ;
        RECT 193.495 24.780 193.665 27.040 ;
        RECT 194.375 24.780 194.545 27.040 ;
        RECT 195.255 24.780 195.425 27.040 ;
        RECT 196.135 24.780 196.305 27.040 ;
        RECT 197.015 24.780 197.185 27.040 ;
        RECT 197.895 24.780 198.065 27.040 ;
        RECT 198.775 24.780 198.945 27.040 ;
        RECT 199.655 24.780 199.825 27.040 ;
        RECT 200.535 24.780 200.705 27.040 ;
        RECT 201.415 24.780 201.585 27.040 ;
        RECT 202.295 24.780 202.465 27.040 ;
        RECT 203.175 24.780 203.345 27.040 ;
        RECT 204.055 24.780 204.225 27.040 ;
        RECT 204.935 24.780 205.105 27.040 ;
        RECT 205.815 24.780 205.985 27.040 ;
        RECT 206.695 24.780 206.865 27.040 ;
        RECT 192.955 24.280 194.205 24.610 ;
        RECT 194.715 24.280 195.965 24.610 ;
        RECT 196.475 24.280 197.725 24.610 ;
        RECT 198.235 24.280 199.485 24.610 ;
        RECT 207.425 23.880 207.595 27.940 ;
        RECT 184.845 23.710 207.595 23.880 ;
        RECT 208.065 27.940 237.855 28.110 ;
        RECT 208.065 23.880 208.235 27.940 ;
        RECT 209.135 27.210 210.385 27.540 ;
        RECT 210.895 27.210 212.145 27.540 ;
        RECT 212.655 27.210 213.905 27.540 ;
        RECT 221.455 27.210 222.705 27.540 ;
        RECT 223.215 27.210 224.465 27.540 ;
        RECT 232.015 27.210 233.265 27.540 ;
        RECT 233.775 27.210 235.025 27.540 ;
        RECT 235.535 27.210 236.785 27.540 ;
        RECT 208.795 24.780 208.965 27.040 ;
        RECT 209.675 24.780 209.845 27.040 ;
        RECT 210.555 24.780 210.725 27.040 ;
        RECT 211.435 24.780 211.605 27.040 ;
        RECT 212.315 24.780 212.485 27.040 ;
        RECT 213.195 24.780 213.365 27.040 ;
        RECT 214.075 24.780 214.245 27.040 ;
        RECT 214.955 24.780 215.125 27.040 ;
        RECT 215.835 24.780 216.005 27.040 ;
        RECT 216.715 24.780 216.885 27.040 ;
        RECT 217.595 24.780 217.765 27.040 ;
        RECT 218.475 24.780 218.645 27.040 ;
        RECT 219.355 24.780 219.525 27.040 ;
        RECT 220.235 24.780 220.405 27.040 ;
        RECT 221.115 24.780 221.285 27.040 ;
        RECT 221.995 24.780 222.165 27.040 ;
        RECT 222.875 24.780 223.045 27.040 ;
        RECT 223.755 24.780 223.925 27.040 ;
        RECT 224.635 24.780 224.805 27.040 ;
        RECT 225.515 24.780 225.685 27.040 ;
        RECT 226.395 24.780 226.565 27.040 ;
        RECT 227.275 24.780 227.445 27.040 ;
        RECT 228.155 24.780 228.325 27.040 ;
        RECT 229.035 24.780 229.205 27.040 ;
        RECT 229.915 24.780 230.085 27.040 ;
        RECT 230.795 24.780 230.965 27.040 ;
        RECT 231.675 24.780 231.845 27.040 ;
        RECT 232.555 24.780 232.725 27.040 ;
        RECT 233.435 24.780 233.605 27.040 ;
        RECT 234.315 24.780 234.485 27.040 ;
        RECT 235.195 24.780 235.365 27.040 ;
        RECT 236.075 24.780 236.245 27.040 ;
        RECT 236.955 24.780 237.125 27.040 ;
        RECT 214.415 24.280 215.665 24.610 ;
        RECT 216.175 24.280 217.425 24.610 ;
        RECT 217.935 24.280 219.185 24.610 ;
        RECT 219.695 24.280 220.945 24.610 ;
        RECT 224.975 24.280 226.225 24.610 ;
        RECT 226.735 24.280 227.985 24.610 ;
        RECT 228.495 24.280 229.745 24.610 ;
        RECT 230.255 24.280 231.505 24.610 ;
        RECT 237.685 23.880 237.855 27.940 ;
        RECT 208.065 23.710 237.855 23.880 ;
        RECT 238.405 27.940 280.510 28.110 ;
        RECT 238.405 23.880 238.575 27.940 ;
        RECT 239.475 27.210 240.725 27.540 ;
        RECT 276.435 27.210 277.685 27.540 ;
        RECT 278.195 27.210 279.445 27.540 ;
        RECT 239.135 24.780 239.305 27.040 ;
        RECT 240.015 24.780 240.185 27.040 ;
        RECT 240.895 24.780 241.065 27.040 ;
        RECT 241.775 24.780 241.945 27.040 ;
        RECT 242.655 24.780 242.825 27.040 ;
        RECT 243.535 24.780 243.705 27.040 ;
        RECT 244.415 24.780 244.585 27.040 ;
        RECT 245.295 24.780 245.465 27.040 ;
        RECT 246.175 24.780 246.345 27.040 ;
        RECT 247.055 24.780 247.225 27.040 ;
        RECT 247.935 24.780 248.105 27.040 ;
        RECT 248.815 24.780 248.985 27.040 ;
        RECT 249.695 24.780 249.865 27.040 ;
        RECT 250.575 24.780 250.745 27.040 ;
        RECT 251.455 24.780 251.625 27.040 ;
        RECT 252.335 24.780 252.505 27.040 ;
        RECT 253.215 24.780 253.385 27.040 ;
        RECT 254.095 24.780 254.265 27.040 ;
        RECT 254.975 24.780 255.145 27.040 ;
        RECT 255.855 24.780 256.025 27.040 ;
        RECT 256.735 24.780 256.905 27.040 ;
        RECT 257.615 24.780 257.785 27.040 ;
        RECT 258.495 24.780 258.665 27.040 ;
        RECT 259.375 24.780 259.545 27.040 ;
        RECT 260.255 24.780 260.425 27.040 ;
        RECT 261.135 24.780 261.305 27.040 ;
        RECT 262.015 24.780 262.185 27.040 ;
        RECT 262.895 24.780 263.065 27.040 ;
        RECT 263.775 24.780 263.945 27.040 ;
        RECT 264.655 24.780 264.825 27.040 ;
        RECT 265.535 24.780 265.705 27.040 ;
        RECT 266.415 24.780 266.585 27.040 ;
        RECT 267.295 24.780 267.465 27.040 ;
        RECT 268.175 24.780 268.345 27.040 ;
        RECT 269.055 24.780 269.225 27.040 ;
        RECT 269.935 24.780 270.105 27.040 ;
        RECT 270.815 24.780 270.985 27.040 ;
        RECT 271.695 24.780 271.865 27.040 ;
        RECT 272.575 24.780 272.745 27.040 ;
        RECT 273.455 24.780 273.625 27.040 ;
        RECT 274.335 24.780 274.505 27.040 ;
        RECT 275.215 24.780 275.385 27.040 ;
        RECT 276.095 24.780 276.265 27.040 ;
        RECT 276.975 24.780 277.145 27.040 ;
        RECT 277.855 24.780 278.025 27.040 ;
        RECT 278.735 24.780 278.905 27.040 ;
        RECT 279.615 24.780 279.785 27.040 ;
        RECT 241.235 24.280 242.485 24.610 ;
        RECT 242.995 24.280 244.245 24.610 ;
        RECT 244.755 24.280 246.005 24.610 ;
        RECT 246.515 24.280 247.765 24.610 ;
        RECT 248.275 24.280 249.525 24.610 ;
        RECT 250.035 24.280 251.285 24.610 ;
        RECT 251.795 24.280 253.045 24.610 ;
        RECT 253.555 24.280 254.805 24.610 ;
        RECT 255.315 24.280 256.565 24.610 ;
        RECT 257.075 24.280 258.325 24.610 ;
        RECT 258.835 24.280 260.085 24.610 ;
        RECT 260.595 24.280 261.845 24.610 ;
        RECT 262.355 24.280 263.605 24.610 ;
        RECT 264.115 24.280 265.365 24.610 ;
        RECT 265.875 24.280 267.125 24.610 ;
        RECT 267.635 24.280 268.885 24.610 ;
        RECT 269.395 24.280 270.645 24.610 ;
        RECT 271.155 24.280 272.405 24.610 ;
        RECT 272.915 24.280 274.165 24.610 ;
        RECT 274.675 24.280 275.925 24.610 ;
        RECT 280.340 23.880 280.510 27.940 ;
        RECT 238.405 23.710 280.510 23.880 ;
        RECT 330.725 27.940 372.830 28.110 ;
        RECT 330.725 23.880 330.895 27.940 ;
        RECT 331.790 27.210 333.040 27.540 ;
        RECT 333.550 27.210 334.800 27.540 ;
        RECT 370.510 27.210 371.760 27.540 ;
        RECT 331.450 24.780 331.620 27.040 ;
        RECT 332.330 24.780 332.500 27.040 ;
        RECT 333.210 24.780 333.380 27.040 ;
        RECT 334.090 24.780 334.260 27.040 ;
        RECT 334.970 24.780 335.140 27.040 ;
        RECT 335.850 24.780 336.020 27.040 ;
        RECT 336.730 24.780 336.900 27.040 ;
        RECT 337.610 24.780 337.780 27.040 ;
        RECT 338.490 24.780 338.660 27.040 ;
        RECT 339.370 24.780 339.540 27.040 ;
        RECT 340.250 24.780 340.420 27.040 ;
        RECT 341.130 24.780 341.300 27.040 ;
        RECT 342.010 24.780 342.180 27.040 ;
        RECT 342.890 24.780 343.060 27.040 ;
        RECT 343.770 24.780 343.940 27.040 ;
        RECT 344.650 24.780 344.820 27.040 ;
        RECT 345.530 24.780 345.700 27.040 ;
        RECT 346.410 24.780 346.580 27.040 ;
        RECT 347.290 24.780 347.460 27.040 ;
        RECT 348.170 24.780 348.340 27.040 ;
        RECT 349.050 24.780 349.220 27.040 ;
        RECT 349.930 24.780 350.100 27.040 ;
        RECT 350.810 24.780 350.980 27.040 ;
        RECT 351.690 24.780 351.860 27.040 ;
        RECT 352.570 24.780 352.740 27.040 ;
        RECT 353.450 24.780 353.620 27.040 ;
        RECT 354.330 24.780 354.500 27.040 ;
        RECT 355.210 24.780 355.380 27.040 ;
        RECT 356.090 24.780 356.260 27.040 ;
        RECT 356.970 24.780 357.140 27.040 ;
        RECT 357.850 24.780 358.020 27.040 ;
        RECT 358.730 24.780 358.900 27.040 ;
        RECT 359.610 24.780 359.780 27.040 ;
        RECT 360.490 24.780 360.660 27.040 ;
        RECT 361.370 24.780 361.540 27.040 ;
        RECT 362.250 24.780 362.420 27.040 ;
        RECT 363.130 24.780 363.300 27.040 ;
        RECT 364.010 24.780 364.180 27.040 ;
        RECT 364.890 24.780 365.060 27.040 ;
        RECT 365.770 24.780 365.940 27.040 ;
        RECT 366.650 24.780 366.820 27.040 ;
        RECT 367.530 24.780 367.700 27.040 ;
        RECT 368.410 24.780 368.580 27.040 ;
        RECT 369.290 24.780 369.460 27.040 ;
        RECT 370.170 24.780 370.340 27.040 ;
        RECT 371.050 24.780 371.220 27.040 ;
        RECT 371.930 24.780 372.100 27.040 ;
        RECT 335.310 24.280 336.560 24.610 ;
        RECT 337.070 24.280 338.320 24.610 ;
        RECT 338.830 24.280 340.080 24.610 ;
        RECT 340.590 24.280 341.840 24.610 ;
        RECT 342.350 24.280 343.600 24.610 ;
        RECT 344.110 24.280 345.360 24.610 ;
        RECT 345.870 24.280 347.120 24.610 ;
        RECT 347.630 24.280 348.880 24.610 ;
        RECT 349.390 24.280 350.640 24.610 ;
        RECT 351.150 24.280 352.400 24.610 ;
        RECT 352.910 24.280 354.160 24.610 ;
        RECT 354.670 24.280 355.920 24.610 ;
        RECT 356.430 24.280 357.680 24.610 ;
        RECT 358.190 24.280 359.440 24.610 ;
        RECT 359.950 24.280 361.200 24.610 ;
        RECT 361.710 24.280 362.960 24.610 ;
        RECT 363.470 24.280 364.720 24.610 ;
        RECT 365.230 24.280 366.480 24.610 ;
        RECT 366.990 24.280 368.240 24.610 ;
        RECT 368.750 24.280 370.000 24.610 ;
        RECT 372.660 23.880 372.830 27.940 ;
        RECT 330.725 23.710 372.830 23.880 ;
        RECT 373.380 27.940 403.170 28.110 ;
        RECT 373.380 23.880 373.550 27.940 ;
        RECT 374.450 27.210 375.700 27.540 ;
        RECT 376.210 27.210 377.460 27.540 ;
        RECT 377.970 27.210 379.220 27.540 ;
        RECT 386.770 27.210 388.020 27.540 ;
        RECT 388.530 27.210 389.780 27.540 ;
        RECT 397.330 27.210 398.580 27.540 ;
        RECT 399.090 27.210 400.340 27.540 ;
        RECT 400.850 27.210 402.100 27.540 ;
        RECT 374.110 24.780 374.280 27.040 ;
        RECT 374.990 24.780 375.160 27.040 ;
        RECT 375.870 24.780 376.040 27.040 ;
        RECT 376.750 24.780 376.920 27.040 ;
        RECT 377.630 24.780 377.800 27.040 ;
        RECT 378.510 24.780 378.680 27.040 ;
        RECT 379.390 24.780 379.560 27.040 ;
        RECT 380.270 24.780 380.440 27.040 ;
        RECT 381.150 24.780 381.320 27.040 ;
        RECT 382.030 24.780 382.200 27.040 ;
        RECT 382.910 24.780 383.080 27.040 ;
        RECT 383.790 24.780 383.960 27.040 ;
        RECT 384.670 24.780 384.840 27.040 ;
        RECT 385.550 24.780 385.720 27.040 ;
        RECT 386.430 24.780 386.600 27.040 ;
        RECT 387.310 24.780 387.480 27.040 ;
        RECT 388.190 24.780 388.360 27.040 ;
        RECT 389.070 24.780 389.240 27.040 ;
        RECT 389.950 24.780 390.120 27.040 ;
        RECT 390.830 24.780 391.000 27.040 ;
        RECT 391.710 24.780 391.880 27.040 ;
        RECT 392.590 24.780 392.760 27.040 ;
        RECT 393.470 24.780 393.640 27.040 ;
        RECT 394.350 24.780 394.520 27.040 ;
        RECT 395.230 24.780 395.400 27.040 ;
        RECT 396.110 24.780 396.280 27.040 ;
        RECT 396.990 24.780 397.160 27.040 ;
        RECT 397.870 24.780 398.040 27.040 ;
        RECT 398.750 24.780 398.920 27.040 ;
        RECT 399.630 24.780 399.800 27.040 ;
        RECT 400.510 24.780 400.680 27.040 ;
        RECT 401.390 24.780 401.560 27.040 ;
        RECT 402.270 24.780 402.440 27.040 ;
        RECT 379.730 24.280 380.980 24.610 ;
        RECT 381.490 24.280 382.740 24.610 ;
        RECT 383.250 24.280 384.500 24.610 ;
        RECT 385.010 24.280 386.260 24.610 ;
        RECT 390.290 24.280 391.540 24.610 ;
        RECT 392.050 24.280 393.300 24.610 ;
        RECT 393.810 24.280 395.060 24.610 ;
        RECT 395.570 24.280 396.820 24.610 ;
        RECT 403.000 23.880 403.170 27.940 ;
        RECT 373.380 23.710 403.170 23.880 ;
        RECT 403.640 27.940 426.390 28.110 ;
        RECT 403.640 23.880 403.810 27.940 ;
        RECT 404.710 27.210 405.960 27.540 ;
        RECT 406.470 27.210 407.720 27.540 ;
        RECT 408.230 27.210 409.480 27.540 ;
        RECT 409.990 27.210 411.240 27.540 ;
        RECT 418.790 27.210 420.040 27.540 ;
        RECT 420.550 27.210 421.800 27.540 ;
        RECT 422.310 27.210 423.560 27.540 ;
        RECT 424.070 27.210 425.320 27.540 ;
        RECT 404.370 24.780 404.540 27.040 ;
        RECT 405.250 24.780 405.420 27.040 ;
        RECT 406.130 24.780 406.300 27.040 ;
        RECT 407.010 24.780 407.180 27.040 ;
        RECT 407.890 24.780 408.060 27.040 ;
        RECT 408.770 24.780 408.940 27.040 ;
        RECT 409.650 24.780 409.820 27.040 ;
        RECT 410.530 24.780 410.700 27.040 ;
        RECT 411.410 24.780 411.580 27.040 ;
        RECT 412.290 24.780 412.460 27.040 ;
        RECT 413.170 24.780 413.340 27.040 ;
        RECT 414.050 24.780 414.220 27.040 ;
        RECT 414.930 24.780 415.100 27.040 ;
        RECT 415.810 24.780 415.980 27.040 ;
        RECT 416.690 24.780 416.860 27.040 ;
        RECT 417.570 24.780 417.740 27.040 ;
        RECT 418.450 24.780 418.620 27.040 ;
        RECT 419.330 24.780 419.500 27.040 ;
        RECT 420.210 24.780 420.380 27.040 ;
        RECT 421.090 24.780 421.260 27.040 ;
        RECT 421.970 24.780 422.140 27.040 ;
        RECT 422.850 24.780 423.020 27.040 ;
        RECT 423.730 24.780 423.900 27.040 ;
        RECT 424.610 24.780 424.780 27.040 ;
        RECT 425.490 24.780 425.660 27.040 ;
        RECT 411.750 24.280 413.000 24.610 ;
        RECT 413.510 24.280 414.760 24.610 ;
        RECT 415.270 24.280 416.520 24.610 ;
        RECT 417.030 24.280 418.280 24.610 ;
        RECT 426.220 23.880 426.390 27.940 ;
        RECT 403.640 23.710 426.390 23.880 ;
        RECT 184.845 21.455 207.595 21.625 ;
        RECT 184.845 17.395 185.015 21.455 ;
        RECT 185.915 20.725 187.165 21.055 ;
        RECT 187.675 20.725 188.925 21.055 ;
        RECT 189.435 20.725 190.685 21.055 ;
        RECT 191.195 20.725 192.445 21.055 ;
        RECT 199.995 20.725 201.245 21.055 ;
        RECT 201.755 20.725 203.005 21.055 ;
        RECT 203.515 20.725 204.765 21.055 ;
        RECT 205.275 20.725 206.525 21.055 ;
        RECT 185.575 18.295 185.745 20.555 ;
        RECT 186.455 18.295 186.625 20.555 ;
        RECT 187.335 18.295 187.505 20.555 ;
        RECT 188.215 18.295 188.385 20.555 ;
        RECT 189.095 18.295 189.265 20.555 ;
        RECT 189.975 18.295 190.145 20.555 ;
        RECT 190.855 18.295 191.025 20.555 ;
        RECT 191.735 18.295 191.905 20.555 ;
        RECT 192.615 18.295 192.785 20.555 ;
        RECT 193.495 18.295 193.665 20.555 ;
        RECT 194.375 18.295 194.545 20.555 ;
        RECT 195.255 18.295 195.425 20.555 ;
        RECT 196.135 18.295 196.305 20.555 ;
        RECT 197.015 18.295 197.185 20.555 ;
        RECT 197.895 18.295 198.065 20.555 ;
        RECT 198.775 18.295 198.945 20.555 ;
        RECT 199.655 18.295 199.825 20.555 ;
        RECT 200.535 18.295 200.705 20.555 ;
        RECT 201.415 18.295 201.585 20.555 ;
        RECT 202.295 18.295 202.465 20.555 ;
        RECT 203.175 18.295 203.345 20.555 ;
        RECT 204.055 18.295 204.225 20.555 ;
        RECT 204.935 18.295 205.105 20.555 ;
        RECT 205.815 18.295 205.985 20.555 ;
        RECT 206.695 18.295 206.865 20.555 ;
        RECT 192.955 17.795 194.205 18.125 ;
        RECT 194.715 17.795 195.965 18.125 ;
        RECT 196.475 17.795 197.725 18.125 ;
        RECT 198.235 17.795 199.485 18.125 ;
        RECT 207.425 17.395 207.595 21.455 ;
        RECT 184.845 17.225 207.595 17.395 ;
        RECT 208.065 21.455 237.855 21.625 ;
        RECT 208.065 17.395 208.235 21.455 ;
        RECT 209.135 20.725 210.385 21.055 ;
        RECT 210.895 20.725 212.145 21.055 ;
        RECT 212.655 20.725 213.905 21.055 ;
        RECT 214.415 20.725 215.665 21.055 ;
        RECT 216.175 20.725 217.425 21.055 ;
        RECT 217.935 20.725 219.185 21.055 ;
        RECT 219.695 20.725 220.945 21.055 ;
        RECT 224.975 20.725 226.225 21.055 ;
        RECT 226.735 20.725 227.985 21.055 ;
        RECT 228.495 20.725 229.745 21.055 ;
        RECT 230.255 20.725 231.505 21.055 ;
        RECT 232.015 20.725 233.265 21.055 ;
        RECT 233.775 20.725 235.025 21.055 ;
        RECT 235.535 20.725 236.785 21.055 ;
        RECT 208.795 18.295 208.965 20.555 ;
        RECT 209.675 18.295 209.845 20.555 ;
        RECT 210.555 18.295 210.725 20.555 ;
        RECT 211.435 18.295 211.605 20.555 ;
        RECT 212.315 18.295 212.485 20.555 ;
        RECT 213.195 18.295 213.365 20.555 ;
        RECT 214.075 18.295 214.245 20.555 ;
        RECT 214.955 18.295 215.125 20.555 ;
        RECT 215.835 18.295 216.005 20.555 ;
        RECT 216.715 18.295 216.885 20.555 ;
        RECT 217.595 18.295 217.765 20.555 ;
        RECT 218.475 18.295 218.645 20.555 ;
        RECT 219.355 18.295 219.525 20.555 ;
        RECT 220.235 18.295 220.405 20.555 ;
        RECT 221.115 18.295 221.285 20.555 ;
        RECT 221.995 18.295 222.165 20.555 ;
        RECT 222.875 18.295 223.045 20.555 ;
        RECT 223.755 18.295 223.925 20.555 ;
        RECT 224.635 18.295 224.805 20.555 ;
        RECT 225.515 18.295 225.685 20.555 ;
        RECT 226.395 18.295 226.565 20.555 ;
        RECT 227.275 18.295 227.445 20.555 ;
        RECT 228.155 18.295 228.325 20.555 ;
        RECT 229.035 18.295 229.205 20.555 ;
        RECT 229.915 18.295 230.085 20.555 ;
        RECT 230.795 18.295 230.965 20.555 ;
        RECT 231.675 18.295 231.845 20.555 ;
        RECT 232.555 18.295 232.725 20.555 ;
        RECT 233.435 18.295 233.605 20.555 ;
        RECT 234.315 18.295 234.485 20.555 ;
        RECT 235.195 18.295 235.365 20.555 ;
        RECT 236.075 18.295 236.245 20.555 ;
        RECT 236.955 18.295 237.125 20.555 ;
        RECT 221.455 17.795 222.705 18.125 ;
        RECT 223.215 17.795 224.465 18.125 ;
        RECT 237.685 17.395 237.855 21.455 ;
        RECT 208.065 17.225 237.855 17.395 ;
        RECT 238.405 21.455 280.510 21.625 ;
        RECT 238.405 17.395 238.575 21.455 ;
        RECT 239.475 20.725 240.725 21.055 ;
        RECT 241.235 20.725 242.485 21.055 ;
        RECT 242.995 20.725 244.245 21.055 ;
        RECT 244.755 20.725 246.005 21.055 ;
        RECT 246.515 20.725 247.765 21.055 ;
        RECT 248.275 20.725 249.525 21.055 ;
        RECT 250.035 20.725 251.285 21.055 ;
        RECT 251.795 20.725 253.045 21.055 ;
        RECT 253.555 20.725 254.805 21.055 ;
        RECT 255.315 20.725 256.565 21.055 ;
        RECT 257.075 20.725 258.325 21.055 ;
        RECT 258.835 20.725 260.085 21.055 ;
        RECT 260.595 20.725 261.845 21.055 ;
        RECT 262.355 20.725 263.605 21.055 ;
        RECT 264.115 20.725 265.365 21.055 ;
        RECT 265.875 20.725 267.125 21.055 ;
        RECT 267.635 20.725 268.885 21.055 ;
        RECT 269.395 20.725 270.645 21.055 ;
        RECT 271.155 20.725 272.405 21.055 ;
        RECT 272.915 20.725 274.165 21.055 ;
        RECT 274.675 20.725 275.925 21.055 ;
        RECT 276.435 20.725 277.685 21.055 ;
        RECT 278.195 20.725 279.445 21.055 ;
        RECT 239.135 18.295 239.305 20.555 ;
        RECT 240.015 18.295 240.185 20.555 ;
        RECT 240.895 18.295 241.065 20.555 ;
        RECT 241.775 18.295 241.945 20.555 ;
        RECT 242.655 18.295 242.825 20.555 ;
        RECT 243.535 18.295 243.705 20.555 ;
        RECT 244.415 18.295 244.585 20.555 ;
        RECT 245.295 18.295 245.465 20.555 ;
        RECT 246.175 18.295 246.345 20.555 ;
        RECT 247.055 18.295 247.225 20.555 ;
        RECT 247.935 18.295 248.105 20.555 ;
        RECT 248.815 18.295 248.985 20.555 ;
        RECT 249.695 18.295 249.865 20.555 ;
        RECT 250.575 18.295 250.745 20.555 ;
        RECT 251.455 18.295 251.625 20.555 ;
        RECT 252.335 18.295 252.505 20.555 ;
        RECT 253.215 18.295 253.385 20.555 ;
        RECT 254.095 18.295 254.265 20.555 ;
        RECT 254.975 18.295 255.145 20.555 ;
        RECT 255.855 18.295 256.025 20.555 ;
        RECT 256.735 18.295 256.905 20.555 ;
        RECT 257.615 18.295 257.785 20.555 ;
        RECT 258.495 18.295 258.665 20.555 ;
        RECT 259.375 18.295 259.545 20.555 ;
        RECT 260.255 18.295 260.425 20.555 ;
        RECT 261.135 18.295 261.305 20.555 ;
        RECT 262.015 18.295 262.185 20.555 ;
        RECT 262.895 18.295 263.065 20.555 ;
        RECT 263.775 18.295 263.945 20.555 ;
        RECT 264.655 18.295 264.825 20.555 ;
        RECT 265.535 18.295 265.705 20.555 ;
        RECT 266.415 18.295 266.585 20.555 ;
        RECT 267.295 18.295 267.465 20.555 ;
        RECT 268.175 18.295 268.345 20.555 ;
        RECT 269.055 18.295 269.225 20.555 ;
        RECT 269.935 18.295 270.105 20.555 ;
        RECT 270.815 18.295 270.985 20.555 ;
        RECT 271.695 18.295 271.865 20.555 ;
        RECT 272.575 18.295 272.745 20.555 ;
        RECT 273.455 18.295 273.625 20.555 ;
        RECT 274.335 18.295 274.505 20.555 ;
        RECT 275.215 18.295 275.385 20.555 ;
        RECT 276.095 18.295 276.265 20.555 ;
        RECT 276.975 18.295 277.145 20.555 ;
        RECT 277.855 18.295 278.025 20.555 ;
        RECT 278.735 18.295 278.905 20.555 ;
        RECT 279.615 18.295 279.785 20.555 ;
        RECT 280.340 17.395 280.510 21.455 ;
        RECT 238.405 17.225 280.510 17.395 ;
        RECT 330.725 21.455 372.830 21.625 ;
        RECT 330.725 17.395 330.895 21.455 ;
        RECT 331.790 20.725 333.040 21.055 ;
        RECT 333.550 20.725 334.800 21.055 ;
        RECT 335.310 20.725 336.560 21.055 ;
        RECT 337.070 20.725 338.320 21.055 ;
        RECT 338.830 20.725 340.080 21.055 ;
        RECT 340.590 20.725 341.840 21.055 ;
        RECT 342.350 20.725 343.600 21.055 ;
        RECT 344.110 20.725 345.360 21.055 ;
        RECT 345.870 20.725 347.120 21.055 ;
        RECT 347.630 20.725 348.880 21.055 ;
        RECT 349.390 20.725 350.640 21.055 ;
        RECT 351.150 20.725 352.400 21.055 ;
        RECT 352.910 20.725 354.160 21.055 ;
        RECT 354.670 20.725 355.920 21.055 ;
        RECT 356.430 20.725 357.680 21.055 ;
        RECT 358.190 20.725 359.440 21.055 ;
        RECT 359.950 20.725 361.200 21.055 ;
        RECT 361.710 20.725 362.960 21.055 ;
        RECT 363.470 20.725 364.720 21.055 ;
        RECT 365.230 20.725 366.480 21.055 ;
        RECT 366.990 20.725 368.240 21.055 ;
        RECT 368.750 20.725 370.000 21.055 ;
        RECT 370.510 20.725 371.760 21.055 ;
        RECT 331.450 18.295 331.620 20.555 ;
        RECT 332.330 18.295 332.500 20.555 ;
        RECT 333.210 18.295 333.380 20.555 ;
        RECT 334.090 18.295 334.260 20.555 ;
        RECT 334.970 18.295 335.140 20.555 ;
        RECT 335.850 18.295 336.020 20.555 ;
        RECT 336.730 18.295 336.900 20.555 ;
        RECT 337.610 18.295 337.780 20.555 ;
        RECT 338.490 18.295 338.660 20.555 ;
        RECT 339.370 18.295 339.540 20.555 ;
        RECT 340.250 18.295 340.420 20.555 ;
        RECT 341.130 18.295 341.300 20.555 ;
        RECT 342.010 18.295 342.180 20.555 ;
        RECT 342.890 18.295 343.060 20.555 ;
        RECT 343.770 18.295 343.940 20.555 ;
        RECT 344.650 18.295 344.820 20.555 ;
        RECT 345.530 18.295 345.700 20.555 ;
        RECT 346.410 18.295 346.580 20.555 ;
        RECT 347.290 18.295 347.460 20.555 ;
        RECT 348.170 18.295 348.340 20.555 ;
        RECT 349.050 18.295 349.220 20.555 ;
        RECT 349.930 18.295 350.100 20.555 ;
        RECT 350.810 18.295 350.980 20.555 ;
        RECT 351.690 18.295 351.860 20.555 ;
        RECT 352.570 18.295 352.740 20.555 ;
        RECT 353.450 18.295 353.620 20.555 ;
        RECT 354.330 18.295 354.500 20.555 ;
        RECT 355.210 18.295 355.380 20.555 ;
        RECT 356.090 18.295 356.260 20.555 ;
        RECT 356.970 18.295 357.140 20.555 ;
        RECT 357.850 18.295 358.020 20.555 ;
        RECT 358.730 18.295 358.900 20.555 ;
        RECT 359.610 18.295 359.780 20.555 ;
        RECT 360.490 18.295 360.660 20.555 ;
        RECT 361.370 18.295 361.540 20.555 ;
        RECT 362.250 18.295 362.420 20.555 ;
        RECT 363.130 18.295 363.300 20.555 ;
        RECT 364.010 18.295 364.180 20.555 ;
        RECT 364.890 18.295 365.060 20.555 ;
        RECT 365.770 18.295 365.940 20.555 ;
        RECT 366.650 18.295 366.820 20.555 ;
        RECT 367.530 18.295 367.700 20.555 ;
        RECT 368.410 18.295 368.580 20.555 ;
        RECT 369.290 18.295 369.460 20.555 ;
        RECT 370.170 18.295 370.340 20.555 ;
        RECT 371.050 18.295 371.220 20.555 ;
        RECT 371.930 18.295 372.100 20.555 ;
        RECT 372.660 17.395 372.830 21.455 ;
        RECT 330.725 17.225 372.830 17.395 ;
        RECT 373.380 21.455 403.170 21.625 ;
        RECT 373.380 17.395 373.550 21.455 ;
        RECT 374.450 20.725 375.700 21.055 ;
        RECT 376.210 20.725 377.460 21.055 ;
        RECT 377.970 20.725 379.220 21.055 ;
        RECT 379.730 20.725 380.980 21.055 ;
        RECT 381.490 20.725 382.740 21.055 ;
        RECT 383.250 20.725 384.500 21.055 ;
        RECT 385.010 20.725 386.260 21.055 ;
        RECT 390.290 20.725 391.540 21.055 ;
        RECT 392.050 20.725 393.300 21.055 ;
        RECT 393.810 20.725 395.060 21.055 ;
        RECT 395.570 20.725 396.820 21.055 ;
        RECT 397.330 20.725 398.580 21.055 ;
        RECT 399.090 20.725 400.340 21.055 ;
        RECT 400.850 20.725 402.100 21.055 ;
        RECT 374.110 18.295 374.280 20.555 ;
        RECT 374.990 18.295 375.160 20.555 ;
        RECT 375.870 18.295 376.040 20.555 ;
        RECT 376.750 18.295 376.920 20.555 ;
        RECT 377.630 18.295 377.800 20.555 ;
        RECT 378.510 18.295 378.680 20.555 ;
        RECT 379.390 18.295 379.560 20.555 ;
        RECT 380.270 18.295 380.440 20.555 ;
        RECT 381.150 18.295 381.320 20.555 ;
        RECT 382.030 18.295 382.200 20.555 ;
        RECT 382.910 18.295 383.080 20.555 ;
        RECT 383.790 18.295 383.960 20.555 ;
        RECT 384.670 18.295 384.840 20.555 ;
        RECT 385.550 18.295 385.720 20.555 ;
        RECT 386.430 18.295 386.600 20.555 ;
        RECT 387.310 18.295 387.480 20.555 ;
        RECT 388.190 18.295 388.360 20.555 ;
        RECT 389.070 18.295 389.240 20.555 ;
        RECT 389.950 18.295 390.120 20.555 ;
        RECT 390.830 18.295 391.000 20.555 ;
        RECT 391.710 18.295 391.880 20.555 ;
        RECT 392.590 18.295 392.760 20.555 ;
        RECT 393.470 18.295 393.640 20.555 ;
        RECT 394.350 18.295 394.520 20.555 ;
        RECT 395.230 18.295 395.400 20.555 ;
        RECT 396.110 18.295 396.280 20.555 ;
        RECT 396.990 18.295 397.160 20.555 ;
        RECT 397.870 18.295 398.040 20.555 ;
        RECT 398.750 18.295 398.920 20.555 ;
        RECT 399.630 18.295 399.800 20.555 ;
        RECT 400.510 18.295 400.680 20.555 ;
        RECT 401.390 18.295 401.560 20.555 ;
        RECT 402.270 18.295 402.440 20.555 ;
        RECT 386.770 17.795 388.020 18.125 ;
        RECT 388.530 17.795 389.780 18.125 ;
        RECT 403.000 17.395 403.170 21.455 ;
        RECT 373.380 17.225 403.170 17.395 ;
        RECT 403.640 21.455 426.390 21.625 ;
        RECT 403.640 17.395 403.810 21.455 ;
        RECT 404.710 20.725 405.960 21.055 ;
        RECT 406.470 20.725 407.720 21.055 ;
        RECT 408.230 20.725 409.480 21.055 ;
        RECT 409.990 20.725 411.240 21.055 ;
        RECT 418.790 20.725 420.040 21.055 ;
        RECT 420.550 20.725 421.800 21.055 ;
        RECT 422.310 20.725 423.560 21.055 ;
        RECT 424.070 20.725 425.320 21.055 ;
        RECT 404.370 18.295 404.540 20.555 ;
        RECT 405.250 18.295 405.420 20.555 ;
        RECT 406.130 18.295 406.300 20.555 ;
        RECT 407.010 18.295 407.180 20.555 ;
        RECT 407.890 18.295 408.060 20.555 ;
        RECT 408.770 18.295 408.940 20.555 ;
        RECT 409.650 18.295 409.820 20.555 ;
        RECT 410.530 18.295 410.700 20.555 ;
        RECT 411.410 18.295 411.580 20.555 ;
        RECT 412.290 18.295 412.460 20.555 ;
        RECT 413.170 18.295 413.340 20.555 ;
        RECT 414.050 18.295 414.220 20.555 ;
        RECT 414.930 18.295 415.100 20.555 ;
        RECT 415.810 18.295 415.980 20.555 ;
        RECT 416.690 18.295 416.860 20.555 ;
        RECT 417.570 18.295 417.740 20.555 ;
        RECT 418.450 18.295 418.620 20.555 ;
        RECT 419.330 18.295 419.500 20.555 ;
        RECT 420.210 18.295 420.380 20.555 ;
        RECT 421.090 18.295 421.260 20.555 ;
        RECT 421.970 18.295 422.140 20.555 ;
        RECT 422.850 18.295 423.020 20.555 ;
        RECT 423.730 18.295 423.900 20.555 ;
        RECT 424.610 18.295 424.780 20.555 ;
        RECT 425.490 18.295 425.660 20.555 ;
        RECT 411.750 17.795 413.000 18.125 ;
        RECT 413.510 17.795 414.760 18.125 ;
        RECT 415.270 17.795 416.520 18.125 ;
        RECT 417.030 17.795 418.280 18.125 ;
        RECT 426.220 17.395 426.390 21.455 ;
        RECT 403.640 17.225 426.390 17.395 ;
      LAYER met1 ;
        RECT 74.400 209.365 116.550 209.655 ;
        RECT 74.400 199.385 74.690 209.365 ;
        RECT 78.980 208.755 113.730 209.085 ;
        RECT 75.095 199.575 75.375 208.605 ;
        RECT 75.975 199.575 76.255 208.605 ;
        RECT 76.855 199.575 77.135 208.605 ;
        RECT 77.735 199.575 78.015 208.605 ;
        RECT 78.615 199.575 78.895 208.605 ;
        RECT 79.495 199.575 79.775 208.605 ;
        RECT 80.375 199.575 80.655 208.605 ;
        RECT 81.255 199.575 81.535 208.605 ;
        RECT 82.135 199.575 82.415 208.605 ;
        RECT 83.015 199.575 83.295 208.605 ;
        RECT 83.895 199.575 84.175 208.605 ;
        RECT 84.775 199.575 85.055 208.605 ;
        RECT 85.655 199.575 85.935 208.605 ;
        RECT 86.535 199.575 86.815 208.605 ;
        RECT 87.415 199.575 87.695 208.605 ;
        RECT 88.295 199.575 88.575 208.605 ;
        RECT 89.175 199.575 89.455 208.605 ;
        RECT 90.055 199.575 90.335 208.605 ;
        RECT 90.935 199.575 91.215 208.605 ;
        RECT 91.815 199.575 92.095 208.605 ;
        RECT 92.695 199.575 92.975 208.605 ;
        RECT 93.575 199.575 93.855 208.605 ;
        RECT 94.455 199.575 94.735 208.605 ;
        RECT 95.335 199.575 95.615 208.605 ;
        RECT 96.215 199.575 96.495 208.605 ;
        RECT 97.095 199.575 97.375 208.605 ;
        RECT 97.975 199.575 98.255 208.605 ;
        RECT 98.855 199.575 99.135 208.605 ;
        RECT 99.735 199.575 100.015 208.605 ;
        RECT 100.615 199.575 100.895 208.605 ;
        RECT 101.495 199.575 101.775 208.605 ;
        RECT 102.375 199.575 102.655 208.605 ;
        RECT 103.255 199.575 103.535 208.605 ;
        RECT 104.135 199.575 104.415 208.605 ;
        RECT 105.015 199.575 105.295 208.605 ;
        RECT 105.895 199.575 106.175 208.605 ;
        RECT 106.775 199.575 107.055 208.605 ;
        RECT 107.655 199.575 107.935 208.605 ;
        RECT 108.535 199.575 108.815 208.605 ;
        RECT 109.415 199.575 109.695 208.605 ;
        RECT 110.295 199.575 110.575 208.605 ;
        RECT 111.175 199.575 111.455 208.605 ;
        RECT 112.055 199.575 112.335 208.605 ;
        RECT 112.935 199.575 113.215 208.605 ;
        RECT 113.815 199.575 114.095 208.605 ;
        RECT 114.695 199.575 114.975 208.605 ;
        RECT 115.575 199.575 115.855 208.605 ;
        RECT 116.260 199.385 116.550 209.365 ;
        RECT 74.400 199.095 78.530 199.385 ;
        RECT 114.180 199.095 116.550 199.385 ;
        RECT 74.400 198.815 74.690 199.095 ;
        RECT 116.260 198.815 116.550 199.095 ;
        RECT 74.400 198.525 116.550 198.815 ;
        RECT 117.060 209.365 146.890 209.655 ;
        RECT 117.060 199.385 117.350 209.365 ;
        RECT 121.640 208.755 142.310 209.085 ;
        RECT 117.755 199.575 118.035 208.605 ;
        RECT 118.635 199.575 118.915 208.605 ;
        RECT 119.515 199.575 119.795 208.605 ;
        RECT 120.395 199.575 120.675 208.605 ;
        RECT 121.275 199.575 121.555 208.605 ;
        RECT 122.155 199.575 122.435 208.605 ;
        RECT 123.035 199.575 123.315 208.605 ;
        RECT 123.915 199.575 124.195 208.605 ;
        RECT 124.795 199.575 125.075 208.605 ;
        RECT 125.675 199.575 125.955 208.605 ;
        RECT 126.555 199.575 126.835 208.605 ;
        RECT 127.435 199.575 127.715 208.605 ;
        RECT 128.315 199.575 128.595 208.605 ;
        RECT 129.195 199.575 129.475 208.605 ;
        RECT 130.075 199.575 130.355 208.605 ;
        RECT 130.955 199.575 131.235 208.605 ;
        RECT 131.835 199.575 132.115 208.605 ;
        RECT 132.715 199.575 132.995 208.605 ;
        RECT 133.595 199.575 133.875 208.605 ;
        RECT 134.475 199.575 134.755 208.605 ;
        RECT 135.355 199.575 135.635 208.605 ;
        RECT 136.235 199.575 136.515 208.605 ;
        RECT 137.115 199.575 137.395 208.605 ;
        RECT 137.995 199.575 138.275 208.605 ;
        RECT 138.875 199.575 139.155 208.605 ;
        RECT 139.755 199.575 140.035 208.605 ;
        RECT 140.635 199.575 140.915 208.605 ;
        RECT 141.515 199.575 141.795 208.605 ;
        RECT 142.395 199.575 142.675 208.605 ;
        RECT 143.275 199.575 143.555 208.605 ;
        RECT 144.155 199.575 144.435 208.605 ;
        RECT 145.035 199.575 145.315 208.605 ;
        RECT 145.915 199.575 146.195 208.605 ;
        RECT 146.600 199.385 146.890 209.365 ;
        RECT 117.060 199.095 121.190 199.385 ;
        RECT 142.760 199.095 146.890 199.385 ;
        RECT 117.060 198.815 117.350 199.095 ;
        RECT 146.600 198.815 146.890 199.095 ;
        RECT 117.060 198.525 146.890 198.815 ;
        RECT 74.400 197.000 116.550 197.290 ;
        RECT 74.400 196.720 74.690 197.000 ;
        RECT 116.260 196.720 116.550 197.000 ;
        RECT 74.400 196.430 78.530 196.720 ;
        RECT 114.180 196.430 116.550 196.720 ;
        RECT 74.400 186.450 74.690 196.430 ;
        RECT 75.095 187.210 75.375 196.240 ;
        RECT 75.975 187.210 76.255 196.240 ;
        RECT 76.855 187.210 77.135 196.240 ;
        RECT 77.735 187.210 78.015 196.240 ;
        RECT 78.615 187.210 78.895 196.240 ;
        RECT 79.495 187.210 79.775 196.240 ;
        RECT 80.375 187.210 80.655 196.240 ;
        RECT 81.255 187.210 81.535 196.240 ;
        RECT 82.135 187.210 82.415 196.240 ;
        RECT 83.015 187.210 83.295 196.240 ;
        RECT 83.895 187.210 84.175 196.240 ;
        RECT 84.775 187.210 85.055 196.240 ;
        RECT 85.655 187.210 85.935 196.240 ;
        RECT 86.535 187.210 86.815 196.240 ;
        RECT 87.415 187.210 87.695 196.240 ;
        RECT 88.295 187.210 88.575 196.240 ;
        RECT 89.175 187.210 89.455 196.240 ;
        RECT 90.055 187.210 90.335 196.240 ;
        RECT 90.935 187.210 91.215 196.240 ;
        RECT 91.815 187.210 92.095 196.240 ;
        RECT 92.695 187.210 92.975 196.240 ;
        RECT 93.575 187.210 93.855 196.240 ;
        RECT 94.455 187.210 94.735 196.240 ;
        RECT 95.335 187.210 95.615 196.240 ;
        RECT 96.215 187.210 96.495 196.240 ;
        RECT 97.095 187.210 97.375 196.240 ;
        RECT 97.975 187.210 98.255 196.240 ;
        RECT 98.855 187.210 99.135 196.240 ;
        RECT 99.735 187.210 100.015 196.240 ;
        RECT 100.615 187.210 100.895 196.240 ;
        RECT 101.495 187.210 101.775 196.240 ;
        RECT 102.375 187.210 102.655 196.240 ;
        RECT 103.255 187.210 103.535 196.240 ;
        RECT 104.135 187.210 104.415 196.240 ;
        RECT 105.015 187.210 105.295 196.240 ;
        RECT 105.895 187.210 106.175 196.240 ;
        RECT 106.775 187.210 107.055 196.240 ;
        RECT 107.655 187.210 107.935 196.240 ;
        RECT 108.535 187.210 108.815 196.240 ;
        RECT 109.415 187.210 109.695 196.240 ;
        RECT 110.295 187.210 110.575 196.240 ;
        RECT 111.175 187.210 111.455 196.240 ;
        RECT 112.055 187.210 112.335 196.240 ;
        RECT 112.935 187.210 113.215 196.240 ;
        RECT 113.815 187.210 114.095 196.240 ;
        RECT 114.695 187.210 114.975 196.240 ;
        RECT 115.575 187.210 115.855 196.240 ;
        RECT 78.980 186.690 113.730 187.020 ;
        RECT 116.260 186.450 116.550 196.430 ;
        RECT 74.400 186.160 116.550 186.450 ;
        RECT 117.060 197.000 146.890 197.290 ;
        RECT 117.060 196.720 117.350 197.000 ;
        RECT 146.600 196.720 146.890 197.000 ;
        RECT 117.060 196.430 122.950 196.720 ;
        RECT 130.440 196.430 133.510 196.720 ;
        RECT 141.000 196.430 146.890 196.720 ;
        RECT 117.060 186.450 117.350 196.430 ;
        RECT 117.755 187.210 118.035 196.240 ;
        RECT 118.635 187.210 118.915 196.240 ;
        RECT 119.515 187.210 119.795 196.240 ;
        RECT 120.395 187.210 120.675 196.240 ;
        RECT 121.275 187.210 121.555 196.240 ;
        RECT 122.155 187.210 122.435 196.240 ;
        RECT 123.035 187.210 123.315 196.240 ;
        RECT 123.915 187.210 124.195 196.240 ;
        RECT 124.795 187.210 125.075 196.240 ;
        RECT 125.675 187.210 125.955 196.240 ;
        RECT 126.555 187.210 126.835 196.240 ;
        RECT 127.435 187.210 127.715 196.240 ;
        RECT 128.315 187.210 128.595 196.240 ;
        RECT 129.195 187.210 129.475 196.240 ;
        RECT 130.075 187.210 130.355 196.240 ;
        RECT 130.955 187.210 131.235 196.430 ;
        RECT 131.835 187.210 132.115 196.430 ;
        RECT 132.715 187.210 132.995 196.430 ;
        RECT 133.595 187.210 133.875 196.240 ;
        RECT 134.475 187.210 134.755 196.240 ;
        RECT 135.355 187.210 135.635 196.240 ;
        RECT 136.235 187.210 136.515 196.240 ;
        RECT 137.115 187.210 137.395 196.240 ;
        RECT 137.995 187.210 138.275 196.240 ;
        RECT 138.875 187.210 139.155 196.240 ;
        RECT 139.755 187.210 140.035 196.240 ;
        RECT 140.635 187.210 140.915 196.240 ;
        RECT 141.515 187.210 141.795 196.240 ;
        RECT 142.395 187.210 142.675 196.240 ;
        RECT 143.275 187.210 143.555 196.240 ;
        RECT 144.155 187.210 144.435 196.240 ;
        RECT 145.035 187.210 145.315 196.240 ;
        RECT 145.915 187.210 146.195 196.240 ;
        RECT 123.345 186.730 129.990 187.020 ;
        RECT 123.345 186.690 129.935 186.730 ;
        RECT 133.960 186.690 140.550 187.020 ;
        RECT 146.600 186.450 146.890 196.430 ;
        RECT 147.280 194.155 170.150 194.445 ;
        RECT 147.280 193.325 147.570 194.155 ;
        RECT 148.380 193.625 152.190 193.915 ;
        RECT 151.900 193.325 152.190 193.625 ;
        RECT 165.240 193.625 169.050 193.915 ;
        RECT 165.240 193.325 165.530 193.625 ;
        RECT 169.860 193.325 170.150 194.155 ;
        RECT 147.280 193.035 151.450 193.325 ;
        RECT 151.900 193.035 165.530 193.325 ;
        RECT 165.980 193.035 170.150 193.325 ;
        RECT 147.280 190.395 147.570 193.035 ;
        RECT 148.015 190.585 148.295 192.845 ;
        RECT 148.895 190.585 149.175 192.845 ;
        RECT 149.775 190.585 150.055 192.845 ;
        RECT 150.655 190.585 150.935 192.845 ;
        RECT 151.535 190.585 151.815 192.845 ;
        RECT 152.415 190.585 152.695 192.845 ;
        RECT 153.295 190.585 153.575 192.845 ;
        RECT 154.175 190.585 154.455 192.845 ;
        RECT 155.055 190.585 155.335 192.845 ;
        RECT 155.935 190.585 156.215 192.845 ;
        RECT 156.815 190.585 157.095 192.845 ;
        RECT 157.695 190.585 157.975 192.845 ;
        RECT 158.575 190.585 158.855 192.845 ;
        RECT 159.455 190.585 159.735 192.845 ;
        RECT 160.335 190.585 160.615 192.845 ;
        RECT 161.215 190.585 161.495 192.845 ;
        RECT 162.095 190.585 162.375 192.845 ;
        RECT 162.975 190.585 163.255 192.845 ;
        RECT 163.855 190.585 164.135 192.845 ;
        RECT 164.735 190.585 165.015 192.845 ;
        RECT 165.615 190.585 165.895 192.845 ;
        RECT 166.495 190.585 166.775 192.845 ;
        RECT 167.375 190.585 167.655 192.845 ;
        RECT 168.255 190.585 168.535 192.845 ;
        RECT 169.135 190.585 169.415 192.845 ;
        RECT 169.860 190.395 170.150 193.035 ;
        RECT 147.280 190.105 151.450 190.395 ;
        RECT 151.900 190.105 165.530 190.395 ;
        RECT 165.980 190.105 170.150 190.395 ;
        RECT 147.280 189.270 147.570 190.105 ;
        RECT 151.900 189.805 152.190 190.105 ;
        RECT 148.380 189.515 152.190 189.805 ;
        RECT 165.240 189.805 165.530 190.105 ;
        RECT 165.240 189.515 169.050 189.805 ;
        RECT 169.860 189.270 170.150 190.105 ;
        RECT 147.280 188.980 170.150 189.270 ;
        RECT 184.785 189.355 207.655 189.645 ;
        RECT 117.060 186.160 146.890 186.450 ;
        RECT 184.785 186.065 185.075 189.355 ;
        RECT 192.925 188.705 199.515 189.035 ;
        RECT 185.520 186.255 185.800 188.515 ;
        RECT 186.400 186.255 186.680 188.515 ;
        RECT 187.280 186.255 187.560 188.515 ;
        RECT 188.160 186.255 188.440 188.515 ;
        RECT 189.040 186.255 189.320 188.515 ;
        RECT 189.920 186.255 190.200 188.515 ;
        RECT 190.800 186.255 191.080 188.515 ;
        RECT 191.680 186.255 191.960 188.515 ;
        RECT 192.560 186.255 192.840 188.515 ;
        RECT 193.440 186.255 193.720 188.515 ;
        RECT 194.320 186.255 194.600 188.515 ;
        RECT 195.200 186.255 195.480 188.515 ;
        RECT 196.080 186.255 196.360 188.515 ;
        RECT 196.960 186.255 197.240 188.515 ;
        RECT 197.840 186.255 198.120 188.515 ;
        RECT 198.720 186.255 199.000 188.515 ;
        RECT 199.600 186.255 199.880 188.515 ;
        RECT 200.480 186.255 200.760 188.515 ;
        RECT 201.360 186.255 201.640 188.515 ;
        RECT 202.240 186.255 202.520 188.515 ;
        RECT 203.120 186.255 203.400 188.515 ;
        RECT 204.000 186.255 204.280 188.515 ;
        RECT 204.880 186.255 205.160 188.515 ;
        RECT 205.760 186.255 206.040 188.515 ;
        RECT 206.640 186.255 206.920 188.515 ;
        RECT 207.365 186.065 207.655 189.355 ;
        RECT 184.785 185.775 192.475 186.065 ;
        RECT 199.965 185.775 207.655 186.065 ;
        RECT 184.785 185.415 185.075 185.775 ;
        RECT 207.365 185.415 207.655 185.775 ;
        RECT 74.365 185.075 116.590 185.365 ;
        RECT 74.365 184.715 74.655 185.075 ;
        RECT 116.300 184.715 116.590 185.075 ;
        RECT 74.365 184.425 78.530 184.715 ;
        RECT 114.180 184.425 116.590 184.715 ;
        RECT 74.365 183.605 74.655 184.425 ;
        RECT 74.360 182.605 74.655 183.605 ;
        RECT 74.365 181.135 74.655 182.605 ;
        RECT 75.095 181.975 75.375 184.235 ;
        RECT 75.975 181.975 76.255 184.235 ;
        RECT 76.855 181.975 77.135 184.235 ;
        RECT 77.735 181.975 78.015 184.235 ;
        RECT 78.615 181.975 78.895 184.235 ;
        RECT 79.495 181.975 79.775 184.235 ;
        RECT 80.375 181.975 80.655 184.235 ;
        RECT 81.255 181.975 81.535 184.235 ;
        RECT 82.135 181.975 82.415 184.235 ;
        RECT 83.015 181.975 83.295 184.235 ;
        RECT 83.895 181.975 84.175 184.235 ;
        RECT 84.775 181.975 85.055 184.235 ;
        RECT 85.655 181.975 85.935 184.235 ;
        RECT 86.535 181.975 86.815 184.235 ;
        RECT 87.415 181.975 87.695 184.235 ;
        RECT 88.295 181.975 88.575 184.235 ;
        RECT 89.175 181.975 89.455 184.235 ;
        RECT 90.055 181.975 90.335 184.235 ;
        RECT 90.935 181.975 91.215 184.235 ;
        RECT 91.815 181.975 92.095 184.235 ;
        RECT 92.695 181.975 92.975 184.235 ;
        RECT 93.575 181.975 93.855 184.235 ;
        RECT 94.455 181.975 94.735 184.235 ;
        RECT 95.335 181.975 95.615 184.235 ;
        RECT 96.215 181.975 96.495 184.235 ;
        RECT 97.095 181.975 97.375 184.235 ;
        RECT 97.975 181.975 98.255 184.235 ;
        RECT 98.855 181.975 99.135 184.235 ;
        RECT 99.735 181.975 100.015 184.235 ;
        RECT 100.615 181.975 100.895 184.235 ;
        RECT 101.495 181.975 101.775 184.235 ;
        RECT 102.375 181.975 102.655 184.235 ;
        RECT 103.255 181.975 103.535 184.235 ;
        RECT 104.135 181.975 104.415 184.235 ;
        RECT 105.015 181.975 105.295 184.235 ;
        RECT 105.895 181.975 106.175 184.235 ;
        RECT 106.775 181.975 107.055 184.235 ;
        RECT 107.655 181.975 107.935 184.235 ;
        RECT 108.535 181.975 108.815 184.235 ;
        RECT 109.415 181.975 109.695 184.235 ;
        RECT 110.295 181.975 110.575 184.235 ;
        RECT 111.175 181.975 111.455 184.235 ;
        RECT 112.055 181.975 112.335 184.235 ;
        RECT 112.935 181.975 113.215 184.235 ;
        RECT 113.815 181.975 114.095 184.235 ;
        RECT 114.695 181.975 114.975 184.235 ;
        RECT 115.575 181.975 115.855 184.235 ;
        RECT 78.980 181.455 115.760 181.785 ;
        RECT 116.300 181.135 116.590 184.425 ;
        RECT 74.365 180.845 116.590 181.135 ;
        RECT 117.020 185.075 146.930 185.365 ;
        RECT 117.020 184.715 117.310 185.075 ;
        RECT 146.640 184.715 146.930 185.075 ;
        RECT 117.020 184.425 122.950 184.715 ;
        RECT 130.440 184.425 133.510 184.715 ;
        RECT 141.000 184.425 146.930 184.715 ;
        RECT 117.020 181.135 117.310 184.425 ;
        RECT 117.755 181.975 118.035 184.235 ;
        RECT 118.635 181.975 118.915 184.235 ;
        RECT 119.515 181.975 119.795 184.235 ;
        RECT 120.395 181.975 120.675 184.235 ;
        RECT 121.275 181.975 121.555 184.235 ;
        RECT 122.155 181.975 122.435 184.235 ;
        RECT 123.035 181.975 123.315 184.235 ;
        RECT 123.915 181.975 124.195 184.235 ;
        RECT 124.795 181.975 125.075 184.235 ;
        RECT 125.675 181.975 125.955 184.235 ;
        RECT 126.555 181.975 126.835 184.235 ;
        RECT 127.435 181.975 127.715 184.235 ;
        RECT 128.315 181.975 128.595 184.235 ;
        RECT 129.195 181.975 129.475 184.235 ;
        RECT 130.075 181.975 130.355 184.235 ;
        RECT 130.955 181.975 131.235 184.425 ;
        RECT 131.835 181.975 132.115 184.425 ;
        RECT 132.715 181.975 132.995 184.425 ;
        RECT 133.595 181.975 133.875 184.235 ;
        RECT 134.475 181.975 134.755 184.235 ;
        RECT 135.355 181.975 135.635 184.235 ;
        RECT 136.235 181.975 136.515 184.235 ;
        RECT 137.115 181.975 137.395 184.235 ;
        RECT 137.995 181.975 138.275 184.235 ;
        RECT 138.875 181.975 139.155 184.235 ;
        RECT 139.755 181.975 140.035 184.235 ;
        RECT 140.635 181.975 140.915 184.235 ;
        RECT 141.515 181.975 141.795 184.235 ;
        RECT 142.395 181.975 142.675 184.235 ;
        RECT 143.275 181.975 143.555 184.235 ;
        RECT 144.155 181.975 144.435 184.235 ;
        RECT 145.035 181.975 145.315 184.235 ;
        RECT 145.915 181.975 146.195 184.235 ;
        RECT 123.400 181.455 143.275 181.785 ;
        RECT 146.640 181.135 146.930 184.425 ;
        RECT 117.020 180.845 146.930 181.135 ;
        RECT 147.280 185.075 170.150 185.365 ;
        RECT 184.785 185.125 207.655 185.415 ;
        RECT 208.005 189.355 237.915 189.645 ;
        RECT 208.005 186.065 208.295 189.355 ;
        RECT 221.425 188.705 224.495 188.995 ;
        RECT 208.740 186.255 209.020 188.515 ;
        RECT 209.620 186.255 209.900 188.515 ;
        RECT 210.500 186.255 210.780 188.515 ;
        RECT 211.380 186.255 211.660 188.515 ;
        RECT 212.260 186.255 212.540 188.515 ;
        RECT 213.140 186.255 213.420 188.515 ;
        RECT 214.020 186.255 214.300 188.515 ;
        RECT 214.900 186.255 215.180 188.515 ;
        RECT 215.780 186.255 216.060 188.515 ;
        RECT 216.660 186.255 216.940 188.515 ;
        RECT 217.540 186.255 217.820 188.515 ;
        RECT 218.420 186.255 218.700 188.515 ;
        RECT 219.300 186.255 219.580 188.515 ;
        RECT 220.180 186.255 220.460 188.515 ;
        RECT 221.060 186.255 221.340 188.515 ;
        RECT 221.940 186.255 222.220 188.705 ;
        RECT 222.820 186.255 223.100 188.515 ;
        RECT 223.700 186.255 223.980 188.705 ;
        RECT 224.580 186.255 224.860 188.515 ;
        RECT 225.460 186.255 225.740 188.515 ;
        RECT 226.340 186.255 226.620 188.515 ;
        RECT 227.220 186.255 227.500 188.515 ;
        RECT 228.100 186.255 228.380 188.515 ;
        RECT 228.980 186.255 229.260 188.515 ;
        RECT 229.860 186.255 230.140 188.515 ;
        RECT 230.740 186.255 231.020 188.515 ;
        RECT 231.620 186.255 231.900 188.515 ;
        RECT 232.500 186.255 232.780 188.515 ;
        RECT 233.380 186.255 233.660 188.515 ;
        RECT 234.260 186.255 234.540 188.515 ;
        RECT 235.140 186.255 235.420 188.515 ;
        RECT 236.020 186.255 236.300 188.515 ;
        RECT 236.900 186.255 237.180 188.515 ;
        RECT 237.625 186.065 237.915 189.355 ;
        RECT 208.005 185.775 213.935 186.065 ;
        RECT 214.385 185.775 231.535 186.065 ;
        RECT 231.985 185.775 237.915 186.065 ;
        RECT 208.005 185.415 208.295 185.775 ;
        RECT 237.625 185.415 237.915 185.775 ;
        RECT 208.005 185.125 237.915 185.415 ;
        RECT 238.345 189.355 280.570 189.645 ;
        RECT 238.345 186.065 238.635 189.355 ;
        RECT 239.080 186.255 239.360 188.515 ;
        RECT 239.960 186.255 240.240 188.515 ;
        RECT 240.840 186.255 241.120 188.515 ;
        RECT 241.720 186.255 242.000 188.515 ;
        RECT 242.600 186.255 242.880 188.515 ;
        RECT 243.480 186.255 243.760 188.515 ;
        RECT 244.360 186.255 244.640 188.515 ;
        RECT 245.240 186.255 245.520 188.515 ;
        RECT 246.120 186.255 246.400 188.515 ;
        RECT 247.000 186.255 247.280 188.515 ;
        RECT 247.880 186.255 248.160 188.515 ;
        RECT 248.760 186.255 249.040 188.515 ;
        RECT 249.640 186.255 249.920 188.515 ;
        RECT 250.520 186.255 250.800 188.515 ;
        RECT 251.400 186.255 251.680 188.515 ;
        RECT 252.280 186.255 252.560 188.515 ;
        RECT 253.160 186.255 253.440 188.515 ;
        RECT 254.040 186.255 254.320 188.515 ;
        RECT 254.920 186.255 255.200 188.515 ;
        RECT 255.800 186.255 256.080 188.515 ;
        RECT 256.680 186.255 256.960 188.515 ;
        RECT 257.560 186.255 257.840 188.515 ;
        RECT 258.440 186.255 258.720 188.515 ;
        RECT 259.320 186.255 259.600 188.515 ;
        RECT 260.200 186.255 260.480 188.515 ;
        RECT 261.080 186.255 261.360 188.515 ;
        RECT 261.960 186.255 262.240 188.515 ;
        RECT 262.840 186.255 263.120 188.515 ;
        RECT 263.720 186.255 264.000 188.515 ;
        RECT 264.600 186.255 264.880 188.515 ;
        RECT 265.480 186.255 265.760 188.515 ;
        RECT 266.360 186.255 266.640 188.515 ;
        RECT 267.240 186.255 267.520 188.515 ;
        RECT 268.120 186.255 268.400 188.515 ;
        RECT 269.000 186.255 269.280 188.515 ;
        RECT 269.880 186.255 270.160 188.515 ;
        RECT 270.760 186.255 271.040 188.515 ;
        RECT 271.640 186.255 271.920 188.515 ;
        RECT 272.520 186.255 272.800 188.515 ;
        RECT 273.400 186.255 273.680 188.515 ;
        RECT 274.280 186.255 274.560 188.515 ;
        RECT 275.160 186.255 275.440 188.515 ;
        RECT 276.040 186.255 276.320 188.515 ;
        RECT 276.920 186.255 277.200 188.515 ;
        RECT 277.800 186.255 278.080 188.515 ;
        RECT 278.680 186.255 278.960 188.515 ;
        RECT 279.560 186.255 279.840 188.515 ;
        RECT 280.280 187.885 280.570 189.355 ;
        RECT 280.280 186.885 280.575 187.885 ;
        RECT 280.280 186.065 280.570 186.885 ;
        RECT 238.345 185.775 240.755 186.065 ;
        RECT 241.205 185.775 275.955 186.065 ;
        RECT 276.405 185.775 280.570 186.065 ;
        RECT 238.345 185.415 238.635 185.775 ;
        RECT 280.280 185.415 280.570 185.775 ;
        RECT 238.345 185.125 280.570 185.415 ;
        RECT 147.280 184.715 147.570 185.075 ;
        RECT 169.860 184.715 170.150 185.075 ;
        RECT 147.280 184.425 154.970 184.715 ;
        RECT 162.460 184.425 170.150 184.715 ;
        RECT 147.280 181.135 147.570 184.425 ;
        RECT 148.015 181.975 148.295 184.235 ;
        RECT 148.895 181.975 149.175 184.235 ;
        RECT 149.775 181.975 150.055 184.235 ;
        RECT 150.655 181.975 150.935 184.235 ;
        RECT 151.535 181.975 151.815 184.235 ;
        RECT 152.415 181.975 152.695 184.235 ;
        RECT 153.295 181.975 153.575 184.235 ;
        RECT 154.175 181.975 154.455 184.235 ;
        RECT 155.055 181.975 155.335 184.235 ;
        RECT 155.935 181.975 156.215 184.235 ;
        RECT 156.815 181.975 157.095 184.235 ;
        RECT 157.695 181.975 157.975 184.235 ;
        RECT 158.575 181.975 158.855 184.235 ;
        RECT 159.455 181.975 159.735 184.235 ;
        RECT 160.335 181.975 160.615 184.235 ;
        RECT 161.215 181.975 161.495 184.235 ;
        RECT 162.095 181.975 162.375 184.235 ;
        RECT 162.975 181.975 163.255 184.235 ;
        RECT 163.855 181.975 164.135 184.235 ;
        RECT 164.735 181.975 165.015 184.235 ;
        RECT 165.615 181.975 165.895 184.235 ;
        RECT 166.495 181.975 166.775 184.235 ;
        RECT 167.375 181.975 167.655 184.235 ;
        RECT 168.255 181.975 168.535 184.235 ;
        RECT 169.135 181.975 169.415 184.235 ;
        RECT 155.420 181.455 162.030 181.785 ;
        RECT 169.860 181.135 170.150 184.425 ;
        RECT 147.280 180.845 170.150 181.135 ;
        RECT 184.785 182.870 207.655 183.160 ;
        RECT 184.785 179.580 185.075 182.870 ;
        RECT 192.905 182.220 199.515 182.550 ;
        RECT 185.520 179.770 185.800 182.030 ;
        RECT 186.400 179.770 186.680 182.030 ;
        RECT 187.280 179.770 187.560 182.030 ;
        RECT 188.160 179.770 188.440 182.030 ;
        RECT 189.040 179.770 189.320 182.030 ;
        RECT 189.920 179.770 190.200 182.030 ;
        RECT 190.800 179.770 191.080 182.030 ;
        RECT 191.680 179.770 191.960 182.030 ;
        RECT 192.560 179.770 192.840 182.030 ;
        RECT 193.440 179.770 193.720 182.030 ;
        RECT 194.320 179.770 194.600 182.030 ;
        RECT 195.200 179.770 195.480 182.030 ;
        RECT 196.080 179.770 196.360 182.030 ;
        RECT 196.960 179.770 197.240 182.030 ;
        RECT 197.840 179.770 198.120 182.030 ;
        RECT 198.720 179.770 199.000 182.030 ;
        RECT 199.600 179.770 199.880 182.030 ;
        RECT 200.480 179.770 200.760 182.030 ;
        RECT 201.360 179.770 201.640 182.030 ;
        RECT 202.240 179.770 202.520 182.030 ;
        RECT 203.120 179.770 203.400 182.030 ;
        RECT 204.000 179.770 204.280 182.030 ;
        RECT 204.880 179.770 205.160 182.030 ;
        RECT 205.760 179.770 206.040 182.030 ;
        RECT 206.640 179.770 206.920 182.030 ;
        RECT 207.365 179.580 207.655 182.870 ;
        RECT 184.785 179.290 192.475 179.580 ;
        RECT 199.965 179.290 207.655 179.580 ;
        RECT 184.785 178.930 185.075 179.290 ;
        RECT 207.365 178.930 207.655 179.290 ;
        RECT 74.365 178.590 116.590 178.880 ;
        RECT 74.365 178.230 74.655 178.590 ;
        RECT 116.300 178.230 116.590 178.590 ;
        RECT 74.365 177.940 78.530 178.230 ;
        RECT 78.980 177.940 113.730 178.230 ;
        RECT 114.180 177.940 116.590 178.230 ;
        RECT 74.365 177.120 74.655 177.940 ;
        RECT 74.360 176.120 74.655 177.120 ;
        RECT 74.365 174.650 74.655 176.120 ;
        RECT 75.095 175.490 75.375 177.750 ;
        RECT 75.975 175.490 76.255 177.750 ;
        RECT 76.855 175.490 77.135 177.750 ;
        RECT 77.735 175.490 78.015 177.750 ;
        RECT 78.615 175.490 78.895 177.750 ;
        RECT 79.495 175.490 79.775 177.750 ;
        RECT 80.375 175.490 80.655 177.750 ;
        RECT 81.255 175.490 81.535 177.750 ;
        RECT 82.135 175.490 82.415 177.750 ;
        RECT 83.015 175.490 83.295 177.750 ;
        RECT 83.895 175.490 84.175 177.750 ;
        RECT 84.775 175.490 85.055 177.750 ;
        RECT 85.655 175.490 85.935 177.750 ;
        RECT 86.535 175.490 86.815 177.750 ;
        RECT 87.415 175.490 87.695 177.750 ;
        RECT 88.295 175.490 88.575 177.750 ;
        RECT 89.175 175.490 89.455 177.750 ;
        RECT 90.055 175.490 90.335 177.750 ;
        RECT 90.935 175.490 91.215 177.750 ;
        RECT 91.815 175.490 92.095 177.750 ;
        RECT 92.695 175.490 92.975 177.750 ;
        RECT 93.575 175.490 93.855 177.750 ;
        RECT 94.455 175.490 94.735 177.750 ;
        RECT 95.335 175.490 95.615 177.750 ;
        RECT 96.215 175.490 96.495 177.750 ;
        RECT 97.095 175.490 97.375 177.750 ;
        RECT 97.975 175.490 98.255 177.750 ;
        RECT 98.855 175.490 99.135 177.750 ;
        RECT 99.735 175.490 100.015 177.750 ;
        RECT 100.615 175.490 100.895 177.750 ;
        RECT 101.495 175.490 101.775 177.750 ;
        RECT 102.375 175.490 102.655 177.750 ;
        RECT 103.255 175.490 103.535 177.750 ;
        RECT 104.135 175.490 104.415 177.750 ;
        RECT 105.015 175.490 105.295 177.750 ;
        RECT 105.895 175.490 106.175 177.750 ;
        RECT 106.775 175.490 107.055 177.750 ;
        RECT 107.655 175.490 107.935 177.750 ;
        RECT 108.535 175.490 108.815 177.750 ;
        RECT 109.415 175.490 109.695 177.750 ;
        RECT 110.295 175.490 110.575 177.750 ;
        RECT 111.175 175.490 111.455 177.750 ;
        RECT 112.055 175.490 112.335 177.750 ;
        RECT 112.935 175.490 113.215 177.750 ;
        RECT 113.815 175.490 114.095 177.750 ;
        RECT 114.695 175.490 114.975 177.750 ;
        RECT 115.575 175.490 115.855 177.750 ;
        RECT 116.300 174.650 116.590 177.940 ;
        RECT 74.365 174.360 116.590 174.650 ;
        RECT 117.020 178.590 146.930 178.880 ;
        RECT 117.020 178.230 117.310 178.590 ;
        RECT 146.640 178.230 146.930 178.590 ;
        RECT 117.020 177.940 122.950 178.230 ;
        RECT 123.400 177.940 140.550 178.230 ;
        RECT 141.000 177.940 146.930 178.230 ;
        RECT 117.020 174.650 117.310 177.940 ;
        RECT 117.755 175.490 118.035 177.750 ;
        RECT 118.635 175.490 118.915 177.750 ;
        RECT 119.515 175.490 119.795 177.750 ;
        RECT 120.395 175.490 120.675 177.750 ;
        RECT 121.275 175.490 121.555 177.750 ;
        RECT 122.155 175.490 122.435 177.750 ;
        RECT 123.035 175.490 123.315 177.750 ;
        RECT 123.915 175.490 124.195 177.750 ;
        RECT 124.795 175.490 125.075 177.750 ;
        RECT 125.675 175.490 125.955 177.750 ;
        RECT 126.555 175.490 126.835 177.750 ;
        RECT 127.435 175.490 127.715 177.750 ;
        RECT 128.315 175.490 128.595 177.750 ;
        RECT 129.195 175.490 129.475 177.750 ;
        RECT 130.075 175.490 130.355 177.750 ;
        RECT 130.955 175.300 131.235 177.750 ;
        RECT 131.835 175.490 132.115 177.750 ;
        RECT 132.715 175.300 132.995 177.750 ;
        RECT 133.595 175.490 133.875 177.750 ;
        RECT 134.475 175.490 134.755 177.750 ;
        RECT 135.355 175.490 135.635 177.750 ;
        RECT 136.235 175.490 136.515 177.750 ;
        RECT 137.115 175.490 137.395 177.750 ;
        RECT 137.995 175.490 138.275 177.750 ;
        RECT 138.875 175.490 139.155 177.750 ;
        RECT 139.755 175.490 140.035 177.750 ;
        RECT 140.635 175.490 140.915 177.750 ;
        RECT 141.515 175.490 141.795 177.750 ;
        RECT 142.395 175.490 142.675 177.750 ;
        RECT 143.275 175.490 143.555 177.750 ;
        RECT 144.155 175.490 144.435 177.750 ;
        RECT 145.035 175.490 145.315 177.750 ;
        RECT 145.915 175.490 146.195 177.750 ;
        RECT 130.440 175.010 133.510 175.300 ;
        RECT 146.640 174.650 146.930 177.940 ;
        RECT 117.020 174.360 146.930 174.650 ;
        RECT 147.280 178.590 170.150 178.880 ;
        RECT 184.785 178.640 207.655 178.930 ;
        RECT 208.005 182.870 237.915 183.160 ;
        RECT 208.005 179.580 208.295 182.870 ;
        RECT 211.660 182.220 231.535 182.550 ;
        RECT 208.740 179.770 209.020 182.030 ;
        RECT 209.620 179.770 209.900 182.030 ;
        RECT 210.500 179.770 210.780 182.030 ;
        RECT 211.380 179.770 211.660 182.030 ;
        RECT 212.260 179.770 212.540 182.030 ;
        RECT 213.140 179.770 213.420 182.030 ;
        RECT 214.020 179.770 214.300 182.030 ;
        RECT 214.900 179.770 215.180 182.030 ;
        RECT 215.780 179.770 216.060 182.030 ;
        RECT 216.660 179.770 216.940 182.030 ;
        RECT 217.540 179.770 217.820 182.030 ;
        RECT 218.420 179.770 218.700 182.030 ;
        RECT 219.300 179.770 219.580 182.030 ;
        RECT 220.180 179.770 220.460 182.030 ;
        RECT 221.060 179.770 221.340 182.030 ;
        RECT 221.940 179.580 222.220 182.030 ;
        RECT 222.820 179.580 223.100 182.030 ;
        RECT 223.700 179.580 223.980 182.030 ;
        RECT 224.580 179.770 224.860 182.030 ;
        RECT 225.460 179.770 225.740 182.030 ;
        RECT 226.340 179.770 226.620 182.030 ;
        RECT 227.220 179.770 227.500 182.030 ;
        RECT 228.100 179.770 228.380 182.030 ;
        RECT 228.980 179.770 229.260 182.030 ;
        RECT 229.860 179.770 230.140 182.030 ;
        RECT 230.740 179.770 231.020 182.030 ;
        RECT 231.620 179.770 231.900 182.030 ;
        RECT 232.500 179.770 232.780 182.030 ;
        RECT 233.380 179.770 233.660 182.030 ;
        RECT 234.260 179.770 234.540 182.030 ;
        RECT 235.140 179.770 235.420 182.030 ;
        RECT 236.020 179.770 236.300 182.030 ;
        RECT 236.900 179.770 237.180 182.030 ;
        RECT 237.625 179.580 237.915 182.870 ;
        RECT 208.005 179.290 213.935 179.580 ;
        RECT 221.425 179.290 224.495 179.580 ;
        RECT 231.985 179.290 237.915 179.580 ;
        RECT 208.005 178.930 208.295 179.290 ;
        RECT 237.625 178.930 237.915 179.290 ;
        RECT 208.005 178.640 237.915 178.930 ;
        RECT 238.345 182.870 280.570 183.160 ;
        RECT 238.345 179.580 238.635 182.870 ;
        RECT 239.175 182.220 275.955 182.550 ;
        RECT 239.080 179.770 239.360 182.030 ;
        RECT 239.960 179.770 240.240 182.030 ;
        RECT 240.840 179.770 241.120 182.030 ;
        RECT 241.720 179.770 242.000 182.030 ;
        RECT 242.600 179.770 242.880 182.030 ;
        RECT 243.480 179.770 243.760 182.030 ;
        RECT 244.360 179.770 244.640 182.030 ;
        RECT 245.240 179.770 245.520 182.030 ;
        RECT 246.120 179.770 246.400 182.030 ;
        RECT 247.000 179.770 247.280 182.030 ;
        RECT 247.880 179.770 248.160 182.030 ;
        RECT 248.760 179.770 249.040 182.030 ;
        RECT 249.640 179.770 249.920 182.030 ;
        RECT 250.520 179.770 250.800 182.030 ;
        RECT 251.400 179.770 251.680 182.030 ;
        RECT 252.280 179.770 252.560 182.030 ;
        RECT 253.160 179.770 253.440 182.030 ;
        RECT 254.040 179.770 254.320 182.030 ;
        RECT 254.920 179.770 255.200 182.030 ;
        RECT 255.800 179.770 256.080 182.030 ;
        RECT 256.680 179.770 256.960 182.030 ;
        RECT 257.560 179.770 257.840 182.030 ;
        RECT 258.440 179.770 258.720 182.030 ;
        RECT 259.320 179.770 259.600 182.030 ;
        RECT 260.200 179.770 260.480 182.030 ;
        RECT 261.080 179.770 261.360 182.030 ;
        RECT 261.960 179.770 262.240 182.030 ;
        RECT 262.840 179.770 263.120 182.030 ;
        RECT 263.720 179.770 264.000 182.030 ;
        RECT 264.600 179.770 264.880 182.030 ;
        RECT 265.480 179.770 265.760 182.030 ;
        RECT 266.360 179.770 266.640 182.030 ;
        RECT 267.240 179.770 267.520 182.030 ;
        RECT 268.120 179.770 268.400 182.030 ;
        RECT 269.000 179.770 269.280 182.030 ;
        RECT 269.880 179.770 270.160 182.030 ;
        RECT 270.760 179.770 271.040 182.030 ;
        RECT 271.640 179.770 271.920 182.030 ;
        RECT 272.520 179.770 272.800 182.030 ;
        RECT 273.400 179.770 273.680 182.030 ;
        RECT 274.280 179.770 274.560 182.030 ;
        RECT 275.160 179.770 275.440 182.030 ;
        RECT 276.040 179.770 276.320 182.030 ;
        RECT 276.920 179.770 277.200 182.030 ;
        RECT 277.800 179.770 278.080 182.030 ;
        RECT 278.680 179.770 278.960 182.030 ;
        RECT 279.560 179.770 279.840 182.030 ;
        RECT 280.280 181.400 280.570 182.870 ;
        RECT 280.280 180.400 280.575 181.400 ;
        RECT 280.280 179.580 280.570 180.400 ;
        RECT 238.345 179.290 240.755 179.580 ;
        RECT 276.405 179.290 280.570 179.580 ;
        RECT 238.345 178.930 238.635 179.290 ;
        RECT 280.280 178.930 280.570 179.290 ;
        RECT 238.345 178.640 280.570 178.930 ;
        RECT 147.280 178.230 147.570 178.590 ;
        RECT 169.860 178.230 170.150 178.590 ;
        RECT 147.280 177.940 154.970 178.230 ;
        RECT 162.460 177.940 170.150 178.230 ;
        RECT 147.280 174.650 147.570 177.940 ;
        RECT 148.015 175.490 148.295 177.750 ;
        RECT 148.895 175.490 149.175 177.750 ;
        RECT 149.775 175.490 150.055 177.750 ;
        RECT 150.655 175.490 150.935 177.750 ;
        RECT 151.535 175.490 151.815 177.750 ;
        RECT 152.415 175.490 152.695 177.750 ;
        RECT 153.295 175.490 153.575 177.750 ;
        RECT 154.175 175.490 154.455 177.750 ;
        RECT 155.055 175.490 155.335 177.750 ;
        RECT 155.935 175.490 156.215 177.750 ;
        RECT 156.815 175.490 157.095 177.750 ;
        RECT 157.695 175.490 157.975 177.750 ;
        RECT 158.575 175.490 158.855 177.750 ;
        RECT 159.455 175.490 159.735 177.750 ;
        RECT 160.335 175.490 160.615 177.750 ;
        RECT 161.215 175.490 161.495 177.750 ;
        RECT 162.095 175.490 162.375 177.750 ;
        RECT 162.975 175.490 163.255 177.750 ;
        RECT 163.855 175.490 164.135 177.750 ;
        RECT 164.735 175.490 165.015 177.750 ;
        RECT 165.615 175.490 165.895 177.750 ;
        RECT 166.495 175.490 166.775 177.750 ;
        RECT 167.375 175.490 167.655 177.750 ;
        RECT 168.255 175.490 168.535 177.750 ;
        RECT 169.135 175.490 169.415 177.750 ;
        RECT 155.420 174.970 162.010 175.300 ;
        RECT 169.860 174.650 170.150 177.940 ;
        RECT 208.045 177.555 237.875 177.845 ;
        RECT 147.280 174.360 170.150 174.650 ;
        RECT 184.785 174.735 207.655 175.025 ;
        RECT 184.785 173.900 185.075 174.735 ;
        RECT 185.885 174.200 189.695 174.490 ;
        RECT 189.405 173.900 189.695 174.200 ;
        RECT 202.745 174.200 206.555 174.490 ;
        RECT 202.745 173.900 203.035 174.200 ;
        RECT 207.365 173.900 207.655 174.735 ;
        RECT 184.785 173.610 188.955 173.900 ;
        RECT 189.405 173.610 203.035 173.900 ;
        RECT 203.485 173.610 207.655 173.900 ;
        RECT 184.785 170.970 185.075 173.610 ;
        RECT 185.520 171.160 185.800 173.420 ;
        RECT 186.400 171.160 186.680 173.420 ;
        RECT 187.280 171.160 187.560 173.420 ;
        RECT 188.160 171.160 188.440 173.420 ;
        RECT 189.040 171.160 189.320 173.420 ;
        RECT 189.920 171.160 190.200 173.420 ;
        RECT 190.800 171.160 191.080 173.420 ;
        RECT 191.680 171.160 191.960 173.420 ;
        RECT 192.560 171.160 192.840 173.420 ;
        RECT 193.440 171.160 193.720 173.420 ;
        RECT 194.320 171.160 194.600 173.420 ;
        RECT 195.200 171.160 195.480 173.420 ;
        RECT 196.080 171.160 196.360 173.420 ;
        RECT 196.960 171.160 197.240 173.420 ;
        RECT 197.840 171.160 198.120 173.420 ;
        RECT 198.720 171.160 199.000 173.420 ;
        RECT 199.600 171.160 199.880 173.420 ;
        RECT 200.480 171.160 200.760 173.420 ;
        RECT 201.360 171.160 201.640 173.420 ;
        RECT 202.240 171.160 202.520 173.420 ;
        RECT 203.120 171.160 203.400 173.420 ;
        RECT 204.000 171.160 204.280 173.420 ;
        RECT 204.880 171.160 205.160 173.420 ;
        RECT 205.760 171.160 206.040 173.420 ;
        RECT 206.640 171.160 206.920 173.420 ;
        RECT 207.365 170.970 207.655 173.610 ;
        RECT 184.785 170.680 188.955 170.970 ;
        RECT 189.405 170.680 203.035 170.970 ;
        RECT 203.485 170.680 207.655 170.970 ;
        RECT 184.785 169.850 185.075 170.680 ;
        RECT 189.405 170.380 189.695 170.680 ;
        RECT 185.885 170.090 189.695 170.380 ;
        RECT 202.745 170.380 203.035 170.680 ;
        RECT 202.745 170.090 206.555 170.380 ;
        RECT 207.365 169.850 207.655 170.680 ;
        RECT 184.785 169.560 207.655 169.850 ;
        RECT 208.045 167.575 208.335 177.555 ;
        RECT 214.385 176.985 220.975 177.315 ;
        RECT 225.000 177.275 231.590 177.315 ;
        RECT 224.945 176.985 231.590 177.275 ;
        RECT 208.740 167.765 209.020 176.795 ;
        RECT 209.620 167.765 209.900 176.795 ;
        RECT 210.500 167.765 210.780 176.795 ;
        RECT 211.380 167.765 211.660 176.795 ;
        RECT 212.260 167.765 212.540 176.795 ;
        RECT 213.140 167.765 213.420 176.795 ;
        RECT 214.020 167.765 214.300 176.795 ;
        RECT 214.900 167.765 215.180 176.795 ;
        RECT 215.780 167.765 216.060 176.795 ;
        RECT 216.660 167.765 216.940 176.795 ;
        RECT 217.540 167.765 217.820 176.795 ;
        RECT 218.420 167.765 218.700 176.795 ;
        RECT 219.300 167.765 219.580 176.795 ;
        RECT 220.180 167.765 220.460 176.795 ;
        RECT 221.060 167.765 221.340 176.795 ;
        RECT 221.940 167.575 222.220 176.795 ;
        RECT 222.820 167.575 223.100 176.795 ;
        RECT 223.700 167.575 223.980 176.795 ;
        RECT 224.580 167.765 224.860 176.795 ;
        RECT 225.460 167.765 225.740 176.795 ;
        RECT 226.340 167.765 226.620 176.795 ;
        RECT 227.220 167.765 227.500 176.795 ;
        RECT 228.100 167.765 228.380 176.795 ;
        RECT 228.980 167.765 229.260 176.795 ;
        RECT 229.860 167.765 230.140 176.795 ;
        RECT 230.740 167.765 231.020 176.795 ;
        RECT 231.620 167.765 231.900 176.795 ;
        RECT 232.500 167.765 232.780 176.795 ;
        RECT 233.380 167.765 233.660 176.795 ;
        RECT 234.260 167.765 234.540 176.795 ;
        RECT 235.140 167.765 235.420 176.795 ;
        RECT 236.020 167.765 236.300 176.795 ;
        RECT 236.900 167.765 237.180 176.795 ;
        RECT 237.585 167.575 237.875 177.555 ;
        RECT 208.045 167.285 213.935 167.575 ;
        RECT 221.425 167.285 224.495 167.575 ;
        RECT 231.985 167.285 237.875 167.575 ;
        RECT 208.045 167.005 208.335 167.285 ;
        RECT 237.585 167.005 237.875 167.285 ;
        RECT 208.045 166.715 237.875 167.005 ;
        RECT 238.385 177.555 280.535 177.845 ;
        RECT 238.385 167.575 238.675 177.555 ;
        RECT 241.205 176.985 275.955 177.315 ;
        RECT 239.080 167.765 239.360 176.795 ;
        RECT 239.960 167.765 240.240 176.795 ;
        RECT 240.840 167.765 241.120 176.795 ;
        RECT 241.720 167.765 242.000 176.795 ;
        RECT 242.600 167.765 242.880 176.795 ;
        RECT 243.480 167.765 243.760 176.795 ;
        RECT 244.360 167.765 244.640 176.795 ;
        RECT 245.240 167.765 245.520 176.795 ;
        RECT 246.120 167.765 246.400 176.795 ;
        RECT 247.000 167.765 247.280 176.795 ;
        RECT 247.880 167.765 248.160 176.795 ;
        RECT 248.760 167.765 249.040 176.795 ;
        RECT 249.640 167.765 249.920 176.795 ;
        RECT 250.520 167.765 250.800 176.795 ;
        RECT 251.400 167.765 251.680 176.795 ;
        RECT 252.280 167.765 252.560 176.795 ;
        RECT 253.160 167.765 253.440 176.795 ;
        RECT 254.040 167.765 254.320 176.795 ;
        RECT 254.920 167.765 255.200 176.795 ;
        RECT 255.800 167.765 256.080 176.795 ;
        RECT 256.680 167.765 256.960 176.795 ;
        RECT 257.560 167.765 257.840 176.795 ;
        RECT 258.440 167.765 258.720 176.795 ;
        RECT 259.320 167.765 259.600 176.795 ;
        RECT 260.200 167.765 260.480 176.795 ;
        RECT 261.080 167.765 261.360 176.795 ;
        RECT 261.960 167.765 262.240 176.795 ;
        RECT 262.840 167.765 263.120 176.795 ;
        RECT 263.720 167.765 264.000 176.795 ;
        RECT 264.600 167.765 264.880 176.795 ;
        RECT 265.480 167.765 265.760 176.795 ;
        RECT 266.360 167.765 266.640 176.795 ;
        RECT 267.240 167.765 267.520 176.795 ;
        RECT 268.120 167.765 268.400 176.795 ;
        RECT 269.000 167.765 269.280 176.795 ;
        RECT 269.880 167.765 270.160 176.795 ;
        RECT 270.760 167.765 271.040 176.795 ;
        RECT 271.640 167.765 271.920 176.795 ;
        RECT 272.520 167.765 272.800 176.795 ;
        RECT 273.400 167.765 273.680 176.795 ;
        RECT 274.280 167.765 274.560 176.795 ;
        RECT 275.160 167.765 275.440 176.795 ;
        RECT 276.040 167.765 276.320 176.795 ;
        RECT 276.920 167.765 277.200 176.795 ;
        RECT 277.800 167.765 278.080 176.795 ;
        RECT 278.680 167.765 278.960 176.795 ;
        RECT 279.560 167.765 279.840 176.795 ;
        RECT 280.245 167.575 280.535 177.555 ;
        RECT 238.385 167.285 240.755 167.575 ;
        RECT 276.405 167.285 280.535 167.575 ;
        RECT 238.385 167.005 238.675 167.285 ;
        RECT 280.245 167.005 280.535 167.285 ;
        RECT 238.385 166.715 280.535 167.005 ;
        RECT 208.045 165.190 237.875 165.480 ;
        RECT 208.045 164.910 208.335 165.190 ;
        RECT 237.585 164.910 237.875 165.190 ;
        RECT 208.045 164.620 212.175 164.910 ;
        RECT 233.745 164.620 237.875 164.910 ;
        RECT 208.045 154.640 208.335 164.620 ;
        RECT 208.740 155.400 209.020 164.430 ;
        RECT 209.620 155.400 209.900 164.430 ;
        RECT 210.500 155.400 210.780 164.430 ;
        RECT 211.380 155.400 211.660 164.430 ;
        RECT 212.260 155.400 212.540 164.430 ;
        RECT 213.140 155.400 213.420 164.430 ;
        RECT 214.020 155.400 214.300 164.430 ;
        RECT 214.900 155.400 215.180 164.430 ;
        RECT 215.780 155.400 216.060 164.430 ;
        RECT 216.660 155.400 216.940 164.430 ;
        RECT 217.540 155.400 217.820 164.430 ;
        RECT 218.420 155.400 218.700 164.430 ;
        RECT 219.300 155.400 219.580 164.430 ;
        RECT 220.180 155.400 220.460 164.430 ;
        RECT 221.060 155.400 221.340 164.430 ;
        RECT 221.940 155.400 222.220 164.430 ;
        RECT 222.820 155.400 223.100 164.430 ;
        RECT 223.700 155.400 223.980 164.430 ;
        RECT 224.580 155.400 224.860 164.430 ;
        RECT 225.460 155.400 225.740 164.430 ;
        RECT 226.340 155.400 226.620 164.430 ;
        RECT 227.220 155.400 227.500 164.430 ;
        RECT 228.100 155.400 228.380 164.430 ;
        RECT 228.980 155.400 229.260 164.430 ;
        RECT 229.860 155.400 230.140 164.430 ;
        RECT 230.740 155.400 231.020 164.430 ;
        RECT 231.620 155.400 231.900 164.430 ;
        RECT 232.500 155.400 232.780 164.430 ;
        RECT 233.380 155.400 233.660 164.430 ;
        RECT 234.260 155.400 234.540 164.430 ;
        RECT 235.140 155.400 235.420 164.430 ;
        RECT 236.020 155.400 236.300 164.430 ;
        RECT 236.900 155.400 237.180 164.430 ;
        RECT 212.625 154.920 233.295 155.250 ;
        RECT 237.585 154.640 237.875 164.620 ;
        RECT 208.045 154.350 237.875 154.640 ;
        RECT 238.385 165.190 280.535 165.480 ;
        RECT 238.385 164.910 238.675 165.190 ;
        RECT 280.245 164.910 280.535 165.190 ;
        RECT 238.385 164.620 240.755 164.910 ;
        RECT 276.405 164.620 280.535 164.910 ;
        RECT 238.385 154.640 238.675 164.620 ;
        RECT 239.080 155.400 239.360 164.430 ;
        RECT 239.960 155.400 240.240 164.430 ;
        RECT 240.840 155.400 241.120 164.430 ;
        RECT 241.720 155.400 242.000 164.430 ;
        RECT 242.600 155.400 242.880 164.430 ;
        RECT 243.480 155.400 243.760 164.430 ;
        RECT 244.360 155.400 244.640 164.430 ;
        RECT 245.240 155.400 245.520 164.430 ;
        RECT 246.120 155.400 246.400 164.430 ;
        RECT 247.000 155.400 247.280 164.430 ;
        RECT 247.880 155.400 248.160 164.430 ;
        RECT 248.760 155.400 249.040 164.430 ;
        RECT 249.640 155.400 249.920 164.430 ;
        RECT 250.520 155.400 250.800 164.430 ;
        RECT 251.400 155.400 251.680 164.430 ;
        RECT 252.280 155.400 252.560 164.430 ;
        RECT 253.160 155.400 253.440 164.430 ;
        RECT 254.040 155.400 254.320 164.430 ;
        RECT 254.920 155.400 255.200 164.430 ;
        RECT 255.800 155.400 256.080 164.430 ;
        RECT 256.680 155.400 256.960 164.430 ;
        RECT 257.560 155.400 257.840 164.430 ;
        RECT 258.440 155.400 258.720 164.430 ;
        RECT 259.320 155.400 259.600 164.430 ;
        RECT 260.200 155.400 260.480 164.430 ;
        RECT 261.080 155.400 261.360 164.430 ;
        RECT 261.960 155.400 262.240 164.430 ;
        RECT 262.840 155.400 263.120 164.430 ;
        RECT 263.720 155.400 264.000 164.430 ;
        RECT 264.600 155.400 264.880 164.430 ;
        RECT 265.480 155.400 265.760 164.430 ;
        RECT 266.360 155.400 266.640 164.430 ;
        RECT 267.240 155.400 267.520 164.430 ;
        RECT 268.120 155.400 268.400 164.430 ;
        RECT 269.000 155.400 269.280 164.430 ;
        RECT 269.880 155.400 270.160 164.430 ;
        RECT 270.760 155.400 271.040 164.430 ;
        RECT 271.640 155.400 271.920 164.430 ;
        RECT 272.520 155.400 272.800 164.430 ;
        RECT 273.400 155.400 273.680 164.430 ;
        RECT 274.280 155.400 274.560 164.430 ;
        RECT 275.160 155.400 275.440 164.430 ;
        RECT 276.040 155.400 276.320 164.430 ;
        RECT 276.920 155.400 277.200 164.430 ;
        RECT 277.800 155.400 278.080 164.430 ;
        RECT 278.680 155.400 278.960 164.430 ;
        RECT 279.560 155.400 279.840 164.430 ;
        RECT 241.205 154.920 275.955 155.250 ;
        RECT 280.245 154.640 280.535 164.620 ;
        RECT 238.385 154.350 280.535 154.640 ;
        RECT 185.685 149.505 186.995 151.610 ;
        RECT 187.695 149.505 189.005 151.610 ;
        RECT 189.705 149.505 191.015 151.610 ;
        RECT 191.715 149.505 193.025 151.610 ;
        RECT 193.725 149.505 195.035 151.610 ;
        RECT 195.735 149.505 197.045 151.610 ;
        RECT 197.745 149.505 199.055 151.610 ;
        RECT 199.755 149.505 201.065 151.610 ;
        RECT 201.765 149.505 203.075 151.610 ;
        RECT 203.775 149.505 205.085 151.610 ;
        RECT 205.785 149.505 207.095 151.610 ;
        RECT 207.795 149.505 209.105 151.610 ;
        RECT 209.805 149.505 211.115 151.610 ;
        RECT 211.815 149.505 213.125 151.610 ;
        RECT 213.825 149.505 215.135 151.610 ;
        RECT 215.835 149.505 217.145 151.610 ;
        RECT 217.845 149.505 219.155 151.610 ;
        RECT 219.855 149.505 221.165 151.610 ;
        RECT 221.865 149.505 223.175 151.610 ;
        RECT 223.875 149.505 225.185 151.610 ;
        RECT 225.885 149.505 227.195 151.610 ;
        RECT 227.895 149.505 229.205 151.610 ;
        RECT 229.905 149.505 231.215 151.610 ;
        RECT 231.915 149.505 233.225 151.610 ;
        RECT 233.925 149.505 235.235 151.610 ;
        RECT 235.935 149.505 237.245 151.610 ;
        RECT 237.945 149.505 239.255 151.610 ;
        RECT 239.955 149.505 241.265 151.610 ;
        RECT 241.965 149.505 243.275 151.610 ;
        RECT 243.975 149.505 245.285 151.610 ;
        RECT 245.985 149.505 247.295 151.610 ;
        RECT 247.995 149.505 249.305 151.610 ;
        RECT 250.005 149.505 251.315 151.610 ;
        RECT 252.015 149.505 253.325 151.610 ;
        RECT 254.025 149.505 255.335 151.610 ;
        RECT 256.035 149.505 257.345 151.610 ;
        RECT 258.045 149.505 259.355 151.610 ;
        RECT 260.055 149.505 261.365 151.610 ;
        RECT 262.065 149.505 263.375 151.610 ;
        RECT 264.075 149.505 265.385 151.610 ;
        RECT 266.085 149.505 267.395 151.610 ;
        RECT 268.095 149.505 269.405 151.610 ;
        RECT 270.105 149.505 271.415 151.610 ;
        RECT 272.115 149.505 273.425 151.610 ;
        RECT 274.125 149.505 275.435 151.610 ;
        RECT 276.135 149.505 277.445 151.610 ;
        RECT 278.145 149.505 279.455 151.610 ;
        RECT 280.155 149.505 281.465 151.610 ;
        RECT 282.165 149.505 283.475 151.610 ;
        RECT 284.175 149.505 285.485 151.610 ;
        RECT 286.185 149.505 287.495 151.610 ;
        RECT 288.195 149.505 289.505 151.610 ;
        RECT 290.205 149.505 291.515 151.610 ;
        RECT 292.215 149.505 293.525 151.610 ;
        RECT 301.220 149.505 302.530 151.610 ;
        RECT 303.230 149.505 304.540 151.610 ;
        RECT 305.240 149.505 306.550 151.610 ;
        RECT 307.250 149.505 308.560 151.610 ;
        RECT 309.260 149.505 310.570 151.610 ;
        RECT 311.270 149.505 312.580 151.610 ;
        RECT 313.280 149.505 314.590 151.610 ;
        RECT 315.290 149.505 316.600 151.610 ;
        RECT 317.300 149.505 318.610 151.610 ;
        RECT 319.310 149.505 320.620 151.610 ;
        RECT 321.320 149.505 322.630 151.610 ;
        RECT 323.330 149.505 324.640 151.610 ;
        RECT 325.340 149.505 326.650 151.610 ;
        RECT 327.350 149.505 328.660 151.610 ;
        RECT 329.360 149.505 330.670 151.610 ;
        RECT 331.370 149.505 332.680 151.610 ;
        RECT 333.380 149.505 334.690 151.610 ;
        RECT 335.390 149.505 336.700 151.610 ;
        RECT 337.400 149.505 338.710 151.610 ;
        RECT 339.410 149.505 340.720 151.610 ;
        RECT 341.420 149.505 342.730 151.610 ;
        RECT 343.430 149.505 344.740 151.610 ;
        RECT 345.440 149.505 346.750 151.610 ;
        RECT 347.450 149.505 348.760 151.610 ;
        RECT 349.460 149.505 350.770 151.610 ;
        RECT 351.470 149.505 352.780 151.610 ;
        RECT 353.480 149.505 354.790 151.610 ;
        RECT 355.490 149.505 356.800 151.610 ;
        RECT 357.500 149.505 358.810 151.610 ;
        RECT 359.510 149.505 360.820 151.610 ;
        RECT 361.520 149.505 362.830 151.610 ;
        RECT 363.530 149.505 364.840 151.610 ;
        RECT 365.540 149.505 366.850 151.610 ;
        RECT 367.550 149.505 368.860 151.610 ;
        RECT 369.560 149.505 370.870 151.610 ;
        RECT 371.570 149.505 372.880 151.610 ;
        RECT 373.580 149.505 374.890 151.610 ;
        RECT 375.590 149.505 376.900 151.610 ;
        RECT 377.600 149.505 378.910 151.610 ;
        RECT 379.610 149.505 380.920 151.610 ;
        RECT 381.620 149.505 382.930 151.610 ;
        RECT 383.630 149.505 384.940 151.610 ;
        RECT 385.640 149.505 386.950 151.610 ;
        RECT 387.650 149.505 388.960 151.610 ;
        RECT 389.660 149.505 390.970 151.610 ;
        RECT 391.670 149.505 392.980 151.610 ;
        RECT 393.680 149.505 394.990 151.610 ;
        RECT 395.690 149.505 397.000 151.610 ;
        RECT 397.700 149.505 399.010 151.610 ;
        RECT 399.710 149.505 401.020 151.610 ;
        RECT 401.720 149.505 403.030 151.610 ;
        RECT 403.730 149.505 405.040 151.610 ;
        RECT 405.740 149.505 407.050 151.610 ;
        RECT 407.750 149.505 409.060 151.610 ;
        RECT 184.800 144.775 185.060 146.775 ;
        RECT 294.150 144.775 294.410 146.775 ;
        RECT 300.335 144.775 300.595 146.775 ;
        RECT 409.685 144.775 409.945 146.775 ;
        RECT 185.685 139.910 186.995 142.015 ;
        RECT 187.695 139.910 189.005 142.015 ;
        RECT 189.705 139.910 191.015 142.015 ;
        RECT 191.715 139.910 193.025 142.015 ;
        RECT 193.725 139.910 195.035 142.015 ;
        RECT 195.735 139.910 197.045 142.015 ;
        RECT 197.745 139.910 199.055 142.015 ;
        RECT 199.755 139.910 201.065 142.015 ;
        RECT 201.765 139.910 203.075 142.015 ;
        RECT 203.775 139.910 205.085 142.015 ;
        RECT 205.785 139.910 207.095 142.015 ;
        RECT 207.795 139.910 209.105 142.015 ;
        RECT 209.805 139.910 211.115 142.015 ;
        RECT 211.815 139.910 213.125 142.015 ;
        RECT 213.825 139.910 215.135 142.015 ;
        RECT 215.835 139.910 217.145 142.015 ;
        RECT 217.845 139.910 219.155 142.015 ;
        RECT 219.855 139.910 221.165 142.015 ;
        RECT 221.865 139.910 223.175 142.015 ;
        RECT 223.875 139.910 225.185 142.015 ;
        RECT 225.885 139.910 227.195 142.015 ;
        RECT 227.895 139.910 229.205 142.015 ;
        RECT 229.905 139.910 231.215 142.015 ;
        RECT 231.915 139.910 233.225 142.015 ;
        RECT 233.925 139.910 235.235 142.015 ;
        RECT 235.935 139.910 237.245 142.015 ;
        RECT 237.945 139.910 239.255 142.015 ;
        RECT 239.955 139.910 241.265 142.015 ;
        RECT 241.965 139.910 243.275 142.015 ;
        RECT 243.975 139.910 245.285 142.015 ;
        RECT 245.985 139.910 247.295 142.015 ;
        RECT 247.995 139.910 249.305 142.015 ;
        RECT 250.005 139.910 251.315 142.015 ;
        RECT 252.015 139.910 253.325 142.015 ;
        RECT 254.025 139.910 255.335 142.015 ;
        RECT 256.035 139.910 257.345 142.015 ;
        RECT 258.045 139.910 259.355 142.015 ;
        RECT 260.055 139.910 261.365 142.015 ;
        RECT 262.065 139.910 263.375 142.015 ;
        RECT 264.075 139.910 265.385 142.015 ;
        RECT 266.085 139.910 267.395 142.015 ;
        RECT 268.095 139.910 269.405 142.015 ;
        RECT 270.105 139.910 271.415 142.015 ;
        RECT 272.115 139.910 273.425 142.015 ;
        RECT 274.125 139.910 275.435 142.015 ;
        RECT 276.135 139.910 277.445 142.015 ;
        RECT 278.145 139.910 279.455 142.015 ;
        RECT 280.155 139.910 281.465 142.015 ;
        RECT 282.165 139.910 283.475 142.015 ;
        RECT 284.175 139.910 285.485 142.015 ;
        RECT 286.185 139.910 287.495 142.015 ;
        RECT 288.195 139.910 289.505 142.015 ;
        RECT 290.205 139.910 291.515 142.015 ;
        RECT 292.215 139.910 293.525 142.015 ;
        RECT 301.220 139.910 302.530 142.015 ;
        RECT 303.230 139.910 304.540 142.015 ;
        RECT 305.240 139.910 306.550 142.015 ;
        RECT 307.250 139.910 308.560 142.015 ;
        RECT 309.260 139.910 310.570 142.015 ;
        RECT 311.270 139.910 312.580 142.015 ;
        RECT 313.280 139.910 314.590 142.015 ;
        RECT 315.290 139.910 316.600 142.015 ;
        RECT 317.300 139.910 318.610 142.015 ;
        RECT 319.310 139.910 320.620 142.015 ;
        RECT 321.320 139.910 322.630 142.015 ;
        RECT 323.330 139.910 324.640 142.015 ;
        RECT 325.340 139.910 326.650 142.015 ;
        RECT 327.350 139.910 328.660 142.015 ;
        RECT 329.360 139.910 330.670 142.015 ;
        RECT 331.370 139.910 332.680 142.015 ;
        RECT 333.380 139.910 334.690 142.015 ;
        RECT 335.390 139.910 336.700 142.015 ;
        RECT 337.400 139.910 338.710 142.015 ;
        RECT 339.410 139.910 340.720 142.015 ;
        RECT 341.420 139.910 342.730 142.015 ;
        RECT 343.430 139.910 344.740 142.015 ;
        RECT 345.440 139.910 346.750 142.015 ;
        RECT 347.450 139.910 348.760 142.015 ;
        RECT 349.460 139.910 350.770 142.015 ;
        RECT 351.470 139.910 352.780 142.015 ;
        RECT 353.480 139.910 354.790 142.015 ;
        RECT 355.490 139.910 356.800 142.015 ;
        RECT 357.500 139.910 358.810 142.015 ;
        RECT 359.510 139.910 360.820 142.015 ;
        RECT 361.520 139.910 362.830 142.015 ;
        RECT 363.530 139.910 364.840 142.015 ;
        RECT 365.540 139.910 366.850 142.015 ;
        RECT 367.550 139.910 368.860 142.015 ;
        RECT 369.560 139.910 370.870 142.015 ;
        RECT 371.570 139.910 372.880 142.015 ;
        RECT 373.580 139.910 374.890 142.015 ;
        RECT 375.590 139.910 376.900 142.015 ;
        RECT 377.600 139.910 378.910 142.015 ;
        RECT 379.610 139.910 380.920 142.015 ;
        RECT 381.620 139.910 382.930 142.015 ;
        RECT 383.630 139.910 384.940 142.015 ;
        RECT 385.640 139.910 386.950 142.015 ;
        RECT 387.650 139.910 388.960 142.015 ;
        RECT 389.660 139.910 390.970 142.015 ;
        RECT 391.670 139.910 392.980 142.015 ;
        RECT 393.680 139.910 394.990 142.015 ;
        RECT 395.690 139.910 397.000 142.015 ;
        RECT 397.700 139.910 399.010 142.015 ;
        RECT 399.710 139.910 401.020 142.015 ;
        RECT 401.720 139.910 403.030 142.015 ;
        RECT 403.730 139.910 405.040 142.015 ;
        RECT 405.740 139.910 407.050 142.015 ;
        RECT 407.750 139.910 409.060 142.015 ;
        RECT 185.685 135.340 186.995 137.445 ;
        RECT 187.695 135.340 189.005 137.445 ;
        RECT 189.705 135.340 191.015 137.445 ;
        RECT 191.715 135.340 193.025 137.445 ;
        RECT 193.725 135.340 195.035 137.445 ;
        RECT 195.735 135.340 197.045 137.445 ;
        RECT 197.745 135.340 199.055 137.445 ;
        RECT 199.755 135.340 201.065 137.445 ;
        RECT 201.765 135.340 203.075 137.445 ;
        RECT 203.775 135.340 205.085 137.445 ;
        RECT 205.785 135.340 207.095 137.445 ;
        RECT 207.795 135.340 209.105 137.445 ;
        RECT 209.805 135.340 211.115 137.445 ;
        RECT 211.815 135.340 213.125 137.445 ;
        RECT 213.825 135.340 215.135 137.445 ;
        RECT 215.835 135.340 217.145 137.445 ;
        RECT 217.845 135.340 219.155 137.445 ;
        RECT 219.855 135.340 221.165 137.445 ;
        RECT 221.865 135.340 223.175 137.445 ;
        RECT 223.875 135.340 225.185 137.445 ;
        RECT 225.885 135.340 227.195 137.445 ;
        RECT 227.895 135.340 229.205 137.445 ;
        RECT 229.905 135.340 231.215 137.445 ;
        RECT 231.915 135.340 233.225 137.445 ;
        RECT 233.925 135.340 235.235 137.445 ;
        RECT 235.935 135.340 237.245 137.445 ;
        RECT 237.945 135.340 239.255 137.445 ;
        RECT 239.955 135.340 241.265 137.445 ;
        RECT 241.965 135.340 243.275 137.445 ;
        RECT 243.975 135.340 245.285 137.445 ;
        RECT 245.985 135.340 247.295 137.445 ;
        RECT 247.995 135.340 249.305 137.445 ;
        RECT 250.005 135.340 251.315 137.445 ;
        RECT 252.015 135.340 253.325 137.445 ;
        RECT 254.025 135.340 255.335 137.445 ;
        RECT 256.035 135.340 257.345 137.445 ;
        RECT 258.045 135.340 259.355 137.445 ;
        RECT 260.055 135.340 261.365 137.445 ;
        RECT 262.065 135.340 263.375 137.445 ;
        RECT 264.075 135.340 265.385 137.445 ;
        RECT 266.085 135.340 267.395 137.445 ;
        RECT 268.095 135.340 269.405 137.445 ;
        RECT 270.105 135.340 271.415 137.445 ;
        RECT 272.115 135.340 273.425 137.445 ;
        RECT 274.125 135.340 275.435 137.445 ;
        RECT 276.135 135.340 277.445 137.445 ;
        RECT 278.145 135.340 279.455 137.445 ;
        RECT 280.155 135.340 281.465 137.445 ;
        RECT 282.165 135.340 283.475 137.445 ;
        RECT 284.175 135.340 285.485 137.445 ;
        RECT 286.185 135.340 287.495 137.445 ;
        RECT 288.195 135.340 289.505 137.445 ;
        RECT 290.205 135.340 291.515 137.445 ;
        RECT 292.215 135.340 293.525 137.445 ;
        RECT 301.220 135.340 302.530 137.445 ;
        RECT 303.230 135.340 304.540 137.445 ;
        RECT 305.240 135.340 306.550 137.445 ;
        RECT 307.250 135.340 308.560 137.445 ;
        RECT 309.260 135.340 310.570 137.445 ;
        RECT 311.270 135.340 312.580 137.445 ;
        RECT 313.280 135.340 314.590 137.445 ;
        RECT 315.290 135.340 316.600 137.445 ;
        RECT 317.300 135.340 318.610 137.445 ;
        RECT 319.310 135.340 320.620 137.445 ;
        RECT 321.320 135.340 322.630 137.445 ;
        RECT 323.330 135.340 324.640 137.445 ;
        RECT 325.340 135.340 326.650 137.445 ;
        RECT 327.350 135.340 328.660 137.445 ;
        RECT 329.360 135.340 330.670 137.445 ;
        RECT 331.370 135.340 332.680 137.445 ;
        RECT 333.380 135.340 334.690 137.445 ;
        RECT 335.390 135.340 336.700 137.445 ;
        RECT 337.400 135.340 338.710 137.445 ;
        RECT 339.410 135.340 340.720 137.445 ;
        RECT 341.420 135.340 342.730 137.445 ;
        RECT 343.430 135.340 344.740 137.445 ;
        RECT 345.440 135.340 346.750 137.445 ;
        RECT 347.450 135.340 348.760 137.445 ;
        RECT 349.460 135.340 350.770 137.445 ;
        RECT 351.470 135.340 352.780 137.445 ;
        RECT 353.480 135.340 354.790 137.445 ;
        RECT 355.490 135.340 356.800 137.445 ;
        RECT 357.500 135.340 358.810 137.445 ;
        RECT 359.510 135.340 360.820 137.445 ;
        RECT 361.520 135.340 362.830 137.445 ;
        RECT 363.530 135.340 364.840 137.445 ;
        RECT 365.540 135.340 366.850 137.445 ;
        RECT 367.550 135.340 368.860 137.445 ;
        RECT 369.560 135.340 370.870 137.445 ;
        RECT 371.570 135.340 372.880 137.445 ;
        RECT 373.580 135.340 374.890 137.445 ;
        RECT 375.590 135.340 376.900 137.445 ;
        RECT 377.600 135.340 378.910 137.445 ;
        RECT 379.610 135.340 380.920 137.445 ;
        RECT 381.620 135.340 382.930 137.445 ;
        RECT 383.630 135.340 384.940 137.445 ;
        RECT 385.640 135.340 386.950 137.445 ;
        RECT 387.650 135.340 388.960 137.445 ;
        RECT 389.660 135.340 390.970 137.445 ;
        RECT 391.670 135.340 392.980 137.445 ;
        RECT 393.680 135.340 394.990 137.445 ;
        RECT 395.690 135.340 397.000 137.445 ;
        RECT 397.700 135.340 399.010 137.445 ;
        RECT 399.710 135.340 401.020 137.445 ;
        RECT 401.720 135.340 403.030 137.445 ;
        RECT 403.730 135.340 405.040 137.445 ;
        RECT 405.740 135.340 407.050 137.445 ;
        RECT 407.750 135.340 409.060 137.445 ;
        RECT 184.800 130.610 185.060 132.610 ;
        RECT 294.150 130.610 294.410 132.610 ;
        RECT 300.335 130.610 300.595 132.610 ;
        RECT 409.685 130.610 409.945 132.610 ;
        RECT 185.685 125.745 186.995 127.850 ;
        RECT 187.695 125.745 189.005 127.850 ;
        RECT 189.705 125.745 191.015 127.850 ;
        RECT 191.715 125.745 193.025 127.850 ;
        RECT 193.725 125.745 195.035 127.850 ;
        RECT 195.735 125.745 197.045 127.850 ;
        RECT 197.745 125.745 199.055 127.850 ;
        RECT 199.755 125.745 201.065 127.850 ;
        RECT 201.765 125.745 203.075 127.850 ;
        RECT 203.775 125.745 205.085 127.850 ;
        RECT 205.785 125.745 207.095 127.850 ;
        RECT 207.795 125.745 209.105 127.850 ;
        RECT 209.805 125.745 211.115 127.850 ;
        RECT 211.815 125.745 213.125 127.850 ;
        RECT 213.825 125.745 215.135 127.850 ;
        RECT 215.835 125.745 217.145 127.850 ;
        RECT 217.845 125.745 219.155 127.850 ;
        RECT 219.855 125.745 221.165 127.850 ;
        RECT 221.865 125.745 223.175 127.850 ;
        RECT 223.875 125.745 225.185 127.850 ;
        RECT 225.885 125.745 227.195 127.850 ;
        RECT 227.895 125.745 229.205 127.850 ;
        RECT 229.905 125.745 231.215 127.850 ;
        RECT 231.915 125.745 233.225 127.850 ;
        RECT 233.925 125.745 235.235 127.850 ;
        RECT 235.935 125.745 237.245 127.850 ;
        RECT 237.945 125.745 239.255 127.850 ;
        RECT 239.955 125.745 241.265 127.850 ;
        RECT 241.965 125.745 243.275 127.850 ;
        RECT 243.975 125.745 245.285 127.850 ;
        RECT 245.985 125.745 247.295 127.850 ;
        RECT 247.995 125.745 249.305 127.850 ;
        RECT 250.005 125.745 251.315 127.850 ;
        RECT 252.015 125.745 253.325 127.850 ;
        RECT 254.025 125.745 255.335 127.850 ;
        RECT 256.035 125.745 257.345 127.850 ;
        RECT 258.045 125.745 259.355 127.850 ;
        RECT 260.055 125.745 261.365 127.850 ;
        RECT 262.065 125.745 263.375 127.850 ;
        RECT 264.075 125.745 265.385 127.850 ;
        RECT 266.085 125.745 267.395 127.850 ;
        RECT 268.095 125.745 269.405 127.850 ;
        RECT 270.105 125.745 271.415 127.850 ;
        RECT 272.115 125.745 273.425 127.850 ;
        RECT 274.125 125.745 275.435 127.850 ;
        RECT 276.135 125.745 277.445 127.850 ;
        RECT 278.145 125.745 279.455 127.850 ;
        RECT 280.155 125.745 281.465 127.850 ;
        RECT 282.165 125.745 283.475 127.850 ;
        RECT 284.175 125.745 285.485 127.850 ;
        RECT 286.185 125.745 287.495 127.850 ;
        RECT 288.195 125.745 289.505 127.850 ;
        RECT 290.205 125.745 291.515 127.850 ;
        RECT 292.215 125.745 293.525 127.850 ;
        RECT 301.220 125.745 302.530 127.850 ;
        RECT 303.230 125.745 304.540 127.850 ;
        RECT 305.240 125.745 306.550 127.850 ;
        RECT 307.250 125.745 308.560 127.850 ;
        RECT 309.260 125.745 310.570 127.850 ;
        RECT 311.270 125.745 312.580 127.850 ;
        RECT 313.280 125.745 314.590 127.850 ;
        RECT 315.290 125.745 316.600 127.850 ;
        RECT 317.300 125.745 318.610 127.850 ;
        RECT 319.310 125.745 320.620 127.850 ;
        RECT 321.320 125.745 322.630 127.850 ;
        RECT 323.330 125.745 324.640 127.850 ;
        RECT 325.340 125.745 326.650 127.850 ;
        RECT 327.350 125.745 328.660 127.850 ;
        RECT 329.360 125.745 330.670 127.850 ;
        RECT 331.370 125.745 332.680 127.850 ;
        RECT 333.380 125.745 334.690 127.850 ;
        RECT 335.390 125.745 336.700 127.850 ;
        RECT 337.400 125.745 338.710 127.850 ;
        RECT 339.410 125.745 340.720 127.850 ;
        RECT 341.420 125.745 342.730 127.850 ;
        RECT 343.430 125.745 344.740 127.850 ;
        RECT 345.440 125.745 346.750 127.850 ;
        RECT 347.450 125.745 348.760 127.850 ;
        RECT 349.460 125.745 350.770 127.850 ;
        RECT 351.470 125.745 352.780 127.850 ;
        RECT 353.480 125.745 354.790 127.850 ;
        RECT 355.490 125.745 356.800 127.850 ;
        RECT 357.500 125.745 358.810 127.850 ;
        RECT 359.510 125.745 360.820 127.850 ;
        RECT 361.520 125.745 362.830 127.850 ;
        RECT 363.530 125.745 364.840 127.850 ;
        RECT 365.540 125.745 366.850 127.850 ;
        RECT 367.550 125.745 368.860 127.850 ;
        RECT 369.560 125.745 370.870 127.850 ;
        RECT 371.570 125.745 372.880 127.850 ;
        RECT 373.580 125.745 374.890 127.850 ;
        RECT 375.590 125.745 376.900 127.850 ;
        RECT 377.600 125.745 378.910 127.850 ;
        RECT 379.610 125.745 380.920 127.850 ;
        RECT 381.620 125.745 382.930 127.850 ;
        RECT 383.630 125.745 384.940 127.850 ;
        RECT 385.640 125.745 386.950 127.850 ;
        RECT 387.650 125.745 388.960 127.850 ;
        RECT 389.660 125.745 390.970 127.850 ;
        RECT 391.670 125.745 392.980 127.850 ;
        RECT 393.680 125.745 394.990 127.850 ;
        RECT 395.690 125.745 397.000 127.850 ;
        RECT 397.700 125.745 399.010 127.850 ;
        RECT 399.710 125.745 401.020 127.850 ;
        RECT 401.720 125.745 403.030 127.850 ;
        RECT 403.730 125.745 405.040 127.850 ;
        RECT 405.740 125.745 407.050 127.850 ;
        RECT 407.750 125.745 409.060 127.850 ;
        RECT 310.855 120.475 333.725 120.765 ;
        RECT 310.855 117.185 311.145 120.475 ;
        RECT 318.995 119.825 325.585 120.155 ;
        RECT 311.590 117.375 311.870 119.635 ;
        RECT 312.470 117.375 312.750 119.635 ;
        RECT 313.350 117.375 313.630 119.635 ;
        RECT 314.230 117.375 314.510 119.635 ;
        RECT 315.110 117.375 315.390 119.635 ;
        RECT 315.990 117.375 316.270 119.635 ;
        RECT 316.870 117.375 317.150 119.635 ;
        RECT 317.750 117.375 318.030 119.635 ;
        RECT 318.630 117.375 318.910 119.635 ;
        RECT 319.510 117.375 319.790 119.635 ;
        RECT 320.390 117.375 320.670 119.635 ;
        RECT 321.270 117.375 321.550 119.635 ;
        RECT 322.150 117.375 322.430 119.635 ;
        RECT 323.030 117.375 323.310 119.635 ;
        RECT 323.910 117.375 324.190 119.635 ;
        RECT 324.790 117.375 325.070 119.635 ;
        RECT 325.670 117.375 325.950 119.635 ;
        RECT 326.550 117.375 326.830 119.635 ;
        RECT 327.430 117.375 327.710 119.635 ;
        RECT 328.310 117.375 328.590 119.635 ;
        RECT 329.190 117.375 329.470 119.635 ;
        RECT 330.070 117.375 330.350 119.635 ;
        RECT 330.950 117.375 331.230 119.635 ;
        RECT 331.830 117.375 332.110 119.635 ;
        RECT 332.710 117.375 332.990 119.635 ;
        RECT 333.435 117.185 333.725 120.475 ;
        RECT 310.855 116.895 318.545 117.185 ;
        RECT 326.035 116.895 333.725 117.185 ;
        RECT 184.740 114.985 198.410 115.275 ;
        RECT 184.740 113.395 185.030 114.985 ;
        RECT 185.425 113.585 185.685 114.585 ;
        RECT 185.855 113.585 186.115 114.585 ;
        RECT 186.285 113.585 186.545 114.585 ;
        RECT 186.700 113.585 186.960 114.585 ;
        RECT 187.145 113.585 187.405 114.585 ;
        RECT 187.560 113.585 187.820 114.585 ;
        RECT 188.005 113.585 188.265 114.585 ;
        RECT 188.420 113.585 188.680 114.585 ;
        RECT 188.865 113.585 189.125 114.585 ;
        RECT 189.280 113.585 189.540 114.585 ;
        RECT 189.725 113.585 189.985 114.585 ;
        RECT 190.155 113.585 190.415 114.585 ;
        RECT 190.585 113.585 190.845 114.585 ;
        RECT 191.030 113.585 191.290 114.585 ;
        RECT 191.445 113.585 191.705 114.585 ;
        RECT 191.890 113.585 192.150 114.585 ;
        RECT 192.305 113.585 192.565 114.585 ;
        RECT 192.750 113.585 193.010 114.585 ;
        RECT 193.165 113.585 193.425 114.585 ;
        RECT 193.610 113.585 193.870 114.585 ;
        RECT 194.025 113.585 194.285 114.585 ;
        RECT 194.470 113.585 194.730 114.585 ;
        RECT 194.885 113.585 195.145 114.585 ;
        RECT 195.330 113.585 195.590 114.585 ;
        RECT 195.745 113.585 196.005 114.585 ;
        RECT 196.190 113.585 196.450 114.585 ;
        RECT 196.605 113.585 196.865 114.585 ;
        RECT 197.035 113.585 197.295 114.585 ;
        RECT 197.465 113.585 197.725 114.585 ;
        RECT 198.120 113.395 198.410 114.985 ;
        RECT 218.010 114.750 219.320 116.855 ;
        RECT 220.020 114.750 221.330 116.855 ;
        RECT 222.030 116.305 223.340 116.855 ;
        RECT 224.040 116.305 225.350 116.855 ;
        RECT 226.050 116.305 227.360 116.855 ;
        RECT 228.060 116.305 229.370 116.855 ;
        RECT 230.070 116.305 231.380 116.855 ;
        RECT 232.080 116.305 233.390 116.855 ;
        RECT 234.090 116.305 235.400 116.855 ;
        RECT 236.100 116.305 237.410 116.855 ;
        RECT 222.030 115.305 237.410 116.305 ;
        RECT 222.030 114.750 223.340 115.305 ;
        RECT 224.040 114.750 225.350 115.305 ;
        RECT 226.050 114.750 227.360 115.305 ;
        RECT 228.060 114.750 229.370 115.305 ;
        RECT 230.070 114.750 231.380 115.305 ;
        RECT 232.080 114.750 233.390 115.305 ;
        RECT 234.090 114.750 235.400 115.305 ;
        RECT 236.100 114.750 237.410 115.305 ;
        RECT 238.110 116.305 239.420 116.855 ;
        RECT 240.120 116.305 241.430 116.855 ;
        RECT 238.110 115.305 241.430 116.305 ;
        RECT 238.110 114.750 239.420 115.305 ;
        RECT 240.120 114.750 241.430 115.305 ;
        RECT 242.130 116.305 243.440 116.855 ;
        RECT 244.140 116.305 245.450 116.855 ;
        RECT 242.130 115.305 245.450 116.305 ;
        RECT 242.130 114.750 243.440 115.305 ;
        RECT 244.140 114.750 245.450 115.305 ;
        RECT 246.150 116.305 247.460 116.855 ;
        RECT 248.160 116.305 249.470 116.855 ;
        RECT 246.150 115.305 249.470 116.305 ;
        RECT 246.150 114.750 247.460 115.305 ;
        RECT 248.160 114.750 249.470 115.305 ;
        RECT 250.170 116.305 251.480 116.855 ;
        RECT 252.180 116.305 253.490 116.855 ;
        RECT 250.170 115.305 253.490 116.305 ;
        RECT 250.170 114.750 251.480 115.305 ;
        RECT 252.180 114.750 253.490 115.305 ;
        RECT 254.190 116.305 255.500 116.855 ;
        RECT 256.200 116.305 257.510 116.855 ;
        RECT 254.190 115.305 257.510 116.305 ;
        RECT 254.190 114.750 255.500 115.305 ;
        RECT 256.200 114.750 257.510 115.305 ;
        RECT 258.210 116.305 259.520 116.855 ;
        RECT 260.220 116.305 261.530 116.855 ;
        RECT 258.210 115.305 261.530 116.305 ;
        RECT 258.210 114.750 259.520 115.305 ;
        RECT 260.220 114.750 261.530 115.305 ;
        RECT 262.230 116.305 263.540 116.855 ;
        RECT 264.240 116.305 265.550 116.855 ;
        RECT 262.230 115.305 265.550 116.305 ;
        RECT 262.230 114.750 263.540 115.305 ;
        RECT 264.240 114.750 265.550 115.305 ;
        RECT 266.250 116.305 267.560 116.855 ;
        RECT 268.260 116.305 269.570 116.855 ;
        RECT 266.250 115.305 269.570 116.305 ;
        RECT 266.250 114.750 267.560 115.305 ;
        RECT 268.260 114.750 269.570 115.305 ;
        RECT 270.270 116.305 271.580 116.855 ;
        RECT 272.280 116.305 273.590 116.855 ;
        RECT 270.270 115.305 273.590 116.305 ;
        RECT 270.270 114.750 271.580 115.305 ;
        RECT 272.280 114.750 273.590 115.305 ;
        RECT 274.290 116.305 275.600 116.855 ;
        RECT 276.300 116.305 277.610 116.855 ;
        RECT 274.290 115.305 277.610 116.305 ;
        RECT 274.290 114.750 275.600 115.305 ;
        RECT 276.300 114.750 277.610 115.305 ;
        RECT 278.310 116.305 279.620 116.855 ;
        RECT 280.320 116.305 281.630 116.855 ;
        RECT 278.310 115.305 281.630 116.305 ;
        RECT 278.310 114.750 279.620 115.305 ;
        RECT 280.320 114.750 281.630 115.305 ;
        RECT 282.330 116.305 283.640 116.855 ;
        RECT 284.340 116.305 285.650 116.855 ;
        RECT 282.330 115.305 285.650 116.305 ;
        RECT 282.330 114.750 283.640 115.305 ;
        RECT 284.340 114.750 285.650 115.305 ;
        RECT 286.350 114.750 287.660 116.855 ;
        RECT 288.360 114.750 289.670 116.855 ;
        RECT 310.855 116.535 311.145 116.895 ;
        RECT 333.435 116.535 333.725 116.895 ;
        RECT 310.855 116.245 333.725 116.535 ;
        RECT 334.075 120.475 363.985 120.765 ;
        RECT 334.075 117.185 334.365 120.475 ;
        RECT 347.495 119.825 350.565 120.115 ;
        RECT 334.810 117.375 335.090 119.635 ;
        RECT 335.690 117.375 335.970 119.635 ;
        RECT 336.570 117.375 336.850 119.635 ;
        RECT 337.450 117.375 337.730 119.635 ;
        RECT 338.330 117.375 338.610 119.635 ;
        RECT 339.210 117.375 339.490 119.635 ;
        RECT 340.090 117.375 340.370 119.635 ;
        RECT 340.970 117.375 341.250 119.635 ;
        RECT 341.850 117.375 342.130 119.635 ;
        RECT 342.730 117.375 343.010 119.635 ;
        RECT 343.610 117.375 343.890 119.635 ;
        RECT 344.490 117.375 344.770 119.635 ;
        RECT 345.370 117.375 345.650 119.635 ;
        RECT 346.250 117.375 346.530 119.635 ;
        RECT 347.130 117.375 347.410 119.635 ;
        RECT 348.010 117.375 348.290 119.825 ;
        RECT 348.890 117.375 349.170 119.635 ;
        RECT 349.770 117.375 350.050 119.825 ;
        RECT 350.650 117.375 350.930 119.635 ;
        RECT 351.530 117.375 351.810 119.635 ;
        RECT 352.410 117.375 352.690 119.635 ;
        RECT 353.290 117.375 353.570 119.635 ;
        RECT 354.170 117.375 354.450 119.635 ;
        RECT 355.050 117.375 355.330 119.635 ;
        RECT 355.930 117.375 356.210 119.635 ;
        RECT 356.810 117.375 357.090 119.635 ;
        RECT 357.690 117.375 357.970 119.635 ;
        RECT 358.570 117.375 358.850 119.635 ;
        RECT 359.450 117.375 359.730 119.635 ;
        RECT 360.330 117.375 360.610 119.635 ;
        RECT 361.210 117.375 361.490 119.635 ;
        RECT 362.090 117.375 362.370 119.635 ;
        RECT 362.970 117.375 363.250 119.635 ;
        RECT 363.695 117.185 363.985 120.475 ;
        RECT 334.075 116.895 340.005 117.185 ;
        RECT 340.455 116.895 357.605 117.185 ;
        RECT 358.055 116.895 363.985 117.185 ;
        RECT 334.075 116.535 334.365 116.895 ;
        RECT 363.695 116.535 363.985 116.895 ;
        RECT 334.075 116.245 363.985 116.535 ;
        RECT 364.415 120.475 406.640 120.765 ;
        RECT 364.415 117.185 364.705 120.475 ;
        RECT 365.150 117.375 365.430 119.635 ;
        RECT 366.030 117.375 366.310 119.635 ;
        RECT 366.910 117.375 367.190 119.635 ;
        RECT 367.790 117.375 368.070 119.635 ;
        RECT 368.670 117.375 368.950 119.635 ;
        RECT 369.550 117.375 369.830 119.635 ;
        RECT 370.430 117.375 370.710 119.635 ;
        RECT 371.310 117.375 371.590 119.635 ;
        RECT 372.190 117.375 372.470 119.635 ;
        RECT 373.070 117.375 373.350 119.635 ;
        RECT 373.950 117.375 374.230 119.635 ;
        RECT 374.830 117.375 375.110 119.635 ;
        RECT 375.710 117.375 375.990 119.635 ;
        RECT 376.590 117.375 376.870 119.635 ;
        RECT 377.470 117.375 377.750 119.635 ;
        RECT 378.350 117.375 378.630 119.635 ;
        RECT 379.230 117.375 379.510 119.635 ;
        RECT 380.110 117.375 380.390 119.635 ;
        RECT 380.990 117.375 381.270 119.635 ;
        RECT 381.870 117.375 382.150 119.635 ;
        RECT 382.750 117.375 383.030 119.635 ;
        RECT 383.630 117.375 383.910 119.635 ;
        RECT 384.510 117.375 384.790 119.635 ;
        RECT 385.390 117.375 385.670 119.635 ;
        RECT 386.270 117.375 386.550 119.635 ;
        RECT 387.150 117.375 387.430 119.635 ;
        RECT 388.030 117.375 388.310 119.635 ;
        RECT 388.910 117.375 389.190 119.635 ;
        RECT 389.790 117.375 390.070 119.635 ;
        RECT 390.670 117.375 390.950 119.635 ;
        RECT 391.550 117.375 391.830 119.635 ;
        RECT 392.430 117.375 392.710 119.635 ;
        RECT 393.310 117.375 393.590 119.635 ;
        RECT 394.190 117.375 394.470 119.635 ;
        RECT 395.070 117.375 395.350 119.635 ;
        RECT 395.950 117.375 396.230 119.635 ;
        RECT 396.830 117.375 397.110 119.635 ;
        RECT 397.710 117.375 397.990 119.635 ;
        RECT 398.590 117.375 398.870 119.635 ;
        RECT 399.470 117.375 399.750 119.635 ;
        RECT 400.350 117.375 400.630 119.635 ;
        RECT 401.230 117.375 401.510 119.635 ;
        RECT 402.110 117.375 402.390 119.635 ;
        RECT 402.990 117.375 403.270 119.635 ;
        RECT 403.870 117.375 404.150 119.635 ;
        RECT 404.750 117.375 405.030 119.635 ;
        RECT 405.630 117.375 405.910 119.635 ;
        RECT 406.350 119.005 406.640 120.475 ;
        RECT 406.350 118.005 406.645 119.005 ;
        RECT 444.015 118.795 452.685 119.085 ;
        RECT 406.350 117.185 406.640 118.005 ;
        RECT 364.415 116.895 366.825 117.185 ;
        RECT 367.275 116.895 402.025 117.185 ;
        RECT 402.475 116.895 406.640 117.185 ;
        RECT 364.415 116.535 364.705 116.895 ;
        RECT 406.350 116.535 406.640 116.895 ;
        RECT 364.415 116.245 406.640 116.535 ;
        RECT 310.855 113.990 333.725 114.280 ;
        RECT 184.740 113.125 186.275 113.395 ;
        RECT 186.555 113.125 196.595 113.395 ;
        RECT 196.875 113.125 198.410 113.395 ;
        RECT 184.740 112.565 185.030 113.125 ;
        RECT 191.410 112.535 191.740 113.125 ;
        RECT 198.120 112.565 198.410 113.125 ;
        RECT 199.820 113.125 213.490 113.415 ;
        RECT 199.820 112.675 200.110 113.125 ;
        RECT 213.200 112.675 213.490 113.125 ;
        RECT 185.490 112.205 191.740 112.535 ;
        RECT 184.740 111.620 185.030 112.180 ;
        RECT 191.410 111.620 191.740 112.205 ;
        RECT 199.820 112.385 201.360 112.675 ;
        RECT 211.950 112.385 213.490 112.675 ;
        RECT 198.120 111.620 198.410 112.180 ;
        RECT 184.740 111.350 189.715 111.620 ;
        RECT 189.995 111.350 193.155 111.620 ;
        RECT 193.435 111.350 198.410 111.620 ;
        RECT 184.740 109.790 185.030 111.350 ;
        RECT 185.425 110.160 185.685 111.160 ;
        RECT 185.855 110.160 186.115 111.160 ;
        RECT 186.285 110.160 186.545 111.160 ;
        RECT 186.715 110.160 186.975 111.160 ;
        RECT 187.145 110.160 187.405 111.160 ;
        RECT 187.575 110.160 187.835 111.160 ;
        RECT 188.005 110.160 188.265 111.160 ;
        RECT 188.435 110.160 188.695 111.160 ;
        RECT 188.865 110.160 189.125 111.160 ;
        RECT 189.295 110.160 189.555 111.160 ;
        RECT 189.725 110.160 189.985 111.160 ;
        RECT 190.155 110.160 190.415 111.160 ;
        RECT 190.585 110.160 190.845 111.160 ;
        RECT 191.030 110.160 191.290 111.160 ;
        RECT 191.445 110.160 191.705 111.160 ;
        RECT 191.890 110.160 192.150 111.160 ;
        RECT 192.305 110.160 192.565 111.160 ;
        RECT 192.750 110.160 193.010 111.160 ;
        RECT 193.165 110.160 193.425 111.160 ;
        RECT 193.595 110.160 193.855 111.160 ;
        RECT 194.025 110.160 194.285 111.160 ;
        RECT 194.455 110.160 194.715 111.160 ;
        RECT 194.885 110.160 195.145 111.160 ;
        RECT 195.315 110.160 195.575 111.160 ;
        RECT 195.745 110.160 196.005 111.160 ;
        RECT 196.175 110.160 196.435 111.160 ;
        RECT 196.605 110.160 196.865 111.160 ;
        RECT 197.035 110.160 197.295 111.160 ;
        RECT 197.480 110.160 197.710 111.350 ;
        RECT 198.120 109.790 198.410 111.350 ;
        RECT 199.820 110.175 200.110 112.385 ;
        RECT 200.505 111.345 200.765 112.195 ;
        RECT 200.935 111.345 201.195 112.195 ;
        RECT 200.520 111.195 200.750 111.345 ;
        RECT 200.950 111.195 201.180 111.345 ;
        RECT 201.365 111.195 201.625 112.195 ;
        RECT 201.795 111.195 202.055 112.195 ;
        RECT 202.240 111.195 202.500 112.195 ;
        RECT 202.670 111.195 202.930 112.195 ;
        RECT 203.100 111.195 203.360 112.195 ;
        RECT 203.530 111.195 203.790 112.195 ;
        RECT 203.960 111.195 204.220 112.195 ;
        RECT 204.390 111.195 204.650 112.195 ;
        RECT 204.820 111.195 205.080 112.195 ;
        RECT 205.250 111.195 205.510 112.195 ;
        RECT 205.680 111.195 205.940 112.195 ;
        RECT 206.110 111.195 206.370 112.195 ;
        RECT 206.540 111.195 206.800 112.195 ;
        RECT 206.970 111.195 207.230 112.195 ;
        RECT 207.400 111.195 207.660 112.195 ;
        RECT 207.830 111.195 208.090 112.195 ;
        RECT 208.260 111.195 208.520 112.195 ;
        RECT 208.690 111.195 208.950 112.195 ;
        RECT 209.120 111.195 209.380 112.195 ;
        RECT 209.550 111.195 209.810 112.195 ;
        RECT 209.980 111.195 210.240 112.195 ;
        RECT 210.410 111.195 210.670 112.195 ;
        RECT 210.840 111.195 211.100 112.195 ;
        RECT 211.270 111.195 211.530 112.195 ;
        RECT 211.700 111.195 211.960 112.195 ;
        RECT 212.115 111.345 212.375 112.195 ;
        RECT 212.545 111.345 212.805 112.195 ;
        RECT 212.130 111.195 212.360 111.345 ;
        RECT 212.560 111.195 212.790 111.345 ;
        RECT 200.310 110.725 211.675 111.005 ;
        RECT 213.200 110.175 213.490 112.385 ;
        RECT 310.855 110.700 311.145 113.990 ;
        RECT 318.975 113.340 325.585 113.670 ;
        RECT 311.590 110.890 311.870 113.150 ;
        RECT 312.470 110.890 312.750 113.150 ;
        RECT 313.350 110.890 313.630 113.150 ;
        RECT 314.230 110.890 314.510 113.150 ;
        RECT 315.110 110.890 315.390 113.150 ;
        RECT 315.990 110.890 316.270 113.150 ;
        RECT 316.870 110.890 317.150 113.150 ;
        RECT 317.750 110.890 318.030 113.150 ;
        RECT 318.630 110.890 318.910 113.150 ;
        RECT 319.510 110.890 319.790 113.150 ;
        RECT 320.390 110.890 320.670 113.150 ;
        RECT 321.270 110.890 321.550 113.150 ;
        RECT 322.150 110.890 322.430 113.150 ;
        RECT 323.030 110.890 323.310 113.150 ;
        RECT 323.910 110.890 324.190 113.150 ;
        RECT 324.790 110.890 325.070 113.150 ;
        RECT 325.670 110.890 325.950 113.150 ;
        RECT 326.550 110.890 326.830 113.150 ;
        RECT 327.430 110.890 327.710 113.150 ;
        RECT 328.310 110.890 328.590 113.150 ;
        RECT 329.190 110.890 329.470 113.150 ;
        RECT 330.070 110.890 330.350 113.150 ;
        RECT 330.950 110.890 331.230 113.150 ;
        RECT 331.830 110.890 332.110 113.150 ;
        RECT 332.710 110.890 332.990 113.150 ;
        RECT 333.435 110.700 333.725 113.990 ;
        RECT 310.855 110.410 318.545 110.700 ;
        RECT 326.035 110.410 333.725 110.700 ;
        RECT 184.740 109.500 198.410 109.790 ;
        RECT 184.740 107.940 185.030 109.500 ;
        RECT 185.425 108.130 185.685 109.130 ;
        RECT 185.855 108.130 186.115 109.130 ;
        RECT 186.285 108.130 186.545 109.130 ;
        RECT 186.715 108.130 186.975 109.130 ;
        RECT 187.145 108.130 187.405 109.130 ;
        RECT 187.575 108.130 187.835 109.130 ;
        RECT 188.005 108.130 188.265 109.130 ;
        RECT 188.435 108.130 188.695 109.130 ;
        RECT 188.865 108.130 189.125 109.130 ;
        RECT 189.295 108.130 189.555 109.130 ;
        RECT 189.725 108.130 189.985 109.130 ;
        RECT 190.155 108.130 190.415 109.130 ;
        RECT 190.585 108.130 190.845 109.130 ;
        RECT 191.030 108.130 191.290 109.130 ;
        RECT 191.445 108.130 191.705 109.130 ;
        RECT 191.890 108.130 192.150 109.130 ;
        RECT 192.305 108.130 192.565 109.130 ;
        RECT 192.750 108.130 193.010 109.130 ;
        RECT 193.165 108.130 193.425 109.130 ;
        RECT 193.595 108.130 193.855 109.130 ;
        RECT 194.025 108.130 194.285 109.130 ;
        RECT 194.455 108.130 194.715 109.130 ;
        RECT 194.885 108.130 195.145 109.130 ;
        RECT 195.315 108.130 195.575 109.130 ;
        RECT 195.745 108.130 196.005 109.130 ;
        RECT 196.175 108.130 196.435 109.130 ;
        RECT 196.605 108.130 196.865 109.130 ;
        RECT 197.035 108.130 197.295 109.130 ;
        RECT 197.480 107.940 197.710 109.130 ;
        RECT 198.120 107.940 198.410 109.500 ;
        RECT 184.740 107.670 189.715 107.940 ;
        RECT 189.995 107.670 193.155 107.940 ;
        RECT 193.435 107.670 198.410 107.940 ;
        RECT 184.740 107.110 185.030 107.670 ;
        RECT 191.410 107.085 191.740 107.670 ;
        RECT 196.775 107.235 197.735 107.515 ;
        RECT 196.775 107.085 197.105 107.235 ;
        RECT 198.120 107.110 198.410 107.670 ;
        RECT 191.410 106.755 197.105 107.085 ;
        RECT 199.820 106.905 200.110 109.415 ;
        RECT 200.310 108.285 211.675 108.565 ;
        RECT 200.520 107.945 200.750 108.095 ;
        RECT 200.950 107.945 201.180 108.095 ;
        RECT 201.380 107.945 201.610 108.095 ;
        RECT 201.810 107.945 202.040 108.095 ;
        RECT 202.240 107.945 202.470 108.095 ;
        RECT 202.670 107.945 202.900 108.095 ;
        RECT 203.100 107.945 203.330 108.095 ;
        RECT 203.530 107.945 203.760 108.095 ;
        RECT 203.960 107.945 204.190 108.095 ;
        RECT 204.390 107.945 204.620 108.095 ;
        RECT 200.505 107.095 200.765 107.945 ;
        RECT 200.935 107.095 201.195 107.945 ;
        RECT 201.365 107.095 201.625 107.945 ;
        RECT 201.795 107.095 202.055 107.945 ;
        RECT 202.225 107.095 202.485 107.945 ;
        RECT 202.655 107.095 202.915 107.945 ;
        RECT 203.085 107.095 203.345 107.945 ;
        RECT 203.515 107.095 203.775 107.945 ;
        RECT 203.945 107.095 204.205 107.945 ;
        RECT 204.375 107.095 204.635 107.945 ;
        RECT 204.820 107.095 205.080 108.095 ;
        RECT 205.250 107.095 205.510 108.095 ;
        RECT 205.680 107.095 205.940 108.095 ;
        RECT 206.110 107.095 206.370 108.095 ;
        RECT 206.540 107.095 206.800 108.095 ;
        RECT 206.970 107.095 207.230 108.095 ;
        RECT 207.400 107.095 207.660 108.095 ;
        RECT 207.830 107.095 208.090 108.095 ;
        RECT 208.260 107.095 208.520 108.095 ;
        RECT 208.690 107.945 208.920 108.095 ;
        RECT 209.120 107.945 209.350 108.095 ;
        RECT 209.550 107.945 209.780 108.095 ;
        RECT 209.980 107.945 210.210 108.095 ;
        RECT 210.410 107.945 210.640 108.095 ;
        RECT 210.840 107.945 211.070 108.095 ;
        RECT 211.270 107.945 211.500 108.095 ;
        RECT 211.700 107.945 211.930 108.095 ;
        RECT 212.130 107.945 212.360 108.095 ;
        RECT 212.560 107.945 212.790 108.095 ;
        RECT 208.675 107.095 208.935 107.945 ;
        RECT 209.105 107.095 209.365 107.945 ;
        RECT 209.535 107.095 209.795 107.945 ;
        RECT 209.965 107.095 210.225 107.945 ;
        RECT 210.395 107.095 210.655 107.945 ;
        RECT 210.825 107.095 211.085 107.945 ;
        RECT 211.255 107.095 211.515 107.945 ;
        RECT 211.685 107.095 211.945 107.945 ;
        RECT 212.115 107.095 212.375 107.945 ;
        RECT 212.545 107.095 212.805 107.945 ;
        RECT 213.200 106.905 213.490 109.415 ;
        RECT 217.110 108.145 217.400 110.145 ;
        RECT 290.280 108.145 290.570 110.145 ;
        RECT 310.855 110.050 311.145 110.410 ;
        RECT 333.435 110.050 333.725 110.410 ;
        RECT 310.855 109.760 333.725 110.050 ;
        RECT 334.075 113.990 363.985 114.280 ;
        RECT 334.075 110.700 334.365 113.990 ;
        RECT 337.730 113.340 357.605 113.670 ;
        RECT 334.810 110.890 335.090 113.150 ;
        RECT 335.690 110.890 335.970 113.150 ;
        RECT 336.570 110.890 336.850 113.150 ;
        RECT 337.450 110.890 337.730 113.150 ;
        RECT 338.330 110.890 338.610 113.150 ;
        RECT 339.210 110.890 339.490 113.150 ;
        RECT 340.090 110.890 340.370 113.150 ;
        RECT 340.970 110.890 341.250 113.150 ;
        RECT 341.850 110.890 342.130 113.150 ;
        RECT 342.730 110.890 343.010 113.150 ;
        RECT 343.610 110.890 343.890 113.150 ;
        RECT 344.490 110.890 344.770 113.150 ;
        RECT 345.370 110.890 345.650 113.150 ;
        RECT 346.250 110.890 346.530 113.150 ;
        RECT 347.130 110.890 347.410 113.150 ;
        RECT 348.010 110.700 348.290 113.150 ;
        RECT 348.890 110.700 349.170 113.150 ;
        RECT 349.770 110.700 350.050 113.150 ;
        RECT 350.650 110.890 350.930 113.150 ;
        RECT 351.530 110.890 351.810 113.150 ;
        RECT 352.410 110.890 352.690 113.150 ;
        RECT 353.290 110.890 353.570 113.150 ;
        RECT 354.170 110.890 354.450 113.150 ;
        RECT 355.050 110.890 355.330 113.150 ;
        RECT 355.930 110.890 356.210 113.150 ;
        RECT 356.810 110.890 357.090 113.150 ;
        RECT 357.690 110.890 357.970 113.150 ;
        RECT 358.570 110.890 358.850 113.150 ;
        RECT 359.450 110.890 359.730 113.150 ;
        RECT 360.330 110.890 360.610 113.150 ;
        RECT 361.210 110.890 361.490 113.150 ;
        RECT 362.090 110.890 362.370 113.150 ;
        RECT 362.970 110.890 363.250 113.150 ;
        RECT 363.695 110.700 363.985 113.990 ;
        RECT 334.075 110.410 340.005 110.700 ;
        RECT 347.495 110.410 350.565 110.700 ;
        RECT 358.055 110.410 363.985 110.700 ;
        RECT 334.075 110.050 334.365 110.410 ;
        RECT 363.695 110.050 363.985 110.410 ;
        RECT 334.075 109.760 363.985 110.050 ;
        RECT 364.415 113.990 406.640 114.280 ;
        RECT 364.415 110.700 364.705 113.990 ;
        RECT 365.245 113.340 402.025 113.670 ;
        RECT 365.150 110.890 365.430 113.150 ;
        RECT 366.030 110.890 366.310 113.150 ;
        RECT 366.910 110.890 367.190 113.150 ;
        RECT 367.790 110.890 368.070 113.150 ;
        RECT 368.670 110.890 368.950 113.150 ;
        RECT 369.550 110.890 369.830 113.150 ;
        RECT 370.430 110.890 370.710 113.150 ;
        RECT 371.310 110.890 371.590 113.150 ;
        RECT 372.190 110.890 372.470 113.150 ;
        RECT 373.070 110.890 373.350 113.150 ;
        RECT 373.950 110.890 374.230 113.150 ;
        RECT 374.830 110.890 375.110 113.150 ;
        RECT 375.710 110.890 375.990 113.150 ;
        RECT 376.590 110.890 376.870 113.150 ;
        RECT 377.470 110.890 377.750 113.150 ;
        RECT 378.350 110.890 378.630 113.150 ;
        RECT 379.230 110.890 379.510 113.150 ;
        RECT 380.110 110.890 380.390 113.150 ;
        RECT 380.990 110.890 381.270 113.150 ;
        RECT 381.870 110.890 382.150 113.150 ;
        RECT 382.750 110.890 383.030 113.150 ;
        RECT 383.630 110.890 383.910 113.150 ;
        RECT 384.510 110.890 384.790 113.150 ;
        RECT 385.390 110.890 385.670 113.150 ;
        RECT 386.270 110.890 386.550 113.150 ;
        RECT 387.150 110.890 387.430 113.150 ;
        RECT 388.030 110.890 388.310 113.150 ;
        RECT 388.910 110.890 389.190 113.150 ;
        RECT 389.790 110.890 390.070 113.150 ;
        RECT 390.670 110.890 390.950 113.150 ;
        RECT 391.550 110.890 391.830 113.150 ;
        RECT 392.430 110.890 392.710 113.150 ;
        RECT 393.310 110.890 393.590 113.150 ;
        RECT 394.190 110.890 394.470 113.150 ;
        RECT 395.070 110.890 395.350 113.150 ;
        RECT 395.950 110.890 396.230 113.150 ;
        RECT 396.830 110.890 397.110 113.150 ;
        RECT 397.710 110.890 397.990 113.150 ;
        RECT 398.590 110.890 398.870 113.150 ;
        RECT 399.470 110.890 399.750 113.150 ;
        RECT 400.350 110.890 400.630 113.150 ;
        RECT 401.230 110.890 401.510 113.150 ;
        RECT 402.110 110.890 402.390 113.150 ;
        RECT 402.990 110.890 403.270 113.150 ;
        RECT 403.870 110.890 404.150 113.150 ;
        RECT 404.750 110.890 405.030 113.150 ;
        RECT 405.630 110.890 405.910 113.150 ;
        RECT 406.350 112.520 406.640 113.990 ;
        RECT 406.350 111.520 406.645 112.520 ;
        RECT 406.350 110.700 406.640 111.520 ;
        RECT 364.415 110.410 366.825 110.700 ;
        RECT 402.475 110.410 406.640 110.700 ;
        RECT 364.415 110.050 364.705 110.410 ;
        RECT 406.350 110.050 406.640 110.410 ;
        RECT 364.415 109.760 406.640 110.050 ;
        RECT 444.015 109.865 444.305 118.795 ;
        RECT 446.815 118.245 449.885 118.575 ;
        RECT 444.715 115.055 444.945 118.055 ;
        RECT 445.595 115.055 445.825 118.055 ;
        RECT 446.475 115.055 446.705 118.055 ;
        RECT 444.700 113.055 444.960 115.055 ;
        RECT 445.580 113.055 445.840 115.055 ;
        RECT 446.460 113.055 446.720 115.055 ;
        RECT 444.715 110.055 444.945 113.055 ;
        RECT 445.595 110.055 445.825 113.055 ;
        RECT 446.475 110.055 446.705 113.055 ;
        RECT 447.340 110.055 447.600 118.055 ;
        RECT 448.235 115.055 448.465 118.055 ;
        RECT 448.220 113.055 448.480 115.055 ;
        RECT 448.235 110.055 448.465 113.055 ;
        RECT 449.100 110.055 449.360 118.055 ;
        RECT 449.995 115.055 450.225 118.055 ;
        RECT 450.875 115.055 451.105 118.055 ;
        RECT 451.755 115.055 451.985 118.055 ;
        RECT 449.980 113.055 450.240 115.055 ;
        RECT 450.860 113.055 451.120 115.055 ;
        RECT 451.740 113.055 452.000 115.055 ;
        RECT 449.995 110.055 450.225 113.055 ;
        RECT 450.875 110.055 451.105 113.055 ;
        RECT 451.755 110.055 451.985 113.055 ;
        RECT 452.395 109.865 452.685 118.795 ;
        RECT 444.015 109.575 446.365 109.865 ;
        RECT 450.335 109.575 452.685 109.865 ;
        RECT 444.015 109.315 444.305 109.575 ;
        RECT 452.395 109.315 452.685 109.575 ;
        RECT 444.015 109.025 452.685 109.315 ;
        RECT 457.835 118.795 466.505 119.085 ;
        RECT 457.835 109.865 458.125 118.795 ;
        RECT 460.635 118.245 463.705 118.575 ;
        RECT 458.535 115.055 458.765 118.055 ;
        RECT 459.415 115.055 459.645 118.055 ;
        RECT 460.295 115.055 460.525 118.055 ;
        RECT 458.520 113.055 458.780 115.055 ;
        RECT 459.400 113.055 459.660 115.055 ;
        RECT 460.280 113.055 460.540 115.055 ;
        RECT 458.535 110.055 458.765 113.055 ;
        RECT 459.415 110.055 459.645 113.055 ;
        RECT 460.295 110.055 460.525 113.055 ;
        RECT 461.160 110.055 461.420 118.055 ;
        RECT 462.055 115.055 462.285 118.055 ;
        RECT 462.040 113.055 462.300 115.055 ;
        RECT 462.055 110.055 462.285 113.055 ;
        RECT 462.935 110.055 463.195 118.055 ;
        RECT 463.815 115.055 464.045 118.055 ;
        RECT 464.695 115.055 464.925 118.055 ;
        RECT 465.575 115.055 465.805 118.055 ;
        RECT 463.800 113.055 464.060 115.055 ;
        RECT 464.680 113.055 464.940 115.055 ;
        RECT 465.560 113.055 465.820 115.055 ;
        RECT 463.815 110.055 464.045 113.055 ;
        RECT 464.695 110.055 464.925 113.055 ;
        RECT 465.575 110.055 465.805 113.055 ;
        RECT 466.215 109.865 466.505 118.795 ;
        RECT 457.835 109.575 460.185 109.865 ;
        RECT 464.155 109.575 466.505 109.865 ;
        RECT 457.835 109.315 458.125 109.575 ;
        RECT 466.215 109.315 466.505 109.575 ;
        RECT 457.835 109.025 466.505 109.315 ;
        RECT 467.575 118.795 486.265 119.085 ;
        RECT 467.575 109.865 467.865 118.795 ;
        RECT 468.275 115.055 468.505 118.055 ;
        RECT 469.555 115.055 469.785 118.055 ;
        RECT 470.835 115.055 471.065 118.055 ;
        RECT 468.260 113.055 468.520 115.055 ;
        RECT 469.540 113.055 469.800 115.055 ;
        RECT 470.820 113.055 471.080 115.055 ;
        RECT 468.275 110.055 468.505 113.055 ;
        RECT 469.555 110.055 469.785 113.055 ;
        RECT 470.835 110.055 471.065 113.055 ;
        RECT 473.805 110.055 474.065 118.055 ;
        RECT 476.805 115.055 477.035 118.055 ;
        RECT 476.790 113.055 477.050 115.055 ;
        RECT 476.805 110.055 477.035 113.055 ;
        RECT 479.775 110.055 480.035 118.055 ;
        RECT 482.775 115.055 483.005 118.055 ;
        RECT 484.055 115.055 484.285 118.055 ;
        RECT 485.335 115.055 485.565 118.055 ;
        RECT 482.760 113.055 483.020 115.055 ;
        RECT 484.040 113.055 484.300 115.055 ;
        RECT 485.320 113.055 485.580 115.055 ;
        RECT 482.775 110.055 483.005 113.055 ;
        RECT 484.055 110.055 484.285 113.055 ;
        RECT 485.335 110.055 485.565 113.055 ;
        RECT 485.975 109.865 486.265 118.795 ;
        RECT 467.575 109.575 470.605 109.865 ;
        RECT 467.575 109.315 467.865 109.575 ;
        RECT 471.120 109.535 482.720 109.865 ;
        RECT 483.235 109.575 486.265 109.865 ;
        RECT 485.975 109.315 486.265 109.575 ;
        RECT 467.575 109.025 486.265 109.315 ;
        RECT 487.050 118.795 495.720 119.085 ;
        RECT 334.115 108.675 363.945 108.965 ;
        RECT 184.740 106.165 185.030 106.725 ;
        RECT 191.410 106.165 191.740 106.755 ;
        RECT 198.120 106.165 198.410 106.725 ;
        RECT 184.740 105.895 186.275 106.165 ;
        RECT 186.555 105.895 196.595 106.165 ;
        RECT 196.875 105.895 198.410 106.165 ;
        RECT 199.820 106.615 204.885 106.905 ;
        RECT 208.425 106.615 213.490 106.905 ;
        RECT 199.820 106.325 200.110 106.615 ;
        RECT 213.200 106.325 213.490 106.615 ;
        RECT 199.820 106.035 213.490 106.325 ;
        RECT 184.740 104.305 185.030 105.895 ;
        RECT 185.425 104.705 185.685 105.705 ;
        RECT 185.855 104.705 186.115 105.705 ;
        RECT 186.285 104.705 186.545 105.705 ;
        RECT 186.700 104.705 186.960 105.705 ;
        RECT 187.145 104.705 187.405 105.705 ;
        RECT 187.560 104.705 187.820 105.705 ;
        RECT 188.005 104.705 188.265 105.705 ;
        RECT 188.420 104.705 188.680 105.705 ;
        RECT 188.865 104.705 189.125 105.705 ;
        RECT 189.280 104.705 189.540 105.705 ;
        RECT 189.725 104.705 189.985 105.705 ;
        RECT 190.155 104.705 190.415 105.705 ;
        RECT 190.585 104.705 190.845 105.705 ;
        RECT 191.030 104.705 191.290 105.705 ;
        RECT 191.445 104.705 191.705 105.705 ;
        RECT 191.890 104.705 192.150 105.705 ;
        RECT 192.305 104.705 192.565 105.705 ;
        RECT 192.750 104.705 193.010 105.705 ;
        RECT 193.165 104.705 193.425 105.705 ;
        RECT 193.610 104.705 193.870 105.705 ;
        RECT 194.025 104.705 194.285 105.705 ;
        RECT 194.470 104.705 194.730 105.705 ;
        RECT 194.885 104.705 195.145 105.705 ;
        RECT 195.330 104.705 195.590 105.705 ;
        RECT 195.745 104.705 196.005 105.705 ;
        RECT 196.190 104.705 196.450 105.705 ;
        RECT 196.605 104.705 196.865 105.705 ;
        RECT 197.035 104.705 197.295 105.705 ;
        RECT 197.465 104.705 197.725 105.705 ;
        RECT 198.120 104.305 198.410 105.895 ;
        RECT 218.010 105.155 219.320 107.260 ;
        RECT 220.020 105.155 221.330 107.260 ;
        RECT 222.030 106.710 223.340 107.260 ;
        RECT 224.040 106.710 225.350 107.260 ;
        RECT 226.050 106.710 227.360 107.260 ;
        RECT 228.060 106.710 229.370 107.260 ;
        RECT 222.030 105.710 229.370 106.710 ;
        RECT 222.030 105.155 223.340 105.710 ;
        RECT 224.040 105.155 225.350 105.710 ;
        RECT 226.050 105.155 227.360 105.710 ;
        RECT 228.060 105.155 229.370 105.710 ;
        RECT 230.070 106.710 231.380 107.260 ;
        RECT 232.080 106.710 233.390 107.260 ;
        RECT 234.090 106.710 235.400 107.260 ;
        RECT 236.100 106.710 237.410 107.260 ;
        RECT 238.110 106.710 239.420 107.260 ;
        RECT 230.070 105.710 239.420 106.710 ;
        RECT 230.070 105.155 231.380 105.710 ;
        RECT 232.080 105.155 233.390 105.710 ;
        RECT 234.090 105.155 235.400 105.710 ;
        RECT 236.100 105.155 237.410 105.710 ;
        RECT 238.110 105.155 239.420 105.710 ;
        RECT 240.120 106.710 241.430 107.260 ;
        RECT 242.130 106.710 243.440 107.260 ;
        RECT 240.120 105.710 243.440 106.710 ;
        RECT 240.120 105.155 241.430 105.710 ;
        RECT 242.130 105.155 243.440 105.710 ;
        RECT 244.140 106.710 245.450 107.260 ;
        RECT 246.150 106.710 247.460 107.260 ;
        RECT 244.140 105.710 247.460 106.710 ;
        RECT 244.140 105.155 245.450 105.710 ;
        RECT 246.150 105.155 247.460 105.710 ;
        RECT 248.160 106.710 249.470 107.260 ;
        RECT 250.170 106.710 251.480 107.260 ;
        RECT 248.160 105.710 251.480 106.710 ;
        RECT 248.160 105.155 249.470 105.710 ;
        RECT 250.170 105.155 251.480 105.710 ;
        RECT 252.180 106.710 253.490 107.260 ;
        RECT 254.190 106.710 255.500 107.260 ;
        RECT 252.180 105.710 255.500 106.710 ;
        RECT 252.180 105.155 253.490 105.710 ;
        RECT 254.190 105.155 255.500 105.710 ;
        RECT 256.200 106.710 257.510 107.260 ;
        RECT 258.210 106.710 259.520 107.260 ;
        RECT 256.200 105.710 259.520 106.710 ;
        RECT 256.200 105.155 257.510 105.710 ;
        RECT 258.210 105.155 259.520 105.710 ;
        RECT 260.220 106.710 261.530 107.260 ;
        RECT 262.230 106.710 263.540 107.260 ;
        RECT 260.220 105.710 263.540 106.710 ;
        RECT 260.220 105.155 261.530 105.710 ;
        RECT 262.230 105.155 263.540 105.710 ;
        RECT 264.240 106.710 265.550 107.260 ;
        RECT 266.250 106.710 267.560 107.260 ;
        RECT 264.240 105.710 267.560 106.710 ;
        RECT 264.240 105.155 265.550 105.710 ;
        RECT 266.250 105.155 267.560 105.710 ;
        RECT 268.260 106.710 269.570 107.260 ;
        RECT 270.270 106.710 271.580 107.260 ;
        RECT 268.260 105.710 271.580 106.710 ;
        RECT 268.260 105.155 269.570 105.710 ;
        RECT 270.270 105.155 271.580 105.710 ;
        RECT 272.280 106.710 273.590 107.260 ;
        RECT 274.290 106.710 275.600 107.260 ;
        RECT 272.280 105.710 275.600 106.710 ;
        RECT 272.280 105.155 273.590 105.710 ;
        RECT 274.290 105.155 275.600 105.710 ;
        RECT 276.300 106.710 277.610 107.260 ;
        RECT 278.310 106.710 279.620 107.260 ;
        RECT 276.300 105.710 279.620 106.710 ;
        RECT 276.300 105.155 277.610 105.710 ;
        RECT 278.310 105.155 279.620 105.710 ;
        RECT 280.320 106.710 281.630 107.260 ;
        RECT 282.330 106.710 283.640 107.260 ;
        RECT 280.320 105.710 283.640 106.710 ;
        RECT 280.320 105.155 281.630 105.710 ;
        RECT 282.330 105.155 283.640 105.710 ;
        RECT 284.340 105.155 285.650 107.260 ;
        RECT 286.350 105.155 287.660 107.260 ;
        RECT 288.360 105.155 289.670 107.260 ;
        RECT 310.855 105.855 333.725 106.145 ;
        RECT 184.740 104.015 198.410 104.305 ;
        RECT 310.855 105.020 311.145 105.855 ;
        RECT 311.955 105.320 315.765 105.610 ;
        RECT 315.475 105.020 315.765 105.320 ;
        RECT 328.815 105.320 332.625 105.610 ;
        RECT 328.815 105.020 329.105 105.320 ;
        RECT 333.435 105.020 333.725 105.855 ;
        RECT 310.855 104.730 315.025 105.020 ;
        RECT 315.475 104.730 329.105 105.020 ;
        RECT 329.555 104.730 333.725 105.020 ;
        RECT 184.740 102.485 198.410 102.775 ;
        RECT 184.740 100.895 185.030 102.485 ;
        RECT 185.425 101.085 185.685 102.085 ;
        RECT 185.855 101.085 186.115 102.085 ;
        RECT 186.285 101.085 186.545 102.085 ;
        RECT 186.700 101.085 186.960 102.085 ;
        RECT 187.145 101.085 187.405 102.085 ;
        RECT 187.560 101.085 187.820 102.085 ;
        RECT 188.005 101.085 188.265 102.085 ;
        RECT 188.420 101.085 188.680 102.085 ;
        RECT 188.865 101.085 189.125 102.085 ;
        RECT 189.280 101.085 189.540 102.085 ;
        RECT 189.725 101.085 189.985 102.085 ;
        RECT 190.155 101.085 190.415 102.085 ;
        RECT 190.585 101.085 190.845 102.085 ;
        RECT 191.030 101.085 191.290 102.085 ;
        RECT 191.445 101.085 191.705 102.085 ;
        RECT 191.890 101.085 192.150 102.085 ;
        RECT 192.305 101.085 192.565 102.085 ;
        RECT 192.750 101.085 193.010 102.085 ;
        RECT 193.165 101.085 193.425 102.085 ;
        RECT 193.610 101.085 193.870 102.085 ;
        RECT 194.025 101.085 194.285 102.085 ;
        RECT 194.470 101.085 194.730 102.085 ;
        RECT 194.885 101.085 195.145 102.085 ;
        RECT 195.330 101.085 195.590 102.085 ;
        RECT 195.745 101.085 196.005 102.085 ;
        RECT 196.190 101.085 196.450 102.085 ;
        RECT 196.605 101.085 196.865 102.085 ;
        RECT 197.035 101.085 197.295 102.085 ;
        RECT 197.465 101.085 197.725 102.085 ;
        RECT 198.120 100.895 198.410 102.485 ;
        RECT 310.855 102.090 311.145 104.730 ;
        RECT 311.590 102.280 311.870 104.540 ;
        RECT 312.470 102.280 312.750 104.540 ;
        RECT 313.350 102.280 313.630 104.540 ;
        RECT 314.230 102.280 314.510 104.540 ;
        RECT 315.110 102.280 315.390 104.540 ;
        RECT 315.990 102.280 316.270 104.540 ;
        RECT 316.870 102.280 317.150 104.540 ;
        RECT 317.750 102.280 318.030 104.540 ;
        RECT 318.630 102.280 318.910 104.540 ;
        RECT 319.510 102.280 319.790 104.540 ;
        RECT 320.390 102.280 320.670 104.540 ;
        RECT 321.270 102.280 321.550 104.540 ;
        RECT 322.150 102.280 322.430 104.540 ;
        RECT 323.030 102.280 323.310 104.540 ;
        RECT 323.910 102.280 324.190 104.540 ;
        RECT 324.790 102.280 325.070 104.540 ;
        RECT 325.670 102.280 325.950 104.540 ;
        RECT 326.550 102.280 326.830 104.540 ;
        RECT 327.430 102.280 327.710 104.540 ;
        RECT 328.310 102.280 328.590 104.540 ;
        RECT 329.190 102.280 329.470 104.540 ;
        RECT 330.070 102.280 330.350 104.540 ;
        RECT 330.950 102.280 331.230 104.540 ;
        RECT 331.830 102.280 332.110 104.540 ;
        RECT 332.710 102.280 332.990 104.540 ;
        RECT 333.435 102.090 333.725 104.730 ;
        RECT 310.855 101.800 315.025 102.090 ;
        RECT 315.475 101.800 329.105 102.090 ;
        RECT 329.555 101.800 333.725 102.090 ;
        RECT 184.740 100.625 186.275 100.895 ;
        RECT 186.555 100.625 196.595 100.895 ;
        RECT 196.875 100.625 198.410 100.895 ;
        RECT 184.740 100.065 185.030 100.625 ;
        RECT 191.410 100.035 191.740 100.625 ;
        RECT 198.120 100.065 198.410 100.625 ;
        RECT 199.820 100.465 213.490 100.755 ;
        RECT 199.820 100.175 200.110 100.465 ;
        RECT 213.200 100.175 213.490 100.465 ;
        RECT 191.410 99.705 197.105 100.035 ;
        RECT 184.740 99.120 185.030 99.680 ;
        RECT 191.410 99.120 191.740 99.705 ;
        RECT 196.775 99.555 197.105 99.705 ;
        RECT 199.820 99.885 204.885 100.175 ;
        RECT 208.425 99.885 213.490 100.175 ;
        RECT 196.775 99.275 197.735 99.555 ;
        RECT 198.120 99.120 198.410 99.680 ;
        RECT 184.740 98.850 189.715 99.120 ;
        RECT 189.995 98.850 193.155 99.120 ;
        RECT 193.435 98.850 198.410 99.120 ;
        RECT 184.740 97.290 185.030 98.850 ;
        RECT 185.425 97.660 185.685 98.660 ;
        RECT 185.855 97.660 186.115 98.660 ;
        RECT 186.285 97.660 186.545 98.660 ;
        RECT 186.715 97.660 186.975 98.660 ;
        RECT 187.145 97.660 187.405 98.660 ;
        RECT 187.575 97.660 187.835 98.660 ;
        RECT 188.005 97.660 188.265 98.660 ;
        RECT 188.435 97.660 188.695 98.660 ;
        RECT 188.865 97.660 189.125 98.660 ;
        RECT 189.295 97.660 189.555 98.660 ;
        RECT 189.725 97.660 189.985 98.660 ;
        RECT 190.155 97.660 190.415 98.660 ;
        RECT 190.585 97.660 190.845 98.660 ;
        RECT 191.030 97.660 191.290 98.660 ;
        RECT 191.445 97.660 191.705 98.660 ;
        RECT 191.890 97.660 192.150 98.660 ;
        RECT 192.305 97.660 192.565 98.660 ;
        RECT 192.750 97.660 193.010 98.660 ;
        RECT 193.165 97.660 193.425 98.660 ;
        RECT 193.595 97.660 193.855 98.660 ;
        RECT 194.025 97.660 194.285 98.660 ;
        RECT 194.455 97.660 194.715 98.660 ;
        RECT 194.885 97.660 195.145 98.660 ;
        RECT 195.315 97.660 195.575 98.660 ;
        RECT 195.745 97.660 196.005 98.660 ;
        RECT 196.175 97.660 196.435 98.660 ;
        RECT 196.605 97.660 196.865 98.660 ;
        RECT 197.035 97.660 197.295 98.660 ;
        RECT 197.480 97.660 197.710 98.850 ;
        RECT 198.120 97.290 198.410 98.850 ;
        RECT 199.820 97.375 200.110 99.885 ;
        RECT 200.505 98.845 200.765 99.695 ;
        RECT 200.935 98.845 201.195 99.695 ;
        RECT 201.365 98.845 201.625 99.695 ;
        RECT 201.795 98.845 202.055 99.695 ;
        RECT 202.225 98.845 202.485 99.695 ;
        RECT 202.655 98.845 202.915 99.695 ;
        RECT 203.085 98.845 203.345 99.695 ;
        RECT 203.515 98.845 203.775 99.695 ;
        RECT 203.945 98.845 204.205 99.695 ;
        RECT 204.375 98.845 204.635 99.695 ;
        RECT 200.520 98.695 200.750 98.845 ;
        RECT 200.950 98.695 201.180 98.845 ;
        RECT 201.380 98.695 201.610 98.845 ;
        RECT 201.810 98.695 202.040 98.845 ;
        RECT 202.240 98.695 202.470 98.845 ;
        RECT 202.670 98.695 202.900 98.845 ;
        RECT 203.100 98.695 203.330 98.845 ;
        RECT 203.530 98.695 203.760 98.845 ;
        RECT 203.960 98.695 204.190 98.845 ;
        RECT 204.390 98.695 204.620 98.845 ;
        RECT 204.820 98.695 205.080 99.695 ;
        RECT 205.250 98.695 205.510 99.695 ;
        RECT 205.680 98.695 205.940 99.695 ;
        RECT 206.110 98.695 206.370 99.695 ;
        RECT 206.540 98.695 206.800 99.695 ;
        RECT 206.970 98.695 207.230 99.695 ;
        RECT 207.400 98.695 207.660 99.695 ;
        RECT 207.830 98.695 208.090 99.695 ;
        RECT 208.260 98.695 208.520 99.695 ;
        RECT 208.675 98.845 208.935 99.695 ;
        RECT 209.105 98.845 209.365 99.695 ;
        RECT 209.535 98.845 209.795 99.695 ;
        RECT 209.965 98.845 210.225 99.695 ;
        RECT 210.395 98.845 210.655 99.695 ;
        RECT 210.825 98.845 211.085 99.695 ;
        RECT 211.255 98.845 211.515 99.695 ;
        RECT 211.685 98.845 211.945 99.695 ;
        RECT 212.115 98.845 212.375 99.695 ;
        RECT 212.545 98.845 212.805 99.695 ;
        RECT 208.690 98.695 208.920 98.845 ;
        RECT 209.120 98.695 209.350 98.845 ;
        RECT 209.550 98.695 209.780 98.845 ;
        RECT 209.980 98.695 210.210 98.845 ;
        RECT 210.410 98.695 210.640 98.845 ;
        RECT 210.840 98.695 211.070 98.845 ;
        RECT 211.270 98.695 211.500 98.845 ;
        RECT 211.700 98.695 211.930 98.845 ;
        RECT 212.130 98.695 212.360 98.845 ;
        RECT 212.560 98.695 212.790 98.845 ;
        RECT 200.310 98.225 211.675 98.505 ;
        RECT 213.200 97.375 213.490 99.885 ;
        RECT 218.010 99.530 219.320 101.635 ;
        RECT 220.020 99.530 221.330 101.635 ;
        RECT 222.030 101.085 223.340 101.635 ;
        RECT 224.040 101.085 225.350 101.635 ;
        RECT 226.050 101.085 227.360 101.635 ;
        RECT 228.060 101.085 229.370 101.635 ;
        RECT 222.030 100.085 229.370 101.085 ;
        RECT 222.030 99.530 223.340 100.085 ;
        RECT 224.040 99.530 225.350 100.085 ;
        RECT 226.050 99.530 227.360 100.085 ;
        RECT 228.060 99.530 229.370 100.085 ;
        RECT 230.070 101.085 231.380 101.635 ;
        RECT 232.080 101.085 233.390 101.635 ;
        RECT 234.090 101.085 235.400 101.635 ;
        RECT 236.100 101.085 237.410 101.635 ;
        RECT 238.110 101.085 239.420 101.635 ;
        RECT 230.070 100.085 239.420 101.085 ;
        RECT 230.070 99.530 231.380 100.085 ;
        RECT 232.080 99.530 233.390 100.085 ;
        RECT 234.090 99.530 235.400 100.085 ;
        RECT 236.100 99.530 237.410 100.085 ;
        RECT 238.110 99.530 239.420 100.085 ;
        RECT 240.120 101.085 241.430 101.635 ;
        RECT 242.130 101.085 243.440 101.635 ;
        RECT 240.120 100.085 243.440 101.085 ;
        RECT 240.120 99.530 241.430 100.085 ;
        RECT 242.130 99.530 243.440 100.085 ;
        RECT 244.140 101.085 245.450 101.635 ;
        RECT 246.150 101.085 247.460 101.635 ;
        RECT 244.140 100.085 247.460 101.085 ;
        RECT 244.140 99.530 245.450 100.085 ;
        RECT 246.150 99.530 247.460 100.085 ;
        RECT 248.160 101.085 249.470 101.635 ;
        RECT 250.170 101.085 251.480 101.635 ;
        RECT 248.160 100.085 251.480 101.085 ;
        RECT 248.160 99.530 249.470 100.085 ;
        RECT 250.170 99.530 251.480 100.085 ;
        RECT 252.180 101.085 253.490 101.635 ;
        RECT 254.190 101.085 255.500 101.635 ;
        RECT 252.180 100.085 255.500 101.085 ;
        RECT 252.180 99.530 253.490 100.085 ;
        RECT 254.190 99.530 255.500 100.085 ;
        RECT 256.200 101.085 257.510 101.635 ;
        RECT 258.210 101.085 259.520 101.635 ;
        RECT 256.200 100.085 259.520 101.085 ;
        RECT 256.200 99.530 257.510 100.085 ;
        RECT 258.210 99.530 259.520 100.085 ;
        RECT 260.220 101.085 261.530 101.635 ;
        RECT 262.230 101.085 263.540 101.635 ;
        RECT 260.220 100.085 263.540 101.085 ;
        RECT 260.220 99.530 261.530 100.085 ;
        RECT 262.230 99.530 263.540 100.085 ;
        RECT 264.240 101.085 265.550 101.635 ;
        RECT 266.250 101.085 267.560 101.635 ;
        RECT 264.240 100.085 267.560 101.085 ;
        RECT 264.240 99.530 265.550 100.085 ;
        RECT 266.250 99.530 267.560 100.085 ;
        RECT 268.260 101.085 269.570 101.635 ;
        RECT 270.270 101.085 271.580 101.635 ;
        RECT 268.260 100.085 271.580 101.085 ;
        RECT 268.260 99.530 269.570 100.085 ;
        RECT 270.270 99.530 271.580 100.085 ;
        RECT 272.280 101.085 273.590 101.635 ;
        RECT 274.290 101.085 275.600 101.635 ;
        RECT 272.280 100.085 275.600 101.085 ;
        RECT 272.280 99.530 273.590 100.085 ;
        RECT 274.290 99.530 275.600 100.085 ;
        RECT 276.300 101.085 277.610 101.635 ;
        RECT 278.310 101.085 279.620 101.635 ;
        RECT 276.300 100.085 279.620 101.085 ;
        RECT 276.300 99.530 277.610 100.085 ;
        RECT 278.310 99.530 279.620 100.085 ;
        RECT 280.320 101.085 281.630 101.635 ;
        RECT 282.330 101.085 283.640 101.635 ;
        RECT 280.320 100.085 283.640 101.085 ;
        RECT 280.320 99.530 281.630 100.085 ;
        RECT 282.330 99.530 283.640 100.085 ;
        RECT 284.340 99.530 285.650 101.635 ;
        RECT 286.350 99.530 287.660 101.635 ;
        RECT 288.360 99.530 289.670 101.635 ;
        RECT 310.855 100.970 311.145 101.800 ;
        RECT 315.475 101.500 315.765 101.800 ;
        RECT 311.955 101.210 315.765 101.500 ;
        RECT 328.815 101.500 329.105 101.800 ;
        RECT 328.815 101.210 332.625 101.500 ;
        RECT 333.435 100.970 333.725 101.800 ;
        RECT 310.855 100.680 333.725 100.970 ;
        RECT 334.115 98.695 334.405 108.675 ;
        RECT 340.455 108.105 347.045 108.435 ;
        RECT 351.070 108.395 357.660 108.435 ;
        RECT 351.015 108.105 357.660 108.395 ;
        RECT 334.810 98.885 335.090 107.915 ;
        RECT 335.690 98.885 335.970 107.915 ;
        RECT 336.570 98.885 336.850 107.915 ;
        RECT 337.450 98.885 337.730 107.915 ;
        RECT 338.330 98.885 338.610 107.915 ;
        RECT 339.210 98.885 339.490 107.915 ;
        RECT 340.090 98.885 340.370 107.915 ;
        RECT 340.970 98.885 341.250 107.915 ;
        RECT 341.850 98.885 342.130 107.915 ;
        RECT 342.730 98.885 343.010 107.915 ;
        RECT 343.610 98.885 343.890 107.915 ;
        RECT 344.490 98.885 344.770 107.915 ;
        RECT 345.370 98.885 345.650 107.915 ;
        RECT 346.250 98.885 346.530 107.915 ;
        RECT 347.130 98.885 347.410 107.915 ;
        RECT 348.010 98.695 348.290 107.915 ;
        RECT 348.890 98.695 349.170 107.915 ;
        RECT 349.770 98.695 350.050 107.915 ;
        RECT 350.650 98.885 350.930 107.915 ;
        RECT 351.530 98.885 351.810 107.915 ;
        RECT 352.410 98.885 352.690 107.915 ;
        RECT 353.290 98.885 353.570 107.915 ;
        RECT 354.170 98.885 354.450 107.915 ;
        RECT 355.050 98.885 355.330 107.915 ;
        RECT 355.930 98.885 356.210 107.915 ;
        RECT 356.810 98.885 357.090 107.915 ;
        RECT 357.690 98.885 357.970 107.915 ;
        RECT 358.570 98.885 358.850 107.915 ;
        RECT 359.450 98.885 359.730 107.915 ;
        RECT 360.330 98.885 360.610 107.915 ;
        RECT 361.210 98.885 361.490 107.915 ;
        RECT 362.090 98.885 362.370 107.915 ;
        RECT 362.970 98.885 363.250 107.915 ;
        RECT 363.655 98.695 363.945 108.675 ;
        RECT 184.740 97.000 198.410 97.290 ;
        RECT 184.740 95.440 185.030 97.000 ;
        RECT 185.425 95.630 185.685 96.630 ;
        RECT 185.855 95.630 186.115 96.630 ;
        RECT 186.285 95.630 186.545 96.630 ;
        RECT 186.715 95.630 186.975 96.630 ;
        RECT 187.145 95.630 187.405 96.630 ;
        RECT 187.575 95.630 187.835 96.630 ;
        RECT 188.005 95.630 188.265 96.630 ;
        RECT 188.435 95.630 188.695 96.630 ;
        RECT 188.865 95.630 189.125 96.630 ;
        RECT 189.295 95.630 189.555 96.630 ;
        RECT 189.725 95.630 189.985 96.630 ;
        RECT 190.155 95.630 190.415 96.630 ;
        RECT 190.585 95.630 190.845 96.630 ;
        RECT 191.030 95.630 191.290 96.630 ;
        RECT 191.445 95.630 191.705 96.630 ;
        RECT 191.890 95.630 192.150 96.630 ;
        RECT 192.305 95.630 192.565 96.630 ;
        RECT 192.750 95.630 193.010 96.630 ;
        RECT 193.165 95.630 193.425 96.630 ;
        RECT 193.595 95.630 193.855 96.630 ;
        RECT 194.025 95.630 194.285 96.630 ;
        RECT 194.455 95.630 194.715 96.630 ;
        RECT 194.885 95.630 195.145 96.630 ;
        RECT 195.315 95.630 195.575 96.630 ;
        RECT 195.745 95.630 196.005 96.630 ;
        RECT 196.175 95.630 196.435 96.630 ;
        RECT 196.605 95.630 196.865 96.630 ;
        RECT 197.035 95.630 197.295 96.630 ;
        RECT 197.480 95.440 197.710 96.630 ;
        RECT 198.120 95.440 198.410 97.000 ;
        RECT 217.110 96.645 217.400 98.645 ;
        RECT 290.280 96.645 290.570 98.645 ;
        RECT 334.115 98.405 340.005 98.695 ;
        RECT 347.495 98.405 350.565 98.695 ;
        RECT 358.055 98.405 363.945 98.695 ;
        RECT 334.115 98.125 334.405 98.405 ;
        RECT 363.655 98.125 363.945 98.405 ;
        RECT 334.115 97.835 363.945 98.125 ;
        RECT 364.455 108.675 406.605 108.965 ;
        RECT 364.455 98.695 364.745 108.675 ;
        RECT 367.275 108.105 402.025 108.435 ;
        RECT 365.150 98.885 365.430 107.915 ;
        RECT 366.030 98.885 366.310 107.915 ;
        RECT 366.910 98.885 367.190 107.915 ;
        RECT 367.790 98.885 368.070 107.915 ;
        RECT 368.670 98.885 368.950 107.915 ;
        RECT 369.550 98.885 369.830 107.915 ;
        RECT 370.430 98.885 370.710 107.915 ;
        RECT 371.310 98.885 371.590 107.915 ;
        RECT 372.190 98.885 372.470 107.915 ;
        RECT 373.070 98.885 373.350 107.915 ;
        RECT 373.950 98.885 374.230 107.915 ;
        RECT 374.830 98.885 375.110 107.915 ;
        RECT 375.710 98.885 375.990 107.915 ;
        RECT 376.590 98.885 376.870 107.915 ;
        RECT 377.470 98.885 377.750 107.915 ;
        RECT 378.350 98.885 378.630 107.915 ;
        RECT 379.230 98.885 379.510 107.915 ;
        RECT 380.110 98.885 380.390 107.915 ;
        RECT 380.990 98.885 381.270 107.915 ;
        RECT 381.870 98.885 382.150 107.915 ;
        RECT 382.750 98.885 383.030 107.915 ;
        RECT 383.630 98.885 383.910 107.915 ;
        RECT 384.510 98.885 384.790 107.915 ;
        RECT 385.390 98.885 385.670 107.915 ;
        RECT 386.270 98.885 386.550 107.915 ;
        RECT 387.150 98.885 387.430 107.915 ;
        RECT 388.030 98.885 388.310 107.915 ;
        RECT 388.910 98.885 389.190 107.915 ;
        RECT 389.790 98.885 390.070 107.915 ;
        RECT 390.670 98.885 390.950 107.915 ;
        RECT 391.550 98.885 391.830 107.915 ;
        RECT 392.430 98.885 392.710 107.915 ;
        RECT 393.310 98.885 393.590 107.915 ;
        RECT 394.190 98.885 394.470 107.915 ;
        RECT 395.070 98.885 395.350 107.915 ;
        RECT 395.950 98.885 396.230 107.915 ;
        RECT 396.830 98.885 397.110 107.915 ;
        RECT 397.710 98.885 397.990 107.915 ;
        RECT 398.590 98.885 398.870 107.915 ;
        RECT 399.470 98.885 399.750 107.915 ;
        RECT 400.350 98.885 400.630 107.915 ;
        RECT 401.230 98.885 401.510 107.915 ;
        RECT 402.110 98.885 402.390 107.915 ;
        RECT 402.990 98.885 403.270 107.915 ;
        RECT 403.870 98.885 404.150 107.915 ;
        RECT 404.750 98.885 405.030 107.915 ;
        RECT 405.630 98.885 405.910 107.915 ;
        RECT 406.315 98.695 406.605 108.675 ;
        RECT 487.050 108.835 487.340 118.795 ;
        RECT 489.850 118.245 492.920 118.575 ;
        RECT 487.750 115.055 487.980 118.055 ;
        RECT 488.630 115.055 488.860 118.055 ;
        RECT 489.510 115.055 489.740 118.055 ;
        RECT 487.735 113.055 487.995 115.055 ;
        RECT 488.615 113.055 488.875 115.055 ;
        RECT 489.495 113.055 489.755 115.055 ;
        RECT 487.750 109.025 487.980 113.055 ;
        RECT 488.630 109.025 488.860 113.055 ;
        RECT 489.510 109.025 489.740 113.055 ;
        RECT 490.375 109.025 490.635 118.055 ;
        RECT 491.270 115.055 491.500 118.055 ;
        RECT 491.255 113.055 491.515 115.055 ;
        RECT 491.270 109.025 491.500 113.055 ;
        RECT 492.135 109.025 492.395 118.055 ;
        RECT 493.030 115.055 493.260 118.055 ;
        RECT 493.910 115.055 494.140 118.055 ;
        RECT 494.790 115.055 495.020 118.055 ;
        RECT 493.015 113.055 493.275 115.055 ;
        RECT 493.895 113.055 494.155 115.055 ;
        RECT 494.775 113.055 495.035 115.055 ;
        RECT 493.030 109.025 493.260 113.055 ;
        RECT 493.910 109.025 494.140 113.055 ;
        RECT 494.790 109.025 495.020 113.055 ;
        RECT 495.430 108.835 495.720 118.795 ;
        RECT 496.780 118.795 505.450 119.085 ;
        RECT 496.780 109.865 497.070 118.795 ;
        RECT 497.480 115.055 497.710 118.055 ;
        RECT 498.360 115.055 498.590 118.055 ;
        RECT 499.240 115.055 499.470 118.055 ;
        RECT 497.465 113.055 497.725 115.055 ;
        RECT 498.345 113.055 498.605 115.055 ;
        RECT 499.225 113.055 499.485 115.055 ;
        RECT 497.480 110.055 497.710 113.055 ;
        RECT 498.360 110.055 498.590 113.055 ;
        RECT 499.240 110.055 499.470 113.055 ;
        RECT 500.105 110.055 500.365 118.055 ;
        RECT 501.000 115.055 501.230 118.055 ;
        RECT 500.985 113.055 501.245 115.055 ;
        RECT 501.000 110.055 501.230 113.055 ;
        RECT 501.865 110.055 502.125 118.055 ;
        RECT 502.760 115.055 502.990 118.055 ;
        RECT 503.640 115.055 503.870 118.055 ;
        RECT 504.520 115.055 504.750 118.055 ;
        RECT 502.745 113.055 503.005 115.055 ;
        RECT 503.625 113.055 503.885 115.055 ;
        RECT 504.505 113.055 504.765 115.055 ;
        RECT 502.760 110.055 502.990 113.055 ;
        RECT 503.640 110.055 503.870 113.055 ;
        RECT 504.520 110.055 504.750 113.055 ;
        RECT 505.160 109.865 505.450 118.795 ;
        RECT 496.780 109.575 499.130 109.865 ;
        RECT 496.780 109.315 497.070 109.575 ;
        RECT 499.580 109.535 502.650 109.865 ;
        RECT 503.100 109.575 505.450 109.865 ;
        RECT 505.160 109.315 505.450 109.575 ;
        RECT 496.780 109.025 505.450 109.315 ;
        RECT 487.050 108.545 489.400 108.835 ;
        RECT 493.370 108.545 495.720 108.835 ;
        RECT 487.050 108.285 487.340 108.545 ;
        RECT 495.430 108.285 495.720 108.545 ;
        RECT 487.050 107.995 495.720 108.285 ;
        RECT 364.455 98.405 366.825 98.695 ;
        RECT 402.475 98.405 406.605 98.695 ;
        RECT 364.455 98.125 364.745 98.405 ;
        RECT 406.315 98.125 406.605 98.405 ;
        RECT 364.455 97.835 406.605 98.125 ;
        RECT 487.050 105.530 495.720 105.820 ;
        RECT 472.625 97.085 481.215 97.375 ;
        RECT 472.625 96.825 472.915 97.085 ;
        RECT 480.925 96.825 481.215 97.085 ;
        RECT 184.740 95.170 189.715 95.440 ;
        RECT 189.995 95.170 193.155 95.440 ;
        RECT 193.435 95.170 198.410 95.440 ;
        RECT 184.740 94.610 185.030 95.170 ;
        RECT 191.410 94.585 191.740 95.170 ;
        RECT 198.120 94.610 198.410 95.170 ;
        RECT 185.490 94.255 191.740 94.585 ;
        RECT 184.740 93.665 185.030 94.225 ;
        RECT 191.410 93.665 191.740 94.255 ;
        RECT 199.820 94.405 200.110 96.615 ;
        RECT 200.310 95.785 211.675 96.065 ;
        RECT 200.520 95.445 200.750 95.595 ;
        RECT 200.950 95.445 201.180 95.595 ;
        RECT 200.505 94.595 200.765 95.445 ;
        RECT 200.935 94.595 201.195 95.445 ;
        RECT 201.365 94.595 201.625 95.595 ;
        RECT 201.795 94.595 202.055 95.595 ;
        RECT 202.240 94.595 202.500 95.595 ;
        RECT 202.670 94.595 202.930 95.595 ;
        RECT 203.100 94.595 203.360 95.595 ;
        RECT 203.530 94.595 203.790 95.595 ;
        RECT 203.960 94.595 204.220 95.595 ;
        RECT 204.390 94.595 204.650 95.595 ;
        RECT 204.820 94.595 205.080 95.595 ;
        RECT 205.250 94.595 205.510 95.595 ;
        RECT 205.680 94.595 205.940 95.595 ;
        RECT 206.110 94.595 206.370 95.595 ;
        RECT 206.540 94.595 206.800 95.595 ;
        RECT 206.970 94.595 207.230 95.595 ;
        RECT 207.400 94.595 207.660 95.595 ;
        RECT 207.830 94.595 208.090 95.595 ;
        RECT 208.260 94.595 208.520 95.595 ;
        RECT 208.690 94.595 208.950 95.595 ;
        RECT 209.120 94.595 209.380 95.595 ;
        RECT 209.550 94.595 209.810 95.595 ;
        RECT 209.980 94.595 210.240 95.595 ;
        RECT 210.410 94.595 210.670 95.595 ;
        RECT 210.840 94.595 211.100 95.595 ;
        RECT 211.270 94.595 211.530 95.595 ;
        RECT 211.700 94.595 211.960 95.595 ;
        RECT 212.130 95.445 212.360 95.595 ;
        RECT 212.560 95.445 212.790 95.595 ;
        RECT 212.115 94.595 212.375 95.445 ;
        RECT 212.545 94.595 212.805 95.445 ;
        RECT 213.200 94.405 213.490 96.615 ;
        RECT 198.120 93.665 198.410 94.225 ;
        RECT 184.740 93.395 186.275 93.665 ;
        RECT 186.555 93.395 196.595 93.665 ;
        RECT 196.875 93.395 198.410 93.665 ;
        RECT 184.740 91.805 185.030 93.395 ;
        RECT 185.425 92.205 185.685 93.205 ;
        RECT 185.855 92.205 186.115 93.205 ;
        RECT 186.285 92.205 186.545 93.205 ;
        RECT 186.700 92.205 186.960 93.205 ;
        RECT 187.145 92.205 187.405 93.205 ;
        RECT 187.560 92.205 187.820 93.205 ;
        RECT 188.005 92.205 188.265 93.205 ;
        RECT 188.420 92.205 188.680 93.205 ;
        RECT 188.865 92.205 189.125 93.205 ;
        RECT 189.280 92.205 189.540 93.205 ;
        RECT 189.725 92.205 189.985 93.205 ;
        RECT 190.155 92.205 190.415 93.205 ;
        RECT 190.585 92.205 190.845 93.205 ;
        RECT 191.030 92.205 191.290 93.205 ;
        RECT 191.445 92.205 191.705 93.205 ;
        RECT 191.890 92.205 192.150 93.205 ;
        RECT 192.305 92.205 192.565 93.205 ;
        RECT 192.750 92.205 193.010 93.205 ;
        RECT 193.165 92.205 193.425 93.205 ;
        RECT 193.610 92.205 193.870 93.205 ;
        RECT 194.025 92.205 194.285 93.205 ;
        RECT 194.470 92.205 194.730 93.205 ;
        RECT 194.885 92.205 195.145 93.205 ;
        RECT 195.330 92.205 195.590 93.205 ;
        RECT 195.745 92.205 196.005 93.205 ;
        RECT 196.190 92.205 196.450 93.205 ;
        RECT 196.605 92.205 196.865 93.205 ;
        RECT 197.035 92.205 197.295 93.205 ;
        RECT 197.465 92.205 197.725 93.205 ;
        RECT 198.120 91.805 198.410 93.395 ;
        RECT 199.820 94.115 201.360 94.405 ;
        RECT 211.950 94.115 213.490 94.405 ;
        RECT 199.820 93.665 200.110 94.115 ;
        RECT 213.200 93.665 213.490 94.115 ;
        RECT 199.820 93.375 213.490 93.665 ;
        RECT 334.115 96.310 363.945 96.600 ;
        RECT 334.115 96.030 334.405 96.310 ;
        RECT 363.655 96.030 363.945 96.310 ;
        RECT 334.115 95.740 338.245 96.030 ;
        RECT 359.815 95.740 363.945 96.030 ;
        RECT 184.740 91.515 198.410 91.805 ;
        RECT 218.010 89.935 219.320 92.040 ;
        RECT 220.020 89.935 221.330 92.040 ;
        RECT 222.030 91.490 223.340 92.040 ;
        RECT 224.040 91.490 225.350 92.040 ;
        RECT 226.050 91.490 227.360 92.040 ;
        RECT 228.060 91.490 229.370 92.040 ;
        RECT 230.070 91.490 231.380 92.040 ;
        RECT 232.080 91.490 233.390 92.040 ;
        RECT 234.090 91.490 235.400 92.040 ;
        RECT 236.100 91.490 237.410 92.040 ;
        RECT 222.030 90.490 237.410 91.490 ;
        RECT 222.030 89.935 223.340 90.490 ;
        RECT 224.040 89.935 225.350 90.490 ;
        RECT 226.050 89.935 227.360 90.490 ;
        RECT 228.060 89.935 229.370 90.490 ;
        RECT 230.070 89.935 231.380 90.490 ;
        RECT 232.080 89.935 233.390 90.490 ;
        RECT 234.090 89.935 235.400 90.490 ;
        RECT 236.100 89.935 237.410 90.490 ;
        RECT 238.110 91.490 239.420 92.040 ;
        RECT 240.120 91.490 241.430 92.040 ;
        RECT 238.110 90.490 241.430 91.490 ;
        RECT 238.110 89.935 239.420 90.490 ;
        RECT 240.120 89.935 241.430 90.490 ;
        RECT 242.130 91.490 243.440 92.040 ;
        RECT 244.140 91.490 245.450 92.040 ;
        RECT 242.130 90.490 245.450 91.490 ;
        RECT 242.130 89.935 243.440 90.490 ;
        RECT 244.140 89.935 245.450 90.490 ;
        RECT 246.150 91.490 247.460 92.040 ;
        RECT 248.160 91.490 249.470 92.040 ;
        RECT 246.150 90.490 249.470 91.490 ;
        RECT 246.150 89.935 247.460 90.490 ;
        RECT 248.160 89.935 249.470 90.490 ;
        RECT 250.170 91.490 251.480 92.040 ;
        RECT 252.180 91.490 253.490 92.040 ;
        RECT 250.170 90.490 253.490 91.490 ;
        RECT 250.170 89.935 251.480 90.490 ;
        RECT 252.180 89.935 253.490 90.490 ;
        RECT 254.190 91.490 255.500 92.040 ;
        RECT 256.200 91.490 257.510 92.040 ;
        RECT 254.190 90.490 257.510 91.490 ;
        RECT 254.190 89.935 255.500 90.490 ;
        RECT 256.200 89.935 257.510 90.490 ;
        RECT 258.210 91.490 259.520 92.040 ;
        RECT 260.220 91.490 261.530 92.040 ;
        RECT 258.210 90.490 261.530 91.490 ;
        RECT 258.210 89.935 259.520 90.490 ;
        RECT 260.220 89.935 261.530 90.490 ;
        RECT 262.230 91.490 263.540 92.040 ;
        RECT 264.240 91.490 265.550 92.040 ;
        RECT 262.230 90.490 265.550 91.490 ;
        RECT 262.230 89.935 263.540 90.490 ;
        RECT 264.240 89.935 265.550 90.490 ;
        RECT 266.250 91.490 267.560 92.040 ;
        RECT 268.260 91.490 269.570 92.040 ;
        RECT 266.250 90.490 269.570 91.490 ;
        RECT 266.250 89.935 267.560 90.490 ;
        RECT 268.260 89.935 269.570 90.490 ;
        RECT 270.270 91.490 271.580 92.040 ;
        RECT 272.280 91.490 273.590 92.040 ;
        RECT 270.270 90.490 273.590 91.490 ;
        RECT 270.270 89.935 271.580 90.490 ;
        RECT 272.280 89.935 273.590 90.490 ;
        RECT 274.290 91.490 275.600 92.040 ;
        RECT 276.300 91.490 277.610 92.040 ;
        RECT 274.290 90.490 277.610 91.490 ;
        RECT 274.290 89.935 275.600 90.490 ;
        RECT 276.300 89.935 277.610 90.490 ;
        RECT 278.310 91.490 279.620 92.040 ;
        RECT 280.320 91.490 281.630 92.040 ;
        RECT 278.310 90.490 281.630 91.490 ;
        RECT 278.310 89.935 279.620 90.490 ;
        RECT 280.320 89.935 281.630 90.490 ;
        RECT 282.330 91.490 283.640 92.040 ;
        RECT 284.340 91.490 285.650 92.040 ;
        RECT 282.330 90.490 285.650 91.490 ;
        RECT 282.330 89.935 283.640 90.490 ;
        RECT 284.340 89.935 285.650 90.490 ;
        RECT 286.350 89.935 287.660 92.040 ;
        RECT 288.360 89.935 289.670 92.040 ;
        RECT 334.115 85.760 334.405 95.740 ;
        RECT 334.810 86.520 335.090 95.550 ;
        RECT 335.690 86.520 335.970 95.550 ;
        RECT 336.570 86.520 336.850 95.550 ;
        RECT 337.450 86.520 337.730 95.550 ;
        RECT 338.330 86.520 338.610 95.550 ;
        RECT 339.210 86.520 339.490 95.550 ;
        RECT 340.090 86.520 340.370 95.550 ;
        RECT 340.970 86.520 341.250 95.550 ;
        RECT 341.850 86.520 342.130 95.550 ;
        RECT 342.730 86.520 343.010 95.550 ;
        RECT 343.610 86.520 343.890 95.550 ;
        RECT 344.490 86.520 344.770 95.550 ;
        RECT 345.370 86.520 345.650 95.550 ;
        RECT 346.250 86.520 346.530 95.550 ;
        RECT 347.130 86.520 347.410 95.550 ;
        RECT 348.010 86.520 348.290 95.550 ;
        RECT 348.890 86.520 349.170 95.550 ;
        RECT 349.770 86.520 350.050 95.550 ;
        RECT 350.650 86.520 350.930 95.550 ;
        RECT 351.530 86.520 351.810 95.550 ;
        RECT 352.410 86.520 352.690 95.550 ;
        RECT 353.290 86.520 353.570 95.550 ;
        RECT 354.170 86.520 354.450 95.550 ;
        RECT 355.050 86.520 355.330 95.550 ;
        RECT 355.930 86.520 356.210 95.550 ;
        RECT 356.810 86.520 357.090 95.550 ;
        RECT 357.690 86.520 357.970 95.550 ;
        RECT 358.570 86.520 358.850 95.550 ;
        RECT 359.450 86.520 359.730 95.550 ;
        RECT 360.330 86.520 360.610 95.550 ;
        RECT 361.210 86.520 361.490 95.550 ;
        RECT 362.090 86.520 362.370 95.550 ;
        RECT 362.970 86.520 363.250 95.550 ;
        RECT 338.695 86.040 359.365 86.370 ;
        RECT 363.655 85.760 363.945 95.740 ;
        RECT 334.115 85.470 363.945 85.760 ;
        RECT 364.455 96.310 406.605 96.600 ;
        RECT 364.455 96.030 364.745 96.310 ;
        RECT 406.315 96.030 406.605 96.310 ;
        RECT 364.455 95.740 366.825 96.030 ;
        RECT 402.475 95.740 406.605 96.030 ;
        RECT 364.455 85.760 364.745 95.740 ;
        RECT 365.150 86.520 365.430 95.550 ;
        RECT 366.030 86.520 366.310 95.550 ;
        RECT 366.910 86.520 367.190 95.550 ;
        RECT 367.790 86.520 368.070 95.550 ;
        RECT 368.670 86.520 368.950 95.550 ;
        RECT 369.550 86.520 369.830 95.550 ;
        RECT 370.430 86.520 370.710 95.550 ;
        RECT 371.310 86.520 371.590 95.550 ;
        RECT 372.190 86.520 372.470 95.550 ;
        RECT 373.070 86.520 373.350 95.550 ;
        RECT 373.950 86.520 374.230 95.550 ;
        RECT 374.830 86.520 375.110 95.550 ;
        RECT 375.710 86.520 375.990 95.550 ;
        RECT 376.590 86.520 376.870 95.550 ;
        RECT 377.470 86.520 377.750 95.550 ;
        RECT 378.350 86.520 378.630 95.550 ;
        RECT 379.230 86.520 379.510 95.550 ;
        RECT 380.110 86.520 380.390 95.550 ;
        RECT 380.990 86.520 381.270 95.550 ;
        RECT 381.870 86.520 382.150 95.550 ;
        RECT 382.750 86.520 383.030 95.550 ;
        RECT 383.630 86.520 383.910 95.550 ;
        RECT 384.510 86.520 384.790 95.550 ;
        RECT 385.390 86.520 385.670 95.550 ;
        RECT 386.270 86.520 386.550 95.550 ;
        RECT 387.150 86.520 387.430 95.550 ;
        RECT 388.030 86.520 388.310 95.550 ;
        RECT 388.910 86.520 389.190 95.550 ;
        RECT 389.790 86.520 390.070 95.550 ;
        RECT 390.670 86.520 390.950 95.550 ;
        RECT 391.550 86.520 391.830 95.550 ;
        RECT 392.430 86.520 392.710 95.550 ;
        RECT 393.310 86.520 393.590 95.550 ;
        RECT 394.190 86.520 394.470 95.550 ;
        RECT 395.070 86.520 395.350 95.550 ;
        RECT 395.950 86.520 396.230 95.550 ;
        RECT 396.830 86.520 397.110 95.550 ;
        RECT 397.710 86.520 397.990 95.550 ;
        RECT 398.590 86.520 398.870 95.550 ;
        RECT 399.470 86.520 399.750 95.550 ;
        RECT 400.350 86.520 400.630 95.550 ;
        RECT 401.230 86.520 401.510 95.550 ;
        RECT 402.110 86.520 402.390 95.550 ;
        RECT 402.990 86.520 403.270 95.550 ;
        RECT 403.870 86.520 404.150 95.550 ;
        RECT 404.750 86.520 405.030 95.550 ;
        RECT 405.630 86.520 405.910 95.550 ;
        RECT 367.275 86.040 402.025 86.370 ;
        RECT 406.315 85.760 406.605 95.740 ;
        RECT 472.625 96.535 474.935 96.825 ;
        RECT 478.905 96.535 481.215 96.825 ;
        RECT 453.275 94.115 471.065 94.405 ;
        RECT 453.275 93.855 453.565 94.115 ;
        RECT 453.275 93.565 456.445 93.855 ;
        RECT 456.935 93.565 467.405 93.895 ;
        RECT 470.775 93.855 471.065 94.115 ;
        RECT 467.895 93.565 471.065 93.855 ;
        RECT 434.835 91.445 443.425 91.735 ;
        RECT 434.835 91.185 435.125 91.445 ;
        RECT 443.135 91.185 443.425 91.445 ;
        RECT 434.835 90.885 437.145 91.185 ;
        RECT 441.115 90.885 443.425 91.185 ;
        RECT 434.835 87.965 435.125 90.885 ;
        RECT 435.495 90.450 435.725 90.705 ;
        RECT 436.375 90.450 436.605 90.705 ;
        RECT 437.255 90.450 437.485 90.705 ;
        RECT 435.480 88.950 435.740 90.450 ;
        RECT 436.360 88.950 436.620 90.450 ;
        RECT 437.240 88.950 437.500 90.450 ;
        RECT 435.495 88.705 435.725 88.950 ;
        RECT 436.375 88.705 436.605 88.950 ;
        RECT 437.255 88.705 437.485 88.950 ;
        RECT 438.085 88.515 438.415 90.705 ;
        RECT 439.015 90.450 439.245 90.705 ;
        RECT 439.000 88.950 439.260 90.450 ;
        RECT 439.015 88.705 439.245 88.950 ;
        RECT 439.845 88.515 440.175 90.705 ;
        RECT 440.775 90.450 441.005 90.705 ;
        RECT 441.655 90.450 441.885 90.705 ;
        RECT 442.535 90.450 442.765 90.705 ;
        RECT 440.760 88.950 441.020 90.450 ;
        RECT 441.640 88.950 441.900 90.450 ;
        RECT 442.520 88.950 442.780 90.450 ;
        RECT 440.775 88.705 441.005 88.950 ;
        RECT 441.655 88.705 441.885 88.950 ;
        RECT 442.535 88.705 442.765 88.950 ;
        RECT 437.595 88.185 440.665 88.515 ;
        RECT 443.135 87.965 443.425 90.885 ;
        RECT 434.835 87.675 443.425 87.965 ;
        RECT 444.055 91.445 452.645 91.735 ;
        RECT 444.055 91.175 444.345 91.445 ;
        RECT 452.355 91.175 452.645 91.445 ;
        RECT 444.055 90.885 446.365 91.175 ;
        RECT 450.335 90.885 452.645 91.175 ;
        RECT 444.055 87.960 444.345 90.885 ;
        RECT 444.715 90.450 444.945 90.695 ;
        RECT 445.595 90.450 445.825 90.695 ;
        RECT 446.475 90.450 446.705 90.695 ;
        RECT 444.700 88.950 444.960 90.450 ;
        RECT 445.580 88.950 445.840 90.450 ;
        RECT 446.460 88.950 446.720 90.450 ;
        RECT 444.715 88.705 444.945 88.950 ;
        RECT 445.595 88.705 445.825 88.950 ;
        RECT 446.475 88.705 446.705 88.950 ;
        RECT 447.340 88.705 447.600 90.695 ;
        RECT 448.235 90.450 448.465 90.695 ;
        RECT 448.220 88.950 448.480 90.450 ;
        RECT 448.235 88.705 448.465 88.950 ;
        RECT 449.100 88.705 449.360 90.695 ;
        RECT 449.995 90.450 450.225 90.695 ;
        RECT 450.875 90.450 451.105 90.695 ;
        RECT 451.755 90.450 451.985 90.695 ;
        RECT 449.980 88.950 450.240 90.450 ;
        RECT 450.860 88.950 451.120 90.450 ;
        RECT 451.740 88.950 452.000 90.450 ;
        RECT 449.995 88.705 450.225 88.950 ;
        RECT 450.875 88.705 451.105 88.950 ;
        RECT 451.755 88.705 451.985 88.950 ;
        RECT 446.815 88.185 449.885 88.515 ;
        RECT 452.355 87.960 452.645 90.885 ;
        RECT 444.055 87.670 452.645 87.960 ;
        RECT 453.275 91.185 453.565 93.565 ;
        RECT 453.935 93.065 454.165 93.375 ;
        RECT 455.215 93.065 455.445 93.375 ;
        RECT 456.495 93.065 456.725 93.375 ;
        RECT 453.920 91.565 454.180 93.065 ;
        RECT 455.200 91.565 455.460 93.065 ;
        RECT 456.480 91.565 456.740 93.065 ;
        RECT 453.935 91.375 454.165 91.565 ;
        RECT 455.215 91.375 455.445 91.565 ;
        RECT 456.495 91.375 456.725 91.565 ;
        RECT 462.040 91.375 462.300 93.375 ;
        RECT 467.615 93.065 467.845 93.375 ;
        RECT 468.895 93.065 469.125 93.375 ;
        RECT 470.175 93.065 470.405 93.375 ;
        RECT 467.600 91.565 467.860 93.065 ;
        RECT 468.880 91.565 469.140 93.065 ;
        RECT 470.160 91.565 470.420 93.065 ;
        RECT 467.615 91.375 467.845 91.565 ;
        RECT 468.895 91.375 469.125 91.565 ;
        RECT 470.175 91.375 470.405 91.565 ;
        RECT 470.775 91.185 471.065 93.565 ;
        RECT 472.625 93.345 472.915 96.535 ;
        RECT 473.285 95.965 473.515 96.345 ;
        RECT 474.165 95.965 474.395 96.345 ;
        RECT 473.270 94.465 473.530 95.965 ;
        RECT 474.150 94.465 474.410 95.965 ;
        RECT 473.285 94.085 473.515 94.465 ;
        RECT 474.165 94.085 474.395 94.465 ;
        RECT 475.030 94.085 475.290 96.345 ;
        RECT 475.910 94.085 476.170 96.345 ;
        RECT 476.790 94.085 477.050 96.345 ;
        RECT 477.685 94.085 477.945 96.345 ;
        RECT 478.550 94.085 478.810 96.345 ;
        RECT 479.445 95.965 479.675 96.345 ;
        RECT 480.325 95.965 480.555 96.345 ;
        RECT 479.430 94.465 479.690 95.965 ;
        RECT 480.310 94.465 480.570 95.965 ;
        RECT 479.445 94.085 479.675 94.465 ;
        RECT 480.325 94.085 480.555 94.465 ;
        RECT 473.940 93.565 478.455 93.895 ;
        RECT 480.925 93.345 481.215 96.535 ;
        RECT 487.050 95.570 487.340 105.530 ;
        RECT 487.540 104.980 492.920 105.310 ;
        RECT 487.750 101.275 487.980 104.790 ;
        RECT 488.630 101.275 488.860 104.790 ;
        RECT 487.735 99.275 487.995 101.275 ;
        RECT 488.615 99.275 488.875 101.275 ;
        RECT 487.750 95.760 487.980 99.275 ;
        RECT 488.630 95.760 488.860 99.275 ;
        RECT 489.495 95.760 489.755 104.790 ;
        RECT 490.375 95.760 490.635 104.790 ;
        RECT 491.255 95.760 491.515 104.790 ;
        RECT 492.135 95.760 492.395 104.790 ;
        RECT 493.015 95.760 493.275 104.790 ;
        RECT 493.910 101.275 494.140 104.790 ;
        RECT 494.790 101.275 495.020 104.790 ;
        RECT 493.895 99.275 494.155 101.275 ;
        RECT 494.775 99.275 495.035 101.275 ;
        RECT 493.910 95.760 494.140 99.275 ;
        RECT 494.790 95.760 495.020 99.275 ;
        RECT 495.430 95.570 495.720 105.530 ;
        RECT 487.050 95.280 489.400 95.570 ;
        RECT 493.370 95.280 495.720 95.570 ;
        RECT 487.050 95.020 487.340 95.280 ;
        RECT 495.430 95.020 495.720 95.280 ;
        RECT 487.050 94.730 495.720 95.020 ;
        RECT 496.820 97.085 505.410 97.375 ;
        RECT 496.820 96.825 497.110 97.085 ;
        RECT 505.120 96.825 505.410 97.085 ;
        RECT 496.820 96.535 499.130 96.825 ;
        RECT 503.100 96.535 505.410 96.825 ;
        RECT 472.625 93.055 481.215 93.345 ;
        RECT 496.820 93.345 497.110 96.535 ;
        RECT 497.480 95.965 497.710 96.345 ;
        RECT 498.360 95.965 498.590 96.345 ;
        RECT 497.465 94.465 497.725 95.965 ;
        RECT 498.345 94.465 498.605 95.965 ;
        RECT 497.480 94.085 497.710 94.465 ;
        RECT 498.360 94.085 498.590 94.465 ;
        RECT 499.225 94.085 499.485 96.345 ;
        RECT 500.105 94.085 500.365 96.345 ;
        RECT 500.985 94.085 501.245 96.345 ;
        RECT 501.865 94.085 502.125 96.345 ;
        RECT 502.745 94.085 503.005 96.345 ;
        RECT 503.640 95.965 503.870 96.345 ;
        RECT 504.520 95.965 504.750 96.345 ;
        RECT 503.625 94.465 503.885 95.965 ;
        RECT 504.505 94.465 504.765 95.965 ;
        RECT 503.640 94.085 503.870 94.465 ;
        RECT 504.520 94.085 504.750 94.465 ;
        RECT 497.630 93.565 502.650 93.895 ;
        RECT 505.120 93.345 505.410 96.535 ;
        RECT 496.820 93.055 505.410 93.345 ;
        RECT 453.275 90.895 456.445 91.185 ;
        RECT 453.275 87.965 453.565 90.895 ;
        RECT 456.935 90.855 467.405 91.185 ;
        RECT 467.895 90.895 471.065 91.185 ;
        RECT 453.935 90.450 454.165 90.705 ;
        RECT 455.215 90.450 455.445 90.705 ;
        RECT 456.495 90.450 456.725 90.705 ;
        RECT 453.920 88.950 454.180 90.450 ;
        RECT 455.200 88.950 455.460 90.450 ;
        RECT 456.480 88.950 456.740 90.450 ;
        RECT 453.935 88.705 454.165 88.950 ;
        RECT 455.215 88.705 455.445 88.950 ;
        RECT 456.495 88.705 456.725 88.950 ;
        RECT 462.040 88.705 462.300 90.705 ;
        RECT 467.615 90.450 467.845 90.705 ;
        RECT 468.895 90.450 469.125 90.705 ;
        RECT 470.175 90.450 470.405 90.705 ;
        RECT 467.600 88.950 467.860 90.450 ;
        RECT 468.880 88.950 469.140 90.450 ;
        RECT 470.160 88.950 470.420 90.450 ;
        RECT 467.615 88.705 467.845 88.950 ;
        RECT 468.895 88.705 469.125 88.950 ;
        RECT 470.175 88.705 470.405 88.950 ;
        RECT 456.935 88.225 461.845 88.515 ;
        RECT 462.495 88.225 467.405 88.515 ;
        RECT 470.775 87.965 471.065 90.895 ;
        RECT 453.275 87.675 471.065 87.965 ;
        RECT 472.625 91.705 481.215 91.995 ;
        RECT 472.625 91.445 472.915 91.705 ;
        RECT 480.925 91.445 481.215 91.705 ;
        RECT 472.625 91.155 474.935 91.445 ;
        RECT 478.905 91.155 481.215 91.445 ;
        RECT 472.625 87.965 472.915 91.155 ;
        RECT 473.285 90.450 473.515 90.965 ;
        RECT 474.165 90.450 474.395 90.965 ;
        RECT 475.045 90.450 475.275 90.965 ;
        RECT 473.270 88.950 473.530 90.450 ;
        RECT 474.150 88.950 474.410 90.450 ;
        RECT 475.030 88.950 475.290 90.450 ;
        RECT 473.285 88.705 473.515 88.950 ;
        RECT 474.165 88.705 474.395 88.950 ;
        RECT 475.045 88.705 475.275 88.950 ;
        RECT 475.910 88.705 476.170 90.965 ;
        RECT 476.805 90.450 477.035 90.965 ;
        RECT 476.790 88.950 477.050 90.450 ;
        RECT 476.805 88.705 477.035 88.950 ;
        RECT 477.685 88.705 477.945 90.965 ;
        RECT 478.565 90.450 478.795 90.965 ;
        RECT 479.445 90.450 479.675 90.965 ;
        RECT 480.325 90.450 480.555 90.965 ;
        RECT 478.550 88.950 478.810 90.450 ;
        RECT 479.430 88.950 479.690 90.450 ;
        RECT 480.310 88.950 480.570 90.450 ;
        RECT 478.565 88.705 478.795 88.950 ;
        RECT 479.445 88.705 479.675 88.950 ;
        RECT 480.325 88.705 480.555 88.950 ;
        RECT 475.385 88.185 478.455 88.515 ;
        RECT 480.925 87.965 481.215 91.155 ;
        RECT 472.625 87.675 481.215 87.965 ;
        RECT 487.090 91.445 495.680 91.735 ;
        RECT 487.090 88.515 487.380 91.445 ;
        RECT 489.850 90.895 492.920 91.225 ;
        RECT 487.750 90.450 487.980 90.705 ;
        RECT 488.630 90.450 488.860 90.705 ;
        RECT 489.510 90.450 489.740 90.705 ;
        RECT 487.735 88.950 487.995 90.450 ;
        RECT 488.615 88.950 488.875 90.450 ;
        RECT 489.495 88.950 489.755 90.450 ;
        RECT 487.750 88.705 487.980 88.950 ;
        RECT 488.630 88.705 488.860 88.950 ;
        RECT 489.510 88.705 489.740 88.950 ;
        RECT 490.375 88.705 490.635 90.705 ;
        RECT 491.270 90.450 491.500 90.705 ;
        RECT 491.255 88.950 491.515 90.450 ;
        RECT 491.270 88.705 491.500 88.950 ;
        RECT 492.135 88.705 492.395 90.705 ;
        RECT 493.030 90.450 493.260 90.705 ;
        RECT 493.910 90.450 494.140 90.705 ;
        RECT 494.790 90.450 495.020 90.705 ;
        RECT 493.015 88.950 493.275 90.450 ;
        RECT 493.895 88.950 494.155 90.450 ;
        RECT 494.775 88.950 495.035 90.450 ;
        RECT 493.030 88.705 493.260 88.950 ;
        RECT 493.910 88.705 494.140 88.950 ;
        RECT 494.790 88.705 495.020 88.950 ;
        RECT 495.390 88.515 495.680 91.445 ;
        RECT 487.090 88.225 489.400 88.515 ;
        RECT 493.370 88.225 495.680 88.515 ;
        RECT 487.090 87.965 487.380 88.225 ;
        RECT 495.390 87.965 495.680 88.225 ;
        RECT 487.090 87.675 495.680 87.965 ;
        RECT 496.820 91.705 505.410 91.995 ;
        RECT 496.820 91.445 497.110 91.705 ;
        RECT 505.120 91.445 505.410 91.705 ;
        RECT 496.820 91.155 499.130 91.445 ;
        RECT 503.100 91.155 505.410 91.445 ;
        RECT 496.820 87.965 497.110 91.155 ;
        RECT 497.480 90.450 497.710 90.965 ;
        RECT 498.360 90.450 498.590 90.965 ;
        RECT 499.240 90.450 499.470 90.965 ;
        RECT 497.465 88.950 497.725 90.450 ;
        RECT 498.345 88.950 498.605 90.450 ;
        RECT 499.225 88.950 499.485 90.450 ;
        RECT 497.480 88.705 497.710 88.950 ;
        RECT 498.360 88.705 498.590 88.950 ;
        RECT 499.240 88.705 499.470 88.950 ;
        RECT 500.105 88.705 500.365 90.965 ;
        RECT 501.000 90.450 501.230 90.965 ;
        RECT 500.985 88.950 501.245 90.450 ;
        RECT 501.000 88.705 501.230 88.950 ;
        RECT 501.865 88.705 502.125 90.965 ;
        RECT 502.760 90.450 502.990 90.965 ;
        RECT 503.640 90.450 503.870 90.965 ;
        RECT 504.520 90.450 504.750 90.965 ;
        RECT 502.745 88.950 503.005 90.450 ;
        RECT 503.625 88.950 503.885 90.450 ;
        RECT 504.505 88.950 504.765 90.450 ;
        RECT 502.760 88.705 502.990 88.950 ;
        RECT 503.640 88.705 503.870 88.950 ;
        RECT 504.520 88.705 504.750 88.950 ;
        RECT 499.580 88.185 502.650 88.515 ;
        RECT 505.120 87.965 505.410 91.155 ;
        RECT 496.820 87.675 505.410 87.965 ;
        RECT 364.455 85.470 406.605 85.760 ;
        RECT 185.685 78.940 186.995 81.045 ;
        RECT 187.695 78.940 189.005 81.045 ;
        RECT 189.705 78.940 191.015 81.045 ;
        RECT 191.715 78.940 193.025 81.045 ;
        RECT 193.725 78.940 195.035 81.045 ;
        RECT 195.735 78.940 197.045 81.045 ;
        RECT 197.745 78.940 199.055 81.045 ;
        RECT 199.755 78.940 201.065 81.045 ;
        RECT 201.765 78.940 203.075 81.045 ;
        RECT 203.775 78.940 205.085 81.045 ;
        RECT 205.785 78.940 207.095 81.045 ;
        RECT 207.795 78.940 209.105 81.045 ;
        RECT 209.805 78.940 211.115 81.045 ;
        RECT 211.815 78.940 213.125 81.045 ;
        RECT 213.825 78.940 215.135 81.045 ;
        RECT 215.835 78.940 217.145 81.045 ;
        RECT 217.845 78.940 219.155 81.045 ;
        RECT 219.855 78.940 221.165 81.045 ;
        RECT 221.865 78.940 223.175 81.045 ;
        RECT 223.875 78.940 225.185 81.045 ;
        RECT 225.885 78.940 227.195 81.045 ;
        RECT 227.895 78.940 229.205 81.045 ;
        RECT 229.905 78.940 231.215 81.045 ;
        RECT 231.915 78.940 233.225 81.045 ;
        RECT 233.925 78.940 235.235 81.045 ;
        RECT 235.935 78.940 237.245 81.045 ;
        RECT 237.945 78.940 239.255 81.045 ;
        RECT 239.955 78.940 241.265 81.045 ;
        RECT 241.965 78.940 243.275 81.045 ;
        RECT 243.975 78.940 245.285 81.045 ;
        RECT 245.985 78.940 247.295 81.045 ;
        RECT 247.995 78.940 249.305 81.045 ;
        RECT 250.005 78.940 251.315 81.045 ;
        RECT 252.015 78.940 253.325 81.045 ;
        RECT 254.025 78.940 255.335 81.045 ;
        RECT 256.035 78.940 257.345 81.045 ;
        RECT 258.045 78.940 259.355 81.045 ;
        RECT 260.055 78.940 261.365 81.045 ;
        RECT 262.065 78.940 263.375 81.045 ;
        RECT 264.075 78.940 265.385 81.045 ;
        RECT 266.085 78.940 267.395 81.045 ;
        RECT 268.095 78.940 269.405 81.045 ;
        RECT 270.105 78.940 271.415 81.045 ;
        RECT 272.115 78.940 273.425 81.045 ;
        RECT 274.125 78.940 275.435 81.045 ;
        RECT 276.135 78.940 277.445 81.045 ;
        RECT 278.145 78.940 279.455 81.045 ;
        RECT 280.155 78.940 281.465 81.045 ;
        RECT 282.165 78.940 283.475 81.045 ;
        RECT 284.175 78.940 285.485 81.045 ;
        RECT 286.185 78.940 287.495 81.045 ;
        RECT 288.195 78.940 289.505 81.045 ;
        RECT 290.205 78.940 291.515 81.045 ;
        RECT 292.215 78.940 293.525 81.045 ;
        RECT 301.220 78.940 302.530 81.045 ;
        RECT 303.230 78.940 304.540 81.045 ;
        RECT 305.240 78.940 306.550 81.045 ;
        RECT 307.250 78.940 308.560 81.045 ;
        RECT 309.260 78.940 310.570 81.045 ;
        RECT 311.270 78.940 312.580 81.045 ;
        RECT 313.280 78.940 314.590 81.045 ;
        RECT 315.290 78.940 316.600 81.045 ;
        RECT 317.300 78.940 318.610 81.045 ;
        RECT 319.310 78.940 320.620 81.045 ;
        RECT 321.320 78.940 322.630 81.045 ;
        RECT 323.330 78.940 324.640 81.045 ;
        RECT 325.340 78.940 326.650 81.045 ;
        RECT 327.350 78.940 328.660 81.045 ;
        RECT 329.360 78.940 330.670 81.045 ;
        RECT 331.370 78.940 332.680 81.045 ;
        RECT 333.380 78.940 334.690 81.045 ;
        RECT 335.390 78.940 336.700 81.045 ;
        RECT 337.400 78.940 338.710 81.045 ;
        RECT 339.410 78.940 340.720 81.045 ;
        RECT 341.420 78.940 342.730 81.045 ;
        RECT 343.430 78.940 344.740 81.045 ;
        RECT 345.440 78.940 346.750 81.045 ;
        RECT 347.450 78.940 348.760 81.045 ;
        RECT 349.460 78.940 350.770 81.045 ;
        RECT 351.470 78.940 352.780 81.045 ;
        RECT 353.480 78.940 354.790 81.045 ;
        RECT 355.490 78.940 356.800 81.045 ;
        RECT 357.500 78.940 358.810 81.045 ;
        RECT 359.510 78.940 360.820 81.045 ;
        RECT 361.520 78.940 362.830 81.045 ;
        RECT 363.530 78.940 364.840 81.045 ;
        RECT 365.540 78.940 366.850 81.045 ;
        RECT 367.550 78.940 368.860 81.045 ;
        RECT 369.560 78.940 370.870 81.045 ;
        RECT 371.570 78.940 372.880 81.045 ;
        RECT 373.580 78.940 374.890 81.045 ;
        RECT 375.590 78.940 376.900 81.045 ;
        RECT 377.600 78.940 378.910 81.045 ;
        RECT 379.610 78.940 380.920 81.045 ;
        RECT 381.620 78.940 382.930 81.045 ;
        RECT 383.630 78.940 384.940 81.045 ;
        RECT 385.640 78.940 386.950 81.045 ;
        RECT 387.650 78.940 388.960 81.045 ;
        RECT 389.660 78.940 390.970 81.045 ;
        RECT 391.670 78.940 392.980 81.045 ;
        RECT 393.680 78.940 394.990 81.045 ;
        RECT 395.690 78.940 397.000 81.045 ;
        RECT 397.700 78.940 399.010 81.045 ;
        RECT 399.710 78.940 401.020 81.045 ;
        RECT 401.720 78.940 403.030 81.045 ;
        RECT 403.730 78.940 405.040 81.045 ;
        RECT 405.740 78.940 407.050 81.045 ;
        RECT 407.750 78.940 409.060 81.045 ;
        RECT 438.410 80.505 439.720 82.610 ;
        RECT 440.420 80.505 441.730 82.610 ;
        RECT 442.430 80.505 443.740 82.610 ;
        RECT 444.440 80.505 445.750 82.610 ;
        RECT 446.450 80.505 447.760 82.610 ;
        RECT 448.460 80.505 449.770 82.610 ;
        RECT 450.470 80.505 451.780 82.610 ;
        RECT 452.480 80.505 453.790 82.610 ;
        RECT 454.490 80.505 455.800 82.610 ;
        RECT 456.500 80.505 457.810 82.610 ;
        RECT 458.510 80.505 459.820 82.610 ;
        RECT 460.520 80.505 461.830 82.610 ;
        RECT 462.530 80.505 463.840 82.610 ;
        RECT 464.540 80.505 465.850 82.610 ;
        RECT 466.550 80.505 467.860 82.610 ;
        RECT 468.560 80.505 469.870 82.610 ;
        RECT 470.570 80.505 471.880 82.610 ;
        RECT 472.580 80.505 473.890 82.610 ;
        RECT 474.590 80.505 475.900 82.610 ;
        RECT 476.600 80.505 477.910 82.610 ;
        RECT 478.610 80.505 479.920 82.610 ;
        RECT 480.620 80.505 481.930 82.610 ;
        RECT 482.630 80.505 483.940 82.610 ;
        RECT 484.640 80.505 485.950 82.610 ;
        RECT 486.650 80.505 487.960 82.610 ;
        RECT 488.660 80.505 489.970 82.610 ;
        RECT 490.670 80.505 491.980 82.610 ;
        RECT 492.680 80.505 493.990 82.610 ;
        RECT 494.690 80.505 496.000 82.610 ;
        RECT 496.700 80.505 498.010 82.610 ;
        RECT 498.710 80.505 500.020 82.610 ;
        RECT 500.720 80.505 502.030 82.610 ;
        RECT 184.800 74.180 185.060 76.180 ;
        RECT 294.150 74.180 294.410 76.180 ;
        RECT 300.335 74.180 300.595 76.180 ;
        RECT 409.685 74.180 409.945 76.180 ;
        RECT 437.510 73.900 437.800 75.900 ;
        RECT 502.640 73.900 502.930 75.900 ;
        RECT 185.685 69.345 186.995 71.450 ;
        RECT 187.695 69.345 189.005 71.450 ;
        RECT 189.705 69.345 191.015 71.450 ;
        RECT 191.715 69.345 193.025 71.450 ;
        RECT 193.725 69.345 195.035 71.450 ;
        RECT 195.735 69.345 197.045 71.450 ;
        RECT 197.745 69.345 199.055 71.450 ;
        RECT 199.755 69.345 201.065 71.450 ;
        RECT 201.765 69.345 203.075 71.450 ;
        RECT 203.775 69.345 205.085 71.450 ;
        RECT 205.785 69.345 207.095 71.450 ;
        RECT 207.795 69.345 209.105 71.450 ;
        RECT 209.805 69.345 211.115 71.450 ;
        RECT 211.815 69.345 213.125 71.450 ;
        RECT 213.825 69.345 215.135 71.450 ;
        RECT 215.835 69.345 217.145 71.450 ;
        RECT 217.845 69.345 219.155 71.450 ;
        RECT 219.855 69.345 221.165 71.450 ;
        RECT 221.865 69.345 223.175 71.450 ;
        RECT 223.875 69.345 225.185 71.450 ;
        RECT 225.885 69.345 227.195 71.450 ;
        RECT 227.895 69.345 229.205 71.450 ;
        RECT 229.905 69.345 231.215 71.450 ;
        RECT 231.915 69.345 233.225 71.450 ;
        RECT 233.925 69.345 235.235 71.450 ;
        RECT 235.935 69.345 237.245 71.450 ;
        RECT 237.945 69.345 239.255 71.450 ;
        RECT 239.955 69.345 241.265 71.450 ;
        RECT 241.965 69.345 243.275 71.450 ;
        RECT 243.975 69.345 245.285 71.450 ;
        RECT 245.985 69.345 247.295 71.450 ;
        RECT 247.995 69.345 249.305 71.450 ;
        RECT 250.005 69.345 251.315 71.450 ;
        RECT 252.015 69.345 253.325 71.450 ;
        RECT 254.025 69.345 255.335 71.450 ;
        RECT 256.035 69.345 257.345 71.450 ;
        RECT 258.045 69.345 259.355 71.450 ;
        RECT 260.055 69.345 261.365 71.450 ;
        RECT 262.065 69.345 263.375 71.450 ;
        RECT 264.075 69.345 265.385 71.450 ;
        RECT 266.085 69.345 267.395 71.450 ;
        RECT 268.095 69.345 269.405 71.450 ;
        RECT 270.105 69.345 271.415 71.450 ;
        RECT 272.115 69.345 273.425 71.450 ;
        RECT 274.125 69.345 275.435 71.450 ;
        RECT 276.135 69.345 277.445 71.450 ;
        RECT 278.145 69.345 279.455 71.450 ;
        RECT 280.155 69.345 281.465 71.450 ;
        RECT 282.165 69.345 283.475 71.450 ;
        RECT 284.175 69.345 285.485 71.450 ;
        RECT 286.185 69.345 287.495 71.450 ;
        RECT 288.195 69.345 289.505 71.450 ;
        RECT 290.205 69.345 291.515 71.450 ;
        RECT 292.215 69.345 293.525 71.450 ;
        RECT 301.220 69.345 302.530 71.450 ;
        RECT 303.230 69.345 304.540 71.450 ;
        RECT 305.240 69.345 306.550 71.450 ;
        RECT 307.250 69.345 308.560 71.450 ;
        RECT 309.260 69.345 310.570 71.450 ;
        RECT 311.270 69.345 312.580 71.450 ;
        RECT 313.280 69.345 314.590 71.450 ;
        RECT 315.290 69.345 316.600 71.450 ;
        RECT 317.300 69.345 318.610 71.450 ;
        RECT 319.310 69.345 320.620 71.450 ;
        RECT 321.320 69.345 322.630 71.450 ;
        RECT 323.330 69.345 324.640 71.450 ;
        RECT 325.340 69.345 326.650 71.450 ;
        RECT 327.350 69.345 328.660 71.450 ;
        RECT 329.360 69.345 330.670 71.450 ;
        RECT 331.370 69.345 332.680 71.450 ;
        RECT 333.380 69.345 334.690 71.450 ;
        RECT 335.390 69.345 336.700 71.450 ;
        RECT 337.400 69.345 338.710 71.450 ;
        RECT 339.410 69.345 340.720 71.450 ;
        RECT 341.420 69.345 342.730 71.450 ;
        RECT 343.430 69.345 344.740 71.450 ;
        RECT 345.440 69.345 346.750 71.450 ;
        RECT 347.450 69.345 348.760 71.450 ;
        RECT 349.460 69.345 350.770 71.450 ;
        RECT 351.470 69.345 352.780 71.450 ;
        RECT 353.480 69.345 354.790 71.450 ;
        RECT 355.490 69.345 356.800 71.450 ;
        RECT 357.500 69.345 358.810 71.450 ;
        RECT 359.510 69.345 360.820 71.450 ;
        RECT 361.520 69.345 362.830 71.450 ;
        RECT 363.530 69.345 364.840 71.450 ;
        RECT 365.540 69.345 366.850 71.450 ;
        RECT 367.550 69.345 368.860 71.450 ;
        RECT 369.560 69.345 370.870 71.450 ;
        RECT 371.570 69.345 372.880 71.450 ;
        RECT 373.580 69.345 374.890 71.450 ;
        RECT 375.590 69.345 376.900 71.450 ;
        RECT 377.600 69.345 378.910 71.450 ;
        RECT 379.610 69.345 380.920 71.450 ;
        RECT 381.620 69.345 382.930 71.450 ;
        RECT 383.630 69.345 384.940 71.450 ;
        RECT 385.640 69.345 386.950 71.450 ;
        RECT 387.650 69.345 388.960 71.450 ;
        RECT 389.660 69.345 390.970 71.450 ;
        RECT 391.670 69.345 392.980 71.450 ;
        RECT 393.680 69.345 394.990 71.450 ;
        RECT 395.690 69.345 397.000 71.450 ;
        RECT 397.700 69.345 399.010 71.450 ;
        RECT 399.710 69.345 401.020 71.450 ;
        RECT 401.720 69.345 403.030 71.450 ;
        RECT 403.730 69.345 405.040 71.450 ;
        RECT 405.740 69.345 407.050 71.450 ;
        RECT 407.750 69.345 409.060 71.450 ;
        RECT 438.410 70.910 439.720 73.015 ;
        RECT 440.420 70.910 441.730 73.015 ;
        RECT 442.430 70.910 443.740 73.015 ;
        RECT 444.440 70.910 445.750 73.015 ;
        RECT 446.450 70.910 447.760 73.015 ;
        RECT 448.460 70.910 449.770 73.015 ;
        RECT 450.470 70.910 451.780 73.015 ;
        RECT 452.480 70.910 453.790 73.015 ;
        RECT 454.490 70.910 455.800 73.015 ;
        RECT 456.500 70.910 457.810 73.015 ;
        RECT 458.510 70.910 459.820 73.015 ;
        RECT 460.520 70.910 461.830 73.015 ;
        RECT 462.530 70.910 463.840 73.015 ;
        RECT 464.540 70.910 465.850 73.015 ;
        RECT 466.550 70.910 467.860 73.015 ;
        RECT 468.560 70.910 469.870 73.015 ;
        RECT 470.570 70.910 471.880 73.015 ;
        RECT 472.580 70.910 473.890 73.015 ;
        RECT 474.590 70.910 475.900 73.015 ;
        RECT 476.600 70.910 477.910 73.015 ;
        RECT 478.610 70.910 479.920 73.015 ;
        RECT 480.620 70.910 481.930 73.015 ;
        RECT 482.630 70.910 483.940 73.015 ;
        RECT 484.640 70.910 485.950 73.015 ;
        RECT 486.650 70.910 487.960 73.015 ;
        RECT 488.660 70.910 489.970 73.015 ;
        RECT 490.670 70.910 491.980 73.015 ;
        RECT 492.680 70.910 493.990 73.015 ;
        RECT 494.690 70.910 496.000 73.015 ;
        RECT 496.700 70.910 498.010 73.015 ;
        RECT 498.710 70.910 500.020 73.015 ;
        RECT 500.720 70.910 502.030 73.015 ;
        RECT 185.685 64.795 186.995 66.900 ;
        RECT 187.695 64.795 189.005 66.900 ;
        RECT 189.705 64.795 191.015 66.900 ;
        RECT 191.715 64.795 193.025 66.900 ;
        RECT 193.725 64.795 195.035 66.900 ;
        RECT 195.735 64.795 197.045 66.900 ;
        RECT 197.745 64.795 199.055 66.900 ;
        RECT 199.755 64.795 201.065 66.900 ;
        RECT 201.765 64.795 203.075 66.900 ;
        RECT 203.775 64.795 205.085 66.900 ;
        RECT 205.785 64.795 207.095 66.900 ;
        RECT 207.795 64.795 209.105 66.900 ;
        RECT 209.805 64.795 211.115 66.900 ;
        RECT 211.815 64.795 213.125 66.900 ;
        RECT 213.825 64.795 215.135 66.900 ;
        RECT 215.835 64.795 217.145 66.900 ;
        RECT 217.845 64.795 219.155 66.900 ;
        RECT 219.855 64.795 221.165 66.900 ;
        RECT 221.865 64.795 223.175 66.900 ;
        RECT 223.875 64.795 225.185 66.900 ;
        RECT 225.885 64.795 227.195 66.900 ;
        RECT 227.895 64.795 229.205 66.900 ;
        RECT 229.905 64.795 231.215 66.900 ;
        RECT 231.915 64.795 233.225 66.900 ;
        RECT 233.925 64.795 235.235 66.900 ;
        RECT 235.935 64.795 237.245 66.900 ;
        RECT 237.945 64.795 239.255 66.900 ;
        RECT 239.955 64.795 241.265 66.900 ;
        RECT 241.965 64.795 243.275 66.900 ;
        RECT 243.975 64.795 245.285 66.900 ;
        RECT 245.985 64.795 247.295 66.900 ;
        RECT 247.995 64.795 249.305 66.900 ;
        RECT 250.005 64.795 251.315 66.900 ;
        RECT 252.015 64.795 253.325 66.900 ;
        RECT 254.025 64.795 255.335 66.900 ;
        RECT 256.035 64.795 257.345 66.900 ;
        RECT 258.045 64.795 259.355 66.900 ;
        RECT 260.055 64.795 261.365 66.900 ;
        RECT 262.065 64.795 263.375 66.900 ;
        RECT 264.075 64.795 265.385 66.900 ;
        RECT 266.085 64.795 267.395 66.900 ;
        RECT 268.095 64.795 269.405 66.900 ;
        RECT 270.105 64.795 271.415 66.900 ;
        RECT 272.115 64.795 273.425 66.900 ;
        RECT 274.125 64.795 275.435 66.900 ;
        RECT 276.135 64.795 277.445 66.900 ;
        RECT 278.145 64.795 279.455 66.900 ;
        RECT 280.155 64.795 281.465 66.900 ;
        RECT 282.165 64.795 283.475 66.900 ;
        RECT 284.175 64.795 285.485 66.900 ;
        RECT 286.185 64.795 287.495 66.900 ;
        RECT 288.195 64.795 289.505 66.900 ;
        RECT 290.205 64.795 291.515 66.900 ;
        RECT 292.215 64.795 293.525 66.900 ;
        RECT 301.220 64.795 302.530 66.900 ;
        RECT 303.230 64.795 304.540 66.900 ;
        RECT 305.240 64.795 306.550 66.900 ;
        RECT 307.250 64.795 308.560 66.900 ;
        RECT 309.260 64.795 310.570 66.900 ;
        RECT 311.270 64.795 312.580 66.900 ;
        RECT 313.280 64.795 314.590 66.900 ;
        RECT 315.290 64.795 316.600 66.900 ;
        RECT 317.300 64.795 318.610 66.900 ;
        RECT 319.310 64.795 320.620 66.900 ;
        RECT 321.320 64.795 322.630 66.900 ;
        RECT 323.330 64.795 324.640 66.900 ;
        RECT 325.340 64.795 326.650 66.900 ;
        RECT 327.350 64.795 328.660 66.900 ;
        RECT 329.360 64.795 330.670 66.900 ;
        RECT 331.370 64.795 332.680 66.900 ;
        RECT 333.380 64.795 334.690 66.900 ;
        RECT 335.390 64.795 336.700 66.900 ;
        RECT 337.400 64.795 338.710 66.900 ;
        RECT 339.410 64.795 340.720 66.900 ;
        RECT 341.420 64.795 342.730 66.900 ;
        RECT 343.430 64.795 344.740 66.900 ;
        RECT 345.440 64.795 346.750 66.900 ;
        RECT 347.450 64.795 348.760 66.900 ;
        RECT 349.460 64.795 350.770 66.900 ;
        RECT 351.470 64.795 352.780 66.900 ;
        RECT 353.480 64.795 354.790 66.900 ;
        RECT 355.490 64.795 356.800 66.900 ;
        RECT 357.500 64.795 358.810 66.900 ;
        RECT 359.510 64.795 360.820 66.900 ;
        RECT 361.520 64.795 362.830 66.900 ;
        RECT 363.530 64.795 364.840 66.900 ;
        RECT 365.540 64.795 366.850 66.900 ;
        RECT 367.550 64.795 368.860 66.900 ;
        RECT 369.560 64.795 370.870 66.900 ;
        RECT 371.570 64.795 372.880 66.900 ;
        RECT 373.580 64.795 374.890 66.900 ;
        RECT 375.590 64.795 376.900 66.900 ;
        RECT 377.600 64.795 378.910 66.900 ;
        RECT 379.610 64.795 380.920 66.900 ;
        RECT 381.620 64.795 382.930 66.900 ;
        RECT 383.630 64.795 384.940 66.900 ;
        RECT 385.640 64.795 386.950 66.900 ;
        RECT 387.650 64.795 388.960 66.900 ;
        RECT 389.660 64.795 390.970 66.900 ;
        RECT 391.670 64.795 392.980 66.900 ;
        RECT 393.680 64.795 394.990 66.900 ;
        RECT 395.690 64.795 397.000 66.900 ;
        RECT 397.700 64.795 399.010 66.900 ;
        RECT 399.710 64.795 401.020 66.900 ;
        RECT 401.720 64.795 403.030 66.900 ;
        RECT 403.730 64.795 405.040 66.900 ;
        RECT 405.740 64.795 407.050 66.900 ;
        RECT 407.750 64.795 409.060 66.900 ;
        RECT 184.800 60.035 185.060 62.035 ;
        RECT 294.150 60.035 294.410 62.035 ;
        RECT 300.335 60.035 300.595 62.035 ;
        RECT 409.685 60.035 409.945 62.035 ;
        RECT 185.685 55.200 186.995 57.305 ;
        RECT 187.695 55.200 189.005 57.305 ;
        RECT 189.705 55.200 191.015 57.305 ;
        RECT 191.715 55.200 193.025 57.305 ;
        RECT 193.725 55.200 195.035 57.305 ;
        RECT 195.735 55.200 197.045 57.305 ;
        RECT 197.745 55.200 199.055 57.305 ;
        RECT 199.755 55.200 201.065 57.305 ;
        RECT 201.765 55.200 203.075 57.305 ;
        RECT 203.775 55.200 205.085 57.305 ;
        RECT 205.785 55.200 207.095 57.305 ;
        RECT 207.795 55.200 209.105 57.305 ;
        RECT 209.805 55.200 211.115 57.305 ;
        RECT 211.815 55.200 213.125 57.305 ;
        RECT 213.825 55.200 215.135 57.305 ;
        RECT 215.835 55.200 217.145 57.305 ;
        RECT 217.845 55.200 219.155 57.305 ;
        RECT 219.855 55.200 221.165 57.305 ;
        RECT 221.865 55.200 223.175 57.305 ;
        RECT 223.875 55.200 225.185 57.305 ;
        RECT 225.885 55.200 227.195 57.305 ;
        RECT 227.895 55.200 229.205 57.305 ;
        RECT 229.905 55.200 231.215 57.305 ;
        RECT 231.915 55.200 233.225 57.305 ;
        RECT 233.925 55.200 235.235 57.305 ;
        RECT 235.935 55.200 237.245 57.305 ;
        RECT 237.945 55.200 239.255 57.305 ;
        RECT 239.955 55.200 241.265 57.305 ;
        RECT 241.965 55.200 243.275 57.305 ;
        RECT 243.975 55.200 245.285 57.305 ;
        RECT 245.985 55.200 247.295 57.305 ;
        RECT 247.995 55.200 249.305 57.305 ;
        RECT 250.005 55.200 251.315 57.305 ;
        RECT 252.015 55.200 253.325 57.305 ;
        RECT 254.025 55.200 255.335 57.305 ;
        RECT 256.035 55.200 257.345 57.305 ;
        RECT 258.045 55.200 259.355 57.305 ;
        RECT 260.055 55.200 261.365 57.305 ;
        RECT 262.065 55.200 263.375 57.305 ;
        RECT 264.075 55.200 265.385 57.305 ;
        RECT 266.085 55.200 267.395 57.305 ;
        RECT 268.095 55.200 269.405 57.305 ;
        RECT 270.105 55.200 271.415 57.305 ;
        RECT 272.115 55.200 273.425 57.305 ;
        RECT 274.125 55.200 275.435 57.305 ;
        RECT 276.135 55.200 277.445 57.305 ;
        RECT 278.145 55.200 279.455 57.305 ;
        RECT 280.155 55.200 281.465 57.305 ;
        RECT 282.165 55.200 283.475 57.305 ;
        RECT 284.175 55.200 285.485 57.305 ;
        RECT 286.185 55.200 287.495 57.305 ;
        RECT 288.195 55.200 289.505 57.305 ;
        RECT 290.205 55.200 291.515 57.305 ;
        RECT 292.215 55.200 293.525 57.305 ;
        RECT 301.220 55.200 302.530 57.305 ;
        RECT 303.230 55.200 304.540 57.305 ;
        RECT 305.240 55.200 306.550 57.305 ;
        RECT 307.250 55.200 308.560 57.305 ;
        RECT 309.260 55.200 310.570 57.305 ;
        RECT 311.270 55.200 312.580 57.305 ;
        RECT 313.280 55.200 314.590 57.305 ;
        RECT 315.290 55.200 316.600 57.305 ;
        RECT 317.300 55.200 318.610 57.305 ;
        RECT 319.310 55.200 320.620 57.305 ;
        RECT 321.320 55.200 322.630 57.305 ;
        RECT 323.330 55.200 324.640 57.305 ;
        RECT 325.340 55.200 326.650 57.305 ;
        RECT 327.350 55.200 328.660 57.305 ;
        RECT 329.360 55.200 330.670 57.305 ;
        RECT 331.370 55.200 332.680 57.305 ;
        RECT 333.380 55.200 334.690 57.305 ;
        RECT 335.390 55.200 336.700 57.305 ;
        RECT 337.400 55.200 338.710 57.305 ;
        RECT 339.410 55.200 340.720 57.305 ;
        RECT 341.420 55.200 342.730 57.305 ;
        RECT 343.430 55.200 344.740 57.305 ;
        RECT 345.440 55.200 346.750 57.305 ;
        RECT 347.450 55.200 348.760 57.305 ;
        RECT 349.460 55.200 350.770 57.305 ;
        RECT 351.470 55.200 352.780 57.305 ;
        RECT 353.480 55.200 354.790 57.305 ;
        RECT 355.490 55.200 356.800 57.305 ;
        RECT 357.500 55.200 358.810 57.305 ;
        RECT 359.510 55.200 360.820 57.305 ;
        RECT 361.520 55.200 362.830 57.305 ;
        RECT 363.530 55.200 364.840 57.305 ;
        RECT 365.540 55.200 366.850 57.305 ;
        RECT 367.550 55.200 368.860 57.305 ;
        RECT 369.560 55.200 370.870 57.305 ;
        RECT 371.570 55.200 372.880 57.305 ;
        RECT 373.580 55.200 374.890 57.305 ;
        RECT 375.590 55.200 376.900 57.305 ;
        RECT 377.600 55.200 378.910 57.305 ;
        RECT 379.610 55.200 380.920 57.305 ;
        RECT 381.620 55.200 382.930 57.305 ;
        RECT 383.630 55.200 384.940 57.305 ;
        RECT 385.640 55.200 386.950 57.305 ;
        RECT 387.650 55.200 388.960 57.305 ;
        RECT 389.660 55.200 390.970 57.305 ;
        RECT 391.670 55.200 392.980 57.305 ;
        RECT 393.680 55.200 394.990 57.305 ;
        RECT 395.690 55.200 397.000 57.305 ;
        RECT 397.700 55.200 399.010 57.305 ;
        RECT 399.710 55.200 401.020 57.305 ;
        RECT 401.720 55.200 403.030 57.305 ;
        RECT 403.730 55.200 405.040 57.305 ;
        RECT 405.740 55.200 407.050 57.305 ;
        RECT 407.750 55.200 409.060 57.305 ;
        RECT 208.045 52.170 237.875 52.460 ;
        RECT 208.045 42.190 208.335 52.170 ;
        RECT 212.625 51.560 233.295 51.890 ;
        RECT 208.740 42.380 209.020 51.410 ;
        RECT 209.620 42.380 209.900 51.410 ;
        RECT 210.500 42.380 210.780 51.410 ;
        RECT 211.380 42.380 211.660 51.410 ;
        RECT 212.260 42.380 212.540 51.410 ;
        RECT 213.140 42.380 213.420 51.410 ;
        RECT 214.020 42.380 214.300 51.410 ;
        RECT 214.900 42.380 215.180 51.410 ;
        RECT 215.780 42.380 216.060 51.410 ;
        RECT 216.660 42.380 216.940 51.410 ;
        RECT 217.540 42.380 217.820 51.410 ;
        RECT 218.420 42.380 218.700 51.410 ;
        RECT 219.300 42.380 219.580 51.410 ;
        RECT 220.180 42.380 220.460 51.410 ;
        RECT 221.060 42.380 221.340 51.410 ;
        RECT 221.940 42.380 222.220 51.410 ;
        RECT 222.820 42.380 223.100 51.410 ;
        RECT 223.700 42.380 223.980 51.410 ;
        RECT 224.580 42.380 224.860 51.410 ;
        RECT 225.460 42.380 225.740 51.410 ;
        RECT 226.340 42.380 226.620 51.410 ;
        RECT 227.220 42.380 227.500 51.410 ;
        RECT 228.100 42.380 228.380 51.410 ;
        RECT 228.980 42.380 229.260 51.410 ;
        RECT 229.860 42.380 230.140 51.410 ;
        RECT 230.740 42.380 231.020 51.410 ;
        RECT 231.620 42.380 231.900 51.410 ;
        RECT 232.500 42.380 232.780 51.410 ;
        RECT 233.380 42.380 233.660 51.410 ;
        RECT 234.260 42.380 234.540 51.410 ;
        RECT 235.140 42.380 235.420 51.410 ;
        RECT 236.020 42.380 236.300 51.410 ;
        RECT 236.900 42.380 237.180 51.410 ;
        RECT 237.585 42.190 237.875 52.170 ;
        RECT 208.045 41.900 212.175 42.190 ;
        RECT 233.745 41.900 237.875 42.190 ;
        RECT 208.045 41.620 208.335 41.900 ;
        RECT 237.585 41.620 237.875 41.900 ;
        RECT 208.045 41.330 237.875 41.620 ;
        RECT 238.385 52.170 280.535 52.460 ;
        RECT 238.385 42.190 238.675 52.170 ;
        RECT 241.205 51.560 275.955 51.890 ;
        RECT 239.080 42.380 239.360 51.410 ;
        RECT 239.960 42.380 240.240 51.410 ;
        RECT 240.840 42.380 241.120 51.410 ;
        RECT 241.720 42.380 242.000 51.410 ;
        RECT 242.600 42.380 242.880 51.410 ;
        RECT 243.480 42.380 243.760 51.410 ;
        RECT 244.360 42.380 244.640 51.410 ;
        RECT 245.240 42.380 245.520 51.410 ;
        RECT 246.120 42.380 246.400 51.410 ;
        RECT 247.000 42.380 247.280 51.410 ;
        RECT 247.880 42.380 248.160 51.410 ;
        RECT 248.760 42.380 249.040 51.410 ;
        RECT 249.640 42.380 249.920 51.410 ;
        RECT 250.520 42.380 250.800 51.410 ;
        RECT 251.400 42.380 251.680 51.410 ;
        RECT 252.280 42.380 252.560 51.410 ;
        RECT 253.160 42.380 253.440 51.410 ;
        RECT 254.040 42.380 254.320 51.410 ;
        RECT 254.920 42.380 255.200 51.410 ;
        RECT 255.800 42.380 256.080 51.410 ;
        RECT 256.680 42.380 256.960 51.410 ;
        RECT 257.560 42.380 257.840 51.410 ;
        RECT 258.440 42.380 258.720 51.410 ;
        RECT 259.320 42.380 259.600 51.410 ;
        RECT 260.200 42.380 260.480 51.410 ;
        RECT 261.080 42.380 261.360 51.410 ;
        RECT 261.960 42.380 262.240 51.410 ;
        RECT 262.840 42.380 263.120 51.410 ;
        RECT 263.720 42.380 264.000 51.410 ;
        RECT 264.600 42.380 264.880 51.410 ;
        RECT 265.480 42.380 265.760 51.410 ;
        RECT 266.360 42.380 266.640 51.410 ;
        RECT 267.240 42.380 267.520 51.410 ;
        RECT 268.120 42.380 268.400 51.410 ;
        RECT 269.000 42.380 269.280 51.410 ;
        RECT 269.880 42.380 270.160 51.410 ;
        RECT 270.760 42.380 271.040 51.410 ;
        RECT 271.640 42.380 271.920 51.410 ;
        RECT 272.520 42.380 272.800 51.410 ;
        RECT 273.400 42.380 273.680 51.410 ;
        RECT 274.280 42.380 274.560 51.410 ;
        RECT 275.160 42.380 275.440 51.410 ;
        RECT 276.040 42.380 276.320 51.410 ;
        RECT 276.920 42.380 277.200 51.410 ;
        RECT 277.800 42.380 278.080 51.410 ;
        RECT 278.680 42.380 278.960 51.410 ;
        RECT 279.560 42.380 279.840 51.410 ;
        RECT 280.245 42.190 280.535 52.170 ;
        RECT 238.385 41.900 240.755 42.190 ;
        RECT 276.405 41.900 280.535 42.190 ;
        RECT 238.385 41.620 238.675 41.900 ;
        RECT 280.245 41.620 280.535 41.900 ;
        RECT 238.385 41.330 280.535 41.620 ;
        RECT 330.700 52.170 372.850 52.460 ;
        RECT 330.700 42.190 330.990 52.170 ;
        RECT 335.280 51.560 370.030 51.890 ;
        RECT 331.395 42.380 331.675 51.410 ;
        RECT 332.275 42.380 332.555 51.410 ;
        RECT 333.155 42.380 333.435 51.410 ;
        RECT 334.035 42.380 334.315 51.410 ;
        RECT 334.915 42.380 335.195 51.410 ;
        RECT 335.795 42.380 336.075 51.410 ;
        RECT 336.675 42.380 336.955 51.410 ;
        RECT 337.555 42.380 337.835 51.410 ;
        RECT 338.435 42.380 338.715 51.410 ;
        RECT 339.315 42.380 339.595 51.410 ;
        RECT 340.195 42.380 340.475 51.410 ;
        RECT 341.075 42.380 341.355 51.410 ;
        RECT 341.955 42.380 342.235 51.410 ;
        RECT 342.835 42.380 343.115 51.410 ;
        RECT 343.715 42.380 343.995 51.410 ;
        RECT 344.595 42.380 344.875 51.410 ;
        RECT 345.475 42.380 345.755 51.410 ;
        RECT 346.355 42.380 346.635 51.410 ;
        RECT 347.235 42.380 347.515 51.410 ;
        RECT 348.115 42.380 348.395 51.410 ;
        RECT 348.995 42.380 349.275 51.410 ;
        RECT 349.875 42.380 350.155 51.410 ;
        RECT 350.755 42.380 351.035 51.410 ;
        RECT 351.635 42.380 351.915 51.410 ;
        RECT 352.515 42.380 352.795 51.410 ;
        RECT 353.395 42.380 353.675 51.410 ;
        RECT 354.275 42.380 354.555 51.410 ;
        RECT 355.155 42.380 355.435 51.410 ;
        RECT 356.035 42.380 356.315 51.410 ;
        RECT 356.915 42.380 357.195 51.410 ;
        RECT 357.795 42.380 358.075 51.410 ;
        RECT 358.675 42.380 358.955 51.410 ;
        RECT 359.555 42.380 359.835 51.410 ;
        RECT 360.435 42.380 360.715 51.410 ;
        RECT 361.315 42.380 361.595 51.410 ;
        RECT 362.195 42.380 362.475 51.410 ;
        RECT 363.075 42.380 363.355 51.410 ;
        RECT 363.955 42.380 364.235 51.410 ;
        RECT 364.835 42.380 365.115 51.410 ;
        RECT 365.715 42.380 365.995 51.410 ;
        RECT 366.595 42.380 366.875 51.410 ;
        RECT 367.475 42.380 367.755 51.410 ;
        RECT 368.355 42.380 368.635 51.410 ;
        RECT 369.235 42.380 369.515 51.410 ;
        RECT 370.115 42.380 370.395 51.410 ;
        RECT 370.995 42.380 371.275 51.410 ;
        RECT 371.875 42.380 372.155 51.410 ;
        RECT 372.560 42.190 372.850 52.170 ;
        RECT 330.700 41.900 334.830 42.190 ;
        RECT 370.480 41.900 372.850 42.190 ;
        RECT 330.700 41.620 330.990 41.900 ;
        RECT 372.560 41.620 372.850 41.900 ;
        RECT 330.700 41.330 372.850 41.620 ;
        RECT 373.360 52.170 403.190 52.460 ;
        RECT 373.360 42.190 373.650 52.170 ;
        RECT 377.940 51.560 398.610 51.890 ;
        RECT 374.055 42.380 374.335 51.410 ;
        RECT 374.935 42.380 375.215 51.410 ;
        RECT 375.815 42.380 376.095 51.410 ;
        RECT 376.695 42.380 376.975 51.410 ;
        RECT 377.575 42.380 377.855 51.410 ;
        RECT 378.455 42.380 378.735 51.410 ;
        RECT 379.335 42.380 379.615 51.410 ;
        RECT 380.215 42.380 380.495 51.410 ;
        RECT 381.095 42.380 381.375 51.410 ;
        RECT 381.975 42.380 382.255 51.410 ;
        RECT 382.855 42.380 383.135 51.410 ;
        RECT 383.735 42.380 384.015 51.410 ;
        RECT 384.615 42.380 384.895 51.410 ;
        RECT 385.495 42.380 385.775 51.410 ;
        RECT 386.375 42.380 386.655 51.410 ;
        RECT 387.255 42.380 387.535 51.410 ;
        RECT 388.135 42.380 388.415 51.410 ;
        RECT 389.015 42.380 389.295 51.410 ;
        RECT 389.895 42.380 390.175 51.410 ;
        RECT 390.775 42.380 391.055 51.410 ;
        RECT 391.655 42.380 391.935 51.410 ;
        RECT 392.535 42.380 392.815 51.410 ;
        RECT 393.415 42.380 393.695 51.410 ;
        RECT 394.295 42.380 394.575 51.410 ;
        RECT 395.175 42.380 395.455 51.410 ;
        RECT 396.055 42.380 396.335 51.410 ;
        RECT 396.935 42.380 397.215 51.410 ;
        RECT 397.815 42.380 398.095 51.410 ;
        RECT 398.695 42.380 398.975 51.410 ;
        RECT 399.575 42.380 399.855 51.410 ;
        RECT 400.455 42.380 400.735 51.410 ;
        RECT 401.335 42.380 401.615 51.410 ;
        RECT 402.215 42.380 402.495 51.410 ;
        RECT 402.900 42.190 403.190 52.170 ;
        RECT 373.360 41.900 377.490 42.190 ;
        RECT 399.060 41.900 403.190 42.190 ;
        RECT 373.360 41.620 373.650 41.900 ;
        RECT 402.900 41.620 403.190 41.900 ;
        RECT 373.360 41.330 403.190 41.620 ;
        RECT 208.045 39.805 237.875 40.095 ;
        RECT 208.045 39.525 208.335 39.805 ;
        RECT 237.585 39.525 237.875 39.805 ;
        RECT 208.045 39.235 213.935 39.525 ;
        RECT 221.425 39.235 224.495 39.525 ;
        RECT 231.985 39.235 237.875 39.525 ;
        RECT 184.785 36.960 207.655 37.250 ;
        RECT 184.785 36.130 185.075 36.960 ;
        RECT 185.885 36.430 189.695 36.720 ;
        RECT 189.405 36.130 189.695 36.430 ;
        RECT 202.745 36.430 206.555 36.720 ;
        RECT 202.745 36.130 203.035 36.430 ;
        RECT 207.365 36.130 207.655 36.960 ;
        RECT 184.785 35.840 188.955 36.130 ;
        RECT 189.405 35.840 203.035 36.130 ;
        RECT 203.485 35.840 207.655 36.130 ;
        RECT 184.785 33.200 185.075 35.840 ;
        RECT 185.520 33.390 185.800 35.650 ;
        RECT 186.400 33.390 186.680 35.650 ;
        RECT 187.280 33.390 187.560 35.650 ;
        RECT 188.160 33.390 188.440 35.650 ;
        RECT 189.040 33.390 189.320 35.650 ;
        RECT 189.920 33.390 190.200 35.650 ;
        RECT 190.800 33.390 191.080 35.650 ;
        RECT 191.680 33.390 191.960 35.650 ;
        RECT 192.560 33.390 192.840 35.650 ;
        RECT 193.440 33.390 193.720 35.650 ;
        RECT 194.320 33.390 194.600 35.650 ;
        RECT 195.200 33.390 195.480 35.650 ;
        RECT 196.080 33.390 196.360 35.650 ;
        RECT 196.960 33.390 197.240 35.650 ;
        RECT 197.840 33.390 198.120 35.650 ;
        RECT 198.720 33.390 199.000 35.650 ;
        RECT 199.600 33.390 199.880 35.650 ;
        RECT 200.480 33.390 200.760 35.650 ;
        RECT 201.360 33.390 201.640 35.650 ;
        RECT 202.240 33.390 202.520 35.650 ;
        RECT 203.120 33.390 203.400 35.650 ;
        RECT 204.000 33.390 204.280 35.650 ;
        RECT 204.880 33.390 205.160 35.650 ;
        RECT 205.760 33.390 206.040 35.650 ;
        RECT 206.640 33.390 206.920 35.650 ;
        RECT 207.365 33.200 207.655 35.840 ;
        RECT 184.785 32.910 188.955 33.200 ;
        RECT 189.405 32.910 203.035 33.200 ;
        RECT 203.485 32.910 207.655 33.200 ;
        RECT 184.785 32.075 185.075 32.910 ;
        RECT 189.405 32.610 189.695 32.910 ;
        RECT 185.885 32.320 189.695 32.610 ;
        RECT 202.745 32.610 203.035 32.910 ;
        RECT 202.745 32.320 206.555 32.610 ;
        RECT 207.365 32.075 207.655 32.910 ;
        RECT 184.785 31.785 207.655 32.075 ;
        RECT 208.045 29.255 208.335 39.235 ;
        RECT 208.740 30.015 209.020 39.045 ;
        RECT 209.620 30.015 209.900 39.045 ;
        RECT 210.500 30.015 210.780 39.045 ;
        RECT 211.380 30.015 211.660 39.045 ;
        RECT 212.260 30.015 212.540 39.045 ;
        RECT 213.140 30.015 213.420 39.045 ;
        RECT 214.020 30.015 214.300 39.045 ;
        RECT 214.900 30.015 215.180 39.045 ;
        RECT 215.780 30.015 216.060 39.045 ;
        RECT 216.660 30.015 216.940 39.045 ;
        RECT 217.540 30.015 217.820 39.045 ;
        RECT 218.420 30.015 218.700 39.045 ;
        RECT 219.300 30.015 219.580 39.045 ;
        RECT 220.180 30.015 220.460 39.045 ;
        RECT 221.060 30.015 221.340 39.045 ;
        RECT 221.940 30.015 222.220 39.235 ;
        RECT 222.820 30.015 223.100 39.235 ;
        RECT 223.700 30.015 223.980 39.235 ;
        RECT 224.580 30.015 224.860 39.045 ;
        RECT 225.460 30.015 225.740 39.045 ;
        RECT 226.340 30.015 226.620 39.045 ;
        RECT 227.220 30.015 227.500 39.045 ;
        RECT 228.100 30.015 228.380 39.045 ;
        RECT 228.980 30.015 229.260 39.045 ;
        RECT 229.860 30.015 230.140 39.045 ;
        RECT 230.740 30.015 231.020 39.045 ;
        RECT 231.620 30.015 231.900 39.045 ;
        RECT 232.500 30.015 232.780 39.045 ;
        RECT 233.380 30.015 233.660 39.045 ;
        RECT 234.260 30.015 234.540 39.045 ;
        RECT 235.140 30.015 235.420 39.045 ;
        RECT 236.020 30.015 236.300 39.045 ;
        RECT 236.900 30.015 237.180 39.045 ;
        RECT 214.385 29.495 220.975 29.825 ;
        RECT 224.945 29.535 231.590 29.825 ;
        RECT 225.000 29.495 231.590 29.535 ;
        RECT 237.585 29.255 237.875 39.235 ;
        RECT 208.045 28.965 237.875 29.255 ;
        RECT 238.385 39.805 280.535 40.095 ;
        RECT 238.385 39.525 238.675 39.805 ;
        RECT 280.245 39.525 280.535 39.805 ;
        RECT 238.385 39.235 240.755 39.525 ;
        RECT 276.405 39.235 280.535 39.525 ;
        RECT 238.385 29.255 238.675 39.235 ;
        RECT 239.080 30.015 239.360 39.045 ;
        RECT 239.960 30.015 240.240 39.045 ;
        RECT 240.840 30.015 241.120 39.045 ;
        RECT 241.720 30.015 242.000 39.045 ;
        RECT 242.600 30.015 242.880 39.045 ;
        RECT 243.480 30.015 243.760 39.045 ;
        RECT 244.360 30.015 244.640 39.045 ;
        RECT 245.240 30.015 245.520 39.045 ;
        RECT 246.120 30.015 246.400 39.045 ;
        RECT 247.000 30.015 247.280 39.045 ;
        RECT 247.880 30.015 248.160 39.045 ;
        RECT 248.760 30.015 249.040 39.045 ;
        RECT 249.640 30.015 249.920 39.045 ;
        RECT 250.520 30.015 250.800 39.045 ;
        RECT 251.400 30.015 251.680 39.045 ;
        RECT 252.280 30.015 252.560 39.045 ;
        RECT 253.160 30.015 253.440 39.045 ;
        RECT 254.040 30.015 254.320 39.045 ;
        RECT 254.920 30.015 255.200 39.045 ;
        RECT 255.800 30.015 256.080 39.045 ;
        RECT 256.680 30.015 256.960 39.045 ;
        RECT 257.560 30.015 257.840 39.045 ;
        RECT 258.440 30.015 258.720 39.045 ;
        RECT 259.320 30.015 259.600 39.045 ;
        RECT 260.200 30.015 260.480 39.045 ;
        RECT 261.080 30.015 261.360 39.045 ;
        RECT 261.960 30.015 262.240 39.045 ;
        RECT 262.840 30.015 263.120 39.045 ;
        RECT 263.720 30.015 264.000 39.045 ;
        RECT 264.600 30.015 264.880 39.045 ;
        RECT 265.480 30.015 265.760 39.045 ;
        RECT 266.360 30.015 266.640 39.045 ;
        RECT 267.240 30.015 267.520 39.045 ;
        RECT 268.120 30.015 268.400 39.045 ;
        RECT 269.000 30.015 269.280 39.045 ;
        RECT 269.880 30.015 270.160 39.045 ;
        RECT 270.760 30.015 271.040 39.045 ;
        RECT 271.640 30.015 271.920 39.045 ;
        RECT 272.520 30.015 272.800 39.045 ;
        RECT 273.400 30.015 273.680 39.045 ;
        RECT 274.280 30.015 274.560 39.045 ;
        RECT 275.160 30.015 275.440 39.045 ;
        RECT 276.040 30.015 276.320 39.045 ;
        RECT 276.920 30.015 277.200 39.045 ;
        RECT 277.800 30.015 278.080 39.045 ;
        RECT 278.680 30.015 278.960 39.045 ;
        RECT 279.560 30.015 279.840 39.045 ;
        RECT 241.205 29.495 275.955 29.825 ;
        RECT 280.245 29.255 280.535 39.235 ;
        RECT 238.385 28.965 280.535 29.255 ;
        RECT 330.700 39.805 372.850 40.095 ;
        RECT 330.700 39.525 330.990 39.805 ;
        RECT 372.560 39.525 372.850 39.805 ;
        RECT 330.700 39.235 334.830 39.525 ;
        RECT 370.480 39.235 372.850 39.525 ;
        RECT 330.700 29.255 330.990 39.235 ;
        RECT 331.395 30.015 331.675 39.045 ;
        RECT 332.275 30.015 332.555 39.045 ;
        RECT 333.155 30.015 333.435 39.045 ;
        RECT 334.035 30.015 334.315 39.045 ;
        RECT 334.915 30.015 335.195 39.045 ;
        RECT 335.795 30.015 336.075 39.045 ;
        RECT 336.675 30.015 336.955 39.045 ;
        RECT 337.555 30.015 337.835 39.045 ;
        RECT 338.435 30.015 338.715 39.045 ;
        RECT 339.315 30.015 339.595 39.045 ;
        RECT 340.195 30.015 340.475 39.045 ;
        RECT 341.075 30.015 341.355 39.045 ;
        RECT 341.955 30.015 342.235 39.045 ;
        RECT 342.835 30.015 343.115 39.045 ;
        RECT 343.715 30.015 343.995 39.045 ;
        RECT 344.595 30.015 344.875 39.045 ;
        RECT 345.475 30.015 345.755 39.045 ;
        RECT 346.355 30.015 346.635 39.045 ;
        RECT 347.235 30.015 347.515 39.045 ;
        RECT 348.115 30.015 348.395 39.045 ;
        RECT 348.995 30.015 349.275 39.045 ;
        RECT 349.875 30.015 350.155 39.045 ;
        RECT 350.755 30.015 351.035 39.045 ;
        RECT 351.635 30.015 351.915 39.045 ;
        RECT 352.515 30.015 352.795 39.045 ;
        RECT 353.395 30.015 353.675 39.045 ;
        RECT 354.275 30.015 354.555 39.045 ;
        RECT 355.155 30.015 355.435 39.045 ;
        RECT 356.035 30.015 356.315 39.045 ;
        RECT 356.915 30.015 357.195 39.045 ;
        RECT 357.795 30.015 358.075 39.045 ;
        RECT 358.675 30.015 358.955 39.045 ;
        RECT 359.555 30.015 359.835 39.045 ;
        RECT 360.435 30.015 360.715 39.045 ;
        RECT 361.315 30.015 361.595 39.045 ;
        RECT 362.195 30.015 362.475 39.045 ;
        RECT 363.075 30.015 363.355 39.045 ;
        RECT 363.955 30.015 364.235 39.045 ;
        RECT 364.835 30.015 365.115 39.045 ;
        RECT 365.715 30.015 365.995 39.045 ;
        RECT 366.595 30.015 366.875 39.045 ;
        RECT 367.475 30.015 367.755 39.045 ;
        RECT 368.355 30.015 368.635 39.045 ;
        RECT 369.235 30.015 369.515 39.045 ;
        RECT 370.115 30.015 370.395 39.045 ;
        RECT 370.995 30.015 371.275 39.045 ;
        RECT 371.875 30.015 372.155 39.045 ;
        RECT 335.280 29.495 370.030 29.825 ;
        RECT 372.560 29.255 372.850 39.235 ;
        RECT 330.700 28.965 372.850 29.255 ;
        RECT 373.360 39.805 403.190 40.095 ;
        RECT 373.360 39.525 373.650 39.805 ;
        RECT 402.900 39.525 403.190 39.805 ;
        RECT 373.360 39.235 379.250 39.525 ;
        RECT 386.740 39.235 389.810 39.525 ;
        RECT 397.300 39.235 403.190 39.525 ;
        RECT 373.360 29.255 373.650 39.235 ;
        RECT 374.055 30.015 374.335 39.045 ;
        RECT 374.935 30.015 375.215 39.045 ;
        RECT 375.815 30.015 376.095 39.045 ;
        RECT 376.695 30.015 376.975 39.045 ;
        RECT 377.575 30.015 377.855 39.045 ;
        RECT 378.455 30.015 378.735 39.045 ;
        RECT 379.335 30.015 379.615 39.045 ;
        RECT 380.215 30.015 380.495 39.045 ;
        RECT 381.095 30.015 381.375 39.045 ;
        RECT 381.975 30.015 382.255 39.045 ;
        RECT 382.855 30.015 383.135 39.045 ;
        RECT 383.735 30.015 384.015 39.045 ;
        RECT 384.615 30.015 384.895 39.045 ;
        RECT 385.495 30.015 385.775 39.045 ;
        RECT 386.375 30.015 386.655 39.045 ;
        RECT 387.255 30.015 387.535 39.235 ;
        RECT 388.135 30.015 388.415 39.235 ;
        RECT 389.015 30.015 389.295 39.235 ;
        RECT 389.895 30.015 390.175 39.045 ;
        RECT 390.775 30.015 391.055 39.045 ;
        RECT 391.655 30.015 391.935 39.045 ;
        RECT 392.535 30.015 392.815 39.045 ;
        RECT 393.415 30.015 393.695 39.045 ;
        RECT 394.295 30.015 394.575 39.045 ;
        RECT 395.175 30.015 395.455 39.045 ;
        RECT 396.055 30.015 396.335 39.045 ;
        RECT 396.935 30.015 397.215 39.045 ;
        RECT 397.815 30.015 398.095 39.045 ;
        RECT 398.695 30.015 398.975 39.045 ;
        RECT 399.575 30.015 399.855 39.045 ;
        RECT 400.455 30.015 400.735 39.045 ;
        RECT 401.335 30.015 401.615 39.045 ;
        RECT 402.215 30.015 402.495 39.045 ;
        RECT 379.645 29.535 386.290 29.825 ;
        RECT 379.645 29.495 386.235 29.535 ;
        RECT 390.260 29.495 396.850 29.825 ;
        RECT 402.900 29.255 403.190 39.235 ;
        RECT 403.580 36.960 426.450 37.250 ;
        RECT 403.580 36.130 403.870 36.960 ;
        RECT 404.680 36.430 408.490 36.720 ;
        RECT 408.200 36.130 408.490 36.430 ;
        RECT 421.540 36.430 425.350 36.720 ;
        RECT 421.540 36.130 421.830 36.430 ;
        RECT 426.160 36.130 426.450 36.960 ;
        RECT 403.580 35.840 407.750 36.130 ;
        RECT 408.200 35.840 421.830 36.130 ;
        RECT 422.280 35.840 426.450 36.130 ;
        RECT 403.580 33.200 403.870 35.840 ;
        RECT 404.315 33.390 404.595 35.650 ;
        RECT 405.195 33.390 405.475 35.650 ;
        RECT 406.075 33.390 406.355 35.650 ;
        RECT 406.955 33.390 407.235 35.650 ;
        RECT 407.835 33.390 408.115 35.650 ;
        RECT 408.715 33.390 408.995 35.650 ;
        RECT 409.595 33.390 409.875 35.650 ;
        RECT 410.475 33.390 410.755 35.650 ;
        RECT 411.355 33.390 411.635 35.650 ;
        RECT 412.235 33.390 412.515 35.650 ;
        RECT 413.115 33.390 413.395 35.650 ;
        RECT 413.995 33.390 414.275 35.650 ;
        RECT 414.875 33.390 415.155 35.650 ;
        RECT 415.755 33.390 416.035 35.650 ;
        RECT 416.635 33.390 416.915 35.650 ;
        RECT 417.515 33.390 417.795 35.650 ;
        RECT 418.395 33.390 418.675 35.650 ;
        RECT 419.275 33.390 419.555 35.650 ;
        RECT 420.155 33.390 420.435 35.650 ;
        RECT 421.035 33.390 421.315 35.650 ;
        RECT 421.915 33.390 422.195 35.650 ;
        RECT 422.795 33.390 423.075 35.650 ;
        RECT 423.675 33.390 423.955 35.650 ;
        RECT 424.555 33.390 424.835 35.650 ;
        RECT 425.435 33.390 425.715 35.650 ;
        RECT 426.160 33.200 426.450 35.840 ;
        RECT 403.580 32.910 407.750 33.200 ;
        RECT 408.200 32.910 421.830 33.200 ;
        RECT 422.280 32.910 426.450 33.200 ;
        RECT 403.580 32.075 403.870 32.910 ;
        RECT 408.200 32.610 408.490 32.910 ;
        RECT 404.680 32.320 408.490 32.610 ;
        RECT 421.540 32.610 421.830 32.910 ;
        RECT 421.540 32.320 425.350 32.610 ;
        RECT 426.160 32.075 426.450 32.910 ;
        RECT 403.580 31.785 426.450 32.075 ;
        RECT 373.360 28.965 403.190 29.255 ;
        RECT 184.785 27.880 207.655 28.170 ;
        RECT 184.785 27.520 185.075 27.880 ;
        RECT 207.365 27.520 207.655 27.880 ;
        RECT 184.785 27.230 192.475 27.520 ;
        RECT 199.965 27.230 207.655 27.520 ;
        RECT 184.785 23.940 185.075 27.230 ;
        RECT 185.520 24.780 185.800 27.040 ;
        RECT 186.400 24.780 186.680 27.040 ;
        RECT 187.280 24.780 187.560 27.040 ;
        RECT 188.160 24.780 188.440 27.040 ;
        RECT 189.040 24.780 189.320 27.040 ;
        RECT 189.920 24.780 190.200 27.040 ;
        RECT 190.800 24.780 191.080 27.040 ;
        RECT 191.680 24.780 191.960 27.040 ;
        RECT 192.560 24.780 192.840 27.040 ;
        RECT 193.440 24.780 193.720 27.040 ;
        RECT 194.320 24.780 194.600 27.040 ;
        RECT 195.200 24.780 195.480 27.040 ;
        RECT 196.080 24.780 196.360 27.040 ;
        RECT 196.960 24.780 197.240 27.040 ;
        RECT 197.840 24.780 198.120 27.040 ;
        RECT 198.720 24.780 199.000 27.040 ;
        RECT 199.600 24.780 199.880 27.040 ;
        RECT 200.480 24.780 200.760 27.040 ;
        RECT 201.360 24.780 201.640 27.040 ;
        RECT 202.240 24.780 202.520 27.040 ;
        RECT 203.120 24.780 203.400 27.040 ;
        RECT 204.000 24.780 204.280 27.040 ;
        RECT 204.880 24.780 205.160 27.040 ;
        RECT 205.760 24.780 206.040 27.040 ;
        RECT 206.640 24.780 206.920 27.040 ;
        RECT 192.905 24.260 199.515 24.590 ;
        RECT 207.365 23.940 207.655 27.230 ;
        RECT 184.785 23.650 207.655 23.940 ;
        RECT 208.005 27.880 237.915 28.170 ;
        RECT 208.005 27.520 208.295 27.880 ;
        RECT 237.625 27.520 237.915 27.880 ;
        RECT 208.005 27.230 213.935 27.520 ;
        RECT 221.425 27.230 224.495 27.520 ;
        RECT 231.985 27.230 237.915 27.520 ;
        RECT 208.005 23.940 208.295 27.230 ;
        RECT 208.740 24.780 209.020 27.040 ;
        RECT 209.620 24.780 209.900 27.040 ;
        RECT 210.500 24.780 210.780 27.040 ;
        RECT 211.380 24.780 211.660 27.040 ;
        RECT 212.260 24.780 212.540 27.040 ;
        RECT 213.140 24.780 213.420 27.040 ;
        RECT 214.020 24.780 214.300 27.040 ;
        RECT 214.900 24.780 215.180 27.040 ;
        RECT 215.780 24.780 216.060 27.040 ;
        RECT 216.660 24.780 216.940 27.040 ;
        RECT 217.540 24.780 217.820 27.040 ;
        RECT 218.420 24.780 218.700 27.040 ;
        RECT 219.300 24.780 219.580 27.040 ;
        RECT 220.180 24.780 220.460 27.040 ;
        RECT 221.060 24.780 221.340 27.040 ;
        RECT 221.940 24.780 222.220 27.230 ;
        RECT 222.820 24.780 223.100 27.230 ;
        RECT 223.700 24.780 223.980 27.230 ;
        RECT 224.580 24.780 224.860 27.040 ;
        RECT 225.460 24.780 225.740 27.040 ;
        RECT 226.340 24.780 226.620 27.040 ;
        RECT 227.220 24.780 227.500 27.040 ;
        RECT 228.100 24.780 228.380 27.040 ;
        RECT 228.980 24.780 229.260 27.040 ;
        RECT 229.860 24.780 230.140 27.040 ;
        RECT 230.740 24.780 231.020 27.040 ;
        RECT 231.620 24.780 231.900 27.040 ;
        RECT 232.500 24.780 232.780 27.040 ;
        RECT 233.380 24.780 233.660 27.040 ;
        RECT 234.260 24.780 234.540 27.040 ;
        RECT 235.140 24.780 235.420 27.040 ;
        RECT 236.020 24.780 236.300 27.040 ;
        RECT 236.900 24.780 237.180 27.040 ;
        RECT 211.660 24.260 231.535 24.590 ;
        RECT 237.625 23.940 237.915 27.230 ;
        RECT 208.005 23.650 237.915 23.940 ;
        RECT 238.345 27.880 280.570 28.170 ;
        RECT 238.345 27.520 238.635 27.880 ;
        RECT 280.280 27.520 280.570 27.880 ;
        RECT 238.345 27.230 240.755 27.520 ;
        RECT 276.405 27.230 280.570 27.520 ;
        RECT 238.345 23.940 238.635 27.230 ;
        RECT 239.080 24.780 239.360 27.040 ;
        RECT 239.960 24.780 240.240 27.040 ;
        RECT 240.840 24.780 241.120 27.040 ;
        RECT 241.720 24.780 242.000 27.040 ;
        RECT 242.600 24.780 242.880 27.040 ;
        RECT 243.480 24.780 243.760 27.040 ;
        RECT 244.360 24.780 244.640 27.040 ;
        RECT 245.240 24.780 245.520 27.040 ;
        RECT 246.120 24.780 246.400 27.040 ;
        RECT 247.000 24.780 247.280 27.040 ;
        RECT 247.880 24.780 248.160 27.040 ;
        RECT 248.760 24.780 249.040 27.040 ;
        RECT 249.640 24.780 249.920 27.040 ;
        RECT 250.520 24.780 250.800 27.040 ;
        RECT 251.400 24.780 251.680 27.040 ;
        RECT 252.280 24.780 252.560 27.040 ;
        RECT 253.160 24.780 253.440 27.040 ;
        RECT 254.040 24.780 254.320 27.040 ;
        RECT 254.920 24.780 255.200 27.040 ;
        RECT 255.800 24.780 256.080 27.040 ;
        RECT 256.680 24.780 256.960 27.040 ;
        RECT 257.560 24.780 257.840 27.040 ;
        RECT 258.440 24.780 258.720 27.040 ;
        RECT 259.320 24.780 259.600 27.040 ;
        RECT 260.200 24.780 260.480 27.040 ;
        RECT 261.080 24.780 261.360 27.040 ;
        RECT 261.960 24.780 262.240 27.040 ;
        RECT 262.840 24.780 263.120 27.040 ;
        RECT 263.720 24.780 264.000 27.040 ;
        RECT 264.600 24.780 264.880 27.040 ;
        RECT 265.480 24.780 265.760 27.040 ;
        RECT 266.360 24.780 266.640 27.040 ;
        RECT 267.240 24.780 267.520 27.040 ;
        RECT 268.120 24.780 268.400 27.040 ;
        RECT 269.000 24.780 269.280 27.040 ;
        RECT 269.880 24.780 270.160 27.040 ;
        RECT 270.760 24.780 271.040 27.040 ;
        RECT 271.640 24.780 271.920 27.040 ;
        RECT 272.520 24.780 272.800 27.040 ;
        RECT 273.400 24.780 273.680 27.040 ;
        RECT 274.280 24.780 274.560 27.040 ;
        RECT 275.160 24.780 275.440 27.040 ;
        RECT 276.040 24.780 276.320 27.040 ;
        RECT 276.920 24.780 277.200 27.040 ;
        RECT 277.800 24.780 278.080 27.040 ;
        RECT 278.680 24.780 278.960 27.040 ;
        RECT 279.560 24.780 279.840 27.040 ;
        RECT 280.280 26.410 280.570 27.230 ;
        RECT 330.665 27.880 372.890 28.170 ;
        RECT 330.665 27.520 330.955 27.880 ;
        RECT 372.600 27.520 372.890 27.880 ;
        RECT 330.665 27.230 334.830 27.520 ;
        RECT 370.480 27.230 372.890 27.520 ;
        RECT 330.665 26.410 330.955 27.230 ;
        RECT 280.280 25.410 280.575 26.410 ;
        RECT 330.660 25.410 330.955 26.410 ;
        RECT 239.175 24.260 275.955 24.590 ;
        RECT 280.280 23.940 280.570 25.410 ;
        RECT 238.345 23.650 280.570 23.940 ;
        RECT 330.665 23.940 330.955 25.410 ;
        RECT 331.395 24.780 331.675 27.040 ;
        RECT 332.275 24.780 332.555 27.040 ;
        RECT 333.155 24.780 333.435 27.040 ;
        RECT 334.035 24.780 334.315 27.040 ;
        RECT 334.915 24.780 335.195 27.040 ;
        RECT 335.795 24.780 336.075 27.040 ;
        RECT 336.675 24.780 336.955 27.040 ;
        RECT 337.555 24.780 337.835 27.040 ;
        RECT 338.435 24.780 338.715 27.040 ;
        RECT 339.315 24.780 339.595 27.040 ;
        RECT 340.195 24.780 340.475 27.040 ;
        RECT 341.075 24.780 341.355 27.040 ;
        RECT 341.955 24.780 342.235 27.040 ;
        RECT 342.835 24.780 343.115 27.040 ;
        RECT 343.715 24.780 343.995 27.040 ;
        RECT 344.595 24.780 344.875 27.040 ;
        RECT 345.475 24.780 345.755 27.040 ;
        RECT 346.355 24.780 346.635 27.040 ;
        RECT 347.235 24.780 347.515 27.040 ;
        RECT 348.115 24.780 348.395 27.040 ;
        RECT 348.995 24.780 349.275 27.040 ;
        RECT 349.875 24.780 350.155 27.040 ;
        RECT 350.755 24.780 351.035 27.040 ;
        RECT 351.635 24.780 351.915 27.040 ;
        RECT 352.515 24.780 352.795 27.040 ;
        RECT 353.395 24.780 353.675 27.040 ;
        RECT 354.275 24.780 354.555 27.040 ;
        RECT 355.155 24.780 355.435 27.040 ;
        RECT 356.035 24.780 356.315 27.040 ;
        RECT 356.915 24.780 357.195 27.040 ;
        RECT 357.795 24.780 358.075 27.040 ;
        RECT 358.675 24.780 358.955 27.040 ;
        RECT 359.555 24.780 359.835 27.040 ;
        RECT 360.435 24.780 360.715 27.040 ;
        RECT 361.315 24.780 361.595 27.040 ;
        RECT 362.195 24.780 362.475 27.040 ;
        RECT 363.075 24.780 363.355 27.040 ;
        RECT 363.955 24.780 364.235 27.040 ;
        RECT 364.835 24.780 365.115 27.040 ;
        RECT 365.715 24.780 365.995 27.040 ;
        RECT 366.595 24.780 366.875 27.040 ;
        RECT 367.475 24.780 367.755 27.040 ;
        RECT 368.355 24.780 368.635 27.040 ;
        RECT 369.235 24.780 369.515 27.040 ;
        RECT 370.115 24.780 370.395 27.040 ;
        RECT 370.995 24.780 371.275 27.040 ;
        RECT 371.875 24.780 372.155 27.040 ;
        RECT 335.280 24.260 372.060 24.590 ;
        RECT 372.600 23.940 372.890 27.230 ;
        RECT 330.665 23.650 372.890 23.940 ;
        RECT 373.320 27.880 403.230 28.170 ;
        RECT 373.320 27.520 373.610 27.880 ;
        RECT 402.940 27.520 403.230 27.880 ;
        RECT 373.320 27.230 379.250 27.520 ;
        RECT 386.740 27.230 389.810 27.520 ;
        RECT 397.300 27.230 403.230 27.520 ;
        RECT 373.320 23.940 373.610 27.230 ;
        RECT 374.055 24.780 374.335 27.040 ;
        RECT 374.935 24.780 375.215 27.040 ;
        RECT 375.815 24.780 376.095 27.040 ;
        RECT 376.695 24.780 376.975 27.040 ;
        RECT 377.575 24.780 377.855 27.040 ;
        RECT 378.455 24.780 378.735 27.040 ;
        RECT 379.335 24.780 379.615 27.040 ;
        RECT 380.215 24.780 380.495 27.040 ;
        RECT 381.095 24.780 381.375 27.040 ;
        RECT 381.975 24.780 382.255 27.040 ;
        RECT 382.855 24.780 383.135 27.040 ;
        RECT 383.735 24.780 384.015 27.040 ;
        RECT 384.615 24.780 384.895 27.040 ;
        RECT 385.495 24.780 385.775 27.040 ;
        RECT 386.375 24.780 386.655 27.040 ;
        RECT 387.255 24.780 387.535 27.230 ;
        RECT 388.135 24.780 388.415 27.230 ;
        RECT 389.015 24.780 389.295 27.230 ;
        RECT 389.895 24.780 390.175 27.040 ;
        RECT 390.775 24.780 391.055 27.040 ;
        RECT 391.655 24.780 391.935 27.040 ;
        RECT 392.535 24.780 392.815 27.040 ;
        RECT 393.415 24.780 393.695 27.040 ;
        RECT 394.295 24.780 394.575 27.040 ;
        RECT 395.175 24.780 395.455 27.040 ;
        RECT 396.055 24.780 396.335 27.040 ;
        RECT 396.935 24.780 397.215 27.040 ;
        RECT 397.815 24.780 398.095 27.040 ;
        RECT 398.695 24.780 398.975 27.040 ;
        RECT 399.575 24.780 399.855 27.040 ;
        RECT 400.455 24.780 400.735 27.040 ;
        RECT 401.335 24.780 401.615 27.040 ;
        RECT 402.215 24.780 402.495 27.040 ;
        RECT 379.700 24.260 399.575 24.590 ;
        RECT 402.940 23.940 403.230 27.230 ;
        RECT 373.320 23.650 403.230 23.940 ;
        RECT 403.580 27.880 426.450 28.170 ;
        RECT 403.580 27.520 403.870 27.880 ;
        RECT 426.160 27.520 426.450 27.880 ;
        RECT 403.580 27.230 411.270 27.520 ;
        RECT 418.760 27.230 426.450 27.520 ;
        RECT 403.580 23.940 403.870 27.230 ;
        RECT 404.315 24.780 404.595 27.040 ;
        RECT 405.195 24.780 405.475 27.040 ;
        RECT 406.075 24.780 406.355 27.040 ;
        RECT 406.955 24.780 407.235 27.040 ;
        RECT 407.835 24.780 408.115 27.040 ;
        RECT 408.715 24.780 408.995 27.040 ;
        RECT 409.595 24.780 409.875 27.040 ;
        RECT 410.475 24.780 410.755 27.040 ;
        RECT 411.355 24.780 411.635 27.040 ;
        RECT 412.235 24.780 412.515 27.040 ;
        RECT 413.115 24.780 413.395 27.040 ;
        RECT 413.995 24.780 414.275 27.040 ;
        RECT 414.875 24.780 415.155 27.040 ;
        RECT 415.755 24.780 416.035 27.040 ;
        RECT 416.635 24.780 416.915 27.040 ;
        RECT 417.515 24.780 417.795 27.040 ;
        RECT 418.395 24.780 418.675 27.040 ;
        RECT 419.275 24.780 419.555 27.040 ;
        RECT 420.155 24.780 420.435 27.040 ;
        RECT 421.035 24.780 421.315 27.040 ;
        RECT 421.915 24.780 422.195 27.040 ;
        RECT 422.795 24.780 423.075 27.040 ;
        RECT 423.675 24.780 423.955 27.040 ;
        RECT 424.555 24.780 424.835 27.040 ;
        RECT 425.435 24.780 425.715 27.040 ;
        RECT 411.720 24.260 418.330 24.590 ;
        RECT 426.160 23.940 426.450 27.230 ;
        RECT 403.580 23.650 426.450 23.940 ;
        RECT 184.785 21.395 207.655 21.685 ;
        RECT 184.785 21.035 185.075 21.395 ;
        RECT 207.365 21.035 207.655 21.395 ;
        RECT 184.785 20.745 192.475 21.035 ;
        RECT 199.965 20.745 207.655 21.035 ;
        RECT 184.785 17.455 185.075 20.745 ;
        RECT 185.520 18.295 185.800 20.555 ;
        RECT 186.400 18.295 186.680 20.555 ;
        RECT 187.280 18.295 187.560 20.555 ;
        RECT 188.160 18.295 188.440 20.555 ;
        RECT 189.040 18.295 189.320 20.555 ;
        RECT 189.920 18.295 190.200 20.555 ;
        RECT 190.800 18.295 191.080 20.555 ;
        RECT 191.680 18.295 191.960 20.555 ;
        RECT 192.560 18.295 192.840 20.555 ;
        RECT 193.440 18.295 193.720 20.555 ;
        RECT 194.320 18.295 194.600 20.555 ;
        RECT 195.200 18.295 195.480 20.555 ;
        RECT 196.080 18.295 196.360 20.555 ;
        RECT 196.960 18.295 197.240 20.555 ;
        RECT 197.840 18.295 198.120 20.555 ;
        RECT 198.720 18.295 199.000 20.555 ;
        RECT 199.600 18.295 199.880 20.555 ;
        RECT 200.480 18.295 200.760 20.555 ;
        RECT 201.360 18.295 201.640 20.555 ;
        RECT 202.240 18.295 202.520 20.555 ;
        RECT 203.120 18.295 203.400 20.555 ;
        RECT 204.000 18.295 204.280 20.555 ;
        RECT 204.880 18.295 205.160 20.555 ;
        RECT 205.760 18.295 206.040 20.555 ;
        RECT 206.640 18.295 206.920 20.555 ;
        RECT 192.925 17.775 199.515 18.105 ;
        RECT 207.365 17.455 207.655 20.745 ;
        RECT 184.785 17.165 207.655 17.455 ;
        RECT 208.005 21.395 237.915 21.685 ;
        RECT 208.005 21.035 208.295 21.395 ;
        RECT 237.625 21.035 237.915 21.395 ;
        RECT 208.005 20.745 213.935 21.035 ;
        RECT 214.385 20.745 231.535 21.035 ;
        RECT 231.985 20.745 237.915 21.035 ;
        RECT 208.005 17.455 208.295 20.745 ;
        RECT 208.740 18.295 209.020 20.555 ;
        RECT 209.620 18.295 209.900 20.555 ;
        RECT 210.500 18.295 210.780 20.555 ;
        RECT 211.380 18.295 211.660 20.555 ;
        RECT 212.260 18.295 212.540 20.555 ;
        RECT 213.140 18.295 213.420 20.555 ;
        RECT 214.020 18.295 214.300 20.555 ;
        RECT 214.900 18.295 215.180 20.555 ;
        RECT 215.780 18.295 216.060 20.555 ;
        RECT 216.660 18.295 216.940 20.555 ;
        RECT 217.540 18.295 217.820 20.555 ;
        RECT 218.420 18.295 218.700 20.555 ;
        RECT 219.300 18.295 219.580 20.555 ;
        RECT 220.180 18.295 220.460 20.555 ;
        RECT 221.060 18.295 221.340 20.555 ;
        RECT 221.940 18.105 222.220 20.555 ;
        RECT 222.820 18.295 223.100 20.555 ;
        RECT 223.700 18.105 223.980 20.555 ;
        RECT 224.580 18.295 224.860 20.555 ;
        RECT 225.460 18.295 225.740 20.555 ;
        RECT 226.340 18.295 226.620 20.555 ;
        RECT 227.220 18.295 227.500 20.555 ;
        RECT 228.100 18.295 228.380 20.555 ;
        RECT 228.980 18.295 229.260 20.555 ;
        RECT 229.860 18.295 230.140 20.555 ;
        RECT 230.740 18.295 231.020 20.555 ;
        RECT 231.620 18.295 231.900 20.555 ;
        RECT 232.500 18.295 232.780 20.555 ;
        RECT 233.380 18.295 233.660 20.555 ;
        RECT 234.260 18.295 234.540 20.555 ;
        RECT 235.140 18.295 235.420 20.555 ;
        RECT 236.020 18.295 236.300 20.555 ;
        RECT 236.900 18.295 237.180 20.555 ;
        RECT 221.425 17.815 224.495 18.105 ;
        RECT 237.625 17.455 237.915 20.745 ;
        RECT 208.005 17.165 237.915 17.455 ;
        RECT 238.345 21.395 280.570 21.685 ;
        RECT 238.345 21.035 238.635 21.395 ;
        RECT 280.280 21.035 280.570 21.395 ;
        RECT 238.345 20.745 240.755 21.035 ;
        RECT 241.205 20.745 275.955 21.035 ;
        RECT 276.405 20.745 280.570 21.035 ;
        RECT 238.345 17.455 238.635 20.745 ;
        RECT 239.080 18.295 239.360 20.555 ;
        RECT 239.960 18.295 240.240 20.555 ;
        RECT 240.840 18.295 241.120 20.555 ;
        RECT 241.720 18.295 242.000 20.555 ;
        RECT 242.600 18.295 242.880 20.555 ;
        RECT 243.480 18.295 243.760 20.555 ;
        RECT 244.360 18.295 244.640 20.555 ;
        RECT 245.240 18.295 245.520 20.555 ;
        RECT 246.120 18.295 246.400 20.555 ;
        RECT 247.000 18.295 247.280 20.555 ;
        RECT 247.880 18.295 248.160 20.555 ;
        RECT 248.760 18.295 249.040 20.555 ;
        RECT 249.640 18.295 249.920 20.555 ;
        RECT 250.520 18.295 250.800 20.555 ;
        RECT 251.400 18.295 251.680 20.555 ;
        RECT 252.280 18.295 252.560 20.555 ;
        RECT 253.160 18.295 253.440 20.555 ;
        RECT 254.040 18.295 254.320 20.555 ;
        RECT 254.920 18.295 255.200 20.555 ;
        RECT 255.800 18.295 256.080 20.555 ;
        RECT 256.680 18.295 256.960 20.555 ;
        RECT 257.560 18.295 257.840 20.555 ;
        RECT 258.440 18.295 258.720 20.555 ;
        RECT 259.320 18.295 259.600 20.555 ;
        RECT 260.200 18.295 260.480 20.555 ;
        RECT 261.080 18.295 261.360 20.555 ;
        RECT 261.960 18.295 262.240 20.555 ;
        RECT 262.840 18.295 263.120 20.555 ;
        RECT 263.720 18.295 264.000 20.555 ;
        RECT 264.600 18.295 264.880 20.555 ;
        RECT 265.480 18.295 265.760 20.555 ;
        RECT 266.360 18.295 266.640 20.555 ;
        RECT 267.240 18.295 267.520 20.555 ;
        RECT 268.120 18.295 268.400 20.555 ;
        RECT 269.000 18.295 269.280 20.555 ;
        RECT 269.880 18.295 270.160 20.555 ;
        RECT 270.760 18.295 271.040 20.555 ;
        RECT 271.640 18.295 271.920 20.555 ;
        RECT 272.520 18.295 272.800 20.555 ;
        RECT 273.400 18.295 273.680 20.555 ;
        RECT 274.280 18.295 274.560 20.555 ;
        RECT 275.160 18.295 275.440 20.555 ;
        RECT 276.040 18.295 276.320 20.555 ;
        RECT 276.920 18.295 277.200 20.555 ;
        RECT 277.800 18.295 278.080 20.555 ;
        RECT 278.680 18.295 278.960 20.555 ;
        RECT 279.560 18.295 279.840 20.555 ;
        RECT 280.280 19.925 280.570 20.745 ;
        RECT 330.665 21.395 372.890 21.685 ;
        RECT 330.665 21.035 330.955 21.395 ;
        RECT 372.600 21.035 372.890 21.395 ;
        RECT 330.665 20.745 334.830 21.035 ;
        RECT 335.280 20.745 370.030 21.035 ;
        RECT 370.480 20.745 372.890 21.035 ;
        RECT 330.665 19.925 330.955 20.745 ;
        RECT 280.280 18.925 280.575 19.925 ;
        RECT 330.660 18.925 330.955 19.925 ;
        RECT 280.280 17.455 280.570 18.925 ;
        RECT 238.345 17.165 280.570 17.455 ;
        RECT 330.665 17.455 330.955 18.925 ;
        RECT 331.395 18.295 331.675 20.555 ;
        RECT 332.275 18.295 332.555 20.555 ;
        RECT 333.155 18.295 333.435 20.555 ;
        RECT 334.035 18.295 334.315 20.555 ;
        RECT 334.915 18.295 335.195 20.555 ;
        RECT 335.795 18.295 336.075 20.555 ;
        RECT 336.675 18.295 336.955 20.555 ;
        RECT 337.555 18.295 337.835 20.555 ;
        RECT 338.435 18.295 338.715 20.555 ;
        RECT 339.315 18.295 339.595 20.555 ;
        RECT 340.195 18.295 340.475 20.555 ;
        RECT 341.075 18.295 341.355 20.555 ;
        RECT 341.955 18.295 342.235 20.555 ;
        RECT 342.835 18.295 343.115 20.555 ;
        RECT 343.715 18.295 343.995 20.555 ;
        RECT 344.595 18.295 344.875 20.555 ;
        RECT 345.475 18.295 345.755 20.555 ;
        RECT 346.355 18.295 346.635 20.555 ;
        RECT 347.235 18.295 347.515 20.555 ;
        RECT 348.115 18.295 348.395 20.555 ;
        RECT 348.995 18.295 349.275 20.555 ;
        RECT 349.875 18.295 350.155 20.555 ;
        RECT 350.755 18.295 351.035 20.555 ;
        RECT 351.635 18.295 351.915 20.555 ;
        RECT 352.515 18.295 352.795 20.555 ;
        RECT 353.395 18.295 353.675 20.555 ;
        RECT 354.275 18.295 354.555 20.555 ;
        RECT 355.155 18.295 355.435 20.555 ;
        RECT 356.035 18.295 356.315 20.555 ;
        RECT 356.915 18.295 357.195 20.555 ;
        RECT 357.795 18.295 358.075 20.555 ;
        RECT 358.675 18.295 358.955 20.555 ;
        RECT 359.555 18.295 359.835 20.555 ;
        RECT 360.435 18.295 360.715 20.555 ;
        RECT 361.315 18.295 361.595 20.555 ;
        RECT 362.195 18.295 362.475 20.555 ;
        RECT 363.075 18.295 363.355 20.555 ;
        RECT 363.955 18.295 364.235 20.555 ;
        RECT 364.835 18.295 365.115 20.555 ;
        RECT 365.715 18.295 365.995 20.555 ;
        RECT 366.595 18.295 366.875 20.555 ;
        RECT 367.475 18.295 367.755 20.555 ;
        RECT 368.355 18.295 368.635 20.555 ;
        RECT 369.235 18.295 369.515 20.555 ;
        RECT 370.115 18.295 370.395 20.555 ;
        RECT 370.995 18.295 371.275 20.555 ;
        RECT 371.875 18.295 372.155 20.555 ;
        RECT 372.600 17.455 372.890 20.745 ;
        RECT 330.665 17.165 372.890 17.455 ;
        RECT 373.320 21.395 403.230 21.685 ;
        RECT 373.320 21.035 373.610 21.395 ;
        RECT 402.940 21.035 403.230 21.395 ;
        RECT 373.320 20.745 379.250 21.035 ;
        RECT 379.700 20.745 396.850 21.035 ;
        RECT 397.300 20.745 403.230 21.035 ;
        RECT 373.320 17.455 373.610 20.745 ;
        RECT 374.055 18.295 374.335 20.555 ;
        RECT 374.935 18.295 375.215 20.555 ;
        RECT 375.815 18.295 376.095 20.555 ;
        RECT 376.695 18.295 376.975 20.555 ;
        RECT 377.575 18.295 377.855 20.555 ;
        RECT 378.455 18.295 378.735 20.555 ;
        RECT 379.335 18.295 379.615 20.555 ;
        RECT 380.215 18.295 380.495 20.555 ;
        RECT 381.095 18.295 381.375 20.555 ;
        RECT 381.975 18.295 382.255 20.555 ;
        RECT 382.855 18.295 383.135 20.555 ;
        RECT 383.735 18.295 384.015 20.555 ;
        RECT 384.615 18.295 384.895 20.555 ;
        RECT 385.495 18.295 385.775 20.555 ;
        RECT 386.375 18.295 386.655 20.555 ;
        RECT 387.255 18.105 387.535 20.555 ;
        RECT 388.135 18.295 388.415 20.555 ;
        RECT 389.015 18.105 389.295 20.555 ;
        RECT 389.895 18.295 390.175 20.555 ;
        RECT 390.775 18.295 391.055 20.555 ;
        RECT 391.655 18.295 391.935 20.555 ;
        RECT 392.535 18.295 392.815 20.555 ;
        RECT 393.415 18.295 393.695 20.555 ;
        RECT 394.295 18.295 394.575 20.555 ;
        RECT 395.175 18.295 395.455 20.555 ;
        RECT 396.055 18.295 396.335 20.555 ;
        RECT 396.935 18.295 397.215 20.555 ;
        RECT 397.815 18.295 398.095 20.555 ;
        RECT 398.695 18.295 398.975 20.555 ;
        RECT 399.575 18.295 399.855 20.555 ;
        RECT 400.455 18.295 400.735 20.555 ;
        RECT 401.335 18.295 401.615 20.555 ;
        RECT 402.215 18.295 402.495 20.555 ;
        RECT 386.740 17.815 389.810 18.105 ;
        RECT 402.940 17.455 403.230 20.745 ;
        RECT 373.320 17.165 403.230 17.455 ;
        RECT 403.580 21.395 426.450 21.685 ;
        RECT 403.580 21.035 403.870 21.395 ;
        RECT 426.160 21.035 426.450 21.395 ;
        RECT 403.580 20.745 411.270 21.035 ;
        RECT 418.760 20.745 426.450 21.035 ;
        RECT 403.580 17.455 403.870 20.745 ;
        RECT 404.315 18.295 404.595 20.555 ;
        RECT 405.195 18.295 405.475 20.555 ;
        RECT 406.075 18.295 406.355 20.555 ;
        RECT 406.955 18.295 407.235 20.555 ;
        RECT 407.835 18.295 408.115 20.555 ;
        RECT 408.715 18.295 408.995 20.555 ;
        RECT 409.595 18.295 409.875 20.555 ;
        RECT 410.475 18.295 410.755 20.555 ;
        RECT 411.355 18.295 411.635 20.555 ;
        RECT 412.235 18.295 412.515 20.555 ;
        RECT 413.115 18.295 413.395 20.555 ;
        RECT 413.995 18.295 414.275 20.555 ;
        RECT 414.875 18.295 415.155 20.555 ;
        RECT 415.755 18.295 416.035 20.555 ;
        RECT 416.635 18.295 416.915 20.555 ;
        RECT 417.515 18.295 417.795 20.555 ;
        RECT 418.395 18.295 418.675 20.555 ;
        RECT 419.275 18.295 419.555 20.555 ;
        RECT 420.155 18.295 420.435 20.555 ;
        RECT 421.035 18.295 421.315 20.555 ;
        RECT 421.915 18.295 422.195 20.555 ;
        RECT 422.795 18.295 423.075 20.555 ;
        RECT 423.675 18.295 423.955 20.555 ;
        RECT 424.555 18.295 424.835 20.555 ;
        RECT 425.435 18.295 425.715 20.555 ;
        RECT 411.720 17.775 418.310 18.105 ;
        RECT 426.160 17.455 426.450 20.745 ;
        RECT 403.580 17.165 426.450 17.455 ;
      LAYER met2 ;
        RECT 180.600 216.490 181.680 217.090 ;
        RECT 179.500 214.890 180.580 215.490 ;
        RECT 73.400 210.510 74.570 210.840 ;
        RECT 73.820 187.020 74.150 210.510 ;
        RECT 78.970 208.755 113.740 209.085 ;
        RECT 121.590 208.755 142.360 209.085 ;
        RECT 170.620 208.755 171.790 209.085 ;
        RECT 74.400 203.085 74.690 205.085 ;
        RECT 75.095 203.085 75.375 205.085 ;
        RECT 75.975 203.085 76.255 205.085 ;
        RECT 76.855 203.085 77.135 205.085 ;
        RECT 77.735 203.085 78.015 205.085 ;
        RECT 78.615 203.085 78.895 205.085 ;
        RECT 79.495 198.305 79.775 208.605 ;
        RECT 80.375 203.085 80.655 205.085 ;
        RECT 81.255 198.305 81.535 208.605 ;
        RECT 82.135 203.085 82.415 205.085 ;
        RECT 83.015 198.305 83.295 208.605 ;
        RECT 83.895 203.085 84.175 205.085 ;
        RECT 84.775 198.305 85.055 208.605 ;
        RECT 85.655 203.085 85.935 205.085 ;
        RECT 86.535 198.305 86.815 208.605 ;
        RECT 87.415 203.085 87.695 205.085 ;
        RECT 88.295 198.305 88.575 208.605 ;
        RECT 89.175 203.085 89.455 205.085 ;
        RECT 90.055 198.305 90.335 208.605 ;
        RECT 90.935 203.085 91.215 205.085 ;
        RECT 91.815 198.305 92.095 208.605 ;
        RECT 92.695 203.085 92.975 205.085 ;
        RECT 93.575 198.305 93.855 208.605 ;
        RECT 94.455 203.085 94.735 205.085 ;
        RECT 95.335 198.305 95.615 208.605 ;
        RECT 96.215 203.085 96.495 205.085 ;
        RECT 97.095 198.305 97.375 208.605 ;
        RECT 97.975 203.085 98.255 205.085 ;
        RECT 98.855 198.305 99.135 208.605 ;
        RECT 99.735 203.085 100.015 205.085 ;
        RECT 100.615 198.305 100.895 208.605 ;
        RECT 101.495 203.085 101.775 205.085 ;
        RECT 102.375 198.305 102.655 208.605 ;
        RECT 103.255 203.085 103.535 205.085 ;
        RECT 104.135 198.305 104.415 208.605 ;
        RECT 105.015 203.085 105.295 205.085 ;
        RECT 105.895 198.305 106.175 208.605 ;
        RECT 106.775 203.085 107.055 205.085 ;
        RECT 107.655 198.305 107.935 208.605 ;
        RECT 108.535 203.085 108.815 205.085 ;
        RECT 109.415 198.305 109.695 208.605 ;
        RECT 110.295 203.085 110.575 205.085 ;
        RECT 111.175 198.305 111.455 208.605 ;
        RECT 112.055 203.085 112.335 205.085 ;
        RECT 112.935 198.305 113.215 208.605 ;
        RECT 113.815 203.085 114.095 205.085 ;
        RECT 114.695 203.085 114.975 205.085 ;
        RECT 115.575 203.085 115.855 205.085 ;
        RECT 116.260 203.085 116.550 205.085 ;
        RECT 117.060 203.085 117.350 205.085 ;
        RECT 117.755 203.085 118.035 205.085 ;
        RECT 118.635 203.085 118.915 205.085 ;
        RECT 119.515 203.085 119.795 205.085 ;
        RECT 120.395 203.085 120.675 205.085 ;
        RECT 121.275 203.085 121.555 205.085 ;
        RECT 122.155 198.420 122.435 208.605 ;
        RECT 123.035 203.085 123.315 205.085 ;
        RECT 123.915 198.420 124.195 208.605 ;
        RECT 124.795 203.085 125.075 205.085 ;
        RECT 125.675 198.420 125.955 208.605 ;
        RECT 126.555 203.085 126.835 205.085 ;
        RECT 127.435 198.420 127.715 208.605 ;
        RECT 128.315 203.085 128.595 205.085 ;
        RECT 129.195 198.420 129.475 208.605 ;
        RECT 130.075 203.085 130.355 205.085 ;
        RECT 130.955 198.420 131.235 208.605 ;
        RECT 131.835 203.085 132.115 205.085 ;
        RECT 79.495 197.505 113.215 198.305 ;
        RECT 121.955 198.050 122.635 198.420 ;
        RECT 123.715 198.050 124.395 198.420 ;
        RECT 125.475 198.050 126.155 198.420 ;
        RECT 127.235 198.050 127.915 198.420 ;
        RECT 128.995 198.050 129.675 198.420 ;
        RECT 130.755 198.050 131.435 198.420 ;
        RECT 74.400 190.725 74.690 192.725 ;
        RECT 75.095 190.725 75.375 192.725 ;
        RECT 75.975 190.725 76.255 192.725 ;
        RECT 76.855 190.725 77.135 192.725 ;
        RECT 77.735 190.725 78.015 192.725 ;
        RECT 73.820 186.690 74.990 187.020 ;
        RECT 78.615 186.165 78.895 196.240 ;
        RECT 79.495 187.210 79.775 197.505 ;
        RECT 79.185 186.690 80.035 187.020 ;
        RECT 80.375 186.165 80.655 196.240 ;
        RECT 81.255 187.210 81.535 197.505 ;
        RECT 80.795 186.690 81.995 187.020 ;
        RECT 82.135 186.165 82.415 196.240 ;
        RECT 83.015 187.210 83.295 197.505 ;
        RECT 82.555 186.690 83.755 187.020 ;
        RECT 83.895 186.165 84.175 196.240 ;
        RECT 84.775 187.210 85.055 197.505 ;
        RECT 84.315 186.690 85.515 187.020 ;
        RECT 85.655 186.165 85.935 196.240 ;
        RECT 86.535 187.210 86.815 197.505 ;
        RECT 86.075 186.690 87.275 187.020 ;
        RECT 87.415 186.165 87.695 196.240 ;
        RECT 88.295 187.210 88.575 197.505 ;
        RECT 87.835 186.690 89.035 187.020 ;
        RECT 89.175 186.165 89.455 196.240 ;
        RECT 90.055 187.210 90.335 197.505 ;
        RECT 89.595 186.690 90.795 187.020 ;
        RECT 90.935 186.165 91.215 196.240 ;
        RECT 91.815 187.210 92.095 197.505 ;
        RECT 91.355 186.690 92.555 187.020 ;
        RECT 92.695 186.165 92.975 196.240 ;
        RECT 93.575 187.210 93.855 197.505 ;
        RECT 93.115 186.690 94.315 187.020 ;
        RECT 94.455 186.165 94.735 196.240 ;
        RECT 95.335 187.210 95.615 197.505 ;
        RECT 94.875 186.690 96.075 187.020 ;
        RECT 96.215 186.165 96.495 196.240 ;
        RECT 97.095 187.210 97.375 197.505 ;
        RECT 96.635 186.690 97.835 187.020 ;
        RECT 97.975 186.165 98.255 196.240 ;
        RECT 98.855 187.210 99.135 197.505 ;
        RECT 98.395 186.690 99.595 187.020 ;
        RECT 99.735 186.165 100.015 196.240 ;
        RECT 100.615 187.210 100.895 197.505 ;
        RECT 100.155 186.690 101.355 187.020 ;
        RECT 101.495 186.165 101.775 196.240 ;
        RECT 102.375 187.210 102.655 197.505 ;
        RECT 101.915 186.690 103.115 187.020 ;
        RECT 103.255 186.165 103.535 196.240 ;
        RECT 104.135 187.210 104.415 197.505 ;
        RECT 103.675 186.690 104.875 187.020 ;
        RECT 105.015 186.165 105.295 196.240 ;
        RECT 105.895 187.210 106.175 197.505 ;
        RECT 105.435 186.690 106.635 187.020 ;
        RECT 106.775 186.165 107.055 196.240 ;
        RECT 107.655 187.210 107.935 197.505 ;
        RECT 107.195 186.690 108.395 187.020 ;
        RECT 108.535 186.165 108.815 196.240 ;
        RECT 109.415 187.210 109.695 197.505 ;
        RECT 108.955 186.690 110.155 187.020 ;
        RECT 110.295 186.165 110.575 196.240 ;
        RECT 111.175 187.210 111.455 197.505 ;
        RECT 110.715 186.690 111.915 187.020 ;
        RECT 112.055 186.165 112.335 196.240 ;
        RECT 112.935 187.210 113.215 197.505 ;
        RECT 122.155 197.440 122.435 198.050 ;
        RECT 112.680 186.690 113.530 187.020 ;
        RECT 113.815 186.165 114.095 196.240 ;
        RECT 114.695 190.725 114.975 192.725 ;
        RECT 115.575 190.725 115.855 192.725 ;
        RECT 116.260 190.725 116.550 192.725 ;
        RECT 117.060 190.725 117.350 192.725 ;
        RECT 117.755 190.725 118.035 192.725 ;
        RECT 118.635 190.725 118.915 192.725 ;
        RECT 119.515 190.725 119.795 192.725 ;
        RECT 120.395 190.725 120.675 192.725 ;
        RECT 121.275 190.725 121.555 192.725 ;
        RECT 122.155 190.725 122.435 192.725 ;
        RECT 72.400 185.365 114.095 186.165 ;
        RECT 72.400 172.150 73.000 185.365 ;
        RECT 74.360 182.605 74.650 183.605 ;
        RECT 75.095 182.605 75.375 183.605 ;
        RECT 75.975 182.605 76.255 183.605 ;
        RECT 76.855 182.605 77.135 183.605 ;
        RECT 77.735 182.605 78.015 183.605 ;
        RECT 78.615 181.975 78.895 185.365 ;
        RECT 73.820 181.785 74.150 181.830 ;
        RECT 73.820 181.455 74.990 181.785 ;
        RECT 73.820 172.780 74.150 181.455 ;
        RECT 79.495 180.410 79.775 184.235 ;
        RECT 80.375 181.975 80.655 185.365 ;
        RECT 81.255 180.410 81.535 184.235 ;
        RECT 82.135 181.975 82.415 185.365 ;
        RECT 83.015 180.410 83.295 184.235 ;
        RECT 83.895 181.975 84.175 185.365 ;
        RECT 84.775 180.410 85.055 184.235 ;
        RECT 85.655 181.975 85.935 185.365 ;
        RECT 86.535 180.410 86.815 184.235 ;
        RECT 87.415 181.975 87.695 185.365 ;
        RECT 88.295 180.410 88.575 184.235 ;
        RECT 89.175 181.975 89.455 185.365 ;
        RECT 90.055 180.410 90.335 184.235 ;
        RECT 90.935 181.975 91.215 185.365 ;
        RECT 91.815 180.410 92.095 184.235 ;
        RECT 92.695 181.975 92.975 185.365 ;
        RECT 93.575 180.410 93.855 184.235 ;
        RECT 94.455 181.975 94.735 185.365 ;
        RECT 95.335 180.410 95.615 184.235 ;
        RECT 96.215 181.975 96.495 185.365 ;
        RECT 97.095 180.410 97.375 184.235 ;
        RECT 97.975 181.975 98.255 185.365 ;
        RECT 98.855 180.410 99.135 184.235 ;
        RECT 99.735 181.975 100.015 185.365 ;
        RECT 100.615 180.410 100.895 184.235 ;
        RECT 101.495 181.975 101.775 185.365 ;
        RECT 102.375 180.410 102.655 184.235 ;
        RECT 103.255 181.975 103.535 185.365 ;
        RECT 104.135 180.410 104.415 184.235 ;
        RECT 105.015 181.975 105.295 185.365 ;
        RECT 105.895 180.410 106.175 184.235 ;
        RECT 106.775 181.975 107.055 185.365 ;
        RECT 107.655 180.410 107.935 184.235 ;
        RECT 108.535 181.975 108.815 185.365 ;
        RECT 109.415 180.410 109.695 184.235 ;
        RECT 110.295 181.975 110.575 185.365 ;
        RECT 111.175 180.410 111.455 184.235 ;
        RECT 112.055 181.975 112.335 185.365 ;
        RECT 112.935 180.410 113.215 184.235 ;
        RECT 113.815 181.975 114.095 185.365 ;
        RECT 114.695 182.605 114.975 183.605 ;
        RECT 115.575 182.605 115.855 183.605 ;
        RECT 116.300 182.605 116.590 183.605 ;
        RECT 117.020 182.605 117.310 183.605 ;
        RECT 117.755 182.605 118.035 183.605 ;
        RECT 118.635 182.605 118.915 183.605 ;
        RECT 119.515 182.605 119.795 183.605 ;
        RECT 120.395 182.605 120.675 183.605 ;
        RECT 121.275 182.605 121.555 183.605 ;
        RECT 122.155 182.605 122.435 183.605 ;
        RECT 114.000 181.455 115.760 181.785 ;
        RECT 79.495 179.610 113.215 180.410 ;
        RECT 123.035 180.055 123.315 196.240 ;
        RECT 123.915 187.210 124.195 198.050 ;
        RECT 123.605 186.690 124.455 187.020 ;
        RECT 74.360 176.120 74.650 177.120 ;
        RECT 75.095 176.120 75.375 177.120 ;
        RECT 75.975 176.120 76.255 177.120 ;
        RECT 76.855 176.120 77.135 177.120 ;
        RECT 77.735 176.120 78.015 177.120 ;
        RECT 78.615 176.120 78.895 177.120 ;
        RECT 79.495 175.490 79.775 179.610 ;
        RECT 80.375 176.120 80.655 177.120 ;
        RECT 81.255 175.490 81.535 179.610 ;
        RECT 82.135 176.120 82.415 177.120 ;
        RECT 83.015 175.490 83.295 179.610 ;
        RECT 83.895 176.120 84.175 177.120 ;
        RECT 84.775 175.490 85.055 179.610 ;
        RECT 85.655 176.120 85.935 177.120 ;
        RECT 86.535 175.490 86.815 179.610 ;
        RECT 87.415 176.120 87.695 177.120 ;
        RECT 88.295 175.490 88.575 179.610 ;
        RECT 89.175 176.120 89.455 177.120 ;
        RECT 90.055 175.490 90.335 179.610 ;
        RECT 90.935 176.120 91.215 177.120 ;
        RECT 91.815 175.490 92.095 179.610 ;
        RECT 92.695 176.120 92.975 177.120 ;
        RECT 93.575 175.490 93.855 179.610 ;
        RECT 94.455 176.120 94.735 177.120 ;
        RECT 95.335 175.490 95.615 179.610 ;
        RECT 96.215 176.120 96.495 177.120 ;
        RECT 97.095 175.490 97.375 179.610 ;
        RECT 97.975 176.120 98.255 177.120 ;
        RECT 98.855 175.490 99.135 179.610 ;
        RECT 99.735 176.120 100.015 177.120 ;
        RECT 100.615 175.490 100.895 179.610 ;
        RECT 101.495 176.120 101.775 177.120 ;
        RECT 102.375 175.490 102.655 179.610 ;
        RECT 103.255 176.120 103.535 177.120 ;
        RECT 104.135 175.490 104.415 179.610 ;
        RECT 105.015 176.120 105.295 177.120 ;
        RECT 105.895 175.490 106.175 179.610 ;
        RECT 106.775 176.120 107.055 177.120 ;
        RECT 107.655 175.490 107.935 179.610 ;
        RECT 108.535 176.120 108.815 177.120 ;
        RECT 109.415 175.490 109.695 179.610 ;
        RECT 110.295 176.120 110.575 177.120 ;
        RECT 111.175 175.490 111.455 179.610 ;
        RECT 111.810 177.940 112.580 178.230 ;
        RECT 112.055 176.120 112.335 177.120 ;
        RECT 112.935 175.490 113.215 179.610 ;
        RECT 113.815 176.120 114.095 177.120 ;
        RECT 114.695 176.120 114.975 177.120 ;
        RECT 115.575 176.120 115.855 177.120 ;
        RECT 116.300 176.120 116.590 177.120 ;
        RECT 117.020 176.120 117.310 177.120 ;
        RECT 117.755 176.120 118.035 177.120 ;
        RECT 118.635 176.120 118.915 177.120 ;
        RECT 119.515 176.120 119.795 177.120 ;
        RECT 120.395 176.120 120.675 177.120 ;
        RECT 121.275 176.120 121.555 177.120 ;
        RECT 122.155 176.120 122.435 177.120 ;
        RECT 123.035 176.120 123.315 177.120 ;
        RECT 123.915 173.440 124.195 184.235 ;
        RECT 124.795 180.055 125.075 196.240 ;
        RECT 125.675 187.210 125.955 198.050 ;
        RECT 125.215 186.690 126.415 187.020 ;
        RECT 124.795 176.120 125.075 177.120 ;
        RECT 125.675 173.440 125.955 184.235 ;
        RECT 126.555 180.055 126.835 196.240 ;
        RECT 127.435 187.210 127.715 198.050 ;
        RECT 126.975 186.690 128.175 187.020 ;
        RECT 126.555 176.120 126.835 177.120 ;
        RECT 127.435 173.440 127.715 184.235 ;
        RECT 128.315 180.055 128.595 196.240 ;
        RECT 129.195 187.210 129.475 198.050 ;
        RECT 130.955 197.440 131.235 198.050 ;
        RECT 132.715 197.790 132.995 208.605 ;
        RECT 133.595 203.085 133.875 205.085 ;
        RECT 134.475 197.790 134.755 208.605 ;
        RECT 135.355 203.085 135.635 205.085 ;
        RECT 136.235 197.790 136.515 208.605 ;
        RECT 137.115 203.085 137.395 205.085 ;
        RECT 137.995 197.790 138.275 208.605 ;
        RECT 138.875 203.085 139.155 205.085 ;
        RECT 139.755 197.790 140.035 208.605 ;
        RECT 140.635 203.085 140.915 205.085 ;
        RECT 141.515 197.790 141.795 208.605 ;
        RECT 142.395 203.085 142.675 205.085 ;
        RECT 143.275 203.085 143.555 205.085 ;
        RECT 144.155 203.085 144.435 205.085 ;
        RECT 145.035 203.085 145.315 205.085 ;
        RECT 145.915 203.085 146.195 205.085 ;
        RECT 146.600 203.085 146.890 205.085 ;
        RECT 152.195 198.050 152.875 198.420 ;
        RECT 132.515 197.420 133.195 197.790 ;
        RECT 134.275 197.420 134.955 197.790 ;
        RECT 136.035 197.420 136.715 197.790 ;
        RECT 137.795 197.420 138.475 197.790 ;
        RECT 139.555 197.420 140.235 197.790 ;
        RECT 141.315 197.420 141.995 197.790 ;
        RECT 128.735 186.690 129.935 187.020 ;
        RECT 128.315 176.120 128.595 177.120 ;
        RECT 129.195 173.440 129.475 184.235 ;
        RECT 130.075 180.055 130.355 196.240 ;
        RECT 130.955 190.725 131.235 192.725 ;
        RECT 131.835 190.725 132.115 192.725 ;
        RECT 132.715 190.725 132.995 192.725 ;
        RECT 130.955 182.605 131.235 183.605 ;
        RECT 131.835 182.605 132.115 183.605 ;
        RECT 132.715 182.605 132.995 183.605 ;
        RECT 133.595 180.055 133.875 196.240 ;
        RECT 134.475 187.210 134.755 197.420 ;
        RECT 134.015 186.690 135.215 187.020 ;
        RECT 130.075 176.120 130.355 177.120 ;
        RECT 130.955 176.120 131.235 177.120 ;
        RECT 131.835 176.120 132.115 177.120 ;
        RECT 132.715 176.120 132.995 177.120 ;
        RECT 133.595 176.120 133.875 177.120 ;
        RECT 134.475 175.490 134.755 184.235 ;
        RECT 135.355 180.055 135.635 196.240 ;
        RECT 136.235 187.210 136.515 197.420 ;
        RECT 135.775 186.690 136.975 187.020 ;
        RECT 135.355 176.120 135.635 177.120 ;
        RECT 136.235 175.490 136.515 184.235 ;
        RECT 137.115 180.575 137.395 196.240 ;
        RECT 137.995 187.210 138.275 197.420 ;
        RECT 137.535 186.690 138.735 187.020 ;
        RECT 137.005 178.245 137.505 180.575 ;
        RECT 136.965 177.925 137.545 178.245 ;
        RECT 137.115 176.120 137.395 177.120 ;
        RECT 137.995 175.490 138.275 184.235 ;
        RECT 138.875 180.055 139.155 196.240 ;
        RECT 139.755 187.210 140.035 197.420 ;
        RECT 139.500 186.690 140.350 187.020 ;
        RECT 138.875 176.120 139.155 177.120 ;
        RECT 139.755 175.490 140.035 184.235 ;
        RECT 140.635 180.055 140.915 196.240 ;
        RECT 141.515 190.725 141.795 192.725 ;
        RECT 142.395 190.725 142.675 192.725 ;
        RECT 143.275 190.725 143.555 192.725 ;
        RECT 144.155 190.725 144.435 192.725 ;
        RECT 145.035 190.725 145.315 192.725 ;
        RECT 145.915 190.725 146.195 192.725 ;
        RECT 146.600 190.725 146.890 192.725 ;
        RECT 147.280 191.215 147.570 192.215 ;
        RECT 148.015 191.215 148.295 192.215 ;
        RECT 148.895 191.215 149.175 192.215 ;
        RECT 149.775 191.215 150.055 192.215 ;
        RECT 150.655 191.215 150.935 192.215 ;
        RECT 151.535 188.240 151.815 192.845 ;
        RECT 152.415 190.585 152.695 198.050 ;
        RECT 154.175 197.790 154.455 198.400 ;
        RECT 155.715 198.050 156.395 198.420 ;
        RECT 153.975 197.420 154.655 197.790 ;
        RECT 153.295 188.240 153.575 192.845 ;
        RECT 154.175 190.585 154.455 197.420 ;
        RECT 155.055 188.240 155.335 192.845 ;
        RECT 155.935 190.585 156.215 198.050 ;
        RECT 157.695 197.790 157.975 198.400 ;
        RECT 159.235 198.050 159.915 198.420 ;
        RECT 157.495 197.420 158.175 197.790 ;
        RECT 156.815 188.240 157.095 192.845 ;
        RECT 157.695 190.585 157.975 197.420 ;
        RECT 158.575 188.240 158.855 192.845 ;
        RECT 159.455 190.585 159.735 198.050 ;
        RECT 161.215 197.790 161.495 198.400 ;
        RECT 162.755 198.050 163.435 198.420 ;
        RECT 161.015 197.420 161.695 197.790 ;
        RECT 160.335 188.240 160.615 192.845 ;
        RECT 161.215 190.585 161.495 197.420 ;
        RECT 162.095 188.240 162.375 192.845 ;
        RECT 162.975 190.585 163.255 198.050 ;
        RECT 164.735 197.790 165.015 198.400 ;
        RECT 164.535 197.420 165.215 197.790 ;
        RECT 163.855 188.240 164.135 192.845 ;
        RECT 164.735 190.585 165.015 197.420 ;
        RECT 167.385 193.625 169.050 193.915 ;
        RECT 165.615 188.240 165.895 192.845 ;
        RECT 166.495 191.215 166.775 192.215 ;
        RECT 167.375 191.215 167.655 192.215 ;
        RECT 168.255 191.215 168.535 192.215 ;
        RECT 169.135 191.215 169.415 192.215 ;
        RECT 169.860 191.215 170.150 192.215 ;
        RECT 167.385 189.515 169.050 189.805 ;
        RECT 151.535 187.740 165.895 188.240 ;
        RECT 141.515 182.605 141.795 183.605 ;
        RECT 142.395 182.605 142.675 183.605 ;
        RECT 143.275 182.605 143.555 183.605 ;
        RECT 144.155 182.605 144.435 183.605 ;
        RECT 145.035 182.605 145.315 183.605 ;
        RECT 145.915 182.605 146.195 183.605 ;
        RECT 146.640 182.605 146.930 183.605 ;
        RECT 147.280 182.605 147.570 183.605 ;
        RECT 148.015 182.605 148.295 183.605 ;
        RECT 148.895 182.605 149.175 183.605 ;
        RECT 149.775 182.605 150.055 183.605 ;
        RECT 150.655 182.605 150.935 183.605 ;
        RECT 151.535 182.605 151.815 183.605 ;
        RECT 152.415 182.605 152.695 183.605 ;
        RECT 153.295 182.605 153.575 183.605 ;
        RECT 154.175 182.605 154.455 183.605 ;
        RECT 155.055 181.975 155.335 187.740 ;
        RECT 141.515 181.455 143.275 181.785 ;
        RECT 155.420 181.455 155.795 181.785 ;
        RECT 155.935 180.110 156.215 184.235 ;
        RECT 156.815 181.975 157.095 187.740 ;
        RECT 156.355 181.455 157.555 181.785 ;
        RECT 157.695 180.110 157.975 184.235 ;
        RECT 158.575 181.975 158.855 187.740 ;
        RECT 158.115 181.455 159.315 181.785 ;
        RECT 159.455 180.110 159.735 184.235 ;
        RECT 160.335 181.975 160.615 187.740 ;
        RECT 159.875 181.455 161.075 181.785 ;
        RECT 161.215 180.110 161.495 184.235 ;
        RECT 162.095 181.975 162.375 187.740 ;
        RECT 162.975 182.605 163.255 183.605 ;
        RECT 163.855 182.605 164.135 183.605 ;
        RECT 164.735 182.605 165.015 183.605 ;
        RECT 165.615 182.605 165.895 183.605 ;
        RECT 166.495 182.605 166.775 183.605 ;
        RECT 167.375 182.605 167.655 183.605 ;
        RECT 168.255 182.605 168.535 183.605 ;
        RECT 169.135 182.605 169.415 183.605 ;
        RECT 169.860 182.605 170.150 183.605 ;
        RECT 161.635 181.455 162.030 181.785 ;
        RECT 155.935 179.610 161.495 180.110 ;
        RECT 140.635 176.120 140.915 177.120 ;
        RECT 141.515 176.120 141.795 177.120 ;
        RECT 142.395 176.120 142.675 177.120 ;
        RECT 143.275 176.120 143.555 177.120 ;
        RECT 144.155 176.120 144.435 177.120 ;
        RECT 145.035 176.120 145.315 177.120 ;
        RECT 145.915 176.120 146.195 177.120 ;
        RECT 146.640 176.120 146.930 177.120 ;
        RECT 147.280 176.120 147.570 177.120 ;
        RECT 148.015 176.120 148.295 177.120 ;
        RECT 148.895 176.120 149.175 177.120 ;
        RECT 149.775 176.120 150.055 177.120 ;
        RECT 150.655 176.120 150.935 177.120 ;
        RECT 151.535 176.120 151.815 177.120 ;
        RECT 152.415 176.120 152.695 177.120 ;
        RECT 153.295 176.120 153.575 177.120 ;
        RECT 154.175 176.120 154.455 177.120 ;
        RECT 155.055 176.120 155.335 177.120 ;
        RECT 155.935 175.490 156.215 179.610 ;
        RECT 156.815 176.120 157.095 177.120 ;
        RECT 157.695 175.490 157.975 179.610 ;
        RECT 158.575 176.120 158.855 177.120 ;
        RECT 159.455 175.490 159.735 179.610 ;
        RECT 160.335 176.120 160.615 177.120 ;
        RECT 161.215 175.490 161.495 179.610 ;
        RECT 162.095 176.120 162.375 177.120 ;
        RECT 162.975 176.120 163.255 177.120 ;
        RECT 163.855 176.120 164.135 177.120 ;
        RECT 164.735 176.120 165.015 177.120 ;
        RECT 165.615 176.120 165.895 177.120 ;
        RECT 166.495 176.120 166.775 177.120 ;
        RECT 167.375 176.120 167.655 177.120 ;
        RECT 168.255 176.120 168.535 177.120 ;
        RECT 169.135 176.120 169.415 177.120 ;
        RECT 169.860 176.120 170.150 177.120 ;
        RECT 160.615 174.970 162.010 175.300 ;
        RECT 123.715 173.070 124.395 173.440 ;
        RECT 125.475 173.070 126.155 173.440 ;
        RECT 127.235 173.070 127.915 173.440 ;
        RECT 128.995 173.070 129.675 173.440 ;
        RECT 73.400 172.450 74.570 172.780 ;
        RECT 72.400 171.550 73.505 172.150 ;
        RECT 171.460 155.250 171.790 208.755 ;
        RECT 172.330 177.315 172.660 187.040 ;
        RECT 172.330 176.985 173.500 177.315 ;
        RECT 171.460 154.920 172.630 155.250 ;
        RECT 46.010 0.890 46.910 151.400 ;
        RECT 68.090 0.890 68.990 151.400 ;
        RECT 175.680 103.005 176.280 189.820 ;
        RECT 176.780 8.125 177.380 193.930 ;
        RECT 178.380 150.800 178.980 174.515 ;
        RECT 178.880 79.825 179.480 126.965 ;
        RECT 179.980 94.255 180.580 214.890 ;
        RECT 181.080 112.205 181.680 216.490 ;
        RECT 280.365 191.225 281.535 191.555 ;
        RECT 430.180 191.225 431.350 191.555 ;
        RECT 225.260 190.565 225.940 190.935 ;
        RECT 227.020 190.565 227.700 190.935 ;
        RECT 228.780 190.565 229.460 190.935 ;
        RECT 230.540 190.565 231.220 190.935 ;
        RECT 183.655 188.705 184.825 189.035 ;
        RECT 192.925 188.705 194.320 189.035 ;
        RECT 183.655 175.300 183.985 188.705 ;
        RECT 184.785 186.885 185.075 187.885 ;
        RECT 185.520 186.885 185.800 187.885 ;
        RECT 186.400 186.885 186.680 187.885 ;
        RECT 187.280 186.885 187.560 187.885 ;
        RECT 188.160 186.885 188.440 187.885 ;
        RECT 189.040 186.885 189.320 187.885 ;
        RECT 189.920 186.885 190.200 187.885 ;
        RECT 190.800 186.885 191.080 187.885 ;
        RECT 191.680 186.885 191.960 187.885 ;
        RECT 192.560 186.885 192.840 187.885 ;
        RECT 193.440 184.395 193.720 188.515 ;
        RECT 194.320 186.885 194.600 187.885 ;
        RECT 195.200 184.395 195.480 188.515 ;
        RECT 196.080 186.885 196.360 187.885 ;
        RECT 196.960 184.395 197.240 188.515 ;
        RECT 197.840 186.885 198.120 187.885 ;
        RECT 198.720 184.395 199.000 188.515 ;
        RECT 199.600 186.885 199.880 187.885 ;
        RECT 200.480 186.885 200.760 187.885 ;
        RECT 201.360 186.885 201.640 187.885 ;
        RECT 202.240 186.885 202.520 187.885 ;
        RECT 203.120 186.885 203.400 187.885 ;
        RECT 204.000 186.885 204.280 187.885 ;
        RECT 204.880 186.885 205.160 187.885 ;
        RECT 205.760 186.885 206.040 187.885 ;
        RECT 206.640 186.885 206.920 187.885 ;
        RECT 207.365 186.885 207.655 187.885 ;
        RECT 208.005 186.885 208.295 187.885 ;
        RECT 208.740 186.885 209.020 187.885 ;
        RECT 209.620 186.885 209.900 187.885 ;
        RECT 210.500 186.885 210.780 187.885 ;
        RECT 211.380 186.885 211.660 187.885 ;
        RECT 212.260 186.885 212.540 187.885 ;
        RECT 213.140 186.885 213.420 187.885 ;
        RECT 214.020 186.885 214.300 187.885 ;
        RECT 193.440 183.895 199.000 184.395 ;
        RECT 192.905 182.220 193.300 182.550 ;
        RECT 184.785 180.400 185.075 181.400 ;
        RECT 185.520 180.400 185.800 181.400 ;
        RECT 186.400 180.400 186.680 181.400 ;
        RECT 187.280 180.400 187.560 181.400 ;
        RECT 188.160 180.400 188.440 181.400 ;
        RECT 189.040 180.400 189.320 181.400 ;
        RECT 189.920 180.400 190.200 181.400 ;
        RECT 190.800 180.400 191.080 181.400 ;
        RECT 191.680 180.400 191.960 181.400 ;
        RECT 192.560 176.265 192.840 182.030 ;
        RECT 193.440 179.770 193.720 183.895 ;
        RECT 193.860 182.220 195.060 182.550 ;
        RECT 194.320 176.265 194.600 182.030 ;
        RECT 195.200 179.770 195.480 183.895 ;
        RECT 195.620 182.220 196.820 182.550 ;
        RECT 196.080 176.265 196.360 182.030 ;
        RECT 196.960 179.770 197.240 183.895 ;
        RECT 197.380 182.220 198.580 182.550 ;
        RECT 197.840 176.265 198.120 182.030 ;
        RECT 198.720 179.770 199.000 183.895 ;
        RECT 199.140 182.220 199.515 182.550 ;
        RECT 211.660 182.220 213.420 182.550 ;
        RECT 199.600 176.265 199.880 182.030 ;
        RECT 200.480 180.400 200.760 181.400 ;
        RECT 201.360 180.400 201.640 181.400 ;
        RECT 202.240 180.400 202.520 181.400 ;
        RECT 203.120 180.400 203.400 181.400 ;
        RECT 204.000 180.400 204.280 181.400 ;
        RECT 204.880 180.400 205.160 181.400 ;
        RECT 205.760 180.400 206.040 181.400 ;
        RECT 206.640 180.400 206.920 181.400 ;
        RECT 207.365 180.400 207.655 181.400 ;
        RECT 208.005 180.400 208.295 181.400 ;
        RECT 208.740 180.400 209.020 181.400 ;
        RECT 209.620 180.400 209.900 181.400 ;
        RECT 210.500 180.400 210.780 181.400 ;
        RECT 211.380 180.400 211.660 181.400 ;
        RECT 212.260 180.400 212.540 181.400 ;
        RECT 213.140 180.400 213.420 181.400 ;
        RECT 182.815 174.970 183.985 175.300 ;
        RECT 189.040 175.765 203.400 176.265 ;
        RECT 185.885 174.200 187.550 174.490 ;
        RECT 184.785 171.790 185.075 172.790 ;
        RECT 185.520 171.790 185.800 172.790 ;
        RECT 186.400 171.790 186.680 172.790 ;
        RECT 187.280 171.790 187.560 172.790 ;
        RECT 188.160 171.790 188.440 172.790 ;
        RECT 189.040 171.160 189.320 175.765 ;
        RECT 183.180 120.945 183.780 170.405 ;
        RECT 185.885 170.090 187.550 170.380 ;
        RECT 189.920 166.585 190.200 173.420 ;
        RECT 190.800 171.160 191.080 175.765 ;
        RECT 189.720 166.215 190.400 166.585 ;
        RECT 189.920 165.605 190.200 166.215 ;
        RECT 191.680 165.955 191.960 173.420 ;
        RECT 192.560 171.160 192.840 175.765 ;
        RECT 193.440 166.585 193.720 173.420 ;
        RECT 194.320 171.160 194.600 175.765 ;
        RECT 193.240 166.215 193.920 166.585 ;
        RECT 191.500 165.585 192.180 165.955 ;
        RECT 193.440 165.605 193.720 166.215 ;
        RECT 195.200 165.955 195.480 173.420 ;
        RECT 196.080 171.160 196.360 175.765 ;
        RECT 196.960 166.585 197.240 173.420 ;
        RECT 197.840 171.160 198.120 175.765 ;
        RECT 196.760 166.215 197.440 166.585 ;
        RECT 195.020 165.585 195.700 165.955 ;
        RECT 196.960 165.605 197.240 166.215 ;
        RECT 198.720 165.955 199.000 173.420 ;
        RECT 199.600 171.160 199.880 175.765 ;
        RECT 200.480 166.585 200.760 173.420 ;
        RECT 201.360 171.160 201.640 175.765 ;
        RECT 200.280 166.215 200.960 166.585 ;
        RECT 198.540 165.585 199.220 165.955 ;
        RECT 200.480 165.605 200.760 166.215 ;
        RECT 202.240 165.955 202.520 173.420 ;
        RECT 203.120 171.160 203.400 175.765 ;
        RECT 204.000 171.790 204.280 172.790 ;
        RECT 204.880 171.790 205.160 172.790 ;
        RECT 205.760 171.790 206.040 172.790 ;
        RECT 206.640 171.790 206.920 172.790 ;
        RECT 207.365 171.790 207.655 172.790 ;
        RECT 208.045 171.280 208.335 173.280 ;
        RECT 208.740 171.280 209.020 173.280 ;
        RECT 209.620 171.280 209.900 173.280 ;
        RECT 210.500 171.280 210.780 173.280 ;
        RECT 211.380 171.280 211.660 173.280 ;
        RECT 212.260 171.280 212.540 173.280 ;
        RECT 213.140 171.280 213.420 173.280 ;
        RECT 214.020 167.765 214.300 183.950 ;
        RECT 214.900 179.770 215.180 188.515 ;
        RECT 215.780 186.885 216.060 187.885 ;
        RECT 214.585 176.985 215.435 177.315 ;
        RECT 214.900 166.585 215.180 176.795 ;
        RECT 215.780 167.765 216.060 183.950 ;
        RECT 216.660 179.770 216.940 188.515 ;
        RECT 217.540 186.885 217.820 187.885 ;
        RECT 217.390 185.760 217.970 186.080 ;
        RECT 217.430 183.430 217.930 185.760 ;
        RECT 216.200 176.985 217.400 177.315 ;
        RECT 216.660 166.585 216.940 176.795 ;
        RECT 217.540 167.765 217.820 183.430 ;
        RECT 218.420 179.770 218.700 188.515 ;
        RECT 219.300 186.885 219.580 187.885 ;
        RECT 217.960 176.985 219.160 177.315 ;
        RECT 218.420 166.585 218.700 176.795 ;
        RECT 219.300 167.765 219.580 183.950 ;
        RECT 220.180 179.770 220.460 188.515 ;
        RECT 221.060 186.885 221.340 187.885 ;
        RECT 221.940 186.885 222.220 187.885 ;
        RECT 222.820 186.885 223.100 187.885 ;
        RECT 223.700 186.885 223.980 187.885 ;
        RECT 224.580 186.885 224.860 187.885 ;
        RECT 219.720 176.985 220.920 177.315 ;
        RECT 220.180 166.585 220.460 176.795 ;
        RECT 221.060 167.765 221.340 183.950 ;
        RECT 221.940 180.400 222.220 181.400 ;
        RECT 222.820 180.400 223.100 181.400 ;
        RECT 223.700 180.400 223.980 181.400 ;
        RECT 221.940 171.280 222.220 173.280 ;
        RECT 222.820 171.280 223.100 173.280 ;
        RECT 223.700 171.280 223.980 173.280 ;
        RECT 224.580 167.765 224.860 183.950 ;
        RECT 225.460 179.770 225.740 190.565 ;
        RECT 226.340 186.885 226.620 187.885 ;
        RECT 225.000 176.985 226.200 177.315 ;
        RECT 212.940 166.215 213.620 166.585 ;
        RECT 214.700 166.215 215.380 166.585 ;
        RECT 216.460 166.215 217.140 166.585 ;
        RECT 218.220 166.215 218.900 166.585 ;
        RECT 219.980 166.215 220.660 166.585 ;
        RECT 221.740 166.215 222.420 166.585 ;
        RECT 202.060 165.585 202.740 165.955 ;
        RECT 208.045 158.920 208.335 160.920 ;
        RECT 208.740 158.920 209.020 160.920 ;
        RECT 209.620 158.920 209.900 160.920 ;
        RECT 210.500 158.920 210.780 160.920 ;
        RECT 211.380 158.920 211.660 160.920 ;
        RECT 212.260 158.920 212.540 160.920 ;
        RECT 213.140 155.400 213.420 166.215 ;
        RECT 214.020 158.920 214.300 160.920 ;
        RECT 214.900 155.400 215.180 166.215 ;
        RECT 215.780 158.920 216.060 160.920 ;
        RECT 216.660 155.400 216.940 166.215 ;
        RECT 217.540 158.920 217.820 160.920 ;
        RECT 218.420 155.400 218.700 166.215 ;
        RECT 219.300 158.920 219.580 160.920 ;
        RECT 220.180 155.400 220.460 166.215 ;
        RECT 221.060 158.920 221.340 160.920 ;
        RECT 221.940 155.400 222.220 166.215 ;
        RECT 223.700 165.955 223.980 166.565 ;
        RECT 225.460 165.955 225.740 176.795 ;
        RECT 226.340 167.765 226.620 183.950 ;
        RECT 227.220 179.770 227.500 190.565 ;
        RECT 228.100 186.885 228.380 187.885 ;
        RECT 226.760 176.985 227.960 177.315 ;
        RECT 227.220 165.955 227.500 176.795 ;
        RECT 228.100 167.765 228.380 183.950 ;
        RECT 228.980 179.770 229.260 190.565 ;
        RECT 229.860 186.885 230.140 187.885 ;
        RECT 228.520 176.985 229.720 177.315 ;
        RECT 228.980 165.955 229.260 176.795 ;
        RECT 229.860 167.765 230.140 183.950 ;
        RECT 230.740 179.770 231.020 190.565 ;
        RECT 231.620 186.885 231.900 187.885 ;
        RECT 232.500 186.885 232.780 187.885 ;
        RECT 233.380 186.885 233.660 187.885 ;
        RECT 234.260 186.885 234.540 187.885 ;
        RECT 235.140 186.885 235.420 187.885 ;
        RECT 236.020 186.885 236.300 187.885 ;
        RECT 236.900 186.885 237.180 187.885 ;
        RECT 237.625 186.885 237.915 187.885 ;
        RECT 238.345 186.885 238.635 187.885 ;
        RECT 239.080 186.885 239.360 187.885 ;
        RECT 239.960 186.885 240.240 187.885 ;
        RECT 240.840 186.885 241.120 187.885 ;
        RECT 241.720 184.395 242.000 188.515 ;
        RECT 242.600 186.885 242.880 187.885 ;
        RECT 242.355 185.775 243.125 186.065 ;
        RECT 243.480 184.395 243.760 188.515 ;
        RECT 244.360 186.885 244.640 187.885 ;
        RECT 245.240 184.395 245.520 188.515 ;
        RECT 246.120 186.885 246.400 187.885 ;
        RECT 247.000 184.395 247.280 188.515 ;
        RECT 247.880 186.885 248.160 187.885 ;
        RECT 248.760 184.395 249.040 188.515 ;
        RECT 249.640 186.885 249.920 187.885 ;
        RECT 250.520 184.395 250.800 188.515 ;
        RECT 251.400 186.885 251.680 187.885 ;
        RECT 252.280 184.395 252.560 188.515 ;
        RECT 253.160 186.885 253.440 187.885 ;
        RECT 254.040 184.395 254.320 188.515 ;
        RECT 254.920 186.885 255.200 187.885 ;
        RECT 255.800 184.395 256.080 188.515 ;
        RECT 256.680 186.885 256.960 187.885 ;
        RECT 257.560 184.395 257.840 188.515 ;
        RECT 258.440 186.885 258.720 187.885 ;
        RECT 259.320 184.395 259.600 188.515 ;
        RECT 260.200 186.885 260.480 187.885 ;
        RECT 261.080 184.395 261.360 188.515 ;
        RECT 261.960 186.885 262.240 187.885 ;
        RECT 262.840 184.395 263.120 188.515 ;
        RECT 263.720 186.885 264.000 187.885 ;
        RECT 264.600 184.395 264.880 188.515 ;
        RECT 265.480 186.885 265.760 187.885 ;
        RECT 266.360 184.395 266.640 188.515 ;
        RECT 267.240 186.885 267.520 187.885 ;
        RECT 268.120 184.395 268.400 188.515 ;
        RECT 269.000 186.885 269.280 187.885 ;
        RECT 269.880 184.395 270.160 188.515 ;
        RECT 270.760 186.885 271.040 187.885 ;
        RECT 271.640 184.395 271.920 188.515 ;
        RECT 272.520 186.885 272.800 187.885 ;
        RECT 273.400 184.395 273.680 188.515 ;
        RECT 274.280 186.885 274.560 187.885 ;
        RECT 275.160 184.395 275.440 188.515 ;
        RECT 276.040 186.885 276.320 187.885 ;
        RECT 276.920 186.885 277.200 187.885 ;
        RECT 277.800 186.885 278.080 187.885 ;
        RECT 278.680 186.885 278.960 187.885 ;
        RECT 279.560 186.885 279.840 187.885 ;
        RECT 280.285 186.885 280.575 187.885 ;
        RECT 230.480 176.985 231.330 177.315 ;
        RECT 230.740 165.955 231.020 176.795 ;
        RECT 231.620 167.765 231.900 183.950 ;
        RECT 241.720 183.595 275.440 184.395 ;
        RECT 239.175 182.220 240.935 182.550 ;
        RECT 232.500 180.400 232.780 181.400 ;
        RECT 233.380 180.400 233.660 181.400 ;
        RECT 234.260 180.400 234.540 181.400 ;
        RECT 235.140 180.400 235.420 181.400 ;
        RECT 236.020 180.400 236.300 181.400 ;
        RECT 236.900 180.400 237.180 181.400 ;
        RECT 237.625 180.400 237.915 181.400 ;
        RECT 238.345 180.400 238.635 181.400 ;
        RECT 239.080 180.400 239.360 181.400 ;
        RECT 239.960 180.400 240.240 181.400 ;
        RECT 240.840 178.640 241.120 182.030 ;
        RECT 241.720 179.770 242.000 183.595 ;
        RECT 242.600 178.640 242.880 182.030 ;
        RECT 243.480 179.770 243.760 183.595 ;
        RECT 244.360 178.640 244.640 182.030 ;
        RECT 245.240 179.770 245.520 183.595 ;
        RECT 246.120 178.640 246.400 182.030 ;
        RECT 247.000 179.770 247.280 183.595 ;
        RECT 247.880 178.640 248.160 182.030 ;
        RECT 248.760 179.770 249.040 183.595 ;
        RECT 249.640 178.640 249.920 182.030 ;
        RECT 250.520 179.770 250.800 183.595 ;
        RECT 251.400 178.640 251.680 182.030 ;
        RECT 252.280 179.770 252.560 183.595 ;
        RECT 253.160 178.640 253.440 182.030 ;
        RECT 254.040 179.770 254.320 183.595 ;
        RECT 254.920 178.640 255.200 182.030 ;
        RECT 255.800 179.770 256.080 183.595 ;
        RECT 256.680 178.640 256.960 182.030 ;
        RECT 257.560 179.770 257.840 183.595 ;
        RECT 258.440 178.640 258.720 182.030 ;
        RECT 259.320 179.770 259.600 183.595 ;
        RECT 260.200 178.640 260.480 182.030 ;
        RECT 261.080 179.770 261.360 183.595 ;
        RECT 261.960 178.640 262.240 182.030 ;
        RECT 262.840 179.770 263.120 183.595 ;
        RECT 263.720 178.640 264.000 182.030 ;
        RECT 264.600 179.770 264.880 183.595 ;
        RECT 265.480 178.640 265.760 182.030 ;
        RECT 266.360 179.770 266.640 183.595 ;
        RECT 267.240 178.640 267.520 182.030 ;
        RECT 268.120 179.770 268.400 183.595 ;
        RECT 269.000 178.640 269.280 182.030 ;
        RECT 269.880 179.770 270.160 183.595 ;
        RECT 270.760 178.640 271.040 182.030 ;
        RECT 271.640 179.770 271.920 183.595 ;
        RECT 272.520 178.640 272.800 182.030 ;
        RECT 273.400 179.770 273.680 183.595 ;
        RECT 274.280 178.640 274.560 182.030 ;
        RECT 275.160 179.770 275.440 183.595 ;
        RECT 280.785 182.550 281.115 191.225 ;
        RECT 429.050 189.825 430.220 190.155 ;
        RECT 279.945 182.220 281.115 182.550 ;
        RECT 280.785 182.175 281.115 182.220 ;
        RECT 276.040 178.640 276.320 182.030 ;
        RECT 276.920 180.400 277.200 181.400 ;
        RECT 277.800 180.400 278.080 181.400 ;
        RECT 278.680 180.400 278.960 181.400 ;
        RECT 279.560 180.400 279.840 181.400 ;
        RECT 280.285 180.400 280.575 181.400 ;
        RECT 240.840 177.840 282.535 178.640 ;
        RECT 232.500 171.280 232.780 173.280 ;
        RECT 233.380 171.280 233.660 173.280 ;
        RECT 234.260 171.280 234.540 173.280 ;
        RECT 235.140 171.280 235.420 173.280 ;
        RECT 236.020 171.280 236.300 173.280 ;
        RECT 236.900 171.280 237.180 173.280 ;
        RECT 237.585 171.280 237.875 173.280 ;
        RECT 238.385 171.280 238.675 173.280 ;
        RECT 239.080 171.280 239.360 173.280 ;
        RECT 239.960 171.280 240.240 173.280 ;
        RECT 240.840 167.765 241.120 177.840 ;
        RECT 241.405 176.985 242.255 177.315 ;
        RECT 232.500 165.955 232.780 166.565 ;
        RECT 241.720 166.500 242.000 176.795 ;
        RECT 242.600 167.765 242.880 177.840 ;
        RECT 243.020 176.985 244.220 177.315 ;
        RECT 243.480 166.500 243.760 176.795 ;
        RECT 244.360 167.765 244.640 177.840 ;
        RECT 244.780 176.985 245.980 177.315 ;
        RECT 245.240 166.500 245.520 176.795 ;
        RECT 246.120 167.765 246.400 177.840 ;
        RECT 246.540 176.985 247.740 177.315 ;
        RECT 247.000 166.500 247.280 176.795 ;
        RECT 247.880 167.765 248.160 177.840 ;
        RECT 248.300 176.985 249.500 177.315 ;
        RECT 248.760 166.500 249.040 176.795 ;
        RECT 249.640 167.765 249.920 177.840 ;
        RECT 250.060 176.985 251.260 177.315 ;
        RECT 250.520 166.500 250.800 176.795 ;
        RECT 251.400 167.765 251.680 177.840 ;
        RECT 251.820 176.985 253.020 177.315 ;
        RECT 252.280 166.500 252.560 176.795 ;
        RECT 253.160 167.765 253.440 177.840 ;
        RECT 253.580 176.985 254.780 177.315 ;
        RECT 254.040 166.500 254.320 176.795 ;
        RECT 254.920 167.765 255.200 177.840 ;
        RECT 255.340 176.985 256.540 177.315 ;
        RECT 255.800 166.500 256.080 176.795 ;
        RECT 256.680 167.765 256.960 177.840 ;
        RECT 257.100 176.985 258.300 177.315 ;
        RECT 257.560 166.500 257.840 176.795 ;
        RECT 258.440 167.765 258.720 177.840 ;
        RECT 258.860 176.985 260.060 177.315 ;
        RECT 259.320 166.500 259.600 176.795 ;
        RECT 260.200 167.765 260.480 177.840 ;
        RECT 260.620 176.985 261.820 177.315 ;
        RECT 261.080 166.500 261.360 176.795 ;
        RECT 261.960 167.765 262.240 177.840 ;
        RECT 262.380 176.985 263.580 177.315 ;
        RECT 262.840 166.500 263.120 176.795 ;
        RECT 263.720 167.765 264.000 177.840 ;
        RECT 264.140 176.985 265.340 177.315 ;
        RECT 264.600 166.500 264.880 176.795 ;
        RECT 265.480 167.765 265.760 177.840 ;
        RECT 265.900 176.985 267.100 177.315 ;
        RECT 266.360 166.500 266.640 176.795 ;
        RECT 267.240 167.765 267.520 177.840 ;
        RECT 267.660 176.985 268.860 177.315 ;
        RECT 268.120 166.500 268.400 176.795 ;
        RECT 269.000 167.765 269.280 177.840 ;
        RECT 269.420 176.985 270.620 177.315 ;
        RECT 269.880 166.500 270.160 176.795 ;
        RECT 270.760 167.765 271.040 177.840 ;
        RECT 271.180 176.985 272.380 177.315 ;
        RECT 271.640 166.500 271.920 176.795 ;
        RECT 272.520 167.765 272.800 177.840 ;
        RECT 272.940 176.985 274.140 177.315 ;
        RECT 273.400 166.500 273.680 176.795 ;
        RECT 274.280 167.765 274.560 177.840 ;
        RECT 274.900 176.985 275.750 177.315 ;
        RECT 275.160 166.500 275.440 176.795 ;
        RECT 276.040 167.765 276.320 177.840 ;
        RECT 279.945 176.985 281.115 177.315 ;
        RECT 276.920 171.280 277.200 173.280 ;
        RECT 277.800 171.280 278.080 173.280 ;
        RECT 278.680 171.280 278.960 173.280 ;
        RECT 279.560 171.280 279.840 173.280 ;
        RECT 280.245 171.280 280.535 173.280 ;
        RECT 223.500 165.585 224.180 165.955 ;
        RECT 225.260 165.585 225.940 165.955 ;
        RECT 227.020 165.585 227.700 165.955 ;
        RECT 228.780 165.585 229.460 165.955 ;
        RECT 230.540 165.585 231.220 165.955 ;
        RECT 232.300 165.585 232.980 165.955 ;
        RECT 241.720 165.700 275.440 166.500 ;
        RECT 222.820 158.920 223.100 160.920 ;
        RECT 223.700 155.400 223.980 165.585 ;
        RECT 224.580 158.920 224.860 160.920 ;
        RECT 225.460 155.400 225.740 165.585 ;
        RECT 226.340 158.920 226.620 160.920 ;
        RECT 227.220 155.400 227.500 165.585 ;
        RECT 228.100 158.920 228.380 160.920 ;
        RECT 228.980 155.400 229.260 165.585 ;
        RECT 229.860 158.920 230.140 160.920 ;
        RECT 230.740 155.400 231.020 165.585 ;
        RECT 231.620 158.920 231.900 160.920 ;
        RECT 232.500 155.400 232.780 165.585 ;
        RECT 233.380 158.920 233.660 160.920 ;
        RECT 234.260 158.920 234.540 160.920 ;
        RECT 235.140 158.920 235.420 160.920 ;
        RECT 236.020 158.920 236.300 160.920 ;
        RECT 236.900 158.920 237.180 160.920 ;
        RECT 237.585 158.920 237.875 160.920 ;
        RECT 238.385 158.920 238.675 160.920 ;
        RECT 239.080 158.920 239.360 160.920 ;
        RECT 239.960 158.920 240.240 160.920 ;
        RECT 240.840 158.920 241.120 160.920 ;
        RECT 241.720 155.400 242.000 165.700 ;
        RECT 242.600 158.920 242.880 160.920 ;
        RECT 243.480 155.400 243.760 165.700 ;
        RECT 244.360 158.920 244.640 160.920 ;
        RECT 245.240 155.400 245.520 165.700 ;
        RECT 246.120 158.920 246.400 160.920 ;
        RECT 247.000 155.400 247.280 165.700 ;
        RECT 247.880 158.920 248.160 160.920 ;
        RECT 248.760 155.400 249.040 165.700 ;
        RECT 249.640 158.920 249.920 160.920 ;
        RECT 250.520 155.400 250.800 165.700 ;
        RECT 251.400 158.920 251.680 160.920 ;
        RECT 252.280 155.400 252.560 165.700 ;
        RECT 253.160 158.920 253.440 160.920 ;
        RECT 254.040 155.400 254.320 165.700 ;
        RECT 254.920 158.920 255.200 160.920 ;
        RECT 255.800 155.400 256.080 165.700 ;
        RECT 256.680 158.920 256.960 160.920 ;
        RECT 257.560 155.400 257.840 165.700 ;
        RECT 258.440 158.920 258.720 160.920 ;
        RECT 259.320 155.400 259.600 165.700 ;
        RECT 260.200 158.920 260.480 160.920 ;
        RECT 261.080 155.400 261.360 165.700 ;
        RECT 261.960 158.920 262.240 160.920 ;
        RECT 262.840 155.400 263.120 165.700 ;
        RECT 263.720 158.920 264.000 160.920 ;
        RECT 264.600 155.400 264.880 165.700 ;
        RECT 265.480 158.920 265.760 160.920 ;
        RECT 266.360 155.400 266.640 165.700 ;
        RECT 267.240 158.920 267.520 160.920 ;
        RECT 268.120 155.400 268.400 165.700 ;
        RECT 269.000 158.920 269.280 160.920 ;
        RECT 269.880 155.400 270.160 165.700 ;
        RECT 270.760 158.920 271.040 160.920 ;
        RECT 271.640 155.400 271.920 165.700 ;
        RECT 272.520 158.920 272.800 160.920 ;
        RECT 273.400 155.400 273.680 165.700 ;
        RECT 274.280 158.920 274.560 160.920 ;
        RECT 275.160 155.400 275.440 165.700 ;
        RECT 276.040 158.920 276.320 160.920 ;
        RECT 276.920 158.920 277.200 160.920 ;
        RECT 277.800 158.920 278.080 160.920 ;
        RECT 278.680 158.920 278.960 160.920 ;
        RECT 279.560 158.920 279.840 160.920 ;
        RECT 280.245 158.920 280.535 160.920 ;
        RECT 212.575 154.920 233.345 155.250 ;
        RECT 241.195 154.920 275.965 155.250 ;
        RECT 280.785 153.495 281.115 176.985 ;
        RECT 280.365 153.165 281.535 153.495 ;
        RECT 281.935 152.865 282.535 177.840 ;
        RECT 281.935 152.265 283.040 152.865 ;
        RECT 189.705 150.060 193.025 151.060 ;
        RECT 193.725 150.060 197.045 151.060 ;
        RECT 197.745 150.060 201.065 151.060 ;
        RECT 201.765 150.060 205.085 151.060 ;
        RECT 205.785 150.060 209.105 151.060 ;
        RECT 209.805 150.060 213.125 151.060 ;
        RECT 213.825 150.060 217.145 151.060 ;
        RECT 217.845 150.060 221.165 151.060 ;
        RECT 221.865 150.060 225.185 151.060 ;
        RECT 225.885 150.060 229.205 151.060 ;
        RECT 229.905 150.060 233.225 151.060 ;
        RECT 233.925 150.060 237.245 151.060 ;
        RECT 237.945 150.060 241.265 151.060 ;
        RECT 241.965 150.060 245.285 151.060 ;
        RECT 245.985 150.060 249.305 151.060 ;
        RECT 250.005 150.060 253.325 151.060 ;
        RECT 254.025 150.060 257.345 151.060 ;
        RECT 258.045 150.060 261.365 151.060 ;
        RECT 262.065 150.060 265.385 151.060 ;
        RECT 266.085 150.060 269.405 151.060 ;
        RECT 270.105 150.060 273.425 151.060 ;
        RECT 274.125 150.060 277.445 151.060 ;
        RECT 278.145 150.060 281.465 151.060 ;
        RECT 282.165 150.060 285.485 151.060 ;
        RECT 286.185 150.060 289.505 151.060 ;
        RECT 184.790 144.775 185.070 146.775 ;
        RECT 294.140 144.775 294.420 146.775 ;
        RECT 189.705 140.465 191.015 141.465 ;
        RECT 191.715 140.465 195.035 141.465 ;
        RECT 195.735 140.465 199.055 141.465 ;
        RECT 199.755 140.465 203.075 141.465 ;
        RECT 203.775 140.465 207.095 141.465 ;
        RECT 207.795 140.465 211.115 141.465 ;
        RECT 211.815 140.465 215.135 141.465 ;
        RECT 215.835 140.465 219.155 141.465 ;
        RECT 219.855 140.465 223.175 141.465 ;
        RECT 223.875 140.465 227.195 141.465 ;
        RECT 227.895 140.465 231.215 141.465 ;
        RECT 231.915 140.465 235.235 141.465 ;
        RECT 235.935 140.465 239.255 141.465 ;
        RECT 239.955 140.465 243.275 141.465 ;
        RECT 243.975 140.465 247.295 141.465 ;
        RECT 247.995 140.465 251.315 141.465 ;
        RECT 252.015 140.465 255.335 141.465 ;
        RECT 256.035 140.465 259.355 141.465 ;
        RECT 260.055 140.465 263.375 141.465 ;
        RECT 264.075 140.465 267.395 141.465 ;
        RECT 268.095 140.465 271.415 141.465 ;
        RECT 272.115 140.465 275.435 141.465 ;
        RECT 276.135 140.465 279.455 141.465 ;
        RECT 280.155 140.465 283.475 141.465 ;
        RECT 284.175 140.465 287.495 141.465 ;
        RECT 288.195 140.465 289.505 141.465 ;
        RECT 297.075 140.465 297.675 152.865 ;
        RECT 305.240 150.060 308.560 151.060 ;
        RECT 309.260 150.060 312.580 151.060 ;
        RECT 313.280 150.060 316.600 151.060 ;
        RECT 317.300 150.060 320.620 151.060 ;
        RECT 321.320 150.060 324.640 151.060 ;
        RECT 325.340 150.060 328.660 151.060 ;
        RECT 329.360 150.060 332.680 151.060 ;
        RECT 333.380 150.060 336.700 151.060 ;
        RECT 337.400 150.060 340.720 151.060 ;
        RECT 341.420 150.060 344.740 151.060 ;
        RECT 345.440 150.060 348.760 151.060 ;
        RECT 349.460 150.060 352.780 151.060 ;
        RECT 353.480 150.060 356.800 151.060 ;
        RECT 357.500 150.060 360.820 151.060 ;
        RECT 361.520 150.060 364.840 151.060 ;
        RECT 365.540 150.060 368.860 151.060 ;
        RECT 369.560 150.060 372.880 151.060 ;
        RECT 373.580 150.060 376.900 151.060 ;
        RECT 377.600 150.060 380.920 151.060 ;
        RECT 381.620 150.060 384.940 151.060 ;
        RECT 385.640 150.060 388.960 151.060 ;
        RECT 389.660 150.060 392.980 151.060 ;
        RECT 393.680 150.060 397.000 151.060 ;
        RECT 397.700 150.060 401.020 151.060 ;
        RECT 401.720 150.060 405.040 151.060 ;
        RECT 300.325 144.775 300.605 146.775 ;
        RECT 409.675 144.775 409.955 146.775 ;
        RECT 305.240 140.465 306.550 141.465 ;
        RECT 307.250 140.465 310.570 141.465 ;
        RECT 311.270 140.465 314.590 141.465 ;
        RECT 315.290 140.465 318.610 141.465 ;
        RECT 319.310 140.465 322.630 141.465 ;
        RECT 323.330 140.465 326.650 141.465 ;
        RECT 327.350 140.465 330.670 141.465 ;
        RECT 331.370 140.465 334.690 141.465 ;
        RECT 335.390 140.465 338.710 141.465 ;
        RECT 339.410 140.465 342.730 141.465 ;
        RECT 343.430 140.465 346.750 141.465 ;
        RECT 347.450 140.465 350.770 141.465 ;
        RECT 351.470 140.465 354.790 141.465 ;
        RECT 355.490 140.465 358.810 141.465 ;
        RECT 359.510 140.465 362.830 141.465 ;
        RECT 363.530 140.465 366.850 141.465 ;
        RECT 367.550 140.465 370.870 141.465 ;
        RECT 371.570 140.465 374.890 141.465 ;
        RECT 375.590 140.465 378.910 141.465 ;
        RECT 379.610 140.465 382.930 141.465 ;
        RECT 383.630 140.465 386.950 141.465 ;
        RECT 387.650 140.465 390.970 141.465 ;
        RECT 391.670 140.465 394.990 141.465 ;
        RECT 395.690 140.465 399.010 141.465 ;
        RECT 399.710 140.465 403.030 141.465 ;
        RECT 403.730 140.465 405.040 141.465 ;
        RECT 410.505 138.960 411.105 141.470 ;
        RECT 299.055 138.360 300.160 138.960 ;
        RECT 410.025 138.360 411.105 138.960 ;
        RECT 189.705 135.895 193.025 136.895 ;
        RECT 193.725 135.895 197.045 136.895 ;
        RECT 197.745 135.895 201.065 136.895 ;
        RECT 201.765 135.895 205.085 136.895 ;
        RECT 205.785 135.895 209.105 136.895 ;
        RECT 209.805 135.895 213.125 136.895 ;
        RECT 213.825 135.895 217.145 136.895 ;
        RECT 217.845 135.895 221.165 136.895 ;
        RECT 221.865 135.895 225.185 136.895 ;
        RECT 225.885 135.895 229.205 136.895 ;
        RECT 229.905 135.895 233.225 136.895 ;
        RECT 233.925 135.895 237.245 136.895 ;
        RECT 237.945 135.895 241.265 136.895 ;
        RECT 241.965 135.895 245.285 136.895 ;
        RECT 245.985 135.895 249.305 136.895 ;
        RECT 250.005 135.895 253.325 136.895 ;
        RECT 254.025 135.895 257.345 136.895 ;
        RECT 258.045 135.895 261.365 136.895 ;
        RECT 262.065 135.895 265.385 136.895 ;
        RECT 266.085 135.895 269.405 136.895 ;
        RECT 270.105 135.895 273.425 136.895 ;
        RECT 274.125 135.895 277.445 136.895 ;
        RECT 278.145 135.895 281.465 136.895 ;
        RECT 282.165 135.895 285.485 136.895 ;
        RECT 286.185 135.895 289.505 136.895 ;
        RECT 184.790 130.610 185.070 132.610 ;
        RECT 294.140 130.610 294.420 132.610 ;
        RECT 189.705 126.300 191.015 127.300 ;
        RECT 191.715 126.300 195.035 127.300 ;
        RECT 195.735 126.300 199.055 127.300 ;
        RECT 199.755 126.300 203.075 127.300 ;
        RECT 203.775 126.300 207.095 127.300 ;
        RECT 207.795 126.300 211.115 127.300 ;
        RECT 211.815 126.300 215.135 127.300 ;
        RECT 215.835 126.300 219.155 127.300 ;
        RECT 219.855 126.300 223.175 127.300 ;
        RECT 223.875 126.300 227.195 127.300 ;
        RECT 227.895 126.300 231.215 127.300 ;
        RECT 231.915 126.300 235.235 127.300 ;
        RECT 235.935 126.300 239.255 127.300 ;
        RECT 239.955 126.300 243.275 127.300 ;
        RECT 243.975 126.300 247.295 127.300 ;
        RECT 247.995 126.300 251.315 127.300 ;
        RECT 252.015 126.300 255.335 127.300 ;
        RECT 256.035 126.300 259.355 127.300 ;
        RECT 260.055 126.300 263.375 127.300 ;
        RECT 264.075 126.300 267.395 127.300 ;
        RECT 268.095 126.300 271.415 127.300 ;
        RECT 272.115 126.300 275.435 127.300 ;
        RECT 276.135 126.300 279.455 127.300 ;
        RECT 280.155 126.300 283.475 127.300 ;
        RECT 284.175 126.300 287.495 127.300 ;
        RECT 288.195 126.300 289.505 127.300 ;
        RECT 295.375 121.545 295.975 127.300 ;
        RECT 225.160 120.945 226.240 121.545 ;
        RECT 294.895 120.945 295.975 121.545 ;
        RECT 184.740 113.585 185.030 114.585 ;
        RECT 185.415 113.585 185.695 114.585 ;
        RECT 185.845 113.585 186.125 114.585 ;
        RECT 186.275 113.585 186.555 114.585 ;
        RECT 186.700 112.535 186.960 114.585 ;
        RECT 187.135 113.585 187.415 114.585 ;
        RECT 187.560 112.535 187.820 114.585 ;
        RECT 187.995 113.585 188.275 114.585 ;
        RECT 188.420 112.535 188.680 114.585 ;
        RECT 188.855 113.585 189.135 114.585 ;
        RECT 189.280 112.535 189.540 114.585 ;
        RECT 189.715 113.585 189.995 114.585 ;
        RECT 190.155 112.535 190.415 114.585 ;
        RECT 190.575 113.585 190.855 114.585 ;
        RECT 191.030 112.535 191.290 114.585 ;
        RECT 191.435 113.585 191.715 114.585 ;
        RECT 191.890 112.535 192.150 114.585 ;
        RECT 192.295 113.585 192.575 114.585 ;
        RECT 192.750 112.535 193.010 114.585 ;
        RECT 193.155 113.585 193.435 114.585 ;
        RECT 193.610 112.535 193.870 114.585 ;
        RECT 194.015 113.585 194.295 114.585 ;
        RECT 194.470 112.535 194.730 114.585 ;
        RECT 194.875 113.585 195.155 114.585 ;
        RECT 195.330 112.535 195.590 114.585 ;
        RECT 195.735 113.585 196.015 114.585 ;
        RECT 196.190 112.535 196.450 114.585 ;
        RECT 196.595 113.585 196.875 114.585 ;
        RECT 197.025 113.585 197.305 114.585 ;
        RECT 197.455 113.585 197.735 114.585 ;
        RECT 198.120 113.585 198.410 114.585 ;
        RECT 185.490 112.205 186.330 112.535 ;
        RECT 186.690 112.205 199.090 112.535 ;
        RECT 184.740 110.160 185.030 111.160 ;
        RECT 185.415 110.160 185.695 111.160 ;
        RECT 185.845 110.160 186.125 111.160 ;
        RECT 186.275 110.160 186.555 111.160 ;
        RECT 186.705 110.160 186.985 111.160 ;
        RECT 187.135 110.160 187.415 111.160 ;
        RECT 187.565 110.160 187.845 111.160 ;
        RECT 187.995 110.160 188.275 111.160 ;
        RECT 188.425 110.160 188.705 111.160 ;
        RECT 188.855 110.160 189.135 111.160 ;
        RECT 189.285 110.160 189.565 111.160 ;
        RECT 189.715 110.160 189.995 111.160 ;
        RECT 190.155 110.160 190.415 112.205 ;
        RECT 190.575 110.160 190.855 111.160 ;
        RECT 191.030 110.160 191.290 112.205 ;
        RECT 191.435 110.160 191.715 111.160 ;
        RECT 191.890 110.160 192.150 112.205 ;
        RECT 192.295 110.160 192.575 111.160 ;
        RECT 192.750 110.160 193.010 112.205 ;
        RECT 193.155 110.160 193.435 111.160 ;
        RECT 193.585 110.160 193.865 111.160 ;
        RECT 194.015 110.160 194.295 111.160 ;
        RECT 194.445 110.160 194.725 111.160 ;
        RECT 194.875 110.160 195.155 111.160 ;
        RECT 195.305 110.160 195.585 111.160 ;
        RECT 195.735 110.160 196.015 111.160 ;
        RECT 196.165 110.160 196.445 111.160 ;
        RECT 196.595 110.160 196.875 111.160 ;
        RECT 197.025 110.160 197.305 111.160 ;
        RECT 184.740 108.130 185.030 109.130 ;
        RECT 185.415 108.130 185.695 109.130 ;
        RECT 185.845 108.130 186.125 109.130 ;
        RECT 186.275 108.130 186.555 109.130 ;
        RECT 186.705 108.130 186.985 109.130 ;
        RECT 187.135 108.130 187.415 109.130 ;
        RECT 187.565 108.130 187.845 109.130 ;
        RECT 187.995 108.130 188.275 109.130 ;
        RECT 188.425 108.130 188.705 109.130 ;
        RECT 188.855 108.130 189.135 109.130 ;
        RECT 189.285 108.130 189.565 109.130 ;
        RECT 189.715 108.130 189.995 109.130 ;
        RECT 190.155 107.085 190.415 109.130 ;
        RECT 190.575 108.130 190.855 109.130 ;
        RECT 191.030 107.085 191.290 109.130 ;
        RECT 191.435 108.130 191.715 109.130 ;
        RECT 191.890 107.085 192.150 109.130 ;
        RECT 192.295 108.130 192.575 109.130 ;
        RECT 192.750 107.085 193.010 109.130 ;
        RECT 193.155 108.130 193.435 109.130 ;
        RECT 193.585 108.130 193.865 109.130 ;
        RECT 194.015 108.130 194.295 109.130 ;
        RECT 194.445 108.130 194.725 109.130 ;
        RECT 194.875 108.130 195.155 109.130 ;
        RECT 195.305 108.130 195.585 109.130 ;
        RECT 195.735 108.130 196.015 109.130 ;
        RECT 196.165 108.130 196.445 109.130 ;
        RECT 196.595 108.130 196.875 109.130 ;
        RECT 197.025 108.130 197.305 109.130 ;
        RECT 197.455 107.515 197.735 112.205 ;
        RECT 198.120 110.160 198.410 111.160 ;
        RECT 198.760 110.680 199.090 112.205 ;
        RECT 199.820 111.345 200.110 112.195 ;
        RECT 200.495 111.345 200.775 112.195 ;
        RECT 200.925 111.345 201.205 112.195 ;
        RECT 200.290 110.680 200.995 111.050 ;
        RECT 201.355 109.840 201.635 112.195 ;
        RECT 198.120 108.130 198.410 109.130 ;
        RECT 201.785 108.705 202.065 112.195 ;
        RECT 202.230 109.860 202.510 112.195 ;
        RECT 202.660 108.705 202.940 112.195 ;
        RECT 203.090 109.860 203.370 112.195 ;
        RECT 203.520 108.705 203.800 112.195 ;
        RECT 203.950 109.860 204.230 112.195 ;
        RECT 204.380 108.705 204.660 112.195 ;
        RECT 196.775 107.235 197.735 107.515 ;
        RECT 198.760 107.085 199.090 108.610 ;
        RECT 200.290 108.240 200.995 108.610 ;
        RECT 199.820 107.095 200.110 107.945 ;
        RECT 200.495 107.095 200.775 107.945 ;
        RECT 200.925 107.095 201.205 107.945 ;
        RECT 201.355 107.095 201.635 107.945 ;
        RECT 201.785 107.095 202.065 107.945 ;
        RECT 202.215 107.095 202.495 107.945 ;
        RECT 202.645 107.095 202.925 107.945 ;
        RECT 203.075 107.095 203.355 107.945 ;
        RECT 203.505 107.095 203.785 107.945 ;
        RECT 203.935 107.095 204.215 107.945 ;
        RECT 204.365 107.095 204.645 107.945 ;
        RECT 204.810 107.095 205.090 112.195 ;
        RECT 205.240 107.095 205.520 112.195 ;
        RECT 205.670 107.095 205.950 112.195 ;
        RECT 206.100 107.095 206.380 112.195 ;
        RECT 206.530 107.095 206.810 112.195 ;
        RECT 206.960 107.095 207.240 112.195 ;
        RECT 207.390 107.095 207.670 112.195 ;
        RECT 207.820 107.095 208.100 112.195 ;
        RECT 208.240 110.610 208.520 112.195 ;
        RECT 208.240 109.840 208.530 110.610 ;
        RECT 208.240 107.095 208.520 109.840 ;
        RECT 208.680 108.705 208.960 112.195 ;
        RECT 209.110 109.860 209.390 112.195 ;
        RECT 209.540 108.705 209.820 112.195 ;
        RECT 209.970 109.860 210.250 112.195 ;
        RECT 210.400 108.705 210.680 112.195 ;
        RECT 210.830 109.860 211.110 112.195 ;
        RECT 211.260 108.705 211.540 112.195 ;
        RECT 211.680 110.630 211.960 112.195 ;
        RECT 212.105 111.345 212.385 112.195 ;
        RECT 212.535 111.345 212.815 112.195 ;
        RECT 213.200 111.345 213.490 112.195 ;
        RECT 211.680 109.860 211.970 110.630 ;
        RECT 208.665 107.095 208.945 107.945 ;
        RECT 209.095 107.095 209.375 107.945 ;
        RECT 209.525 107.095 209.805 107.945 ;
        RECT 209.955 107.095 210.235 107.945 ;
        RECT 210.385 107.095 210.665 107.945 ;
        RECT 210.815 107.095 211.095 107.945 ;
        RECT 211.245 107.095 211.525 107.945 ;
        RECT 211.675 107.095 211.955 107.945 ;
        RECT 212.105 107.095 212.385 107.945 ;
        RECT 212.535 107.095 212.815 107.945 ;
        RECT 213.200 107.095 213.490 107.945 ;
        RECT 186.690 106.755 199.090 107.085 ;
        RECT 184.740 104.705 185.030 105.705 ;
        RECT 185.415 104.705 185.695 105.705 ;
        RECT 185.845 104.705 186.125 105.705 ;
        RECT 186.275 104.705 186.555 105.705 ;
        RECT 186.700 104.705 186.960 106.755 ;
        RECT 187.135 104.705 187.415 105.705 ;
        RECT 187.560 104.705 187.820 106.755 ;
        RECT 187.995 104.705 188.275 105.705 ;
        RECT 188.420 104.705 188.680 106.755 ;
        RECT 188.855 104.705 189.135 105.705 ;
        RECT 189.280 104.705 189.540 106.755 ;
        RECT 189.715 104.705 189.995 105.705 ;
        RECT 190.155 104.705 190.415 106.755 ;
        RECT 190.575 104.705 190.855 105.705 ;
        RECT 191.030 104.705 191.290 106.755 ;
        RECT 191.435 104.705 191.715 105.705 ;
        RECT 191.890 104.705 192.150 106.755 ;
        RECT 192.295 104.705 192.575 105.705 ;
        RECT 192.750 104.705 193.010 106.755 ;
        RECT 193.155 104.705 193.435 105.705 ;
        RECT 193.610 104.705 193.870 106.755 ;
        RECT 194.015 104.705 194.295 105.705 ;
        RECT 194.470 104.705 194.730 106.755 ;
        RECT 194.875 104.705 195.155 105.705 ;
        RECT 195.330 104.705 195.590 106.755 ;
        RECT 195.735 104.705 196.015 105.705 ;
        RECT 196.190 104.705 196.450 106.755 ;
        RECT 196.595 104.705 196.875 105.705 ;
        RECT 197.025 104.705 197.305 105.705 ;
        RECT 197.455 104.705 197.735 105.705 ;
        RECT 198.120 104.705 198.410 105.705 ;
        RECT 184.740 101.085 185.030 102.085 ;
        RECT 185.415 101.085 185.695 102.085 ;
        RECT 185.845 101.085 186.125 102.085 ;
        RECT 186.275 101.085 186.555 102.085 ;
        RECT 186.700 100.035 186.960 102.085 ;
        RECT 187.135 101.085 187.415 102.085 ;
        RECT 187.560 100.035 187.820 102.085 ;
        RECT 187.995 101.085 188.275 102.085 ;
        RECT 188.420 100.035 188.680 102.085 ;
        RECT 188.855 101.085 189.135 102.085 ;
        RECT 189.280 100.035 189.540 102.085 ;
        RECT 189.715 101.085 189.995 102.085 ;
        RECT 190.155 100.035 190.415 102.085 ;
        RECT 190.575 101.085 190.855 102.085 ;
        RECT 191.030 100.035 191.290 102.085 ;
        RECT 191.435 101.085 191.715 102.085 ;
        RECT 191.890 100.035 192.150 102.085 ;
        RECT 192.295 101.085 192.575 102.085 ;
        RECT 192.750 100.035 193.010 102.085 ;
        RECT 193.155 101.085 193.435 102.085 ;
        RECT 193.610 100.035 193.870 102.085 ;
        RECT 194.015 101.085 194.295 102.085 ;
        RECT 194.470 100.035 194.730 102.085 ;
        RECT 194.875 101.085 195.155 102.085 ;
        RECT 195.330 100.035 195.590 102.085 ;
        RECT 195.735 101.085 196.015 102.085 ;
        RECT 196.190 100.035 196.450 102.085 ;
        RECT 196.595 101.085 196.875 102.085 ;
        RECT 197.025 101.085 197.305 102.085 ;
        RECT 197.455 101.085 197.735 102.085 ;
        RECT 198.120 101.085 198.410 102.085 ;
        RECT 186.690 99.705 199.090 100.035 ;
        RECT 184.740 97.660 185.030 98.660 ;
        RECT 185.415 97.660 185.695 98.660 ;
        RECT 185.845 97.660 186.125 98.660 ;
        RECT 186.275 97.660 186.555 98.660 ;
        RECT 186.705 97.660 186.985 98.660 ;
        RECT 187.135 97.660 187.415 98.660 ;
        RECT 187.565 97.660 187.845 98.660 ;
        RECT 187.995 97.660 188.275 98.660 ;
        RECT 188.425 97.660 188.705 98.660 ;
        RECT 188.855 97.660 189.135 98.660 ;
        RECT 189.285 97.660 189.565 98.660 ;
        RECT 189.715 97.660 189.995 98.660 ;
        RECT 190.155 97.660 190.415 99.705 ;
        RECT 190.575 97.660 190.855 98.660 ;
        RECT 191.030 97.660 191.290 99.705 ;
        RECT 191.435 97.660 191.715 98.660 ;
        RECT 191.890 97.660 192.150 99.705 ;
        RECT 192.295 97.660 192.575 98.660 ;
        RECT 192.750 97.660 193.010 99.705 ;
        RECT 196.775 99.275 197.735 99.555 ;
        RECT 193.155 97.660 193.435 98.660 ;
        RECT 193.585 97.660 193.865 98.660 ;
        RECT 194.015 97.660 194.295 98.660 ;
        RECT 194.445 97.660 194.725 98.660 ;
        RECT 194.875 97.660 195.155 98.660 ;
        RECT 195.305 97.660 195.585 98.660 ;
        RECT 195.735 97.660 196.015 98.660 ;
        RECT 196.165 97.660 196.445 98.660 ;
        RECT 196.595 97.660 196.875 98.660 ;
        RECT 197.025 97.660 197.305 98.660 ;
        RECT 184.740 95.630 185.030 96.630 ;
        RECT 185.415 95.630 185.695 96.630 ;
        RECT 185.845 95.630 186.125 96.630 ;
        RECT 186.275 95.630 186.555 96.630 ;
        RECT 186.705 95.630 186.985 96.630 ;
        RECT 187.135 95.630 187.415 96.630 ;
        RECT 187.565 95.630 187.845 96.630 ;
        RECT 187.995 95.630 188.275 96.630 ;
        RECT 188.425 95.630 188.705 96.630 ;
        RECT 188.855 95.630 189.135 96.630 ;
        RECT 189.285 95.630 189.565 96.630 ;
        RECT 189.715 95.630 189.995 96.630 ;
        RECT 190.155 94.585 190.415 96.630 ;
        RECT 190.575 95.630 190.855 96.630 ;
        RECT 191.030 94.585 191.290 96.630 ;
        RECT 191.435 95.630 191.715 96.630 ;
        RECT 191.890 94.585 192.150 96.630 ;
        RECT 192.295 95.630 192.575 96.630 ;
        RECT 192.750 94.585 193.010 96.630 ;
        RECT 193.155 95.630 193.435 96.630 ;
        RECT 193.585 95.630 193.865 96.630 ;
        RECT 194.015 95.630 194.295 96.630 ;
        RECT 194.445 95.630 194.725 96.630 ;
        RECT 194.875 95.630 195.155 96.630 ;
        RECT 195.305 95.630 195.585 96.630 ;
        RECT 195.735 95.630 196.015 96.630 ;
        RECT 196.165 95.630 196.445 96.630 ;
        RECT 196.595 95.630 196.875 96.630 ;
        RECT 197.025 95.630 197.305 96.630 ;
        RECT 197.455 94.585 197.735 99.275 ;
        RECT 198.120 97.660 198.410 98.660 ;
        RECT 198.760 98.180 199.090 99.705 ;
        RECT 199.820 98.845 200.110 99.695 ;
        RECT 200.495 98.845 200.775 99.695 ;
        RECT 200.925 98.845 201.205 99.695 ;
        RECT 201.355 98.845 201.635 99.695 ;
        RECT 201.785 98.845 202.065 99.695 ;
        RECT 202.215 98.845 202.495 99.695 ;
        RECT 202.645 98.845 202.925 99.695 ;
        RECT 203.075 98.845 203.355 99.695 ;
        RECT 203.505 98.845 203.785 99.695 ;
        RECT 203.935 98.845 204.215 99.695 ;
        RECT 204.365 98.845 204.645 99.695 ;
        RECT 200.290 98.180 200.995 98.550 ;
        RECT 198.120 95.630 198.410 96.630 ;
        RECT 198.760 94.585 199.090 96.110 ;
        RECT 200.290 95.740 200.995 96.110 ;
        RECT 199.820 94.595 200.110 95.445 ;
        RECT 200.495 94.595 200.775 95.445 ;
        RECT 200.925 94.595 201.205 95.445 ;
        RECT 201.355 94.595 201.635 96.950 ;
        RECT 201.785 94.595 202.065 98.085 ;
        RECT 202.230 94.595 202.510 96.930 ;
        RECT 202.660 94.595 202.940 98.085 ;
        RECT 203.090 94.595 203.370 96.930 ;
        RECT 203.520 94.595 203.800 98.085 ;
        RECT 203.950 94.595 204.230 96.930 ;
        RECT 204.380 94.595 204.660 98.085 ;
        RECT 204.810 94.595 205.090 99.695 ;
        RECT 205.240 94.595 205.520 99.695 ;
        RECT 205.670 94.595 205.950 99.695 ;
        RECT 206.100 94.595 206.380 99.695 ;
        RECT 206.530 94.595 206.810 99.695 ;
        RECT 206.960 94.595 207.240 99.695 ;
        RECT 207.390 94.595 207.670 99.695 ;
        RECT 207.820 94.595 208.100 99.695 ;
        RECT 208.240 96.950 208.520 99.695 ;
        RECT 208.665 98.845 208.945 99.695 ;
        RECT 209.095 98.845 209.375 99.695 ;
        RECT 209.525 98.845 209.805 99.695 ;
        RECT 209.955 98.845 210.235 99.695 ;
        RECT 210.385 98.845 210.665 99.695 ;
        RECT 210.815 98.845 211.095 99.695 ;
        RECT 211.245 98.845 211.525 99.695 ;
        RECT 211.675 98.845 211.955 99.695 ;
        RECT 212.105 98.845 212.385 99.695 ;
        RECT 212.535 98.845 212.815 99.695 ;
        RECT 213.200 98.845 213.490 99.695 ;
        RECT 208.240 96.180 208.530 96.950 ;
        RECT 208.240 94.595 208.520 96.180 ;
        RECT 208.680 94.595 208.960 98.085 ;
        RECT 209.110 94.595 209.390 96.930 ;
        RECT 209.540 94.595 209.820 98.085 ;
        RECT 209.970 94.595 210.250 96.930 ;
        RECT 210.400 94.595 210.680 98.085 ;
        RECT 210.830 94.595 211.110 96.930 ;
        RECT 211.260 94.595 211.540 98.085 ;
        RECT 214.090 97.335 214.420 116.325 ;
        RECT 222.030 115.305 223.340 116.305 ;
        RECT 214.820 105.690 215.150 109.455 ;
        RECT 215.550 100.065 215.880 110.190 ;
        RECT 217.110 108.145 217.400 110.145 ;
        RECT 225.200 106.675 226.200 120.945 ;
        RECT 290.280 108.145 290.570 110.145 ;
        RECT 225.060 105.745 226.340 106.675 ;
        RECT 240.120 105.710 243.440 106.710 ;
        RECT 225.060 100.120 226.340 101.050 ;
        RECT 211.680 96.160 211.970 96.930 ;
        RECT 211.680 94.595 211.960 96.160 ;
        RECT 212.105 94.595 212.385 95.445 ;
        RECT 212.535 94.595 212.815 95.445 ;
        RECT 213.200 94.595 213.490 95.445 ;
        RECT 185.490 94.255 186.330 94.585 ;
        RECT 186.690 94.255 199.090 94.585 ;
        RECT 184.740 92.205 185.030 93.205 ;
        RECT 185.415 92.205 185.695 93.205 ;
        RECT 185.845 92.205 186.125 93.205 ;
        RECT 186.275 92.205 186.555 93.205 ;
        RECT 186.700 92.205 186.960 94.255 ;
        RECT 187.135 92.205 187.415 93.205 ;
        RECT 187.560 92.205 187.820 94.255 ;
        RECT 187.995 92.205 188.275 93.205 ;
        RECT 188.420 92.205 188.680 94.255 ;
        RECT 188.855 92.205 189.135 93.205 ;
        RECT 189.280 92.205 189.540 94.255 ;
        RECT 189.715 92.205 189.995 93.205 ;
        RECT 190.155 92.205 190.415 94.255 ;
        RECT 190.575 92.205 190.855 93.205 ;
        RECT 191.030 92.205 191.290 94.255 ;
        RECT 191.435 92.205 191.715 93.205 ;
        RECT 191.890 92.205 192.150 94.255 ;
        RECT 192.295 92.205 192.575 93.205 ;
        RECT 192.750 92.205 193.010 94.255 ;
        RECT 193.155 92.205 193.435 93.205 ;
        RECT 193.610 92.205 193.870 94.255 ;
        RECT 194.015 92.205 194.295 93.205 ;
        RECT 194.470 92.205 194.730 94.255 ;
        RECT 194.875 92.205 195.155 93.205 ;
        RECT 195.330 92.205 195.590 94.255 ;
        RECT 195.735 92.205 196.015 93.205 ;
        RECT 196.190 92.205 196.450 94.255 ;
        RECT 196.595 92.205 196.875 93.205 ;
        RECT 197.025 92.205 197.305 93.205 ;
        RECT 197.455 92.205 197.735 93.205 ;
        RECT 198.120 92.205 198.410 93.205 ;
        RECT 214.090 90.470 214.420 96.930 ;
        RECT 217.110 96.645 217.400 98.645 ;
        RECT 222.030 90.490 223.340 91.490 ;
        RECT 225.200 85.845 226.200 100.120 ;
        RECT 240.120 100.085 243.440 101.085 ;
        RECT 284.495 100.085 285.495 106.710 ;
        RECT 299.055 105.680 299.655 138.360 ;
        RECT 305.240 135.895 308.560 136.895 ;
        RECT 309.260 135.895 312.580 136.895 ;
        RECT 313.280 135.895 316.600 136.895 ;
        RECT 317.300 135.895 320.620 136.895 ;
        RECT 321.320 135.895 324.640 136.895 ;
        RECT 325.340 135.895 328.660 136.895 ;
        RECT 329.360 135.895 332.680 136.895 ;
        RECT 333.380 135.895 336.700 136.895 ;
        RECT 337.400 135.895 340.720 136.895 ;
        RECT 341.420 135.895 344.740 136.895 ;
        RECT 345.440 135.895 348.760 136.895 ;
        RECT 349.460 135.895 352.780 136.895 ;
        RECT 353.480 135.895 356.800 136.895 ;
        RECT 357.500 135.895 360.820 136.895 ;
        RECT 361.520 135.895 364.840 136.895 ;
        RECT 365.540 135.895 368.860 136.895 ;
        RECT 369.560 135.895 372.880 136.895 ;
        RECT 373.580 135.895 376.900 136.895 ;
        RECT 377.600 135.895 380.920 136.895 ;
        RECT 381.620 135.895 384.940 136.895 ;
        RECT 385.640 135.895 388.960 136.895 ;
        RECT 389.660 135.895 392.980 136.895 ;
        RECT 393.680 135.895 397.000 136.895 ;
        RECT 397.700 135.895 401.020 136.895 ;
        RECT 401.720 135.895 405.040 136.895 ;
        RECT 300.325 130.610 300.605 132.610 ;
        RECT 409.675 130.610 409.955 132.610 ;
        RECT 305.240 126.300 306.550 127.300 ;
        RECT 307.250 126.300 310.570 127.300 ;
        RECT 311.270 126.300 314.590 127.300 ;
        RECT 315.290 126.300 318.610 127.300 ;
        RECT 319.310 126.300 322.630 127.300 ;
        RECT 323.330 126.300 326.650 127.300 ;
        RECT 327.350 126.300 330.670 127.300 ;
        RECT 331.370 126.300 334.690 127.300 ;
        RECT 335.390 126.300 338.710 127.300 ;
        RECT 339.410 126.300 342.730 127.300 ;
        RECT 343.430 126.300 346.750 127.300 ;
        RECT 347.450 126.300 350.770 127.300 ;
        RECT 351.470 126.300 354.790 127.300 ;
        RECT 355.490 126.300 358.810 127.300 ;
        RECT 359.510 126.300 362.830 127.300 ;
        RECT 363.530 126.300 366.850 127.300 ;
        RECT 367.550 126.300 370.870 127.300 ;
        RECT 371.570 126.300 374.890 127.300 ;
        RECT 375.590 126.300 378.910 127.300 ;
        RECT 379.610 126.300 382.930 127.300 ;
        RECT 383.630 126.300 386.950 127.300 ;
        RECT 387.650 126.300 390.970 127.300 ;
        RECT 391.670 126.300 394.990 127.300 ;
        RECT 395.690 126.300 399.010 127.300 ;
        RECT 399.710 126.300 403.030 127.300 ;
        RECT 403.730 126.300 405.040 127.300 ;
        RECT 410.770 124.385 411.370 127.300 ;
        RECT 410.290 123.785 411.370 124.385 ;
        RECT 406.435 122.345 407.605 122.675 ;
        RECT 351.330 121.685 352.010 122.055 ;
        RECT 353.090 121.685 353.770 122.055 ;
        RECT 354.850 121.685 355.530 122.055 ;
        RECT 356.610 121.685 357.290 122.055 ;
        RECT 318.995 119.825 320.390 120.155 ;
        RECT 310.855 118.005 311.145 119.005 ;
        RECT 311.590 118.005 311.870 119.005 ;
        RECT 312.470 118.005 312.750 119.005 ;
        RECT 313.350 118.005 313.630 119.005 ;
        RECT 314.230 118.005 314.510 119.005 ;
        RECT 315.110 118.005 315.390 119.005 ;
        RECT 315.990 118.005 316.270 119.005 ;
        RECT 316.870 118.005 317.150 119.005 ;
        RECT 317.750 118.005 318.030 119.005 ;
        RECT 318.630 118.005 318.910 119.005 ;
        RECT 319.510 115.515 319.790 119.635 ;
        RECT 320.390 118.005 320.670 119.005 ;
        RECT 321.270 115.515 321.550 119.635 ;
        RECT 322.150 118.005 322.430 119.005 ;
        RECT 323.030 115.515 323.310 119.635 ;
        RECT 323.910 118.005 324.190 119.005 ;
        RECT 324.790 115.515 325.070 119.635 ;
        RECT 325.670 118.005 325.950 119.005 ;
        RECT 326.550 118.005 326.830 119.005 ;
        RECT 327.430 118.005 327.710 119.005 ;
        RECT 328.310 118.005 328.590 119.005 ;
        RECT 329.190 118.005 329.470 119.005 ;
        RECT 330.070 118.005 330.350 119.005 ;
        RECT 330.950 118.005 331.230 119.005 ;
        RECT 331.830 118.005 332.110 119.005 ;
        RECT 332.710 118.005 332.990 119.005 ;
        RECT 333.435 118.005 333.725 119.005 ;
        RECT 334.075 118.005 334.365 119.005 ;
        RECT 334.810 118.005 335.090 119.005 ;
        RECT 335.690 118.005 335.970 119.005 ;
        RECT 336.570 118.005 336.850 119.005 ;
        RECT 337.450 118.005 337.730 119.005 ;
        RECT 338.330 118.005 338.610 119.005 ;
        RECT 339.210 118.005 339.490 119.005 ;
        RECT 340.090 118.005 340.370 119.005 ;
        RECT 319.510 115.015 325.070 115.515 ;
        RECT 318.975 113.340 319.370 113.670 ;
        RECT 310.855 111.520 311.145 112.520 ;
        RECT 311.590 111.520 311.870 112.520 ;
        RECT 312.470 111.520 312.750 112.520 ;
        RECT 313.350 111.520 313.630 112.520 ;
        RECT 314.230 111.520 314.510 112.520 ;
        RECT 315.110 111.520 315.390 112.520 ;
        RECT 315.990 111.520 316.270 112.520 ;
        RECT 316.870 111.520 317.150 112.520 ;
        RECT 317.750 111.520 318.030 112.520 ;
        RECT 318.630 107.385 318.910 113.150 ;
        RECT 319.510 110.890 319.790 115.015 ;
        RECT 319.930 113.340 321.130 113.670 ;
        RECT 320.390 107.385 320.670 113.150 ;
        RECT 321.270 110.890 321.550 115.015 ;
        RECT 321.690 113.340 322.890 113.670 ;
        RECT 322.150 107.385 322.430 113.150 ;
        RECT 323.030 110.890 323.310 115.015 ;
        RECT 323.450 113.340 324.650 113.670 ;
        RECT 323.910 107.385 324.190 113.150 ;
        RECT 324.790 110.890 325.070 115.015 ;
        RECT 325.210 113.340 325.585 113.670 ;
        RECT 337.730 113.340 339.490 113.670 ;
        RECT 325.670 107.385 325.950 113.150 ;
        RECT 326.550 111.520 326.830 112.520 ;
        RECT 327.430 111.520 327.710 112.520 ;
        RECT 328.310 111.520 328.590 112.520 ;
        RECT 329.190 111.520 329.470 112.520 ;
        RECT 330.070 111.520 330.350 112.520 ;
        RECT 330.950 111.520 331.230 112.520 ;
        RECT 331.830 111.520 332.110 112.520 ;
        RECT 332.710 111.520 332.990 112.520 ;
        RECT 333.435 111.520 333.725 112.520 ;
        RECT 334.075 111.520 334.365 112.520 ;
        RECT 334.810 111.520 335.090 112.520 ;
        RECT 335.690 111.520 335.970 112.520 ;
        RECT 336.570 111.520 336.850 112.520 ;
        RECT 337.450 111.520 337.730 112.520 ;
        RECT 338.330 111.520 338.610 112.520 ;
        RECT 339.210 111.520 339.490 112.520 ;
        RECT 315.110 106.885 329.470 107.385 ;
        RECT 299.055 105.310 300.160 105.680 ;
        RECT 311.955 105.320 313.620 105.610 ;
        RECT 310.855 102.910 311.145 103.910 ;
        RECT 311.590 102.910 311.870 103.910 ;
        RECT 312.470 102.910 312.750 103.910 ;
        RECT 313.350 102.910 313.630 103.910 ;
        RECT 314.230 102.910 314.510 103.910 ;
        RECT 315.110 102.280 315.390 106.885 ;
        RECT 299.055 101.130 300.160 101.500 ;
        RECT 311.955 101.210 313.620 101.500 ;
        RECT 290.280 96.645 290.570 98.645 ;
        RECT 178.380 32.295 178.980 56.010 ;
        RECT 183.180 36.385 183.780 85.845 ;
        RECT 225.160 85.245 226.240 85.845 ;
        RECT 294.895 85.245 295.975 85.845 ;
        RECT 189.705 79.490 191.015 80.490 ;
        RECT 191.715 79.490 195.035 80.490 ;
        RECT 195.735 79.490 199.055 80.490 ;
        RECT 199.755 79.490 203.075 80.490 ;
        RECT 203.775 79.490 207.095 80.490 ;
        RECT 207.795 79.490 211.115 80.490 ;
        RECT 211.815 79.490 215.135 80.490 ;
        RECT 215.835 79.490 219.155 80.490 ;
        RECT 219.855 79.490 223.175 80.490 ;
        RECT 223.875 79.490 227.195 80.490 ;
        RECT 227.895 79.490 231.215 80.490 ;
        RECT 231.915 79.490 235.235 80.490 ;
        RECT 235.935 79.490 239.255 80.490 ;
        RECT 239.955 79.490 243.275 80.490 ;
        RECT 243.975 79.490 247.295 80.490 ;
        RECT 247.995 79.490 251.315 80.490 ;
        RECT 252.015 79.490 255.335 80.490 ;
        RECT 256.035 79.490 259.355 80.490 ;
        RECT 260.055 79.490 263.375 80.490 ;
        RECT 264.075 79.490 267.395 80.490 ;
        RECT 268.095 79.490 271.415 80.490 ;
        RECT 272.115 79.490 275.435 80.490 ;
        RECT 276.135 79.490 279.455 80.490 ;
        RECT 280.155 79.490 283.475 80.490 ;
        RECT 284.175 79.490 287.495 80.490 ;
        RECT 288.195 79.490 289.505 80.490 ;
        RECT 295.375 79.490 295.975 85.245 ;
        RECT 184.790 74.180 185.070 76.180 ;
        RECT 294.140 74.180 294.420 76.180 ;
        RECT 189.705 69.895 193.025 70.895 ;
        RECT 193.725 69.895 197.045 70.895 ;
        RECT 197.745 69.895 201.065 70.895 ;
        RECT 201.765 69.895 205.085 70.895 ;
        RECT 205.785 69.895 209.105 70.895 ;
        RECT 209.805 69.895 213.125 70.895 ;
        RECT 213.825 69.895 217.145 70.895 ;
        RECT 217.845 69.895 221.165 70.895 ;
        RECT 221.865 69.895 225.185 70.895 ;
        RECT 225.885 69.895 229.205 70.895 ;
        RECT 229.905 69.895 233.225 70.895 ;
        RECT 233.925 69.895 237.245 70.895 ;
        RECT 237.945 69.895 241.265 70.895 ;
        RECT 241.965 69.895 245.285 70.895 ;
        RECT 245.985 69.895 249.305 70.895 ;
        RECT 250.005 69.895 253.325 70.895 ;
        RECT 254.025 69.895 257.345 70.895 ;
        RECT 258.045 69.895 261.365 70.895 ;
        RECT 262.065 69.895 265.385 70.895 ;
        RECT 266.085 69.895 269.405 70.895 ;
        RECT 270.105 69.895 273.425 70.895 ;
        RECT 274.125 69.895 277.445 70.895 ;
        RECT 278.145 69.895 281.465 70.895 ;
        RECT 282.165 69.895 285.485 70.895 ;
        RECT 286.185 69.895 289.505 70.895 ;
        RECT 299.055 68.430 299.655 101.130 ;
        RECT 315.990 97.705 316.270 104.540 ;
        RECT 316.870 102.280 317.150 106.885 ;
        RECT 315.790 97.335 316.470 97.705 ;
        RECT 315.990 96.725 316.270 97.335 ;
        RECT 317.750 97.075 318.030 104.540 ;
        RECT 318.630 102.280 318.910 106.885 ;
        RECT 319.510 97.705 319.790 104.540 ;
        RECT 320.390 102.280 320.670 106.885 ;
        RECT 319.310 97.335 319.990 97.705 ;
        RECT 317.570 96.705 318.250 97.075 ;
        RECT 319.510 96.725 319.790 97.335 ;
        RECT 321.270 97.075 321.550 104.540 ;
        RECT 322.150 102.280 322.430 106.885 ;
        RECT 323.030 97.705 323.310 104.540 ;
        RECT 323.910 102.280 324.190 106.885 ;
        RECT 322.830 97.335 323.510 97.705 ;
        RECT 321.090 96.705 321.770 97.075 ;
        RECT 323.030 96.725 323.310 97.335 ;
        RECT 324.790 97.075 325.070 104.540 ;
        RECT 325.670 102.280 325.950 106.885 ;
        RECT 326.550 97.705 326.830 104.540 ;
        RECT 327.430 102.280 327.710 106.885 ;
        RECT 326.350 97.335 327.030 97.705 ;
        RECT 324.610 96.705 325.290 97.075 ;
        RECT 326.550 96.725 326.830 97.335 ;
        RECT 328.310 97.075 328.590 104.540 ;
        RECT 329.190 102.280 329.470 106.885 ;
        RECT 330.070 102.910 330.350 103.910 ;
        RECT 330.950 102.910 331.230 103.910 ;
        RECT 331.830 102.910 332.110 103.910 ;
        RECT 332.710 102.910 332.990 103.910 ;
        RECT 333.435 102.910 333.725 103.910 ;
        RECT 334.115 102.400 334.405 104.400 ;
        RECT 334.810 102.400 335.090 104.400 ;
        RECT 335.690 102.400 335.970 104.400 ;
        RECT 336.570 102.400 336.850 104.400 ;
        RECT 337.450 102.400 337.730 104.400 ;
        RECT 338.330 102.400 338.610 104.400 ;
        RECT 339.210 102.400 339.490 104.400 ;
        RECT 340.090 98.885 340.370 115.070 ;
        RECT 340.970 110.890 341.250 119.635 ;
        RECT 341.850 118.005 342.130 119.005 ;
        RECT 340.655 108.105 341.505 108.435 ;
        RECT 340.970 97.705 341.250 107.915 ;
        RECT 341.850 98.885 342.130 115.070 ;
        RECT 342.730 110.890 343.010 119.635 ;
        RECT 343.610 118.005 343.890 119.005 ;
        RECT 343.460 116.880 344.040 117.200 ;
        RECT 343.500 114.550 344.000 116.880 ;
        RECT 342.270 108.105 343.470 108.435 ;
        RECT 342.730 97.705 343.010 107.915 ;
        RECT 343.610 98.885 343.890 114.550 ;
        RECT 344.490 110.890 344.770 119.635 ;
        RECT 345.370 118.005 345.650 119.005 ;
        RECT 344.030 108.105 345.230 108.435 ;
        RECT 344.490 97.705 344.770 107.915 ;
        RECT 345.370 98.885 345.650 115.070 ;
        RECT 346.250 110.890 346.530 119.635 ;
        RECT 347.130 118.005 347.410 119.005 ;
        RECT 348.010 118.005 348.290 119.005 ;
        RECT 348.890 118.005 349.170 119.005 ;
        RECT 349.770 118.005 350.050 119.005 ;
        RECT 350.650 118.005 350.930 119.005 ;
        RECT 345.790 108.105 346.990 108.435 ;
        RECT 346.250 97.705 346.530 107.915 ;
        RECT 347.130 98.885 347.410 115.070 ;
        RECT 348.010 111.520 348.290 112.520 ;
        RECT 348.890 111.520 349.170 112.520 ;
        RECT 349.770 111.520 350.050 112.520 ;
        RECT 348.010 102.400 348.290 104.400 ;
        RECT 348.890 102.400 349.170 104.400 ;
        RECT 349.770 102.400 350.050 104.400 ;
        RECT 350.650 98.885 350.930 115.070 ;
        RECT 351.530 110.890 351.810 121.685 ;
        RECT 352.410 118.005 352.690 119.005 ;
        RECT 351.070 108.105 352.270 108.435 ;
        RECT 339.010 97.335 339.690 97.705 ;
        RECT 340.770 97.335 341.450 97.705 ;
        RECT 342.530 97.335 343.210 97.705 ;
        RECT 344.290 97.335 344.970 97.705 ;
        RECT 346.050 97.335 346.730 97.705 ;
        RECT 347.810 97.335 348.490 97.705 ;
        RECT 328.130 96.705 328.810 97.075 ;
        RECT 334.115 90.040 334.405 92.040 ;
        RECT 334.810 90.040 335.090 92.040 ;
        RECT 335.690 90.040 335.970 92.040 ;
        RECT 336.570 90.040 336.850 92.040 ;
        RECT 337.450 90.040 337.730 92.040 ;
        RECT 338.330 90.040 338.610 92.040 ;
        RECT 339.210 86.520 339.490 97.335 ;
        RECT 340.090 90.040 340.370 92.040 ;
        RECT 340.970 86.520 341.250 97.335 ;
        RECT 341.850 90.040 342.130 92.040 ;
        RECT 342.730 86.520 343.010 97.335 ;
        RECT 343.610 90.040 343.890 92.040 ;
        RECT 344.490 86.520 344.770 97.335 ;
        RECT 345.370 90.040 345.650 92.040 ;
        RECT 346.250 86.520 346.530 97.335 ;
        RECT 347.130 90.040 347.410 92.040 ;
        RECT 348.010 86.520 348.290 97.335 ;
        RECT 349.770 97.075 350.050 97.685 ;
        RECT 351.530 97.075 351.810 107.915 ;
        RECT 352.410 98.885 352.690 115.070 ;
        RECT 353.290 110.890 353.570 121.685 ;
        RECT 354.170 118.005 354.450 119.005 ;
        RECT 352.830 108.105 354.030 108.435 ;
        RECT 353.290 97.075 353.570 107.915 ;
        RECT 354.170 98.885 354.450 115.070 ;
        RECT 355.050 110.890 355.330 121.685 ;
        RECT 355.930 118.005 356.210 119.005 ;
        RECT 354.590 108.105 355.790 108.435 ;
        RECT 355.050 97.075 355.330 107.915 ;
        RECT 355.930 98.885 356.210 115.070 ;
        RECT 356.810 110.890 357.090 121.685 ;
        RECT 357.690 118.005 357.970 119.005 ;
        RECT 358.570 118.005 358.850 119.005 ;
        RECT 359.450 118.005 359.730 119.005 ;
        RECT 360.330 118.005 360.610 119.005 ;
        RECT 361.210 118.005 361.490 119.005 ;
        RECT 362.090 118.005 362.370 119.005 ;
        RECT 362.970 118.005 363.250 119.005 ;
        RECT 363.695 118.005 363.985 119.005 ;
        RECT 364.415 118.005 364.705 119.005 ;
        RECT 365.150 118.005 365.430 119.005 ;
        RECT 366.030 118.005 366.310 119.005 ;
        RECT 366.910 118.005 367.190 119.005 ;
        RECT 367.790 115.515 368.070 119.635 ;
        RECT 368.670 118.005 368.950 119.005 ;
        RECT 368.425 116.895 369.195 117.185 ;
        RECT 369.550 115.515 369.830 119.635 ;
        RECT 370.430 118.005 370.710 119.005 ;
        RECT 371.310 115.515 371.590 119.635 ;
        RECT 372.190 118.005 372.470 119.005 ;
        RECT 373.070 115.515 373.350 119.635 ;
        RECT 373.950 118.005 374.230 119.005 ;
        RECT 374.830 115.515 375.110 119.635 ;
        RECT 375.710 118.005 375.990 119.005 ;
        RECT 376.590 115.515 376.870 119.635 ;
        RECT 377.470 118.005 377.750 119.005 ;
        RECT 378.350 115.515 378.630 119.635 ;
        RECT 379.230 118.005 379.510 119.005 ;
        RECT 380.110 115.515 380.390 119.635 ;
        RECT 380.990 118.005 381.270 119.005 ;
        RECT 381.870 115.515 382.150 119.635 ;
        RECT 382.750 118.005 383.030 119.005 ;
        RECT 383.630 115.515 383.910 119.635 ;
        RECT 384.510 118.005 384.790 119.005 ;
        RECT 385.390 115.515 385.670 119.635 ;
        RECT 386.270 118.005 386.550 119.005 ;
        RECT 387.150 115.515 387.430 119.635 ;
        RECT 388.030 118.005 388.310 119.005 ;
        RECT 388.910 115.515 389.190 119.635 ;
        RECT 389.790 118.005 390.070 119.005 ;
        RECT 390.670 115.515 390.950 119.635 ;
        RECT 391.550 118.005 391.830 119.005 ;
        RECT 392.430 115.515 392.710 119.635 ;
        RECT 393.310 118.005 393.590 119.005 ;
        RECT 394.190 115.515 394.470 119.635 ;
        RECT 395.070 118.005 395.350 119.005 ;
        RECT 395.950 115.515 396.230 119.635 ;
        RECT 396.830 118.005 397.110 119.005 ;
        RECT 397.710 115.515 397.990 119.635 ;
        RECT 398.590 118.005 398.870 119.005 ;
        RECT 399.470 115.515 399.750 119.635 ;
        RECT 400.350 118.005 400.630 119.005 ;
        RECT 401.230 115.515 401.510 119.635 ;
        RECT 402.110 118.005 402.390 119.005 ;
        RECT 402.990 118.005 403.270 119.005 ;
        RECT 403.870 118.005 404.150 119.005 ;
        RECT 404.750 118.005 405.030 119.005 ;
        RECT 405.630 118.005 405.910 119.005 ;
        RECT 406.355 118.005 406.645 119.005 ;
        RECT 356.550 108.105 357.400 108.435 ;
        RECT 356.810 97.075 357.090 107.915 ;
        RECT 357.690 98.885 357.970 115.070 ;
        RECT 367.790 114.715 401.510 115.515 ;
        RECT 365.245 113.340 367.005 113.670 ;
        RECT 358.570 111.520 358.850 112.520 ;
        RECT 359.450 111.520 359.730 112.520 ;
        RECT 360.330 111.520 360.610 112.520 ;
        RECT 361.210 111.520 361.490 112.520 ;
        RECT 362.090 111.520 362.370 112.520 ;
        RECT 362.970 111.520 363.250 112.520 ;
        RECT 363.695 111.520 363.985 112.520 ;
        RECT 364.415 111.520 364.705 112.520 ;
        RECT 365.150 111.520 365.430 112.520 ;
        RECT 366.030 111.520 366.310 112.520 ;
        RECT 366.910 109.760 367.190 113.150 ;
        RECT 367.790 110.890 368.070 114.715 ;
        RECT 368.670 109.760 368.950 113.150 ;
        RECT 369.550 110.890 369.830 114.715 ;
        RECT 370.430 109.760 370.710 113.150 ;
        RECT 371.310 110.890 371.590 114.715 ;
        RECT 372.190 109.760 372.470 113.150 ;
        RECT 373.070 110.890 373.350 114.715 ;
        RECT 373.950 109.760 374.230 113.150 ;
        RECT 374.830 110.890 375.110 114.715 ;
        RECT 375.710 109.760 375.990 113.150 ;
        RECT 376.590 110.890 376.870 114.715 ;
        RECT 377.470 109.760 377.750 113.150 ;
        RECT 378.350 110.890 378.630 114.715 ;
        RECT 379.230 109.760 379.510 113.150 ;
        RECT 380.110 110.890 380.390 114.715 ;
        RECT 380.990 109.760 381.270 113.150 ;
        RECT 381.870 110.890 382.150 114.715 ;
        RECT 382.750 109.760 383.030 113.150 ;
        RECT 383.630 110.890 383.910 114.715 ;
        RECT 384.510 109.760 384.790 113.150 ;
        RECT 385.390 110.890 385.670 114.715 ;
        RECT 386.270 109.760 386.550 113.150 ;
        RECT 387.150 110.890 387.430 114.715 ;
        RECT 388.030 109.760 388.310 113.150 ;
        RECT 388.910 110.890 389.190 114.715 ;
        RECT 389.790 109.760 390.070 113.150 ;
        RECT 390.670 110.890 390.950 114.715 ;
        RECT 391.550 109.760 391.830 113.150 ;
        RECT 392.430 110.890 392.710 114.715 ;
        RECT 393.310 109.760 393.590 113.150 ;
        RECT 394.190 110.890 394.470 114.715 ;
        RECT 395.070 109.760 395.350 113.150 ;
        RECT 395.950 110.890 396.230 114.715 ;
        RECT 396.830 109.760 397.110 113.150 ;
        RECT 397.710 110.890 397.990 114.715 ;
        RECT 398.590 109.760 398.870 113.150 ;
        RECT 399.470 110.890 399.750 114.715 ;
        RECT 400.350 109.760 400.630 113.150 ;
        RECT 401.230 110.890 401.510 114.715 ;
        RECT 406.855 113.670 407.185 122.345 ;
        RECT 406.015 113.340 407.185 113.670 ;
        RECT 406.855 113.295 407.185 113.340 ;
        RECT 402.110 109.760 402.390 113.150 ;
        RECT 402.990 111.520 403.270 112.520 ;
        RECT 403.870 111.520 404.150 112.520 ;
        RECT 404.750 111.520 405.030 112.520 ;
        RECT 405.630 111.520 405.910 112.520 ;
        RECT 406.355 111.520 406.645 112.520 ;
        RECT 366.910 108.960 408.605 109.760 ;
        RECT 358.570 102.400 358.850 104.400 ;
        RECT 359.450 102.400 359.730 104.400 ;
        RECT 360.330 102.400 360.610 104.400 ;
        RECT 361.210 102.400 361.490 104.400 ;
        RECT 362.090 102.400 362.370 104.400 ;
        RECT 362.970 102.400 363.250 104.400 ;
        RECT 363.655 102.400 363.945 104.400 ;
        RECT 364.455 102.400 364.745 104.400 ;
        RECT 365.150 102.400 365.430 104.400 ;
        RECT 366.030 102.400 366.310 104.400 ;
        RECT 366.910 98.885 367.190 108.960 ;
        RECT 367.475 108.105 368.325 108.435 ;
        RECT 358.570 97.075 358.850 97.685 ;
        RECT 367.790 97.620 368.070 107.915 ;
        RECT 368.670 98.885 368.950 108.960 ;
        RECT 369.090 108.105 370.290 108.435 ;
        RECT 369.550 97.620 369.830 107.915 ;
        RECT 370.430 98.885 370.710 108.960 ;
        RECT 370.850 108.105 372.050 108.435 ;
        RECT 371.310 97.620 371.590 107.915 ;
        RECT 372.190 98.885 372.470 108.960 ;
        RECT 372.610 108.105 373.810 108.435 ;
        RECT 373.070 97.620 373.350 107.915 ;
        RECT 373.950 98.885 374.230 108.960 ;
        RECT 374.370 108.105 375.570 108.435 ;
        RECT 374.830 97.620 375.110 107.915 ;
        RECT 375.710 98.885 375.990 108.960 ;
        RECT 376.130 108.105 377.330 108.435 ;
        RECT 376.590 97.620 376.870 107.915 ;
        RECT 377.470 98.885 377.750 108.960 ;
        RECT 377.890 108.105 379.090 108.435 ;
        RECT 378.350 97.620 378.630 107.915 ;
        RECT 379.230 98.885 379.510 108.960 ;
        RECT 379.650 108.105 380.850 108.435 ;
        RECT 380.110 97.620 380.390 107.915 ;
        RECT 380.990 98.885 381.270 108.960 ;
        RECT 381.410 108.105 382.610 108.435 ;
        RECT 381.870 97.620 382.150 107.915 ;
        RECT 382.750 98.885 383.030 108.960 ;
        RECT 383.170 108.105 384.370 108.435 ;
        RECT 383.630 97.620 383.910 107.915 ;
        RECT 384.510 98.885 384.790 108.960 ;
        RECT 384.930 108.105 386.130 108.435 ;
        RECT 385.390 97.620 385.670 107.915 ;
        RECT 386.270 98.885 386.550 108.960 ;
        RECT 386.690 108.105 387.890 108.435 ;
        RECT 387.150 97.620 387.430 107.915 ;
        RECT 388.030 98.885 388.310 108.960 ;
        RECT 388.450 108.105 389.650 108.435 ;
        RECT 388.910 97.620 389.190 107.915 ;
        RECT 389.790 98.885 390.070 108.960 ;
        RECT 390.210 108.105 391.410 108.435 ;
        RECT 390.670 97.620 390.950 107.915 ;
        RECT 391.550 98.885 391.830 108.960 ;
        RECT 391.970 108.105 393.170 108.435 ;
        RECT 392.430 97.620 392.710 107.915 ;
        RECT 393.310 98.885 393.590 108.960 ;
        RECT 393.730 108.105 394.930 108.435 ;
        RECT 394.190 97.620 394.470 107.915 ;
        RECT 395.070 98.885 395.350 108.960 ;
        RECT 395.490 108.105 396.690 108.435 ;
        RECT 395.950 97.620 396.230 107.915 ;
        RECT 396.830 98.885 397.110 108.960 ;
        RECT 397.250 108.105 398.450 108.435 ;
        RECT 397.710 97.620 397.990 107.915 ;
        RECT 398.590 98.885 398.870 108.960 ;
        RECT 399.010 108.105 400.210 108.435 ;
        RECT 399.470 97.620 399.750 107.915 ;
        RECT 400.350 98.885 400.630 108.960 ;
        RECT 400.970 108.105 401.820 108.435 ;
        RECT 401.230 97.620 401.510 107.915 ;
        RECT 402.110 98.885 402.390 108.960 ;
        RECT 406.015 108.105 407.185 108.435 ;
        RECT 402.990 102.400 403.270 104.400 ;
        RECT 403.870 102.400 404.150 104.400 ;
        RECT 404.750 102.400 405.030 104.400 ;
        RECT 405.630 102.400 405.910 104.400 ;
        RECT 406.315 102.400 406.605 104.400 ;
        RECT 349.570 96.705 350.250 97.075 ;
        RECT 351.330 96.705 352.010 97.075 ;
        RECT 353.090 96.705 353.770 97.075 ;
        RECT 354.850 96.705 355.530 97.075 ;
        RECT 356.610 96.705 357.290 97.075 ;
        RECT 358.370 96.705 359.050 97.075 ;
        RECT 367.790 96.820 401.510 97.620 ;
        RECT 348.890 90.040 349.170 92.040 ;
        RECT 349.770 86.520 350.050 96.705 ;
        RECT 350.650 90.040 350.930 92.040 ;
        RECT 351.530 86.520 351.810 96.705 ;
        RECT 352.410 90.040 352.690 92.040 ;
        RECT 353.290 86.520 353.570 96.705 ;
        RECT 354.170 90.040 354.450 92.040 ;
        RECT 355.050 86.520 355.330 96.705 ;
        RECT 355.930 90.040 356.210 92.040 ;
        RECT 356.810 86.520 357.090 96.705 ;
        RECT 357.690 90.040 357.970 92.040 ;
        RECT 358.570 86.520 358.850 96.705 ;
        RECT 359.450 90.040 359.730 92.040 ;
        RECT 360.330 90.040 360.610 92.040 ;
        RECT 361.210 90.040 361.490 92.040 ;
        RECT 362.090 90.040 362.370 92.040 ;
        RECT 362.970 90.040 363.250 92.040 ;
        RECT 363.655 90.040 363.945 92.040 ;
        RECT 364.455 90.040 364.745 92.040 ;
        RECT 365.150 90.040 365.430 92.040 ;
        RECT 366.030 90.040 366.310 92.040 ;
        RECT 366.910 90.040 367.190 92.040 ;
        RECT 367.790 86.520 368.070 96.820 ;
        RECT 368.670 90.040 368.950 92.040 ;
        RECT 369.550 86.520 369.830 96.820 ;
        RECT 370.430 90.040 370.710 92.040 ;
        RECT 371.310 86.520 371.590 96.820 ;
        RECT 372.190 90.040 372.470 92.040 ;
        RECT 373.070 86.520 373.350 96.820 ;
        RECT 373.950 90.040 374.230 92.040 ;
        RECT 374.830 86.520 375.110 96.820 ;
        RECT 375.710 90.040 375.990 92.040 ;
        RECT 376.590 86.520 376.870 96.820 ;
        RECT 377.470 90.040 377.750 92.040 ;
        RECT 378.350 86.520 378.630 96.820 ;
        RECT 379.230 90.040 379.510 92.040 ;
        RECT 380.110 86.520 380.390 96.820 ;
        RECT 380.990 90.040 381.270 92.040 ;
        RECT 381.870 86.520 382.150 96.820 ;
        RECT 382.750 90.040 383.030 92.040 ;
        RECT 383.630 86.520 383.910 96.820 ;
        RECT 384.510 90.040 384.790 92.040 ;
        RECT 385.390 86.520 385.670 96.820 ;
        RECT 386.270 90.040 386.550 92.040 ;
        RECT 387.150 86.520 387.430 96.820 ;
        RECT 388.030 90.040 388.310 92.040 ;
        RECT 388.910 86.520 389.190 96.820 ;
        RECT 389.790 90.040 390.070 92.040 ;
        RECT 390.670 86.520 390.950 96.820 ;
        RECT 391.550 90.040 391.830 92.040 ;
        RECT 392.430 86.520 392.710 96.820 ;
        RECT 393.310 90.040 393.590 92.040 ;
        RECT 394.190 86.520 394.470 96.820 ;
        RECT 395.070 90.040 395.350 92.040 ;
        RECT 395.950 86.520 396.230 96.820 ;
        RECT 396.830 90.040 397.110 92.040 ;
        RECT 397.710 86.520 397.990 96.820 ;
        RECT 398.590 90.040 398.870 92.040 ;
        RECT 399.470 86.520 399.750 96.820 ;
        RECT 400.350 90.040 400.630 92.040 ;
        RECT 401.230 86.520 401.510 96.820 ;
        RECT 402.110 90.040 402.390 92.040 ;
        RECT 402.990 90.040 403.270 92.040 ;
        RECT 403.870 90.040 404.150 92.040 ;
        RECT 404.750 90.040 405.030 92.040 ;
        RECT 405.630 90.040 405.910 92.040 ;
        RECT 406.315 90.040 406.605 92.040 ;
        RECT 338.645 86.040 359.415 86.370 ;
        RECT 367.265 86.040 402.035 86.370 ;
        RECT 406.855 84.615 407.185 108.105 ;
        RECT 406.435 84.285 407.605 84.615 ;
        RECT 305.240 79.490 306.550 80.490 ;
        RECT 307.250 79.490 310.570 80.490 ;
        RECT 311.270 79.490 314.590 80.490 ;
        RECT 315.290 79.490 318.610 80.490 ;
        RECT 319.310 79.490 322.630 80.490 ;
        RECT 323.330 79.490 326.650 80.490 ;
        RECT 327.350 79.490 330.670 80.490 ;
        RECT 331.370 79.490 334.690 80.490 ;
        RECT 335.390 79.490 338.710 80.490 ;
        RECT 339.410 79.490 342.730 80.490 ;
        RECT 343.430 79.490 346.750 80.490 ;
        RECT 347.450 79.490 350.770 80.490 ;
        RECT 351.470 79.490 354.790 80.490 ;
        RECT 355.490 79.490 358.810 80.490 ;
        RECT 359.510 79.490 362.830 80.490 ;
        RECT 363.530 79.490 366.850 80.490 ;
        RECT 367.550 79.490 370.870 80.490 ;
        RECT 371.570 79.490 374.890 80.490 ;
        RECT 375.590 79.490 378.910 80.490 ;
        RECT 379.610 79.490 382.930 80.490 ;
        RECT 383.630 79.490 386.950 80.490 ;
        RECT 387.650 79.490 390.970 80.490 ;
        RECT 391.670 79.490 394.990 80.490 ;
        RECT 395.690 79.490 399.010 80.490 ;
        RECT 399.710 79.490 403.030 80.490 ;
        RECT 403.730 79.490 405.040 80.490 ;
        RECT 408.005 80.290 408.605 108.960 ;
        RECT 408.005 79.690 429.280 80.290 ;
        RECT 300.325 74.180 300.605 76.180 ;
        RECT 409.675 74.180 409.955 76.180 ;
        RECT 305.240 69.895 308.560 70.895 ;
        RECT 309.260 69.895 312.580 70.895 ;
        RECT 313.280 69.895 316.600 70.895 ;
        RECT 317.300 69.895 320.620 70.895 ;
        RECT 321.320 69.895 324.640 70.895 ;
        RECT 325.340 69.895 328.660 70.895 ;
        RECT 329.360 69.895 332.680 70.895 ;
        RECT 333.380 69.895 336.700 70.895 ;
        RECT 337.400 69.895 340.720 70.895 ;
        RECT 341.420 69.895 344.740 70.895 ;
        RECT 345.440 69.895 348.760 70.895 ;
        RECT 349.460 69.895 352.780 70.895 ;
        RECT 353.480 69.895 356.800 70.895 ;
        RECT 357.500 69.895 360.820 70.895 ;
        RECT 361.520 69.895 364.840 70.895 ;
        RECT 365.540 69.895 368.860 70.895 ;
        RECT 369.560 69.895 372.880 70.895 ;
        RECT 373.580 69.895 376.900 70.895 ;
        RECT 377.600 69.895 380.920 70.895 ;
        RECT 381.620 69.895 384.940 70.895 ;
        RECT 385.640 69.895 388.960 70.895 ;
        RECT 389.660 69.895 392.980 70.895 ;
        RECT 393.680 69.895 397.000 70.895 ;
        RECT 397.700 69.895 401.020 70.895 ;
        RECT 401.720 69.895 405.040 70.895 ;
        RECT 299.055 67.830 300.160 68.430 ;
        RECT 410.025 67.830 411.105 68.430 ;
        RECT 189.705 65.345 191.015 66.345 ;
        RECT 191.715 65.345 195.035 66.345 ;
        RECT 195.735 65.345 199.055 66.345 ;
        RECT 199.755 65.345 203.075 66.345 ;
        RECT 203.775 65.345 207.095 66.345 ;
        RECT 207.795 65.345 211.115 66.345 ;
        RECT 211.815 65.345 215.135 66.345 ;
        RECT 215.835 65.345 219.155 66.345 ;
        RECT 219.855 65.345 223.175 66.345 ;
        RECT 223.875 65.345 227.195 66.345 ;
        RECT 227.895 65.345 231.215 66.345 ;
        RECT 231.915 65.345 235.235 66.345 ;
        RECT 235.935 65.345 239.255 66.345 ;
        RECT 239.955 65.345 243.275 66.345 ;
        RECT 243.975 65.345 247.295 66.345 ;
        RECT 247.995 65.345 251.315 66.345 ;
        RECT 252.015 65.345 255.335 66.345 ;
        RECT 256.035 65.345 259.355 66.345 ;
        RECT 260.055 65.345 263.375 66.345 ;
        RECT 264.075 65.345 267.395 66.345 ;
        RECT 268.095 65.345 271.415 66.345 ;
        RECT 272.115 65.345 275.435 66.345 ;
        RECT 276.135 65.345 279.455 66.345 ;
        RECT 280.155 65.345 283.475 66.345 ;
        RECT 284.175 65.345 287.495 66.345 ;
        RECT 288.195 65.345 289.505 66.345 ;
        RECT 184.790 60.035 185.070 62.035 ;
        RECT 294.140 60.035 294.420 62.035 ;
        RECT 189.705 55.750 193.025 56.750 ;
        RECT 193.725 55.750 197.045 56.750 ;
        RECT 197.745 55.750 201.065 56.750 ;
        RECT 201.765 55.750 205.085 56.750 ;
        RECT 205.785 55.750 209.105 56.750 ;
        RECT 209.805 55.750 213.125 56.750 ;
        RECT 213.825 55.750 217.145 56.750 ;
        RECT 217.845 55.750 221.165 56.750 ;
        RECT 221.865 55.750 225.185 56.750 ;
        RECT 225.885 55.750 229.205 56.750 ;
        RECT 229.905 55.750 233.225 56.750 ;
        RECT 233.925 55.750 237.245 56.750 ;
        RECT 237.945 55.750 241.265 56.750 ;
        RECT 241.965 55.750 245.285 56.750 ;
        RECT 245.985 55.750 249.305 56.750 ;
        RECT 250.005 55.750 253.325 56.750 ;
        RECT 254.025 55.750 257.345 56.750 ;
        RECT 258.045 55.750 261.365 56.750 ;
        RECT 262.065 55.750 265.385 56.750 ;
        RECT 266.085 55.750 269.405 56.750 ;
        RECT 270.105 55.750 273.425 56.750 ;
        RECT 274.125 55.750 277.445 56.750 ;
        RECT 278.145 55.750 281.465 56.750 ;
        RECT 282.165 55.750 285.485 56.750 ;
        RECT 286.185 55.750 289.505 56.750 ;
        RECT 281.935 53.945 283.040 54.545 ;
        RECT 297.075 53.945 297.675 66.345 ;
        RECT 305.240 65.345 306.550 66.345 ;
        RECT 307.250 65.345 310.570 66.345 ;
        RECT 311.270 65.345 314.590 66.345 ;
        RECT 315.290 65.345 318.610 66.345 ;
        RECT 319.310 65.345 322.630 66.345 ;
        RECT 323.330 65.345 326.650 66.345 ;
        RECT 327.350 65.345 330.670 66.345 ;
        RECT 331.370 65.345 334.690 66.345 ;
        RECT 335.390 65.345 338.710 66.345 ;
        RECT 339.410 65.345 342.730 66.345 ;
        RECT 343.430 65.345 346.750 66.345 ;
        RECT 347.450 65.345 350.770 66.345 ;
        RECT 351.470 65.345 354.790 66.345 ;
        RECT 355.490 65.345 358.810 66.345 ;
        RECT 359.510 65.345 362.830 66.345 ;
        RECT 363.530 65.345 366.850 66.345 ;
        RECT 367.550 65.345 370.870 66.345 ;
        RECT 371.570 65.345 374.890 66.345 ;
        RECT 375.590 65.345 378.910 66.345 ;
        RECT 379.610 65.345 382.930 66.345 ;
        RECT 383.630 65.345 386.950 66.345 ;
        RECT 387.650 65.345 390.970 66.345 ;
        RECT 391.670 65.345 394.990 66.345 ;
        RECT 395.690 65.345 399.010 66.345 ;
        RECT 399.710 65.345 403.030 66.345 ;
        RECT 403.730 65.345 405.040 66.345 ;
        RECT 410.505 65.345 411.105 67.830 ;
        RECT 300.325 60.035 300.605 62.035 ;
        RECT 409.675 60.035 409.955 62.035 ;
        RECT 305.240 55.750 308.560 56.750 ;
        RECT 309.260 55.750 312.580 56.750 ;
        RECT 313.280 55.750 316.600 56.750 ;
        RECT 317.300 55.750 320.620 56.750 ;
        RECT 321.320 55.750 324.640 56.750 ;
        RECT 325.340 55.750 328.660 56.750 ;
        RECT 329.360 55.750 332.680 56.750 ;
        RECT 333.380 55.750 336.700 56.750 ;
        RECT 337.400 55.750 340.720 56.750 ;
        RECT 341.420 55.750 344.740 56.750 ;
        RECT 345.440 55.750 348.760 56.750 ;
        RECT 349.460 55.750 352.780 56.750 ;
        RECT 353.480 55.750 356.800 56.750 ;
        RECT 357.500 55.750 360.820 56.750 ;
        RECT 361.520 55.750 364.840 56.750 ;
        RECT 365.540 55.750 368.860 56.750 ;
        RECT 369.560 55.750 372.880 56.750 ;
        RECT 373.580 55.750 376.900 56.750 ;
        RECT 377.600 55.750 380.920 56.750 ;
        RECT 381.620 55.750 384.940 56.750 ;
        RECT 385.640 55.750 388.960 56.750 ;
        RECT 389.660 55.750 392.980 56.750 ;
        RECT 393.680 55.750 397.000 56.750 ;
        RECT 397.700 55.750 401.020 56.750 ;
        RECT 401.720 55.750 405.040 56.750 ;
        RECT 280.365 53.315 281.535 53.645 ;
        RECT 212.575 51.560 233.345 51.890 ;
        RECT 241.195 51.560 275.965 51.890 ;
        RECT 208.045 45.890 208.335 47.890 ;
        RECT 208.740 45.890 209.020 47.890 ;
        RECT 209.620 45.890 209.900 47.890 ;
        RECT 210.500 45.890 210.780 47.890 ;
        RECT 211.380 45.890 211.660 47.890 ;
        RECT 212.260 45.890 212.540 47.890 ;
        RECT 189.920 40.595 190.200 41.205 ;
        RECT 191.500 40.855 192.180 41.225 ;
        RECT 189.720 40.225 190.400 40.595 ;
        RECT 185.885 36.430 187.550 36.720 ;
        RECT 184.785 34.020 185.075 35.020 ;
        RECT 185.520 34.020 185.800 35.020 ;
        RECT 186.400 34.020 186.680 35.020 ;
        RECT 187.280 34.020 187.560 35.020 ;
        RECT 188.160 34.020 188.440 35.020 ;
        RECT 185.885 32.320 187.550 32.610 ;
        RECT 189.040 31.045 189.320 35.650 ;
        RECT 189.920 33.390 190.200 40.225 ;
        RECT 190.800 31.045 191.080 35.650 ;
        RECT 191.680 33.390 191.960 40.855 ;
        RECT 193.440 40.595 193.720 41.205 ;
        RECT 195.020 40.855 195.700 41.225 ;
        RECT 193.240 40.225 193.920 40.595 ;
        RECT 192.560 31.045 192.840 35.650 ;
        RECT 193.440 33.390 193.720 40.225 ;
        RECT 194.320 31.045 194.600 35.650 ;
        RECT 195.200 33.390 195.480 40.855 ;
        RECT 196.960 40.595 197.240 41.205 ;
        RECT 198.540 40.855 199.220 41.225 ;
        RECT 196.760 40.225 197.440 40.595 ;
        RECT 196.080 31.045 196.360 35.650 ;
        RECT 196.960 33.390 197.240 40.225 ;
        RECT 197.840 31.045 198.120 35.650 ;
        RECT 198.720 33.390 199.000 40.855 ;
        RECT 200.480 40.595 200.760 41.205 ;
        RECT 202.060 40.855 202.740 41.225 ;
        RECT 200.280 40.225 200.960 40.595 ;
        RECT 199.600 31.045 199.880 35.650 ;
        RECT 200.480 33.390 200.760 40.225 ;
        RECT 201.360 31.045 201.640 35.650 ;
        RECT 202.240 33.390 202.520 40.855 ;
        RECT 213.140 40.595 213.420 51.410 ;
        RECT 214.020 45.890 214.300 47.890 ;
        RECT 214.900 40.595 215.180 51.410 ;
        RECT 215.780 45.890 216.060 47.890 ;
        RECT 216.660 40.595 216.940 51.410 ;
        RECT 217.540 45.890 217.820 47.890 ;
        RECT 218.420 40.595 218.700 51.410 ;
        RECT 219.300 45.890 219.580 47.890 ;
        RECT 220.180 40.595 220.460 51.410 ;
        RECT 221.060 45.890 221.340 47.890 ;
        RECT 221.940 40.595 222.220 51.410 ;
        RECT 222.820 45.890 223.100 47.890 ;
        RECT 223.700 41.225 223.980 51.410 ;
        RECT 224.580 45.890 224.860 47.890 ;
        RECT 225.460 41.225 225.740 51.410 ;
        RECT 226.340 45.890 226.620 47.890 ;
        RECT 227.220 41.225 227.500 51.410 ;
        RECT 228.100 45.890 228.380 47.890 ;
        RECT 228.980 41.225 229.260 51.410 ;
        RECT 229.860 45.890 230.140 47.890 ;
        RECT 230.740 41.225 231.020 51.410 ;
        RECT 231.620 45.890 231.900 47.890 ;
        RECT 232.500 41.225 232.780 51.410 ;
        RECT 233.380 45.890 233.660 47.890 ;
        RECT 234.260 45.890 234.540 47.890 ;
        RECT 235.140 45.890 235.420 47.890 ;
        RECT 236.020 45.890 236.300 47.890 ;
        RECT 236.900 45.890 237.180 47.890 ;
        RECT 237.585 45.890 237.875 47.890 ;
        RECT 238.385 45.890 238.675 47.890 ;
        RECT 239.080 45.890 239.360 47.890 ;
        RECT 239.960 45.890 240.240 47.890 ;
        RECT 240.840 45.890 241.120 47.890 ;
        RECT 223.500 40.855 224.180 41.225 ;
        RECT 225.260 40.855 225.940 41.225 ;
        RECT 227.020 40.855 227.700 41.225 ;
        RECT 228.780 40.855 229.460 41.225 ;
        RECT 230.540 40.855 231.220 41.225 ;
        RECT 232.300 40.855 232.980 41.225 ;
        RECT 241.720 41.110 242.000 51.410 ;
        RECT 242.600 45.890 242.880 47.890 ;
        RECT 243.480 41.110 243.760 51.410 ;
        RECT 244.360 45.890 244.640 47.890 ;
        RECT 245.240 41.110 245.520 51.410 ;
        RECT 246.120 45.890 246.400 47.890 ;
        RECT 247.000 41.110 247.280 51.410 ;
        RECT 247.880 45.890 248.160 47.890 ;
        RECT 248.760 41.110 249.040 51.410 ;
        RECT 249.640 45.890 249.920 47.890 ;
        RECT 250.520 41.110 250.800 51.410 ;
        RECT 251.400 45.890 251.680 47.890 ;
        RECT 252.280 41.110 252.560 51.410 ;
        RECT 253.160 45.890 253.440 47.890 ;
        RECT 254.040 41.110 254.320 51.410 ;
        RECT 254.920 45.890 255.200 47.890 ;
        RECT 255.800 41.110 256.080 51.410 ;
        RECT 256.680 45.890 256.960 47.890 ;
        RECT 257.560 41.110 257.840 51.410 ;
        RECT 258.440 45.890 258.720 47.890 ;
        RECT 259.320 41.110 259.600 51.410 ;
        RECT 260.200 45.890 260.480 47.890 ;
        RECT 261.080 41.110 261.360 51.410 ;
        RECT 261.960 45.890 262.240 47.890 ;
        RECT 262.840 41.110 263.120 51.410 ;
        RECT 263.720 45.890 264.000 47.890 ;
        RECT 264.600 41.110 264.880 51.410 ;
        RECT 265.480 45.890 265.760 47.890 ;
        RECT 266.360 41.110 266.640 51.410 ;
        RECT 267.240 45.890 267.520 47.890 ;
        RECT 268.120 41.110 268.400 51.410 ;
        RECT 269.000 45.890 269.280 47.890 ;
        RECT 269.880 41.110 270.160 51.410 ;
        RECT 270.760 45.890 271.040 47.890 ;
        RECT 271.640 41.110 271.920 51.410 ;
        RECT 272.520 45.890 272.800 47.890 ;
        RECT 273.400 41.110 273.680 51.410 ;
        RECT 274.280 45.890 274.560 47.890 ;
        RECT 275.160 41.110 275.440 51.410 ;
        RECT 276.040 45.890 276.320 47.890 ;
        RECT 276.920 45.890 277.200 47.890 ;
        RECT 277.800 45.890 278.080 47.890 ;
        RECT 278.680 45.890 278.960 47.890 ;
        RECT 279.560 45.890 279.840 47.890 ;
        RECT 280.245 45.890 280.535 47.890 ;
        RECT 212.940 40.225 213.620 40.595 ;
        RECT 214.700 40.225 215.380 40.595 ;
        RECT 216.460 40.225 217.140 40.595 ;
        RECT 218.220 40.225 218.900 40.595 ;
        RECT 219.980 40.225 220.660 40.595 ;
        RECT 221.740 40.225 222.420 40.595 ;
        RECT 223.700 40.245 223.980 40.855 ;
        RECT 203.120 31.045 203.400 35.650 ;
        RECT 204.000 34.020 204.280 35.020 ;
        RECT 204.880 34.020 205.160 35.020 ;
        RECT 205.760 34.020 206.040 35.020 ;
        RECT 206.640 34.020 206.920 35.020 ;
        RECT 207.365 34.020 207.655 35.020 ;
        RECT 208.045 33.530 208.335 35.530 ;
        RECT 208.740 33.530 209.020 35.530 ;
        RECT 209.620 33.530 209.900 35.530 ;
        RECT 210.500 33.530 210.780 35.530 ;
        RECT 211.380 33.530 211.660 35.530 ;
        RECT 212.260 33.530 212.540 35.530 ;
        RECT 213.140 33.530 213.420 35.530 ;
        RECT 189.040 30.545 203.400 31.045 ;
        RECT 184.785 25.410 185.075 26.410 ;
        RECT 185.520 25.410 185.800 26.410 ;
        RECT 186.400 25.410 186.680 26.410 ;
        RECT 187.280 25.410 187.560 26.410 ;
        RECT 188.160 25.410 188.440 26.410 ;
        RECT 189.040 25.410 189.320 26.410 ;
        RECT 189.920 25.410 190.200 26.410 ;
        RECT 190.800 25.410 191.080 26.410 ;
        RECT 191.680 25.410 191.960 26.410 ;
        RECT 192.560 24.780 192.840 30.545 ;
        RECT 192.905 24.260 193.300 24.590 ;
        RECT 193.440 22.915 193.720 27.040 ;
        RECT 194.320 24.780 194.600 30.545 ;
        RECT 193.860 24.260 195.060 24.590 ;
        RECT 195.200 22.915 195.480 27.040 ;
        RECT 196.080 24.780 196.360 30.545 ;
        RECT 195.620 24.260 196.820 24.590 ;
        RECT 196.960 22.915 197.240 27.040 ;
        RECT 197.840 24.780 198.120 30.545 ;
        RECT 197.380 24.260 198.580 24.590 ;
        RECT 198.720 22.915 199.000 27.040 ;
        RECT 199.600 24.780 199.880 30.545 ;
        RECT 200.480 25.410 200.760 26.410 ;
        RECT 201.360 25.410 201.640 26.410 ;
        RECT 202.240 25.410 202.520 26.410 ;
        RECT 203.120 25.410 203.400 26.410 ;
        RECT 204.000 25.410 204.280 26.410 ;
        RECT 204.880 25.410 205.160 26.410 ;
        RECT 205.760 25.410 206.040 26.410 ;
        RECT 206.640 25.410 206.920 26.410 ;
        RECT 207.365 25.410 207.655 26.410 ;
        RECT 208.005 25.410 208.295 26.410 ;
        RECT 208.740 25.410 209.020 26.410 ;
        RECT 209.620 25.410 209.900 26.410 ;
        RECT 210.500 25.410 210.780 26.410 ;
        RECT 211.380 25.410 211.660 26.410 ;
        RECT 212.260 25.410 212.540 26.410 ;
        RECT 213.140 25.410 213.420 26.410 ;
        RECT 199.140 24.260 199.515 24.590 ;
        RECT 211.660 24.260 213.420 24.590 ;
        RECT 193.440 22.415 199.000 22.915 ;
        RECT 214.020 22.860 214.300 39.045 ;
        RECT 214.900 30.015 215.180 40.225 ;
        RECT 214.585 29.495 215.435 29.825 ;
        RECT 184.785 18.925 185.075 19.925 ;
        RECT 185.520 18.925 185.800 19.925 ;
        RECT 186.400 18.925 186.680 19.925 ;
        RECT 187.280 18.925 187.560 19.925 ;
        RECT 188.160 18.925 188.440 19.925 ;
        RECT 189.040 18.925 189.320 19.925 ;
        RECT 189.920 18.925 190.200 19.925 ;
        RECT 190.800 18.925 191.080 19.925 ;
        RECT 191.680 18.925 191.960 19.925 ;
        RECT 192.560 18.925 192.840 19.925 ;
        RECT 193.440 18.295 193.720 22.415 ;
        RECT 194.320 18.925 194.600 19.925 ;
        RECT 195.200 18.295 195.480 22.415 ;
        RECT 196.080 18.925 196.360 19.925 ;
        RECT 196.960 18.295 197.240 22.415 ;
        RECT 197.840 18.925 198.120 19.925 ;
        RECT 198.720 18.295 199.000 22.415 ;
        RECT 199.600 18.925 199.880 19.925 ;
        RECT 200.480 18.925 200.760 19.925 ;
        RECT 201.360 18.925 201.640 19.925 ;
        RECT 202.240 18.925 202.520 19.925 ;
        RECT 203.120 18.925 203.400 19.925 ;
        RECT 204.000 18.925 204.280 19.925 ;
        RECT 204.880 18.925 205.160 19.925 ;
        RECT 205.760 18.925 206.040 19.925 ;
        RECT 206.640 18.925 206.920 19.925 ;
        RECT 207.365 18.925 207.655 19.925 ;
        RECT 208.005 18.925 208.295 19.925 ;
        RECT 208.740 18.925 209.020 19.925 ;
        RECT 209.620 18.925 209.900 19.925 ;
        RECT 210.500 18.925 210.780 19.925 ;
        RECT 211.380 18.925 211.660 19.925 ;
        RECT 212.260 18.925 212.540 19.925 ;
        RECT 213.140 18.925 213.420 19.925 ;
        RECT 214.020 18.925 214.300 19.925 ;
        RECT 214.900 18.295 215.180 27.040 ;
        RECT 215.780 22.860 216.060 39.045 ;
        RECT 216.660 30.015 216.940 40.225 ;
        RECT 216.200 29.495 217.400 29.825 ;
        RECT 215.780 18.925 216.060 19.925 ;
        RECT 216.660 18.295 216.940 27.040 ;
        RECT 217.540 23.380 217.820 39.045 ;
        RECT 218.420 30.015 218.700 40.225 ;
        RECT 217.960 29.495 219.160 29.825 ;
        RECT 217.430 21.050 217.930 23.380 ;
        RECT 217.390 20.730 217.970 21.050 ;
        RECT 217.540 18.925 217.820 19.925 ;
        RECT 218.420 18.295 218.700 27.040 ;
        RECT 219.300 22.860 219.580 39.045 ;
        RECT 220.180 30.015 220.460 40.225 ;
        RECT 219.720 29.495 220.920 29.825 ;
        RECT 219.300 18.925 219.580 19.925 ;
        RECT 220.180 18.295 220.460 27.040 ;
        RECT 221.060 22.860 221.340 39.045 ;
        RECT 221.940 33.530 222.220 35.530 ;
        RECT 222.820 33.530 223.100 35.530 ;
        RECT 223.700 33.530 223.980 35.530 ;
        RECT 221.940 25.410 222.220 26.410 ;
        RECT 222.820 25.410 223.100 26.410 ;
        RECT 223.700 25.410 223.980 26.410 ;
        RECT 224.580 22.860 224.860 39.045 ;
        RECT 225.460 30.015 225.740 40.855 ;
        RECT 225.000 29.495 226.200 29.825 ;
        RECT 221.060 18.925 221.340 19.925 ;
        RECT 221.940 18.925 222.220 19.925 ;
        RECT 222.820 18.925 223.100 19.925 ;
        RECT 223.700 18.925 223.980 19.925 ;
        RECT 224.580 18.925 224.860 19.925 ;
        RECT 192.925 17.775 194.320 18.105 ;
        RECT 225.460 16.245 225.740 27.040 ;
        RECT 226.340 22.860 226.620 39.045 ;
        RECT 227.220 30.015 227.500 40.855 ;
        RECT 226.760 29.495 227.960 29.825 ;
        RECT 226.340 18.925 226.620 19.925 ;
        RECT 227.220 16.245 227.500 27.040 ;
        RECT 228.100 22.860 228.380 39.045 ;
        RECT 228.980 30.015 229.260 40.855 ;
        RECT 228.520 29.495 229.720 29.825 ;
        RECT 228.100 18.925 228.380 19.925 ;
        RECT 228.980 16.245 229.260 27.040 ;
        RECT 229.860 22.860 230.140 39.045 ;
        RECT 230.740 30.015 231.020 40.855 ;
        RECT 232.500 40.245 232.780 40.855 ;
        RECT 241.720 40.310 275.440 41.110 ;
        RECT 230.480 29.495 231.330 29.825 ;
        RECT 229.860 18.925 230.140 19.925 ;
        RECT 230.740 16.245 231.020 27.040 ;
        RECT 231.620 22.860 231.900 39.045 ;
        RECT 232.500 33.530 232.780 35.530 ;
        RECT 233.380 33.530 233.660 35.530 ;
        RECT 234.260 33.530 234.540 35.530 ;
        RECT 235.140 33.530 235.420 35.530 ;
        RECT 236.020 33.530 236.300 35.530 ;
        RECT 236.900 33.530 237.180 35.530 ;
        RECT 237.585 33.530 237.875 35.530 ;
        RECT 238.385 33.530 238.675 35.530 ;
        RECT 239.080 33.530 239.360 35.530 ;
        RECT 239.960 33.530 240.240 35.530 ;
        RECT 240.840 28.970 241.120 39.045 ;
        RECT 241.720 30.015 242.000 40.310 ;
        RECT 241.405 29.495 242.255 29.825 ;
        RECT 242.600 28.970 242.880 39.045 ;
        RECT 243.480 30.015 243.760 40.310 ;
        RECT 243.020 29.495 244.220 29.825 ;
        RECT 244.360 28.970 244.640 39.045 ;
        RECT 245.240 30.015 245.520 40.310 ;
        RECT 244.780 29.495 245.980 29.825 ;
        RECT 246.120 28.970 246.400 39.045 ;
        RECT 247.000 30.015 247.280 40.310 ;
        RECT 246.540 29.495 247.740 29.825 ;
        RECT 247.880 28.970 248.160 39.045 ;
        RECT 248.760 30.015 249.040 40.310 ;
        RECT 248.300 29.495 249.500 29.825 ;
        RECT 249.640 28.970 249.920 39.045 ;
        RECT 250.520 30.015 250.800 40.310 ;
        RECT 250.060 29.495 251.260 29.825 ;
        RECT 251.400 28.970 251.680 39.045 ;
        RECT 252.280 30.015 252.560 40.310 ;
        RECT 251.820 29.495 253.020 29.825 ;
        RECT 253.160 28.970 253.440 39.045 ;
        RECT 254.040 30.015 254.320 40.310 ;
        RECT 253.580 29.495 254.780 29.825 ;
        RECT 254.920 28.970 255.200 39.045 ;
        RECT 255.800 30.015 256.080 40.310 ;
        RECT 255.340 29.495 256.540 29.825 ;
        RECT 256.680 28.970 256.960 39.045 ;
        RECT 257.560 30.015 257.840 40.310 ;
        RECT 257.100 29.495 258.300 29.825 ;
        RECT 258.440 28.970 258.720 39.045 ;
        RECT 259.320 30.015 259.600 40.310 ;
        RECT 258.860 29.495 260.060 29.825 ;
        RECT 260.200 28.970 260.480 39.045 ;
        RECT 261.080 30.015 261.360 40.310 ;
        RECT 260.620 29.495 261.820 29.825 ;
        RECT 261.960 28.970 262.240 39.045 ;
        RECT 262.840 30.015 263.120 40.310 ;
        RECT 262.380 29.495 263.580 29.825 ;
        RECT 263.720 28.970 264.000 39.045 ;
        RECT 264.600 30.015 264.880 40.310 ;
        RECT 264.140 29.495 265.340 29.825 ;
        RECT 265.480 28.970 265.760 39.045 ;
        RECT 266.360 30.015 266.640 40.310 ;
        RECT 265.900 29.495 267.100 29.825 ;
        RECT 267.240 28.970 267.520 39.045 ;
        RECT 268.120 30.015 268.400 40.310 ;
        RECT 267.660 29.495 268.860 29.825 ;
        RECT 269.000 28.970 269.280 39.045 ;
        RECT 269.880 30.015 270.160 40.310 ;
        RECT 269.420 29.495 270.620 29.825 ;
        RECT 270.760 28.970 271.040 39.045 ;
        RECT 271.640 30.015 271.920 40.310 ;
        RECT 271.180 29.495 272.380 29.825 ;
        RECT 272.520 28.970 272.800 39.045 ;
        RECT 273.400 30.015 273.680 40.310 ;
        RECT 272.940 29.495 274.140 29.825 ;
        RECT 274.280 28.970 274.560 39.045 ;
        RECT 275.160 30.015 275.440 40.310 ;
        RECT 274.900 29.495 275.750 29.825 ;
        RECT 276.040 28.970 276.320 39.045 ;
        RECT 276.920 33.530 277.200 35.530 ;
        RECT 277.800 33.530 278.080 35.530 ;
        RECT 278.680 33.530 278.960 35.530 ;
        RECT 279.560 33.530 279.840 35.530 ;
        RECT 280.245 33.530 280.535 35.530 ;
        RECT 280.785 29.825 281.115 53.315 ;
        RECT 279.945 29.495 281.115 29.825 ;
        RECT 281.935 28.970 282.535 53.945 ;
        RECT 240.840 28.170 282.535 28.970 ;
        RECT 328.700 53.925 329.805 54.295 ;
        RECT 426.915 53.925 427.995 54.295 ;
        RECT 328.700 28.970 329.300 53.925 ;
        RECT 329.700 53.315 330.870 53.645 ;
        RECT 330.120 29.825 330.450 53.315 ;
        RECT 335.270 51.560 370.040 51.890 ;
        RECT 377.890 51.560 398.660 51.890 ;
        RECT 330.700 45.890 330.990 47.890 ;
        RECT 331.395 45.890 331.675 47.890 ;
        RECT 332.275 45.890 332.555 47.890 ;
        RECT 333.155 45.890 333.435 47.890 ;
        RECT 334.035 45.890 334.315 47.890 ;
        RECT 334.915 45.890 335.195 47.890 ;
        RECT 335.795 41.110 336.075 51.410 ;
        RECT 336.675 45.890 336.955 47.890 ;
        RECT 337.555 41.110 337.835 51.410 ;
        RECT 338.435 45.890 338.715 47.890 ;
        RECT 339.315 41.110 339.595 51.410 ;
        RECT 340.195 45.890 340.475 47.890 ;
        RECT 341.075 41.110 341.355 51.410 ;
        RECT 341.955 45.890 342.235 47.890 ;
        RECT 342.835 41.110 343.115 51.410 ;
        RECT 343.715 45.890 343.995 47.890 ;
        RECT 344.595 41.110 344.875 51.410 ;
        RECT 345.475 45.890 345.755 47.890 ;
        RECT 346.355 41.110 346.635 51.410 ;
        RECT 347.235 45.890 347.515 47.890 ;
        RECT 348.115 41.110 348.395 51.410 ;
        RECT 348.995 45.890 349.275 47.890 ;
        RECT 349.875 41.110 350.155 51.410 ;
        RECT 350.755 45.890 351.035 47.890 ;
        RECT 351.635 41.110 351.915 51.410 ;
        RECT 352.515 45.890 352.795 47.890 ;
        RECT 353.395 41.110 353.675 51.410 ;
        RECT 354.275 45.890 354.555 47.890 ;
        RECT 355.155 41.110 355.435 51.410 ;
        RECT 356.035 45.890 356.315 47.890 ;
        RECT 356.915 41.110 357.195 51.410 ;
        RECT 357.795 45.890 358.075 47.890 ;
        RECT 358.675 41.110 358.955 51.410 ;
        RECT 359.555 45.890 359.835 47.890 ;
        RECT 360.435 41.110 360.715 51.410 ;
        RECT 361.315 45.890 361.595 47.890 ;
        RECT 362.195 41.110 362.475 51.410 ;
        RECT 363.075 45.890 363.355 47.890 ;
        RECT 363.955 41.110 364.235 51.410 ;
        RECT 364.835 45.890 365.115 47.890 ;
        RECT 365.715 41.110 365.995 51.410 ;
        RECT 366.595 45.890 366.875 47.890 ;
        RECT 367.475 41.110 367.755 51.410 ;
        RECT 368.355 45.890 368.635 47.890 ;
        RECT 369.235 41.110 369.515 51.410 ;
        RECT 370.115 45.890 370.395 47.890 ;
        RECT 370.995 45.890 371.275 47.890 ;
        RECT 371.875 45.890 372.155 47.890 ;
        RECT 372.560 45.890 372.850 47.890 ;
        RECT 373.360 45.890 373.650 47.890 ;
        RECT 374.055 45.890 374.335 47.890 ;
        RECT 374.935 45.890 375.215 47.890 ;
        RECT 375.815 45.890 376.095 47.890 ;
        RECT 376.695 45.890 376.975 47.890 ;
        RECT 377.575 45.890 377.855 47.890 ;
        RECT 378.455 41.225 378.735 51.410 ;
        RECT 379.335 45.890 379.615 47.890 ;
        RECT 380.215 41.225 380.495 51.410 ;
        RECT 381.095 45.890 381.375 47.890 ;
        RECT 381.975 41.225 382.255 51.410 ;
        RECT 382.855 45.890 383.135 47.890 ;
        RECT 383.735 41.225 384.015 51.410 ;
        RECT 384.615 45.890 384.895 47.890 ;
        RECT 385.495 41.225 385.775 51.410 ;
        RECT 386.375 45.890 386.655 47.890 ;
        RECT 387.255 41.225 387.535 51.410 ;
        RECT 388.135 45.890 388.415 47.890 ;
        RECT 335.795 40.310 369.515 41.110 ;
        RECT 378.255 40.855 378.935 41.225 ;
        RECT 380.015 40.855 380.695 41.225 ;
        RECT 381.775 40.855 382.455 41.225 ;
        RECT 383.535 40.855 384.215 41.225 ;
        RECT 385.295 40.855 385.975 41.225 ;
        RECT 387.055 40.855 387.735 41.225 ;
        RECT 330.700 33.530 330.990 35.530 ;
        RECT 331.395 33.530 331.675 35.530 ;
        RECT 332.275 33.530 332.555 35.530 ;
        RECT 333.155 33.530 333.435 35.530 ;
        RECT 334.035 33.530 334.315 35.530 ;
        RECT 330.120 29.495 331.290 29.825 ;
        RECT 334.915 28.970 335.195 39.045 ;
        RECT 335.795 30.015 336.075 40.310 ;
        RECT 335.485 29.495 336.335 29.825 ;
        RECT 336.675 28.970 336.955 39.045 ;
        RECT 337.555 30.015 337.835 40.310 ;
        RECT 337.095 29.495 338.295 29.825 ;
        RECT 338.435 28.970 338.715 39.045 ;
        RECT 339.315 30.015 339.595 40.310 ;
        RECT 338.855 29.495 340.055 29.825 ;
        RECT 340.195 28.970 340.475 39.045 ;
        RECT 341.075 30.015 341.355 40.310 ;
        RECT 340.615 29.495 341.815 29.825 ;
        RECT 341.955 28.970 342.235 39.045 ;
        RECT 342.835 30.015 343.115 40.310 ;
        RECT 342.375 29.495 343.575 29.825 ;
        RECT 343.715 28.970 343.995 39.045 ;
        RECT 344.595 30.015 344.875 40.310 ;
        RECT 344.135 29.495 345.335 29.825 ;
        RECT 345.475 28.970 345.755 39.045 ;
        RECT 346.355 30.015 346.635 40.310 ;
        RECT 345.895 29.495 347.095 29.825 ;
        RECT 347.235 28.970 347.515 39.045 ;
        RECT 348.115 30.015 348.395 40.310 ;
        RECT 347.655 29.495 348.855 29.825 ;
        RECT 348.995 28.970 349.275 39.045 ;
        RECT 349.875 30.015 350.155 40.310 ;
        RECT 349.415 29.495 350.615 29.825 ;
        RECT 350.755 28.970 351.035 39.045 ;
        RECT 351.635 30.015 351.915 40.310 ;
        RECT 351.175 29.495 352.375 29.825 ;
        RECT 352.515 28.970 352.795 39.045 ;
        RECT 353.395 30.015 353.675 40.310 ;
        RECT 352.935 29.495 354.135 29.825 ;
        RECT 354.275 28.970 354.555 39.045 ;
        RECT 355.155 30.015 355.435 40.310 ;
        RECT 354.695 29.495 355.895 29.825 ;
        RECT 356.035 28.970 356.315 39.045 ;
        RECT 356.915 30.015 357.195 40.310 ;
        RECT 356.455 29.495 357.655 29.825 ;
        RECT 357.795 28.970 358.075 39.045 ;
        RECT 358.675 30.015 358.955 40.310 ;
        RECT 358.215 29.495 359.415 29.825 ;
        RECT 359.555 28.970 359.835 39.045 ;
        RECT 360.435 30.015 360.715 40.310 ;
        RECT 359.975 29.495 361.175 29.825 ;
        RECT 361.315 28.970 361.595 39.045 ;
        RECT 362.195 30.015 362.475 40.310 ;
        RECT 361.735 29.495 362.935 29.825 ;
        RECT 363.075 28.970 363.355 39.045 ;
        RECT 363.955 30.015 364.235 40.310 ;
        RECT 363.495 29.495 364.695 29.825 ;
        RECT 364.835 28.970 365.115 39.045 ;
        RECT 365.715 30.015 365.995 40.310 ;
        RECT 365.255 29.495 366.455 29.825 ;
        RECT 366.595 28.970 366.875 39.045 ;
        RECT 367.475 30.015 367.755 40.310 ;
        RECT 367.015 29.495 368.215 29.825 ;
        RECT 368.355 28.970 368.635 39.045 ;
        RECT 369.235 30.015 369.515 40.310 ;
        RECT 378.455 40.245 378.735 40.855 ;
        RECT 368.980 29.495 369.830 29.825 ;
        RECT 370.115 28.970 370.395 39.045 ;
        RECT 370.995 33.530 371.275 35.530 ;
        RECT 371.875 33.530 372.155 35.530 ;
        RECT 372.560 33.530 372.850 35.530 ;
        RECT 373.360 33.530 373.650 35.530 ;
        RECT 374.055 33.530 374.335 35.530 ;
        RECT 374.935 33.530 375.215 35.530 ;
        RECT 375.815 33.530 376.095 35.530 ;
        RECT 376.695 33.530 376.975 35.530 ;
        RECT 377.575 33.530 377.855 35.530 ;
        RECT 378.455 33.530 378.735 35.530 ;
        RECT 328.700 28.170 370.395 28.970 ;
        RECT 232.500 25.410 232.780 26.410 ;
        RECT 233.380 25.410 233.660 26.410 ;
        RECT 234.260 25.410 234.540 26.410 ;
        RECT 235.140 25.410 235.420 26.410 ;
        RECT 236.020 25.410 236.300 26.410 ;
        RECT 236.900 25.410 237.180 26.410 ;
        RECT 237.625 25.410 237.915 26.410 ;
        RECT 238.345 25.410 238.635 26.410 ;
        RECT 239.080 25.410 239.360 26.410 ;
        RECT 239.960 25.410 240.240 26.410 ;
        RECT 240.840 24.780 241.120 28.170 ;
        RECT 239.175 24.260 240.935 24.590 ;
        RECT 241.720 23.215 242.000 27.040 ;
        RECT 242.600 24.780 242.880 28.170 ;
        RECT 243.480 23.215 243.760 27.040 ;
        RECT 244.360 24.780 244.640 28.170 ;
        RECT 245.240 23.215 245.520 27.040 ;
        RECT 246.120 24.780 246.400 28.170 ;
        RECT 247.000 23.215 247.280 27.040 ;
        RECT 247.880 24.780 248.160 28.170 ;
        RECT 248.760 23.215 249.040 27.040 ;
        RECT 249.640 24.780 249.920 28.170 ;
        RECT 250.520 23.215 250.800 27.040 ;
        RECT 251.400 24.780 251.680 28.170 ;
        RECT 252.280 23.215 252.560 27.040 ;
        RECT 253.160 24.780 253.440 28.170 ;
        RECT 254.040 23.215 254.320 27.040 ;
        RECT 254.920 24.780 255.200 28.170 ;
        RECT 255.800 23.215 256.080 27.040 ;
        RECT 256.680 24.780 256.960 28.170 ;
        RECT 257.560 23.215 257.840 27.040 ;
        RECT 258.440 24.780 258.720 28.170 ;
        RECT 259.320 23.215 259.600 27.040 ;
        RECT 260.200 24.780 260.480 28.170 ;
        RECT 261.080 23.215 261.360 27.040 ;
        RECT 261.960 24.780 262.240 28.170 ;
        RECT 262.840 23.215 263.120 27.040 ;
        RECT 263.720 24.780 264.000 28.170 ;
        RECT 264.600 23.215 264.880 27.040 ;
        RECT 265.480 24.780 265.760 28.170 ;
        RECT 266.360 23.215 266.640 27.040 ;
        RECT 267.240 24.780 267.520 28.170 ;
        RECT 268.120 23.215 268.400 27.040 ;
        RECT 269.000 24.780 269.280 28.170 ;
        RECT 269.880 23.215 270.160 27.040 ;
        RECT 270.760 24.780 271.040 28.170 ;
        RECT 271.640 23.215 271.920 27.040 ;
        RECT 272.520 24.780 272.800 28.170 ;
        RECT 273.400 23.215 273.680 27.040 ;
        RECT 274.280 24.780 274.560 28.170 ;
        RECT 275.160 23.215 275.440 27.040 ;
        RECT 276.040 24.780 276.320 28.170 ;
        RECT 276.920 25.410 277.200 26.410 ;
        RECT 277.800 25.410 278.080 26.410 ;
        RECT 278.680 25.410 278.960 26.410 ;
        RECT 279.560 25.410 279.840 26.410 ;
        RECT 280.285 25.410 280.575 26.410 ;
        RECT 280.785 24.590 281.115 24.635 ;
        RECT 279.945 24.260 281.115 24.590 ;
        RECT 241.720 22.415 275.440 23.215 ;
        RECT 231.620 18.925 231.900 19.925 ;
        RECT 232.500 18.925 232.780 19.925 ;
        RECT 233.380 18.925 233.660 19.925 ;
        RECT 234.260 18.925 234.540 19.925 ;
        RECT 235.140 18.925 235.420 19.925 ;
        RECT 236.020 18.925 236.300 19.925 ;
        RECT 236.900 18.925 237.180 19.925 ;
        RECT 237.625 18.925 237.915 19.925 ;
        RECT 238.345 18.925 238.635 19.925 ;
        RECT 239.080 18.925 239.360 19.925 ;
        RECT 239.960 18.925 240.240 19.925 ;
        RECT 240.840 18.925 241.120 19.925 ;
        RECT 241.720 18.295 242.000 22.415 ;
        RECT 242.355 20.745 243.125 21.035 ;
        RECT 242.600 18.925 242.880 19.925 ;
        RECT 243.480 18.295 243.760 22.415 ;
        RECT 244.360 18.925 244.640 19.925 ;
        RECT 245.240 18.295 245.520 22.415 ;
        RECT 246.120 18.925 246.400 19.925 ;
        RECT 247.000 18.295 247.280 22.415 ;
        RECT 247.880 18.925 248.160 19.925 ;
        RECT 248.760 18.295 249.040 22.415 ;
        RECT 249.640 18.925 249.920 19.925 ;
        RECT 250.520 18.295 250.800 22.415 ;
        RECT 251.400 18.925 251.680 19.925 ;
        RECT 252.280 18.295 252.560 22.415 ;
        RECT 253.160 18.925 253.440 19.925 ;
        RECT 254.040 18.295 254.320 22.415 ;
        RECT 254.920 18.925 255.200 19.925 ;
        RECT 255.800 18.295 256.080 22.415 ;
        RECT 256.680 18.925 256.960 19.925 ;
        RECT 257.560 18.295 257.840 22.415 ;
        RECT 258.440 18.925 258.720 19.925 ;
        RECT 259.320 18.295 259.600 22.415 ;
        RECT 260.200 18.925 260.480 19.925 ;
        RECT 261.080 18.295 261.360 22.415 ;
        RECT 261.960 18.925 262.240 19.925 ;
        RECT 262.840 18.295 263.120 22.415 ;
        RECT 263.720 18.925 264.000 19.925 ;
        RECT 264.600 18.295 264.880 22.415 ;
        RECT 265.480 18.925 265.760 19.925 ;
        RECT 266.360 18.295 266.640 22.415 ;
        RECT 267.240 18.925 267.520 19.925 ;
        RECT 268.120 18.295 268.400 22.415 ;
        RECT 269.000 18.925 269.280 19.925 ;
        RECT 269.880 18.295 270.160 22.415 ;
        RECT 270.760 18.925 271.040 19.925 ;
        RECT 271.640 18.295 271.920 22.415 ;
        RECT 272.520 18.925 272.800 19.925 ;
        RECT 273.400 18.295 273.680 22.415 ;
        RECT 274.280 18.925 274.560 19.925 ;
        RECT 275.160 18.295 275.440 22.415 ;
        RECT 276.040 18.925 276.320 19.925 ;
        RECT 276.920 18.925 277.200 19.925 ;
        RECT 277.800 18.925 278.080 19.925 ;
        RECT 278.680 18.925 278.960 19.925 ;
        RECT 279.560 18.925 279.840 19.925 ;
        RECT 280.285 18.925 280.575 19.925 ;
        RECT 225.260 15.875 225.940 16.245 ;
        RECT 227.020 15.875 227.700 16.245 ;
        RECT 228.780 15.875 229.460 16.245 ;
        RECT 230.540 15.875 231.220 16.245 ;
        RECT 280.785 15.585 281.115 24.260 ;
        RECT 280.365 15.255 281.535 15.585 ;
        RECT 328.700 7.125 329.300 28.170 ;
        RECT 330.660 25.410 330.950 26.410 ;
        RECT 331.395 25.410 331.675 26.410 ;
        RECT 332.275 25.410 332.555 26.410 ;
        RECT 333.155 25.410 333.435 26.410 ;
        RECT 334.035 25.410 334.315 26.410 ;
        RECT 334.915 24.780 335.195 28.170 ;
        RECT 330.120 24.590 330.450 24.635 ;
        RECT 330.120 24.260 331.290 24.590 ;
        RECT 330.120 15.585 330.450 24.260 ;
        RECT 335.795 23.215 336.075 27.040 ;
        RECT 336.675 24.780 336.955 28.170 ;
        RECT 337.555 23.215 337.835 27.040 ;
        RECT 338.435 24.780 338.715 28.170 ;
        RECT 339.315 23.215 339.595 27.040 ;
        RECT 340.195 24.780 340.475 28.170 ;
        RECT 341.075 23.215 341.355 27.040 ;
        RECT 341.955 24.780 342.235 28.170 ;
        RECT 342.835 23.215 343.115 27.040 ;
        RECT 343.715 24.780 343.995 28.170 ;
        RECT 344.595 23.215 344.875 27.040 ;
        RECT 345.475 24.780 345.755 28.170 ;
        RECT 346.355 23.215 346.635 27.040 ;
        RECT 347.235 24.780 347.515 28.170 ;
        RECT 348.115 23.215 348.395 27.040 ;
        RECT 348.995 24.780 349.275 28.170 ;
        RECT 349.875 23.215 350.155 27.040 ;
        RECT 350.755 24.780 351.035 28.170 ;
        RECT 351.635 23.215 351.915 27.040 ;
        RECT 352.515 24.780 352.795 28.170 ;
        RECT 353.395 23.215 353.675 27.040 ;
        RECT 354.275 24.780 354.555 28.170 ;
        RECT 355.155 23.215 355.435 27.040 ;
        RECT 356.035 24.780 356.315 28.170 ;
        RECT 356.915 23.215 357.195 27.040 ;
        RECT 357.795 24.780 358.075 28.170 ;
        RECT 358.675 23.215 358.955 27.040 ;
        RECT 359.555 24.780 359.835 28.170 ;
        RECT 360.435 23.215 360.715 27.040 ;
        RECT 361.315 24.780 361.595 28.170 ;
        RECT 362.195 23.215 362.475 27.040 ;
        RECT 363.075 24.780 363.355 28.170 ;
        RECT 363.955 23.215 364.235 27.040 ;
        RECT 364.835 24.780 365.115 28.170 ;
        RECT 365.715 23.215 365.995 27.040 ;
        RECT 366.595 24.780 366.875 28.170 ;
        RECT 367.475 23.215 367.755 27.040 ;
        RECT 368.355 24.780 368.635 28.170 ;
        RECT 369.235 23.215 369.515 27.040 ;
        RECT 370.115 24.780 370.395 28.170 ;
        RECT 370.995 25.410 371.275 26.410 ;
        RECT 371.875 25.410 372.155 26.410 ;
        RECT 372.600 25.410 372.890 26.410 ;
        RECT 373.320 25.410 373.610 26.410 ;
        RECT 374.055 25.410 374.335 26.410 ;
        RECT 374.935 25.410 375.215 26.410 ;
        RECT 375.815 25.410 376.095 26.410 ;
        RECT 376.695 25.410 376.975 26.410 ;
        RECT 377.575 25.410 377.855 26.410 ;
        RECT 378.455 25.410 378.735 26.410 ;
        RECT 370.300 24.260 372.060 24.590 ;
        RECT 335.795 22.415 369.515 23.215 ;
        RECT 379.335 22.860 379.615 39.045 ;
        RECT 380.215 30.015 380.495 40.855 ;
        RECT 379.905 29.495 380.755 29.825 ;
        RECT 330.660 18.925 330.950 19.925 ;
        RECT 331.395 18.925 331.675 19.925 ;
        RECT 332.275 18.925 332.555 19.925 ;
        RECT 333.155 18.925 333.435 19.925 ;
        RECT 334.035 18.925 334.315 19.925 ;
        RECT 334.915 18.925 335.195 19.925 ;
        RECT 335.795 18.295 336.075 22.415 ;
        RECT 336.675 18.925 336.955 19.925 ;
        RECT 337.555 18.295 337.835 22.415 ;
        RECT 338.435 18.925 338.715 19.925 ;
        RECT 339.315 18.295 339.595 22.415 ;
        RECT 340.195 18.925 340.475 19.925 ;
        RECT 341.075 18.295 341.355 22.415 ;
        RECT 341.955 18.925 342.235 19.925 ;
        RECT 342.835 18.295 343.115 22.415 ;
        RECT 343.715 18.925 343.995 19.925 ;
        RECT 344.595 18.295 344.875 22.415 ;
        RECT 345.475 18.925 345.755 19.925 ;
        RECT 346.355 18.295 346.635 22.415 ;
        RECT 347.235 18.925 347.515 19.925 ;
        RECT 348.115 18.295 348.395 22.415 ;
        RECT 348.995 18.925 349.275 19.925 ;
        RECT 349.875 18.295 350.155 22.415 ;
        RECT 350.755 18.925 351.035 19.925 ;
        RECT 351.635 18.295 351.915 22.415 ;
        RECT 352.515 18.925 352.795 19.925 ;
        RECT 353.395 18.295 353.675 22.415 ;
        RECT 354.275 18.925 354.555 19.925 ;
        RECT 355.155 18.295 355.435 22.415 ;
        RECT 356.035 18.925 356.315 19.925 ;
        RECT 356.915 18.295 357.195 22.415 ;
        RECT 357.795 18.925 358.075 19.925 ;
        RECT 358.675 18.295 358.955 22.415 ;
        RECT 359.555 18.925 359.835 19.925 ;
        RECT 360.435 18.295 360.715 22.415 ;
        RECT 361.315 18.925 361.595 19.925 ;
        RECT 362.195 18.295 362.475 22.415 ;
        RECT 363.075 18.925 363.355 19.925 ;
        RECT 363.955 18.295 364.235 22.415 ;
        RECT 364.835 18.925 365.115 19.925 ;
        RECT 365.715 18.295 365.995 22.415 ;
        RECT 366.595 18.925 366.875 19.925 ;
        RECT 367.475 18.295 367.755 22.415 ;
        RECT 368.110 20.745 368.880 21.035 ;
        RECT 368.355 18.925 368.635 19.925 ;
        RECT 369.235 18.295 369.515 22.415 ;
        RECT 370.115 18.925 370.395 19.925 ;
        RECT 370.995 18.925 371.275 19.925 ;
        RECT 371.875 18.925 372.155 19.925 ;
        RECT 372.600 18.925 372.890 19.925 ;
        RECT 373.320 18.925 373.610 19.925 ;
        RECT 374.055 18.925 374.335 19.925 ;
        RECT 374.935 18.925 375.215 19.925 ;
        RECT 375.815 18.925 376.095 19.925 ;
        RECT 376.695 18.925 376.975 19.925 ;
        RECT 377.575 18.925 377.855 19.925 ;
        RECT 378.455 18.925 378.735 19.925 ;
        RECT 379.335 18.925 379.615 19.925 ;
        RECT 380.215 16.245 380.495 27.040 ;
        RECT 381.095 22.860 381.375 39.045 ;
        RECT 381.975 30.015 382.255 40.855 ;
        RECT 381.515 29.495 382.715 29.825 ;
        RECT 381.095 18.925 381.375 19.925 ;
        RECT 381.975 16.245 382.255 27.040 ;
        RECT 382.855 22.860 383.135 39.045 ;
        RECT 383.735 30.015 384.015 40.855 ;
        RECT 383.275 29.495 384.475 29.825 ;
        RECT 382.855 18.925 383.135 19.925 ;
        RECT 383.735 16.245 384.015 27.040 ;
        RECT 384.615 22.860 384.895 39.045 ;
        RECT 385.495 30.015 385.775 40.855 ;
        RECT 387.255 40.245 387.535 40.855 ;
        RECT 389.015 40.595 389.295 51.410 ;
        RECT 389.895 45.890 390.175 47.890 ;
        RECT 390.775 40.595 391.055 51.410 ;
        RECT 391.655 45.890 391.935 47.890 ;
        RECT 392.535 40.595 392.815 51.410 ;
        RECT 393.415 45.890 393.695 47.890 ;
        RECT 394.295 40.595 394.575 51.410 ;
        RECT 395.175 45.890 395.455 47.890 ;
        RECT 396.055 40.595 396.335 51.410 ;
        RECT 396.935 45.890 397.215 47.890 ;
        RECT 397.815 40.595 398.095 51.410 ;
        RECT 398.695 45.890 398.975 47.890 ;
        RECT 399.575 45.890 399.855 47.890 ;
        RECT 400.455 45.890 400.735 47.890 ;
        RECT 401.335 45.890 401.615 47.890 ;
        RECT 402.215 45.890 402.495 47.890 ;
        RECT 402.900 45.890 403.190 47.890 ;
        RECT 408.495 40.855 409.175 41.225 ;
        RECT 388.815 40.225 389.495 40.595 ;
        RECT 390.575 40.225 391.255 40.595 ;
        RECT 392.335 40.225 393.015 40.595 ;
        RECT 394.095 40.225 394.775 40.595 ;
        RECT 395.855 40.225 396.535 40.595 ;
        RECT 397.615 40.225 398.295 40.595 ;
        RECT 385.035 29.495 386.235 29.825 ;
        RECT 384.615 18.925 384.895 19.925 ;
        RECT 385.495 16.245 385.775 27.040 ;
        RECT 386.375 22.860 386.655 39.045 ;
        RECT 387.255 33.530 387.535 35.530 ;
        RECT 388.135 33.530 388.415 35.530 ;
        RECT 389.015 33.530 389.295 35.530 ;
        RECT 387.255 25.410 387.535 26.410 ;
        RECT 388.135 25.410 388.415 26.410 ;
        RECT 389.015 25.410 389.295 26.410 ;
        RECT 389.895 22.860 390.175 39.045 ;
        RECT 390.775 30.015 391.055 40.225 ;
        RECT 390.315 29.495 391.515 29.825 ;
        RECT 386.375 18.925 386.655 19.925 ;
        RECT 387.255 18.925 387.535 19.925 ;
        RECT 388.135 18.925 388.415 19.925 ;
        RECT 389.015 18.925 389.295 19.925 ;
        RECT 389.895 18.925 390.175 19.925 ;
        RECT 390.775 18.295 391.055 27.040 ;
        RECT 391.655 22.860 391.935 39.045 ;
        RECT 392.535 30.015 392.815 40.225 ;
        RECT 392.075 29.495 393.275 29.825 ;
        RECT 391.655 18.925 391.935 19.925 ;
        RECT 392.535 18.295 392.815 27.040 ;
        RECT 393.415 23.380 393.695 39.045 ;
        RECT 394.295 30.015 394.575 40.225 ;
        RECT 393.835 29.495 395.035 29.825 ;
        RECT 393.305 21.050 393.805 23.380 ;
        RECT 393.265 20.730 393.845 21.050 ;
        RECT 393.415 18.925 393.695 19.925 ;
        RECT 394.295 18.295 394.575 27.040 ;
        RECT 395.175 22.860 395.455 39.045 ;
        RECT 396.055 30.015 396.335 40.225 ;
        RECT 395.800 29.495 396.650 29.825 ;
        RECT 395.175 18.925 395.455 19.925 ;
        RECT 396.055 18.295 396.335 27.040 ;
        RECT 396.935 22.860 397.215 39.045 ;
        RECT 397.815 33.530 398.095 35.530 ;
        RECT 398.695 33.530 398.975 35.530 ;
        RECT 399.575 33.530 399.855 35.530 ;
        RECT 400.455 33.530 400.735 35.530 ;
        RECT 401.335 33.530 401.615 35.530 ;
        RECT 402.215 33.530 402.495 35.530 ;
        RECT 402.900 33.530 403.190 35.530 ;
        RECT 403.580 34.020 403.870 35.020 ;
        RECT 404.315 34.020 404.595 35.020 ;
        RECT 405.195 34.020 405.475 35.020 ;
        RECT 406.075 34.020 406.355 35.020 ;
        RECT 406.955 34.020 407.235 35.020 ;
        RECT 407.835 31.045 408.115 35.650 ;
        RECT 408.715 33.390 408.995 40.855 ;
        RECT 410.475 40.595 410.755 41.205 ;
        RECT 412.015 40.855 412.695 41.225 ;
        RECT 410.275 40.225 410.955 40.595 ;
        RECT 409.595 31.045 409.875 35.650 ;
        RECT 410.475 33.390 410.755 40.225 ;
        RECT 411.355 31.045 411.635 35.650 ;
        RECT 412.235 33.390 412.515 40.855 ;
        RECT 413.995 40.595 414.275 41.205 ;
        RECT 415.535 40.855 416.215 41.225 ;
        RECT 413.795 40.225 414.475 40.595 ;
        RECT 413.115 31.045 413.395 35.650 ;
        RECT 413.995 33.390 414.275 40.225 ;
        RECT 414.875 31.045 415.155 35.650 ;
        RECT 415.755 33.390 416.035 40.855 ;
        RECT 417.515 40.595 417.795 41.205 ;
        RECT 419.055 40.855 419.735 41.225 ;
        RECT 417.315 40.225 417.995 40.595 ;
        RECT 416.635 31.045 416.915 35.650 ;
        RECT 417.515 33.390 417.795 40.225 ;
        RECT 418.395 31.045 418.675 35.650 ;
        RECT 419.275 33.390 419.555 40.855 ;
        RECT 421.035 40.595 421.315 41.205 ;
        RECT 420.835 40.225 421.515 40.595 ;
        RECT 420.155 31.045 420.435 35.650 ;
        RECT 421.035 33.390 421.315 40.225 ;
        RECT 423.685 36.430 425.350 36.720 ;
        RECT 427.395 36.405 427.995 53.925 ;
        RECT 421.915 31.045 422.195 35.650 ;
        RECT 422.795 34.020 423.075 35.020 ;
        RECT 423.675 34.020 423.955 35.020 ;
        RECT 424.555 34.020 424.835 35.020 ;
        RECT 425.435 34.020 425.715 35.020 ;
        RECT 426.160 34.020 426.450 35.020 ;
        RECT 423.685 32.320 425.350 32.610 ;
        RECT 428.680 32.295 429.280 79.690 ;
        RECT 407.835 30.545 422.195 31.045 ;
        RECT 397.815 25.410 398.095 26.410 ;
        RECT 398.695 25.410 398.975 26.410 ;
        RECT 399.575 25.410 399.855 26.410 ;
        RECT 400.455 25.410 400.735 26.410 ;
        RECT 401.335 25.410 401.615 26.410 ;
        RECT 402.215 25.410 402.495 26.410 ;
        RECT 402.940 25.410 403.230 26.410 ;
        RECT 403.580 25.410 403.870 26.410 ;
        RECT 404.315 25.410 404.595 26.410 ;
        RECT 405.195 25.410 405.475 26.410 ;
        RECT 406.075 25.410 406.355 26.410 ;
        RECT 406.955 25.410 407.235 26.410 ;
        RECT 407.835 25.410 408.115 26.410 ;
        RECT 408.715 25.410 408.995 26.410 ;
        RECT 409.595 25.410 409.875 26.410 ;
        RECT 410.475 25.410 410.755 26.410 ;
        RECT 411.355 24.780 411.635 30.545 ;
        RECT 397.815 24.260 399.575 24.590 ;
        RECT 411.720 24.260 412.095 24.590 ;
        RECT 412.235 22.915 412.515 27.040 ;
        RECT 413.115 24.780 413.395 30.545 ;
        RECT 412.655 24.260 413.855 24.590 ;
        RECT 413.995 22.915 414.275 27.040 ;
        RECT 414.875 24.780 415.155 30.545 ;
        RECT 414.415 24.260 415.615 24.590 ;
        RECT 415.755 22.915 416.035 27.040 ;
        RECT 416.635 24.780 416.915 30.545 ;
        RECT 416.175 24.260 417.375 24.590 ;
        RECT 417.515 22.915 417.795 27.040 ;
        RECT 418.395 24.780 418.675 30.545 ;
        RECT 419.275 25.410 419.555 26.410 ;
        RECT 420.155 25.410 420.435 26.410 ;
        RECT 421.035 25.410 421.315 26.410 ;
        RECT 421.915 25.410 422.195 26.410 ;
        RECT 422.795 25.410 423.075 26.410 ;
        RECT 423.675 25.410 423.955 26.410 ;
        RECT 424.555 25.410 424.835 26.410 ;
        RECT 425.435 25.410 425.715 26.410 ;
        RECT 426.160 25.410 426.450 26.410 ;
        RECT 417.935 24.260 418.330 24.590 ;
        RECT 412.235 22.415 417.795 22.915 ;
        RECT 396.935 18.925 397.215 19.925 ;
        RECT 397.815 18.925 398.095 19.925 ;
        RECT 398.695 18.925 398.975 19.925 ;
        RECT 399.575 18.925 399.855 19.925 ;
        RECT 400.455 18.925 400.735 19.925 ;
        RECT 401.335 18.925 401.615 19.925 ;
        RECT 402.215 18.925 402.495 19.925 ;
        RECT 402.940 18.925 403.230 19.925 ;
        RECT 403.580 18.925 403.870 19.925 ;
        RECT 404.315 18.925 404.595 19.925 ;
        RECT 405.195 18.925 405.475 19.925 ;
        RECT 406.075 18.925 406.355 19.925 ;
        RECT 406.955 18.925 407.235 19.925 ;
        RECT 407.835 18.925 408.115 19.925 ;
        RECT 408.715 18.925 408.995 19.925 ;
        RECT 409.595 18.925 409.875 19.925 ;
        RECT 410.475 18.925 410.755 19.925 ;
        RECT 411.355 18.925 411.635 19.925 ;
        RECT 412.235 18.295 412.515 22.415 ;
        RECT 413.115 18.925 413.395 19.925 ;
        RECT 413.995 18.295 414.275 22.415 ;
        RECT 414.875 18.925 415.155 19.925 ;
        RECT 415.755 18.295 416.035 22.415 ;
        RECT 416.635 18.925 416.915 19.925 ;
        RECT 417.515 18.295 417.795 22.415 ;
        RECT 418.395 18.925 418.675 19.925 ;
        RECT 419.275 18.925 419.555 19.925 ;
        RECT 420.155 18.925 420.435 19.925 ;
        RECT 421.035 18.925 421.315 19.925 ;
        RECT 421.915 18.925 422.195 19.925 ;
        RECT 422.795 18.925 423.075 19.925 ;
        RECT 423.675 18.925 423.955 19.925 ;
        RECT 424.555 18.925 424.835 19.925 ;
        RECT 425.435 18.925 425.715 19.925 ;
        RECT 426.160 18.925 426.450 19.925 ;
        RECT 416.915 17.775 418.310 18.105 ;
        RECT 429.890 17.755 430.220 189.825 ;
        RECT 380.015 15.875 380.695 16.245 ;
        RECT 381.775 15.875 382.455 16.245 ;
        RECT 383.535 15.875 384.215 16.245 ;
        RECT 385.295 15.875 385.975 16.245 ;
        RECT 431.020 15.585 431.350 191.225 ;
        RECT 432.150 53.295 432.480 153.515 ;
        RECT 433.280 51.540 433.610 154.145 ;
        RECT 446.765 118.245 449.935 118.575 ;
        RECT 460.585 118.245 463.755 118.575 ;
        RECT 489.800 118.245 492.970 118.575 ;
        RECT 444.015 113.055 444.305 115.055 ;
        RECT 444.690 113.055 444.970 115.055 ;
        RECT 445.570 113.055 445.850 115.055 ;
        RECT 446.450 113.055 446.730 115.055 ;
        RECT 434.835 88.950 435.125 90.450 ;
        RECT 435.470 88.950 435.750 90.450 ;
        RECT 436.350 88.950 436.630 90.450 ;
        RECT 437.230 88.950 437.510 90.450 ;
        RECT 438.990 88.950 439.270 90.450 ;
        RECT 440.750 88.950 441.030 90.450 ;
        RECT 441.630 88.950 441.910 90.450 ;
        RECT 442.510 88.950 442.790 90.450 ;
        RECT 443.135 88.950 443.425 90.450 ;
        RECT 444.055 88.950 444.345 90.450 ;
        RECT 444.690 88.950 444.970 90.450 ;
        RECT 445.570 88.950 445.850 90.450 ;
        RECT 446.450 88.950 446.730 90.450 ;
        RECT 447.325 88.705 447.615 118.245 ;
        RECT 448.210 113.055 448.490 115.055 ;
        RECT 448.210 88.950 448.490 90.450 ;
        RECT 449.085 88.705 449.375 118.245 ;
        RECT 449.970 113.055 450.250 115.055 ;
        RECT 450.850 113.055 451.130 115.055 ;
        RECT 451.730 113.055 452.010 115.055 ;
        RECT 452.395 113.055 452.685 115.055 ;
        RECT 457.835 113.055 458.125 115.055 ;
        RECT 458.510 113.055 458.790 115.055 ;
        RECT 459.390 113.055 459.670 115.055 ;
        RECT 460.270 113.055 460.550 115.055 ;
        RECT 461.145 93.895 461.435 118.055 ;
        RECT 462.030 113.055 462.310 115.055 ;
        RECT 462.920 93.895 463.210 118.055 ;
        RECT 463.790 113.055 464.070 115.055 ;
        RECT 464.670 113.055 464.950 115.055 ;
        RECT 465.550 113.055 465.830 115.055 ;
        RECT 466.215 113.055 466.505 115.055 ;
        RECT 467.575 113.055 467.865 115.055 ;
        RECT 468.250 113.055 468.530 115.055 ;
        RECT 469.530 113.055 469.810 115.055 ;
        RECT 470.810 113.055 471.090 115.055 ;
        RECT 473.790 109.865 474.080 118.055 ;
        RECT 476.780 113.055 477.060 115.055 ;
        RECT 479.760 109.865 480.050 118.055 ;
        RECT 482.750 113.055 483.030 115.055 ;
        RECT 484.030 113.055 484.310 115.055 ;
        RECT 485.310 113.055 485.590 115.055 ;
        RECT 485.975 113.055 486.265 115.055 ;
        RECT 487.050 113.055 487.340 115.055 ;
        RECT 487.725 113.055 488.005 115.055 ;
        RECT 488.605 113.055 488.885 115.055 ;
        RECT 489.485 113.055 489.765 115.055 ;
        RECT 473.485 109.535 474.385 109.865 ;
        RECT 479.455 109.535 480.355 109.865 ;
        RECT 473.790 105.310 474.080 109.535 ;
        RECT 479.760 105.310 480.050 109.535 ;
        RECT 490.360 107.055 490.650 118.055 ;
        RECT 491.245 113.055 491.525 115.055 ;
        RECT 492.120 107.055 492.410 118.055 ;
        RECT 493.005 113.055 493.285 115.055 ;
        RECT 493.885 113.055 494.165 115.055 ;
        RECT 494.765 113.055 495.045 115.055 ;
        RECT 495.430 113.055 495.720 115.055 ;
        RECT 496.780 113.055 497.070 115.055 ;
        RECT 497.455 113.055 497.735 115.055 ;
        RECT 498.335 113.055 498.615 115.055 ;
        RECT 499.215 113.055 499.495 115.055 ;
        RECT 500.090 109.865 500.380 118.055 ;
        RECT 500.975 113.055 501.255 115.055 ;
        RECT 501.850 109.865 502.140 118.055 ;
        RECT 502.735 113.055 503.015 115.055 ;
        RECT 503.615 113.055 503.895 115.055 ;
        RECT 504.495 113.055 504.775 115.055 ;
        RECT 505.160 113.055 505.450 115.055 ;
        RECT 500.090 109.535 502.140 109.865 ;
        RECT 500.090 107.705 500.380 109.535 ;
        RECT 501.850 107.705 502.140 109.535 ;
        RECT 499.210 107.375 503.020 107.705 ;
        RECT 489.480 106.725 493.290 107.055 ;
        RECT 473.790 104.980 480.050 105.310 ;
        RECT 487.540 104.980 488.870 105.310 ;
        RECT 472.625 94.465 472.915 95.965 ;
        RECT 473.260 94.465 473.540 95.965 ;
        RECT 474.140 94.465 474.420 95.965 ;
        RECT 475.015 94.085 475.305 104.980 ;
        RECT 456.935 93.565 467.405 93.895 ;
        RECT 473.940 93.565 475.350 93.895 ;
        RECT 453.275 91.565 453.565 93.065 ;
        RECT 453.910 91.565 454.190 93.065 ;
        RECT 455.190 91.565 455.470 93.065 ;
        RECT 456.470 91.565 456.750 93.065 ;
        RECT 449.970 88.950 450.250 90.450 ;
        RECT 450.850 88.950 451.130 90.450 ;
        RECT 451.730 88.950 452.010 90.450 ;
        RECT 452.355 88.950 452.645 90.450 ;
        RECT 453.275 88.950 453.565 90.450 ;
        RECT 453.910 88.950 454.190 90.450 ;
        RECT 455.190 88.950 455.470 90.450 ;
        RECT 456.470 88.950 456.750 90.450 ;
        RECT 462.025 88.705 462.315 93.565 ;
        RECT 467.590 91.565 467.870 93.065 ;
        RECT 468.870 91.565 469.150 93.065 ;
        RECT 470.150 91.565 470.430 93.065 ;
        RECT 470.775 91.565 471.065 93.065 ;
        RECT 475.895 92.670 476.185 96.345 ;
        RECT 476.775 94.085 477.065 104.980 ;
        RECT 477.670 92.670 477.960 96.345 ;
        RECT 478.535 94.085 478.825 104.980 ;
        RECT 487.050 99.275 487.340 101.275 ;
        RECT 487.725 99.275 488.005 101.275 ;
        RECT 488.605 99.275 488.885 101.275 ;
        RECT 479.420 94.465 479.700 95.965 ;
        RECT 480.300 94.465 480.580 95.965 ;
        RECT 480.925 94.465 481.215 95.965 ;
        RECT 489.480 95.760 489.770 106.725 ;
        RECT 475.895 92.380 477.960 92.670 ;
        RECT 467.590 88.950 467.870 90.450 ;
        RECT 468.870 88.950 469.150 90.450 ;
        RECT 470.150 88.950 470.430 90.450 ;
        RECT 470.775 88.950 471.065 90.450 ;
        RECT 472.625 88.950 472.915 90.450 ;
        RECT 473.260 88.950 473.540 90.450 ;
        RECT 474.140 88.950 474.420 90.450 ;
        RECT 475.020 88.950 475.300 90.450 ;
        RECT 475.895 88.705 476.185 92.380 ;
        RECT 476.780 88.950 477.060 90.450 ;
        RECT 477.670 88.705 477.960 92.380 ;
        RECT 490.360 91.225 490.650 104.790 ;
        RECT 491.240 95.760 491.530 106.725 ;
        RECT 492.120 91.225 492.410 104.790 ;
        RECT 493.000 95.760 493.290 106.725 ;
        RECT 493.885 99.275 494.165 101.275 ;
        RECT 494.765 99.275 495.045 101.275 ;
        RECT 495.430 99.275 495.720 101.275 ;
        RECT 496.820 94.465 497.110 95.965 ;
        RECT 497.455 94.465 497.735 95.965 ;
        RECT 498.335 94.465 498.615 95.965 ;
        RECT 499.210 94.085 499.500 107.375 ;
        RECT 497.640 93.565 498.850 93.895 ;
        RECT 490.360 90.895 492.410 91.225 ;
        RECT 478.540 88.950 478.820 90.450 ;
        RECT 479.420 88.950 479.700 90.450 ;
        RECT 480.300 88.950 480.580 90.450 ;
        RECT 480.925 88.950 481.215 90.450 ;
        RECT 487.090 88.950 487.380 90.450 ;
        RECT 487.725 88.950 488.005 90.450 ;
        RECT 488.605 88.950 488.885 90.450 ;
        RECT 489.485 88.950 489.765 90.450 ;
        RECT 490.360 88.705 490.650 90.895 ;
        RECT 491.245 88.950 491.525 90.450 ;
        RECT 492.120 88.705 492.410 90.895 ;
        RECT 500.090 92.670 500.380 96.345 ;
        RECT 500.970 94.085 501.260 107.375 ;
        RECT 501.850 92.670 502.140 96.345 ;
        RECT 502.730 94.085 503.020 107.375 ;
        RECT 503.615 94.465 503.895 95.965 ;
        RECT 504.495 94.465 504.775 95.965 ;
        RECT 505.120 94.465 505.410 95.965 ;
        RECT 500.090 92.380 502.140 92.670 ;
        RECT 493.005 88.950 493.285 90.450 ;
        RECT 493.885 88.950 494.165 90.450 ;
        RECT 494.765 88.950 495.045 90.450 ;
        RECT 495.390 88.950 495.680 90.450 ;
        RECT 496.820 88.950 497.110 90.450 ;
        RECT 497.455 88.950 497.735 90.450 ;
        RECT 498.335 88.950 498.615 90.450 ;
        RECT 499.215 88.950 499.495 90.450 ;
        RECT 500.090 88.705 500.380 92.380 ;
        RECT 500.975 88.950 501.255 90.450 ;
        RECT 501.850 88.705 502.140 92.380 ;
        RECT 502.735 88.950 503.015 90.450 ;
        RECT 503.615 88.950 503.895 90.450 ;
        RECT 504.495 88.950 504.775 90.450 ;
        RECT 505.120 88.950 505.410 90.450 ;
        RECT 437.545 88.185 440.715 88.515 ;
        RECT 446.765 88.185 449.935 88.515 ;
        RECT 475.335 88.185 478.505 88.515 ;
        RECT 499.530 88.185 502.700 88.515 ;
        RECT 442.430 81.060 445.750 82.060 ;
        RECT 446.450 81.060 449.770 82.060 ;
        RECT 450.470 81.060 453.790 82.060 ;
        RECT 454.490 81.060 457.810 82.060 ;
        RECT 458.510 81.060 461.830 82.060 ;
        RECT 462.530 81.060 465.850 82.060 ;
        RECT 466.550 81.060 469.870 82.060 ;
        RECT 470.570 81.060 473.890 82.060 ;
        RECT 474.590 81.060 477.910 82.060 ;
        RECT 478.610 81.060 481.930 82.060 ;
        RECT 482.630 81.060 485.950 82.060 ;
        RECT 486.650 81.060 489.970 82.060 ;
        RECT 490.670 81.060 493.990 82.060 ;
        RECT 494.690 81.060 498.010 82.060 ;
        RECT 437.510 73.900 437.800 75.900 ;
        RECT 502.640 73.900 502.930 75.900 ;
        RECT 442.430 71.465 447.760 72.465 ;
        RECT 448.460 71.465 451.780 72.465 ;
        RECT 452.480 71.465 455.800 72.465 ;
        RECT 456.500 71.465 459.820 72.465 ;
        RECT 460.520 71.465 463.840 72.465 ;
        RECT 464.540 71.465 467.860 72.465 ;
        RECT 468.560 71.465 471.880 72.465 ;
        RECT 472.580 71.465 475.900 72.465 ;
        RECT 476.600 71.465 479.920 72.465 ;
        RECT 480.620 71.465 483.940 72.465 ;
        RECT 484.640 71.465 487.960 72.465 ;
        RECT 488.660 71.465 491.980 72.465 ;
        RECT 492.680 71.465 496.000 72.465 ;
        RECT 496.700 71.465 498.010 72.465 ;
        RECT 329.700 15.255 330.870 15.585 ;
        RECT 430.180 15.255 431.350 15.585 ;
        RECT 328.195 6.525 329.300 7.125 ;
      LAYER met3 ;
        RECT 3.980 219.260 88.940 220.760 ;
        RECT 147.500 217.090 147.820 217.670 ;
        RECT 147.500 216.490 181.705 217.090 ;
        RECT 143.820 215.490 144.140 216.045 ;
        RECT 143.820 214.890 180.605 215.490 ;
        RECT 143.820 214.865 144.140 214.890 ;
        RECT 49.000 211.340 503.815 214.340 ;
        RECT 73.420 210.510 74.550 210.840 ;
        RECT 74.545 209.880 75.345 210.210 ;
        RECT 75.015 209.085 75.345 209.880 ;
        RECT 75.015 208.755 171.790 209.085 ;
        RECT 54.490 192.630 72.000 208.680 ;
        RECT 74.380 203.085 272.340 205.085 ;
        RECT 121.930 198.070 165.240 198.400 ;
        RECT 121.930 197.440 165.240 197.770 ;
        RECT 167.390 193.930 169.050 193.935 ;
        RECT 167.385 193.600 177.380 193.930 ;
        RECT 176.780 192.800 177.380 193.600 ;
        RECT 54.490 175.380 72.000 191.430 ;
        RECT 74.380 190.725 146.910 192.725 ;
        RECT 147.260 191.215 170.170 192.215 ;
        RECT 280.385 191.225 431.350 191.555 ;
        RECT 225.235 190.575 292.705 190.925 ;
        RECT 279.750 189.825 430.220 190.155 ;
        RECT 167.390 189.820 169.050 189.825 ;
        RECT 167.385 189.490 176.280 189.820 ;
        RECT 175.680 188.690 176.280 189.490 ;
        RECT 279.750 189.035 280.080 189.825 ;
        RECT 183.655 188.705 280.080 189.035 ;
        RECT 73.820 186.690 172.660 187.020 ;
        RECT 184.765 186.885 280.595 187.885 ;
        RECT 74.240 185.365 75.045 186.165 ;
        RECT 172.330 185.890 172.660 186.690 ;
        RECT 242.375 185.755 243.105 186.085 ;
        RECT 214.875 184.855 215.205 185.085 ;
        RECT 216.635 184.855 216.965 185.085 ;
        RECT 218.395 184.855 218.725 185.085 ;
        RECT 220.155 184.855 220.485 185.085 ;
        RECT 214.875 184.355 220.485 184.855 ;
        RECT 225.435 184.855 225.765 185.085 ;
        RECT 227.195 184.855 227.525 185.085 ;
        RECT 228.955 184.855 229.285 185.085 ;
        RECT 230.715 184.855 231.045 185.085 ;
        RECT 225.435 184.355 231.045 184.855 ;
        RECT 242.490 183.930 242.990 185.755 ;
        RECT 74.340 182.605 170.170 183.605 ;
        RECT 213.995 183.430 221.365 183.930 ;
        RECT 213.995 183.200 214.325 183.430 ;
        RECT 215.755 183.200 216.085 183.430 ;
        RECT 217.515 183.200 217.845 183.430 ;
        RECT 219.275 183.200 219.605 183.430 ;
        RECT 221.035 183.200 221.365 183.430 ;
        RECT 224.555 183.430 242.990 183.930 ;
        RECT 224.555 183.200 224.885 183.430 ;
        RECT 226.315 183.200 226.645 183.430 ;
        RECT 228.075 183.200 228.405 183.430 ;
        RECT 229.835 183.200 230.165 183.430 ;
        RECT 231.595 183.200 231.925 183.430 ;
        RECT 182.495 182.220 281.115 182.550 ;
        RECT 182.495 181.785 182.825 182.220 ;
        RECT 73.820 181.455 182.825 181.785 ;
        RECT 123.010 180.575 123.340 180.805 ;
        RECT 124.770 180.575 125.100 180.805 ;
        RECT 126.530 180.575 126.860 180.805 ;
        RECT 128.290 180.575 128.620 180.805 ;
        RECT 130.050 180.575 130.380 180.805 ;
        RECT 111.945 180.075 130.380 180.575 ;
        RECT 133.570 180.575 133.900 180.805 ;
        RECT 135.330 180.575 135.660 180.805 ;
        RECT 137.090 180.575 137.420 180.805 ;
        RECT 138.850 180.575 139.180 180.805 ;
        RECT 140.610 180.575 140.940 180.805 ;
        RECT 133.570 180.075 140.940 180.575 ;
        RECT 184.765 180.400 280.595 181.400 ;
        RECT 111.945 178.250 112.445 180.075 ;
        RECT 123.890 179.150 129.500 179.650 ;
        RECT 123.890 178.920 124.220 179.150 ;
        RECT 125.650 178.920 125.980 179.150 ;
        RECT 127.410 178.920 127.740 179.150 ;
        RECT 129.170 178.920 129.500 179.150 ;
        RECT 134.450 179.150 140.060 179.650 ;
        RECT 134.450 178.920 134.780 179.150 ;
        RECT 136.210 178.920 136.540 179.150 ;
        RECT 137.970 178.920 138.300 179.150 ;
        RECT 139.730 178.920 140.060 179.150 ;
        RECT 111.830 177.920 112.560 178.250 ;
        RECT 279.890 177.840 280.695 178.640 ;
        RECT 74.340 176.120 170.170 177.120 ;
        RECT 172.330 176.985 281.115 177.315 ;
        RECT 74.855 174.970 183.985 175.300 ;
        RECT 74.855 174.180 75.185 174.970 ;
        RECT 74.510 173.850 75.185 174.180 ;
        RECT 178.380 174.185 187.550 174.515 ;
        RECT 62.230 173.080 129.700 173.430 ;
        RECT 178.380 173.385 178.980 174.185 ;
        RECT 185.885 174.180 187.545 174.185 ;
        RECT 73.420 172.450 74.550 172.780 ;
        RECT 72.400 171.550 91.065 172.150 ;
        RECT 184.765 171.790 207.675 172.790 ;
        RECT 208.025 171.280 280.555 173.280 ;
        RECT 282.935 172.575 300.445 188.625 ;
        RECT 183.180 170.075 187.550 170.405 ;
        RECT 183.180 169.275 183.780 170.075 ;
        RECT 185.885 170.070 187.545 170.075 ;
        RECT 189.695 166.235 233.005 166.565 ;
        RECT 189.695 165.605 233.005 165.935 ;
        RECT 208.025 158.920 280.555 160.920 ;
        RECT 282.935 155.325 300.445 171.375 ;
        RECT 171.460 154.920 279.920 155.250 ;
        RECT 279.590 154.125 279.920 154.920 ;
        RECT 279.590 153.795 433.610 154.125 ;
        RECT 280.385 153.165 432.480 153.495 ;
        RECT 281.935 152.265 297.675 152.865 ;
        RECT 432.150 152.365 432.480 153.165 ;
        RECT 433.280 152.995 433.610 153.795 ;
        RECT 178.380 151.400 178.980 151.930 ;
        RECT 297.075 151.735 297.675 152.265 ;
        RECT 46.010 150.800 178.980 151.400 ;
        RECT 184.765 144.775 294.445 146.775 ;
        RECT 300.300 144.775 409.980 146.775 ;
        RECT 183.180 141.465 183.780 141.530 ;
        RECT 297.075 141.465 297.675 141.595 ;
        RECT 410.505 141.465 411.105 141.470 ;
        RECT 183.180 140.465 191.020 141.465 ;
        RECT 288.195 140.465 306.555 141.465 ;
        RECT 403.730 140.465 411.105 141.465 ;
        RECT 183.180 140.400 183.780 140.465 ;
        RECT 410.505 140.340 411.105 140.465 ;
        RECT 299.055 138.360 411.130 138.960 ;
        RECT 184.765 130.610 294.445 132.610 ;
        RECT 300.300 130.610 409.980 132.610 ;
        RECT 299.055 127.300 299.655 127.365 ;
        RECT 184.930 126.965 191.020 127.300 ;
        RECT 178.880 126.635 191.020 126.965 ;
        RECT 178.880 125.835 179.480 126.635 ;
        RECT 184.930 126.300 191.020 126.635 ;
        RECT 288.195 126.300 295.975 127.300 ;
        RECT 295.375 126.170 295.975 126.300 ;
        RECT 299.055 126.300 306.555 127.300 ;
        RECT 403.730 126.300 411.370 127.300 ;
        RECT 299.055 126.235 299.655 126.300 ;
        RECT 410.770 126.170 411.370 126.300 ;
        RECT 175.680 124.385 176.280 124.650 ;
        RECT 175.680 123.785 411.395 124.385 ;
        RECT 175.680 123.520 176.280 123.785 ;
        RECT 431.020 122.675 431.350 123.475 ;
        RECT 406.455 122.345 431.350 122.675 ;
        RECT 183.180 121.545 183.780 122.075 ;
        RECT 351.305 121.695 418.775 122.045 ;
        RECT 183.180 120.945 296.000 121.545 ;
        RECT 405.820 120.945 430.220 121.275 ;
        RECT 405.820 120.155 406.150 120.945 ;
        RECT 311.000 119.825 406.150 120.155 ;
        RECT 429.890 120.145 430.220 120.945 ;
        RECT 310.835 118.005 406.665 119.005 ;
        RECT 368.445 116.875 369.175 117.205 ;
        RECT 214.090 115.305 223.340 116.305 ;
        RECT 340.945 115.975 341.275 116.205 ;
        RECT 342.705 115.975 343.035 116.205 ;
        RECT 344.465 115.975 344.795 116.205 ;
        RECT 346.225 115.975 346.555 116.205 ;
        RECT 340.945 115.475 346.555 115.975 ;
        RECT 351.505 115.975 351.835 116.205 ;
        RECT 353.265 115.975 353.595 116.205 ;
        RECT 355.025 115.975 355.355 116.205 ;
        RECT 356.785 115.975 357.115 116.205 ;
        RECT 351.505 115.475 357.115 115.975 ;
        RECT 214.090 115.175 214.420 115.305 ;
        RECT 368.560 115.050 369.060 116.875 ;
        RECT 184.620 113.585 290.545 114.585 ;
        RECT 340.065 114.550 347.435 115.050 ;
        RECT 340.065 114.320 340.395 114.550 ;
        RECT 341.825 114.320 342.155 114.550 ;
        RECT 343.585 114.320 343.915 114.550 ;
        RECT 345.345 114.320 345.675 114.550 ;
        RECT 347.105 114.320 347.435 114.550 ;
        RECT 350.625 114.550 369.060 115.050 ;
        RECT 350.625 114.320 350.955 114.550 ;
        RECT 352.385 114.320 352.715 114.550 ;
        RECT 354.145 114.320 354.475 114.550 ;
        RECT 355.905 114.320 356.235 114.550 ;
        RECT 357.665 114.320 357.995 114.550 ;
        RECT 311.085 113.340 407.185 113.670 ;
        RECT 181.080 112.535 181.680 113.335 ;
        RECT 181.080 112.205 186.430 112.535 ;
        RECT 184.720 110.160 198.430 111.160 ;
        RECT 198.760 111.030 199.090 111.830 ;
        RECT 199.800 111.345 213.510 112.195 ;
        RECT 310.835 111.520 406.665 112.520 ;
        RECT 198.760 110.700 200.995 111.030 ;
        RECT 201.330 110.190 201.660 110.590 ;
        RECT 202.205 110.190 202.535 110.610 ;
        RECT 203.065 110.190 203.395 110.610 ;
        RECT 203.925 110.190 204.255 110.610 ;
        RECT 204.785 110.190 205.115 110.590 ;
        RECT 205.645 110.190 205.975 110.590 ;
        RECT 206.505 110.190 206.835 110.590 ;
        RECT 207.365 110.190 207.695 110.590 ;
        RECT 208.225 110.190 208.555 110.590 ;
        RECT 209.085 110.190 209.415 110.610 ;
        RECT 209.945 110.190 210.275 110.610 ;
        RECT 210.805 110.190 211.135 110.610 ;
        RECT 211.665 110.190 211.995 110.610 ;
        RECT 199.965 109.860 215.880 110.190 ;
        RECT 184.720 108.130 198.430 109.130 ;
        RECT 199.965 109.125 215.150 109.455 ;
        RECT 201.760 108.725 202.090 109.125 ;
        RECT 202.635 108.725 202.965 109.125 ;
        RECT 203.495 108.725 203.825 109.125 ;
        RECT 204.355 108.725 204.685 109.125 ;
        RECT 205.215 108.725 205.545 109.125 ;
        RECT 206.075 108.725 206.405 109.125 ;
        RECT 206.935 108.725 207.265 109.125 ;
        RECT 207.795 108.725 208.125 109.125 ;
        RECT 208.655 108.725 208.985 109.125 ;
        RECT 209.515 108.725 209.845 109.125 ;
        RECT 210.375 108.725 210.705 109.125 ;
        RECT 211.235 108.725 211.565 109.125 ;
        RECT 198.760 108.260 200.995 108.590 ;
        RECT 214.820 108.305 215.150 109.125 ;
        RECT 215.550 109.040 215.880 109.860 ;
        RECT 198.760 107.460 199.090 108.260 ;
        RECT 217.090 108.145 290.590 110.145 ;
        RECT 405.960 108.960 406.765 109.760 ;
        RECT 311.000 108.105 407.185 108.435 ;
        RECT 199.800 107.095 213.510 107.945 ;
        RECT 214.820 106.710 215.150 106.840 ;
        RECT 214.820 105.710 243.440 106.710 ;
        RECT 184.720 104.705 213.245 105.705 ;
        RECT 299.055 105.635 311.330 105.660 ;
        RECT 299.055 105.330 313.620 105.635 ;
        RECT 311.000 105.305 313.620 105.330 ;
        RECT 311.955 105.300 313.615 105.305 ;
        RECT 175.680 103.805 176.280 104.135 ;
        RECT 112.260 103.005 176.280 103.805 ;
        RECT 176.780 103.710 177.380 104.240 ;
        RECT 178.880 103.710 179.480 104.175 ;
        RECT 176.780 103.110 179.480 103.710 ;
        RECT 178.880 102.645 179.480 103.110 ;
        RECT 184.620 102.895 290.545 103.895 ;
        RECT 310.835 102.910 333.745 103.910 ;
        RECT 334.095 102.400 406.625 104.400 ;
        RECT 409.005 103.695 426.515 119.745 ;
        RECT 446.785 118.245 492.950 118.575 ;
        RECT 434.770 113.055 505.570 115.055 ;
        RECT 433.280 107.705 433.610 108.105 ;
        RECT 433.280 107.375 505.190 107.705 ;
        RECT 433.280 106.975 433.610 107.375 ;
        RECT 432.150 105.310 432.480 105.710 ;
        RECT 432.150 104.980 505.190 105.310 ;
        RECT 432.150 104.580 432.480 104.980 ;
        RECT 184.720 101.085 213.245 102.085 ;
        RECT 311.000 101.480 313.620 101.525 ;
        RECT 215.550 101.085 215.880 101.215 ;
        RECT 299.055 101.195 313.620 101.480 ;
        RECT 299.055 101.150 311.330 101.195 ;
        RECT 311.955 101.190 313.615 101.195 ;
        RECT 215.550 100.085 243.440 101.085 ;
        RECT 184.720 97.660 198.430 98.660 ;
        RECT 198.760 98.530 199.090 99.330 ;
        RECT 199.800 98.845 213.510 99.695 ;
        RECT 198.760 98.200 200.995 98.530 ;
        RECT 201.760 97.665 202.090 98.065 ;
        RECT 202.635 97.665 202.965 98.065 ;
        RECT 203.495 97.665 203.825 98.065 ;
        RECT 204.355 97.665 204.685 98.065 ;
        RECT 205.215 97.665 205.545 98.065 ;
        RECT 206.075 97.665 206.405 98.065 ;
        RECT 206.935 97.665 207.265 98.065 ;
        RECT 207.795 97.665 208.125 98.065 ;
        RECT 208.655 97.665 208.985 98.065 ;
        RECT 209.515 97.665 209.845 98.065 ;
        RECT 210.375 97.665 210.705 98.065 ;
        RECT 211.235 97.665 211.565 98.065 ;
        RECT 214.090 97.665 214.420 98.485 ;
        RECT 199.965 97.335 214.420 97.665 ;
        RECT 184.720 95.630 198.430 96.630 ;
        RECT 199.965 96.600 214.420 96.930 ;
        RECT 217.090 96.645 290.590 98.645 ;
        RECT 315.765 97.355 359.075 97.685 ;
        RECT 315.765 96.725 359.075 97.055 ;
        RECT 201.330 96.200 201.660 96.600 ;
        RECT 202.205 96.180 202.535 96.600 ;
        RECT 203.065 96.180 203.395 96.600 ;
        RECT 203.925 96.180 204.255 96.600 ;
        RECT 204.785 96.200 205.115 96.600 ;
        RECT 205.645 96.200 205.975 96.600 ;
        RECT 206.505 96.200 206.835 96.600 ;
        RECT 207.365 96.200 207.695 96.600 ;
        RECT 208.225 96.200 208.555 96.600 ;
        RECT 209.085 96.180 209.415 96.600 ;
        RECT 209.945 96.180 210.275 96.600 ;
        RECT 210.805 96.180 211.135 96.600 ;
        RECT 211.665 96.180 211.995 96.600 ;
        RECT 198.760 95.760 200.995 96.090 ;
        RECT 214.090 95.780 214.420 96.600 ;
        RECT 179.980 94.585 180.580 95.385 ;
        RECT 198.760 94.960 199.090 95.760 ;
        RECT 199.800 94.595 213.510 95.445 ;
        RECT 179.980 94.255 186.430 94.585 ;
        RECT 184.620 92.205 290.545 93.205 ;
        RECT 214.090 91.490 214.420 91.620 ;
        RECT 214.090 90.490 223.340 91.490 ;
        RECT 334.095 90.040 406.625 92.040 ;
        RECT 409.005 86.445 426.515 102.495 ;
        RECT 486.930 99.275 503.815 101.275 ;
        RECT 472.330 94.465 505.570 95.965 ;
        RECT 431.020 93.895 431.350 94.295 ;
        RECT 431.020 93.565 505.270 93.895 ;
        RECT 431.020 93.165 431.350 93.565 ;
        RECT 429.890 91.225 430.220 91.625 ;
        RECT 453.250 91.565 471.085 93.065 ;
        RECT 429.890 90.895 505.270 91.225 ;
        RECT 429.890 90.495 430.220 90.895 ;
        RECT 434.770 88.950 505.570 90.450 ;
        RECT 434.980 88.185 505.270 88.515 ;
        RECT 311.000 86.040 405.990 86.370 ;
        RECT 183.180 85.245 296.000 85.845 ;
        RECT 405.660 85.245 405.990 86.040 ;
        RECT 433.280 85.245 433.610 85.645 ;
        RECT 183.180 84.715 183.780 85.245 ;
        RECT 405.660 84.915 433.610 85.245 ;
        RECT 406.455 84.285 432.480 84.615 ;
        RECT 433.280 84.515 433.610 84.915 ;
        RECT 432.150 83.485 432.480 84.285 ;
        RECT 442.430 81.060 443.740 88.185 ;
        RECT 178.880 80.155 179.480 80.955 ;
        RECT 295.375 80.490 295.975 80.620 ;
        RECT 184.930 80.155 191.020 80.490 ;
        RECT 178.880 79.825 191.020 80.155 ;
        RECT 184.930 79.490 191.020 79.825 ;
        RECT 288.195 79.490 295.975 80.490 ;
        RECT 299.055 80.490 299.655 80.555 ;
        RECT 299.055 79.490 306.555 80.490 ;
        RECT 403.730 79.490 409.815 80.490 ;
        RECT 299.055 79.425 299.655 79.490 ;
        RECT 184.765 74.180 294.445 76.180 ;
        RECT 300.300 74.180 419.895 76.180 ;
        RECT 437.490 73.900 502.950 75.900 ;
        RECT 496.700 71.465 498.010 72.465 ;
        RECT 299.055 67.830 411.130 68.430 ;
        RECT 183.180 66.345 183.780 66.410 ;
        RECT 410.505 66.345 411.105 66.475 ;
        RECT 183.180 65.345 191.020 66.345 ;
        RECT 288.195 65.345 306.555 66.345 ;
        RECT 403.730 65.345 411.105 66.345 ;
        RECT 183.180 65.280 183.780 65.345 ;
        RECT 297.075 65.215 297.675 65.345 ;
        RECT 184.765 60.035 294.445 62.035 ;
        RECT 300.300 60.035 419.895 62.035 ;
        RECT 46.160 55.410 178.980 56.010 ;
        RECT 178.380 54.880 178.980 55.410 ;
        RECT 297.075 54.545 297.675 55.075 ;
        RECT 281.935 53.945 297.675 54.545 ;
        RECT 328.700 53.945 428.020 54.275 ;
        RECT 432.150 53.645 432.480 54.445 ;
        RECT 280.385 53.315 432.480 53.645 ;
        RECT 279.590 52.685 331.645 53.015 ;
        RECT 279.590 51.890 279.920 52.685 ;
        RECT 184.930 51.560 279.920 51.890 ;
        RECT 331.315 51.890 331.645 52.685 ;
        RECT 433.280 51.890 433.610 52.690 ;
        RECT 331.315 51.560 433.610 51.890 ;
        RECT 208.025 45.890 280.555 47.890 ;
        RECT 189.695 40.875 233.005 41.205 ;
        RECT 189.695 40.245 233.005 40.575 ;
        RECT 183.180 36.715 183.780 37.515 ;
        RECT 185.885 36.735 187.545 36.740 ;
        RECT 184.930 36.715 187.550 36.735 ;
        RECT 183.180 36.405 187.550 36.715 ;
        RECT 183.180 36.385 185.260 36.405 ;
        RECT 184.765 34.020 207.675 35.020 ;
        RECT 208.025 33.530 280.555 35.530 ;
        RECT 282.935 35.435 300.445 51.485 ;
        RECT 310.790 35.435 328.300 51.485 ;
        RECT 330.680 45.890 403.210 47.890 ;
        RECT 378.230 40.875 421.540 41.205 ;
        RECT 378.230 40.245 421.540 40.575 ;
        RECT 423.690 36.735 425.350 36.740 ;
        RECT 427.395 36.735 427.995 37.535 ;
        RECT 423.685 36.405 427.995 36.735 ;
        RECT 178.380 32.625 178.980 33.425 ;
        RECT 185.885 32.625 187.545 32.630 ;
        RECT 178.380 32.295 187.550 32.625 ;
        RECT 184.930 29.495 281.115 29.825 ;
        RECT 279.890 28.170 280.695 28.970 ;
        RECT 184.765 25.410 280.595 26.410 ;
        RECT 185.015 24.260 281.115 24.590 ;
        RECT 213.995 23.380 214.325 23.610 ;
        RECT 215.755 23.380 216.085 23.610 ;
        RECT 217.515 23.380 217.845 23.610 ;
        RECT 219.275 23.380 219.605 23.610 ;
        RECT 221.035 23.380 221.365 23.610 ;
        RECT 213.995 22.880 221.365 23.380 ;
        RECT 224.555 23.380 224.885 23.610 ;
        RECT 226.315 23.380 226.645 23.610 ;
        RECT 228.075 23.380 228.405 23.610 ;
        RECT 229.835 23.380 230.165 23.610 ;
        RECT 231.595 23.380 231.925 23.610 ;
        RECT 224.555 22.880 242.990 23.380 ;
        RECT 214.875 21.955 220.485 22.455 ;
        RECT 214.875 21.725 215.205 21.955 ;
        RECT 216.635 21.725 216.965 21.955 ;
        RECT 218.395 21.725 218.725 21.955 ;
        RECT 220.155 21.725 220.485 21.955 ;
        RECT 225.435 21.955 231.045 22.455 ;
        RECT 225.435 21.725 225.765 21.955 ;
        RECT 227.195 21.725 227.525 21.955 ;
        RECT 228.955 21.725 229.285 21.955 ;
        RECT 230.715 21.725 231.045 21.955 ;
        RECT 242.490 21.055 242.990 22.880 ;
        RECT 242.375 20.725 243.105 21.055 ;
        RECT 184.765 18.925 280.595 19.925 ;
        RECT 282.935 18.185 300.445 34.235 ;
        RECT 310.790 18.185 328.300 34.235 ;
        RECT 330.680 33.530 403.210 35.530 ;
        RECT 403.560 34.020 426.470 35.020 ;
        RECT 423.690 32.625 425.350 32.630 ;
        RECT 428.680 32.625 429.280 33.425 ;
        RECT 423.685 32.295 429.280 32.625 ;
        RECT 330.120 29.495 426.305 29.825 ;
        RECT 330.540 28.170 331.345 28.970 ;
        RECT 330.640 25.410 426.470 26.410 ;
        RECT 330.120 24.260 426.220 24.590 ;
        RECT 379.310 23.380 379.640 23.610 ;
        RECT 381.070 23.380 381.400 23.610 ;
        RECT 382.830 23.380 383.160 23.610 ;
        RECT 384.590 23.380 384.920 23.610 ;
        RECT 386.350 23.380 386.680 23.610 ;
        RECT 368.245 22.880 386.680 23.380 ;
        RECT 389.870 23.380 390.200 23.610 ;
        RECT 391.630 23.380 391.960 23.610 ;
        RECT 393.390 23.380 393.720 23.610 ;
        RECT 395.150 23.380 395.480 23.610 ;
        RECT 396.910 23.380 397.240 23.610 ;
        RECT 389.870 22.880 397.240 23.380 ;
        RECT 368.245 21.055 368.745 22.880 ;
        RECT 380.190 21.955 385.800 22.455 ;
        RECT 380.190 21.725 380.520 21.955 ;
        RECT 381.950 21.725 382.280 21.955 ;
        RECT 383.710 21.725 384.040 21.955 ;
        RECT 385.470 21.725 385.800 21.955 ;
        RECT 390.750 21.955 396.360 22.455 ;
        RECT 390.750 21.725 391.080 21.955 ;
        RECT 392.510 21.725 392.840 21.955 ;
        RECT 394.270 21.725 394.600 21.955 ;
        RECT 396.030 21.725 396.360 21.955 ;
        RECT 368.130 20.725 368.860 21.055 ;
        RECT 330.640 18.925 426.470 19.925 ;
        RECT 429.890 18.105 430.220 18.905 ;
        RECT 184.930 17.775 280.080 18.105 ;
        RECT 279.750 16.985 280.080 17.775 ;
        RECT 331.155 17.775 430.220 18.105 ;
        RECT 331.155 16.985 331.485 17.775 ;
        RECT 279.750 16.655 331.485 16.985 ;
        RECT 225.235 15.885 292.705 16.235 ;
        RECT 318.530 15.885 386.000 16.235 ;
        RECT 280.385 15.255 431.350 15.585 ;
        RECT 1.000 10.570 503.815 13.570 ;
        RECT 176.780 8.725 177.380 9.255 ;
        RECT 134.330 8.125 177.380 8.725 ;
        RECT 156.410 6.525 329.300 7.125 ;
        RECT 46.010 0.890 46.910 2.325 ;
        RECT 68.090 0.890 68.990 2.325 ;
      LAYER met4 ;
        RECT 3.990 220.760 4.290 224.760 ;
        RECT 7.670 220.760 7.970 224.760 ;
        RECT 11.350 220.760 11.650 224.760 ;
        RECT 15.030 220.760 15.330 224.760 ;
        RECT 18.710 220.760 19.010 224.760 ;
        RECT 22.390 220.760 22.690 224.760 ;
        RECT 26.070 220.760 26.370 224.760 ;
        RECT 29.750 220.760 30.050 224.760 ;
        RECT 33.430 220.760 33.730 224.760 ;
        RECT 37.110 220.760 37.410 224.760 ;
        RECT 40.790 220.760 41.090 224.760 ;
        RECT 44.470 220.760 44.770 224.760 ;
        RECT 48.150 220.760 48.450 224.760 ;
        RECT 51.830 220.760 52.130 224.760 ;
        RECT 55.510 220.760 55.810 224.760 ;
        RECT 59.190 220.760 59.490 224.760 ;
        RECT 62.870 220.760 63.170 224.760 ;
        RECT 66.550 220.760 66.850 224.760 ;
        RECT 70.230 220.760 70.530 224.760 ;
        RECT 73.910 220.760 74.210 224.760 ;
        RECT 77.590 220.760 77.890 224.760 ;
        RECT 81.270 220.760 81.570 224.760 ;
        RECT 84.950 220.760 85.250 224.760 ;
        RECT 88.630 220.760 88.930 224.760 ;
        RECT 3.975 219.260 4.305 220.760 ;
        RECT 7.655 219.260 7.985 220.760 ;
        RECT 11.335 219.260 11.665 220.760 ;
        RECT 15.015 219.260 15.345 220.760 ;
        RECT 18.695 219.260 19.025 220.760 ;
        RECT 22.375 219.260 22.705 220.760 ;
        RECT 26.055 219.260 26.385 220.760 ;
        RECT 29.735 219.260 30.065 220.760 ;
        RECT 33.415 219.260 33.745 220.760 ;
        RECT 37.095 219.260 37.425 220.760 ;
        RECT 40.775 219.260 41.105 220.760 ;
        RECT 44.455 219.260 44.785 220.760 ;
        RECT 48.135 219.260 48.465 220.760 ;
        RECT 51.815 219.260 52.145 220.760 ;
        RECT 55.495 219.260 55.825 220.760 ;
        RECT 59.175 219.260 59.505 220.760 ;
        RECT 62.855 219.260 63.185 220.760 ;
        RECT 66.535 219.260 66.865 220.760 ;
        RECT 70.215 219.260 70.545 220.760 ;
        RECT 73.895 219.260 74.225 220.760 ;
        RECT 77.575 219.260 77.905 220.760 ;
        RECT 81.255 219.260 81.585 220.760 ;
        RECT 84.935 219.260 85.265 220.760 ;
        RECT 88.615 219.260 88.945 220.760 ;
        RECT 143.830 216.045 144.130 224.760 ;
        RECT 147.510 217.670 147.810 224.760 ;
        RECT 147.495 216.490 147.825 217.670 ;
        RECT 143.815 214.865 144.145 216.045 ;
        RECT 62.255 208.285 62.775 208.635 ;
        RECT 54.885 193.025 70.145 208.285 ;
        RECT 62.430 191.035 62.950 193.025 ;
        RECT 54.885 175.775 70.145 191.035 ;
        RECT 71.480 186.165 72.000 208.680 ;
        RECT 71.480 185.365 75.045 186.165 ;
        RECT 62.255 173.430 62.775 175.775 ;
        RECT 71.480 175.380 72.000 185.365 ;
        RECT 82.595 174.320 84.095 209.775 ;
        RECT 109.095 174.320 110.595 214.340 ;
        RECT 135.595 174.320 137.095 209.775 ;
        RECT 139.095 190.725 157.470 192.725 ;
        RECT 62.255 173.080 62.985 173.430 ;
        RECT 89.140 171.550 91.070 172.150 ;
        RECT 46.010 1.000 46.910 2.325 ;
        RECT 68.090 1.000 68.990 2.325 ;
        RECT 90.170 1.000 91.070 171.550 ;
        RECT 112.255 103.005 113.785 103.805 ;
        RECT 112.255 1.000 113.155 103.005 ;
        RECT 155.470 10.570 157.470 190.725 ;
        RECT 162.095 174.320 163.595 214.340 ;
        RECT 185.245 91.395 186.245 214.340 ;
        RECT 191.340 14.970 192.840 214.340 ;
        RECT 194.245 10.570 195.245 115.395 ;
        RECT 203.245 91.395 204.245 214.340 ;
        RECT 212.245 10.570 213.245 115.395 ;
        RECT 217.840 10.570 219.340 205.085 ;
        RECT 221.245 91.395 222.245 214.340 ;
        RECT 230.245 10.570 231.245 115.395 ;
        RECT 239.245 91.395 240.245 214.340 ;
        RECT 244.340 14.970 245.840 214.340 ;
        RECT 248.245 10.570 249.245 115.395 ;
        RECT 257.245 91.395 258.245 214.340 ;
        RECT 266.245 10.570 267.245 115.395 ;
        RECT 270.840 10.570 272.340 205.085 ;
        RECT 275.245 91.395 276.245 214.340 ;
        RECT 291.950 190.575 292.680 190.925 ;
        RECT 282.935 178.640 283.455 188.625 ;
        RECT 292.160 188.230 292.680 190.575 ;
        RECT 279.890 177.840 283.455 178.640 ;
        RECT 282.935 155.325 283.455 177.840 ;
        RECT 284.790 172.970 300.050 188.230 ;
        RECT 291.985 170.980 292.505 172.970 ;
        RECT 284.790 155.720 300.050 170.980 ;
        RECT 292.160 155.370 292.680 155.720 ;
        RECT 284.245 91.395 285.245 115.395 ;
        RECT 317.410 60.035 318.910 214.340 ;
        RECT 282.935 28.970 283.455 51.485 ;
        RECT 292.160 51.090 292.680 51.440 ;
        RECT 318.555 51.090 319.075 51.440 ;
        RECT 284.790 35.830 300.050 51.090 ;
        RECT 311.185 35.830 326.445 51.090 ;
        RECT 291.985 33.840 292.505 35.830 ;
        RECT 318.730 33.840 319.250 35.830 ;
        RECT 279.890 28.170 283.455 28.970 ;
        RECT 282.935 18.185 283.455 28.170 ;
        RECT 284.790 18.580 300.050 33.840 ;
        RECT 311.185 18.580 326.445 33.840 ;
        RECT 327.780 28.970 328.300 51.485 ;
        RECT 327.780 28.170 331.345 28.970 ;
        RECT 292.160 16.235 292.680 18.580 ;
        RECT 291.950 15.885 292.680 16.235 ;
        RECT 318.555 16.235 319.075 18.580 ;
        RECT 327.780 18.185 328.300 28.170 ;
        RECT 318.555 15.885 319.285 16.235 ;
        RECT 338.895 10.570 340.395 52.580 ;
        RECT 343.910 10.570 345.410 120.805 ;
        RECT 365.395 14.970 366.895 76.180 ;
        RECT 370.410 60.035 371.910 214.340 ;
        RECT 418.020 121.695 418.750 122.045 ;
        RECT 391.895 10.570 393.395 52.580 ;
        RECT 396.910 10.570 398.410 120.805 ;
        RECT 409.005 109.760 409.525 119.745 ;
        RECT 418.230 119.350 418.750 121.695 ;
        RECT 405.960 108.960 409.525 109.760 ;
        RECT 409.005 86.445 409.525 108.960 ;
        RECT 410.860 104.090 426.120 119.350 ;
        RECT 418.055 102.100 418.575 104.090 ;
        RECT 410.860 86.840 426.120 102.100 ;
        RECT 435.815 87.610 437.815 214.340 ;
        RECT 418.230 86.490 418.750 86.840 ;
        RECT 418.395 14.970 419.895 76.180 ;
        RECT 457.815 10.570 459.815 119.205 ;
        RECT 479.815 73.900 481.815 214.340 ;
        RECT 501.815 72.465 503.815 119.205 ;
        RECT 496.700 71.465 503.815 72.465 ;
        RECT 501.815 10.570 503.815 71.465 ;
        RECT 134.330 8.125 135.460 8.725 ;
        RECT 134.330 1.000 135.230 8.125 ;
        RECT 156.410 6.525 157.540 7.125 ;
        RECT 156.410 1.000 157.310 6.525 ;
        RECT 113.150 0.135 113.155 1.000 ;
  END
END tt_um_CktA_InstAmp
END LIBRARY

