VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_KolosKoblasz_mixer
  CLASS BLOCK ;
  FOREIGN tt_um_KolosKoblasz_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.736000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.736000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.088000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.088000 ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1223.933350 ;
    ANTENNADIFFAREA 164.215347 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 57.000 202.085 131.440 203.690 ;
      LAYER pwell ;
        RECT 57.195 200.885 58.565 201.695 ;
        RECT 58.575 200.885 60.405 201.695 ;
        RECT 60.875 200.885 62.245 201.665 ;
        RECT 62.255 200.885 67.765 201.695 ;
        RECT 67.775 200.885 69.605 201.695 ;
        RECT 70.085 200.970 70.515 201.755 ;
        RECT 70.535 200.885 72.365 201.565 ;
        RECT 72.375 200.885 75.125 201.695 ;
        RECT 75.195 200.885 76.965 201.795 ;
        RECT 76.975 200.885 79.725 201.695 ;
        RECT 80.195 200.885 81.565 201.665 ;
        RECT 81.575 200.885 82.945 201.695 ;
        RECT 82.965 200.970 83.395 201.755 ;
        RECT 83.415 200.885 85.245 201.695 ;
        RECT 85.265 200.885 86.615 201.795 ;
        RECT 86.730 201.565 87.650 201.795 ;
        RECT 86.730 200.885 90.195 201.565 ;
        RECT 90.315 200.885 91.685 201.665 ;
        RECT 91.695 200.885 95.365 201.695 ;
        RECT 95.845 200.970 96.275 201.755 ;
        RECT 97.215 200.885 98.585 201.665 ;
        RECT 99.080 201.595 100.435 201.795 ;
        RECT 99.080 201.565 101.760 201.595 ;
        RECT 105.390 201.565 106.310 201.795 ;
        RECT 98.595 200.915 101.760 201.565 ;
        RECT 98.595 200.885 100.435 200.915 ;
        RECT 102.845 200.885 106.310 201.565 ;
        RECT 106.415 200.885 108.245 201.695 ;
        RECT 108.725 200.970 109.155 201.755 ;
        RECT 109.835 201.565 113.765 201.795 ;
        RECT 109.350 200.885 113.765 201.565 ;
        RECT 115.155 200.885 118.825 201.695 ;
        RECT 118.835 200.885 120.205 201.665 ;
        RECT 120.215 200.885 121.585 201.695 ;
        RECT 121.605 200.970 122.035 201.755 ;
        RECT 122.055 200.885 127.565 201.695 ;
        RECT 127.575 200.885 129.405 201.695 ;
        RECT 129.875 200.885 131.245 201.695 ;
        RECT 57.335 200.675 57.505 200.885 ;
        RECT 58.715 200.675 58.885 200.885 ;
        RECT 60.550 200.725 60.670 200.835 ;
        RECT 61.025 200.695 61.195 200.885 ;
        RECT 62.395 200.695 62.565 200.885 ;
        RECT 64.235 200.675 64.405 200.865 ;
        RECT 67.915 200.695 68.085 200.885 ;
        RECT 69.755 200.835 69.925 200.865 ;
        RECT 69.750 200.725 69.925 200.835 ;
        RECT 69.755 200.675 69.925 200.725 ;
        RECT 70.675 200.695 70.845 200.885 ;
        RECT 71.590 200.725 71.710 200.835 ;
        RECT 72.055 200.675 72.225 200.865 ;
        RECT 72.515 200.695 72.685 200.885 ;
        RECT 76.650 200.695 76.820 200.885 ;
        RECT 77.115 200.695 77.285 200.885 ;
        RECT 78.500 200.695 78.670 200.865 ;
        RECT 79.875 200.835 80.045 200.865 ;
        RECT 78.965 200.720 79.125 200.830 ;
        RECT 79.870 200.725 80.045 200.835 ;
        RECT 78.500 200.675 78.635 200.695 ;
        RECT 79.875 200.675 80.045 200.725 ;
        RECT 80.345 200.695 80.515 200.885 ;
        RECT 81.715 200.695 81.885 200.885 ;
        RECT 83.555 200.695 83.725 200.885 ;
        RECT 84.930 200.675 85.100 200.865 ;
        RECT 85.390 200.725 85.510 200.835 ;
        RECT 86.315 200.695 86.485 200.885 ;
        RECT 89.995 200.695 90.165 200.885 ;
        RECT 90.455 200.695 90.625 200.885 ;
        RECT 91.835 200.695 92.005 200.885 ;
        RECT 92.755 200.675 92.925 200.865 ;
        RECT 93.215 200.675 93.385 200.865 ;
        RECT 95.510 200.725 95.630 200.835 ;
        RECT 96.445 200.730 96.605 200.840 ;
        RECT 97.355 200.695 97.525 200.885 ;
        RECT 98.735 200.695 98.905 200.885 ;
        RECT 101.965 200.730 102.125 200.840 ;
        RECT 102.875 200.695 103.045 200.885 ;
        RECT 103.980 200.675 104.150 200.865 ;
        RECT 105.635 200.675 105.805 200.865 ;
        RECT 106.095 200.675 106.265 200.865 ;
        RECT 106.555 200.695 106.725 200.885 ;
        RECT 109.350 200.865 109.460 200.885 ;
        RECT 108.390 200.725 108.510 200.835 ;
        RECT 109.290 200.695 109.485 200.865 ;
        RECT 111.150 200.725 111.270 200.835 ;
        RECT 109.315 200.675 109.485 200.695 ;
        RECT 111.615 200.675 111.785 200.865 ;
        RECT 113.915 200.695 114.085 200.865 ;
        RECT 115.295 200.695 115.465 200.885 ;
        RECT 118.975 200.695 119.145 200.885 ;
        RECT 120.355 200.695 120.525 200.885 ;
        RECT 122.195 200.695 122.365 200.885 ;
        RECT 124.035 200.675 124.205 200.865 ;
        RECT 124.495 200.675 124.665 200.865 ;
        RECT 125.875 200.675 126.045 200.865 ;
        RECT 127.715 200.695 127.885 200.885 ;
        RECT 129.550 200.725 129.670 200.835 ;
        RECT 130.935 200.675 131.105 200.885 ;
        RECT 57.195 199.865 58.565 200.675 ;
        RECT 58.575 199.865 64.085 200.675 ;
        RECT 64.095 199.865 69.605 200.675 ;
        RECT 69.615 199.865 71.445 200.675 ;
        RECT 71.955 199.765 75.125 200.675 ;
        RECT 75.135 199.765 78.635 200.675 ;
        RECT 79.735 199.765 82.945 200.675 ;
        RECT 82.965 199.805 83.395 200.590 ;
        RECT 83.415 199.765 85.245 200.675 ;
        RECT 85.755 199.995 93.065 200.675 ;
        RECT 93.075 199.995 100.385 200.675 ;
        RECT 100.665 199.995 104.565 200.675 ;
        RECT 85.755 199.765 87.105 199.995 ;
        RECT 88.640 199.775 89.550 199.995 ;
        RECT 96.590 199.775 97.500 199.995 ;
        RECT 99.035 199.765 100.385 199.995 ;
        RECT 103.635 199.765 104.565 199.995 ;
        RECT 104.585 199.765 105.935 200.675 ;
        RECT 105.955 199.865 108.705 200.675 ;
        RECT 108.725 199.805 109.155 200.590 ;
        RECT 109.175 199.865 111.005 200.675 ;
        RECT 111.475 199.995 120.665 200.675 ;
        RECT 115.985 199.775 116.915 199.995 ;
        RECT 119.745 199.765 120.665 199.995 ;
        RECT 120.770 199.995 124.235 200.675 ;
        RECT 120.770 199.765 121.690 199.995 ;
        RECT 124.365 199.765 125.715 200.675 ;
        RECT 125.735 199.865 129.405 200.675 ;
        RECT 129.875 199.865 131.245 200.675 ;
      LAYER nwell ;
        RECT 57.000 196.645 131.440 199.475 ;
      LAYER pwell ;
        RECT 57.195 195.445 58.565 196.255 ;
        RECT 58.575 195.445 64.085 196.255 ;
        RECT 64.095 195.445 69.605 196.255 ;
        RECT 70.085 195.530 70.515 196.315 ;
        RECT 70.535 195.445 74.205 196.255 ;
        RECT 74.215 195.445 75.585 196.255 ;
        RECT 75.595 195.445 78.345 196.355 ;
        RECT 78.355 195.445 82.025 196.255 ;
        RECT 82.495 196.125 83.420 196.355 ;
        RECT 82.495 195.445 86.165 196.125 ;
        RECT 87.095 195.445 88.910 196.355 ;
        RECT 92.050 196.125 92.970 196.355 ;
        RECT 89.505 195.445 92.970 196.125 ;
        RECT 93.095 195.445 94.445 196.355 ;
        RECT 94.455 195.445 95.825 196.255 ;
        RECT 95.845 195.530 96.275 196.315 ;
        RECT 96.375 195.445 99.825 196.355 ;
        RECT 99.975 195.445 103.185 196.355 ;
        RECT 103.195 195.445 104.565 196.255 ;
        RECT 113.775 196.125 114.705 196.355 ;
        RECT 119.720 196.155 120.665 196.355 ;
        RECT 104.660 195.445 113.765 196.125 ;
        RECT 113.775 195.445 117.675 196.125 ;
        RECT 117.915 195.475 120.665 196.155 ;
        RECT 121.605 195.530 122.035 196.315 ;
        RECT 57.335 195.235 57.505 195.445 ;
        RECT 58.715 195.235 58.885 195.445 ;
        RECT 64.235 195.235 64.405 195.445 ;
        RECT 69.755 195.395 69.925 195.425 ;
        RECT 69.750 195.285 69.925 195.395 ;
        RECT 69.755 195.235 69.925 195.285 ;
        RECT 70.675 195.255 70.845 195.445 ;
        RECT 74.355 195.255 74.525 195.445 ;
        RECT 75.275 195.235 75.445 195.425 ;
        RECT 78.035 195.255 78.205 195.445 ;
        RECT 78.310 195.235 78.480 195.425 ;
        RECT 78.495 195.255 78.665 195.445 ;
        RECT 82.170 195.390 82.290 195.395 ;
        RECT 82.170 195.285 82.345 195.390 ;
        RECT 82.185 195.280 82.345 195.285 ;
        RECT 82.640 195.255 82.810 195.445 ;
        RECT 86.325 195.290 86.485 195.400 ;
        RECT 88.615 195.255 88.785 195.445 ;
        RECT 89.070 195.285 89.190 195.395 ;
        RECT 89.535 195.255 89.705 195.445 ;
        RECT 92.295 195.235 92.465 195.425 ;
        RECT 92.755 195.235 92.925 195.425 ;
        RECT 93.210 195.255 93.380 195.445 ;
        RECT 94.135 195.235 94.305 195.425 ;
        RECT 94.595 195.255 94.765 195.445 ;
        RECT 96.435 195.255 96.605 195.445 ;
        RECT 99.655 195.235 99.825 195.425 ;
        RECT 100.105 195.255 100.275 195.445 ;
        RECT 103.335 195.255 103.505 195.445 ;
        RECT 104.255 195.255 104.425 195.425 ;
        RECT 104.275 195.235 104.425 195.255 ;
        RECT 106.560 195.235 106.730 195.425 ;
        RECT 107.945 195.280 108.105 195.390 ;
        RECT 109.315 195.235 109.485 195.425 ;
        RECT 113.455 195.255 113.625 195.445 ;
        RECT 114.190 195.255 114.360 195.445 ;
        RECT 118.060 195.255 118.230 195.475 ;
        RECT 119.720 195.445 120.665 195.475 ;
        RECT 122.055 195.445 123.425 196.225 ;
        RECT 123.435 195.445 128.945 196.255 ;
        RECT 129.875 195.445 131.245 196.255 ;
        RECT 118.515 195.235 118.685 195.425 ;
        RECT 120.825 195.290 120.985 195.400 ;
        RECT 123.115 195.255 123.285 195.445 ;
        RECT 123.575 195.255 123.745 195.445 ;
        RECT 124.035 195.235 124.205 195.425 ;
        RECT 129.105 195.290 129.265 195.400 ;
        RECT 129.550 195.285 129.670 195.395 ;
        RECT 130.935 195.235 131.105 195.445 ;
        RECT 57.195 194.425 58.565 195.235 ;
        RECT 58.575 194.425 64.085 195.235 ;
        RECT 64.095 194.425 69.605 195.235 ;
        RECT 69.615 194.425 75.125 195.235 ;
        RECT 75.135 194.425 77.885 195.235 ;
        RECT 77.895 194.555 81.795 195.235 ;
        RECT 77.895 194.325 78.825 194.555 ;
        RECT 82.965 194.365 83.395 195.150 ;
        RECT 83.500 194.555 92.605 195.235 ;
        RECT 92.615 194.455 93.985 195.235 ;
        RECT 93.995 194.425 99.505 195.235 ;
        RECT 99.515 194.425 103.185 195.235 ;
        RECT 104.275 194.415 106.205 195.235 ;
        RECT 105.255 194.325 106.205 194.415 ;
        RECT 106.415 194.325 107.765 195.235 ;
        RECT 108.725 194.365 109.155 195.150 ;
        RECT 109.175 194.555 118.280 195.235 ;
        RECT 118.375 194.425 123.885 195.235 ;
        RECT 123.895 194.425 129.405 195.235 ;
        RECT 129.875 194.425 131.245 195.235 ;
      LAYER nwell ;
        RECT 57.000 191.205 131.440 194.035 ;
      LAYER pwell ;
        RECT 57.195 190.005 58.565 190.815 ;
        RECT 58.575 190.005 64.085 190.815 ;
        RECT 64.095 190.005 69.605 190.815 ;
        RECT 70.085 190.090 70.515 190.875 ;
        RECT 70.535 190.005 76.045 190.815 ;
        RECT 76.055 190.005 77.885 190.815 ;
        RECT 78.355 190.005 81.525 190.915 ;
        RECT 81.575 190.715 82.520 190.915 ;
        RECT 81.575 190.035 84.325 190.715 ;
        RECT 81.575 190.005 82.520 190.035 ;
        RECT 57.335 189.795 57.505 190.005 ;
        RECT 58.715 189.795 58.885 190.005 ;
        RECT 64.235 189.795 64.405 190.005 ;
        RECT 69.755 189.955 69.925 189.985 ;
        RECT 69.750 189.845 69.925 189.955 ;
        RECT 69.755 189.795 69.925 189.845 ;
        RECT 70.675 189.815 70.845 190.005 ;
        RECT 75.275 189.795 75.445 189.985 ;
        RECT 76.195 189.815 76.365 190.005 ;
        RECT 78.030 189.845 78.150 189.955 ;
        RECT 57.195 188.985 58.565 189.795 ;
        RECT 58.575 188.985 64.085 189.795 ;
        RECT 64.095 188.985 69.605 189.795 ;
        RECT 69.615 188.985 75.125 189.795 ;
        RECT 75.135 188.985 78.805 189.795 ;
        RECT 78.960 189.765 79.130 189.985 ;
        RECT 81.255 189.815 81.425 190.005 ;
        RECT 81.715 189.795 81.885 189.985 ;
        RECT 83.555 189.795 83.725 189.985 ;
        RECT 84.010 189.815 84.180 190.035 ;
        RECT 84.335 190.005 85.705 190.815 ;
        RECT 86.765 190.685 87.695 190.915 ;
        RECT 85.860 190.005 87.695 190.685 ;
        RECT 88.055 190.685 89.405 190.915 ;
        RECT 90.940 190.685 91.850 190.905 ;
        RECT 88.055 190.005 95.365 190.685 ;
        RECT 95.845 190.090 96.275 190.875 ;
        RECT 96.335 190.685 97.685 190.915 ;
        RECT 99.220 190.685 100.130 190.905 ;
        RECT 96.335 190.005 103.645 190.685 ;
        RECT 103.655 190.005 109.165 190.815 ;
        RECT 109.215 190.685 110.565 190.915 ;
        RECT 112.100 190.685 113.010 190.905 ;
        RECT 109.215 190.005 116.525 190.685 ;
        RECT 116.535 190.005 120.205 190.815 ;
        RECT 120.215 190.005 121.585 190.815 ;
        RECT 121.605 190.090 122.035 190.875 ;
        RECT 122.055 190.005 127.565 190.815 ;
        RECT 127.575 190.005 129.405 190.815 ;
        RECT 129.875 190.005 131.245 190.815 ;
        RECT 84.475 189.815 84.645 190.005 ;
        RECT 85.860 189.985 86.025 190.005 ;
        RECT 85.855 189.815 86.025 189.985 ;
        RECT 87.230 189.845 87.350 189.955 ;
        RECT 80.620 189.765 81.565 189.795 ;
        RECT 78.815 189.085 81.565 189.765 ;
        RECT 80.620 188.885 81.565 189.085 ;
        RECT 81.575 188.985 82.945 189.795 ;
        RECT 82.965 188.925 83.395 189.710 ;
        RECT 83.415 188.985 87.085 189.795 ;
        RECT 87.700 189.765 87.870 189.985 ;
        RECT 90.915 189.795 91.085 189.985 ;
        RECT 95.055 189.815 95.225 190.005 ;
        RECT 95.510 189.845 95.630 189.955 ;
        RECT 96.430 189.845 96.550 189.955 ;
        RECT 96.895 189.795 97.065 189.985 ;
        RECT 101.490 189.795 101.660 189.985 ;
        RECT 101.955 189.795 102.125 189.985 ;
        RECT 103.335 189.815 103.505 190.005 ;
        RECT 103.795 189.815 103.965 190.005 ;
        RECT 107.475 189.795 107.645 189.985 ;
        RECT 109.315 189.795 109.485 189.985 ;
        RECT 114.835 189.795 115.005 189.985 ;
        RECT 116.215 189.815 116.385 190.005 ;
        RECT 116.675 189.815 116.845 190.005 ;
        RECT 120.355 189.795 120.525 190.005 ;
        RECT 122.195 189.815 122.365 190.005 ;
        RECT 125.875 189.795 126.045 189.985 ;
        RECT 127.255 189.795 127.425 189.985 ;
        RECT 127.715 189.815 127.885 190.005 ;
        RECT 129.105 189.840 129.265 189.950 ;
        RECT 129.550 189.845 129.670 189.955 ;
        RECT 130.935 189.795 131.105 190.005 ;
        RECT 89.830 189.765 90.765 189.795 ;
        RECT 87.700 189.565 90.765 189.765 ;
        RECT 87.555 189.085 90.765 189.565 ;
        RECT 87.555 188.885 88.485 189.085 ;
        RECT 89.815 188.885 90.765 189.085 ;
        RECT 90.775 188.985 96.285 189.795 ;
        RECT 96.865 189.115 100.330 189.795 ;
        RECT 99.410 188.885 100.330 189.115 ;
        RECT 100.455 188.885 101.805 189.795 ;
        RECT 101.815 188.985 107.325 189.795 ;
        RECT 107.335 188.985 108.705 189.795 ;
        RECT 108.725 188.925 109.155 189.710 ;
        RECT 109.175 188.985 114.685 189.795 ;
        RECT 114.695 188.985 120.205 189.795 ;
        RECT 120.215 188.985 125.725 189.795 ;
        RECT 125.735 188.985 127.105 189.795 ;
        RECT 127.115 189.115 128.945 189.795 ;
        RECT 127.600 188.885 128.945 189.115 ;
        RECT 129.875 188.985 131.245 189.795 ;
      LAYER nwell ;
        RECT 57.000 185.765 131.440 188.595 ;
      LAYER pwell ;
        RECT 57.195 184.565 58.565 185.375 ;
        RECT 58.575 184.565 64.085 185.375 ;
        RECT 64.095 184.565 69.605 185.375 ;
        RECT 70.085 184.650 70.515 185.435 ;
        RECT 70.535 184.565 76.045 185.375 ;
        RECT 76.055 184.565 81.565 185.375 ;
        RECT 81.575 184.565 87.085 185.375 ;
        RECT 87.095 184.565 92.605 185.375 ;
        RECT 92.615 184.565 95.365 185.375 ;
        RECT 95.845 184.650 96.275 185.435 ;
        RECT 96.295 184.565 101.805 185.375 ;
        RECT 101.815 184.565 107.325 185.375 ;
        RECT 107.335 184.565 112.845 185.375 ;
        RECT 112.855 184.565 118.365 185.375 ;
        RECT 118.375 184.565 121.125 185.375 ;
        RECT 121.605 184.650 122.035 185.435 ;
        RECT 122.055 184.565 127.565 185.375 ;
        RECT 127.575 184.565 129.405 185.375 ;
        RECT 129.875 184.565 131.245 185.375 ;
        RECT 57.335 184.355 57.505 184.565 ;
        RECT 58.715 184.355 58.885 184.565 ;
        RECT 64.235 184.355 64.405 184.565 ;
        RECT 69.755 184.515 69.925 184.545 ;
        RECT 69.750 184.405 69.925 184.515 ;
        RECT 69.755 184.355 69.925 184.405 ;
        RECT 70.675 184.375 70.845 184.565 ;
        RECT 75.275 184.355 75.445 184.545 ;
        RECT 76.195 184.375 76.365 184.565 ;
        RECT 80.795 184.355 80.965 184.545 ;
        RECT 81.715 184.375 81.885 184.565 ;
        RECT 82.630 184.405 82.750 184.515 ;
        RECT 83.555 184.355 83.725 184.545 ;
        RECT 87.235 184.375 87.405 184.565 ;
        RECT 89.075 184.355 89.245 184.545 ;
        RECT 92.755 184.375 92.925 184.565 ;
        RECT 94.595 184.355 94.765 184.545 ;
        RECT 95.510 184.405 95.630 184.515 ;
        RECT 96.435 184.375 96.605 184.565 ;
        RECT 100.115 184.355 100.285 184.545 ;
        RECT 101.955 184.375 102.125 184.565 ;
        RECT 105.635 184.355 105.805 184.545 ;
        RECT 107.475 184.375 107.645 184.565 ;
        RECT 108.390 184.405 108.510 184.515 ;
        RECT 109.315 184.355 109.485 184.545 ;
        RECT 112.995 184.375 113.165 184.565 ;
        RECT 114.835 184.355 115.005 184.545 ;
        RECT 118.515 184.375 118.685 184.565 ;
        RECT 120.355 184.355 120.525 184.545 ;
        RECT 121.270 184.405 121.390 184.515 ;
        RECT 122.195 184.375 122.365 184.565 ;
        RECT 125.875 184.355 126.045 184.545 ;
        RECT 127.715 184.375 127.885 184.565 ;
        RECT 129.550 184.405 129.670 184.515 ;
        RECT 130.935 184.355 131.105 184.565 ;
        RECT 57.195 183.545 58.565 184.355 ;
        RECT 58.575 183.545 64.085 184.355 ;
        RECT 64.095 183.545 69.605 184.355 ;
        RECT 69.615 183.545 75.125 184.355 ;
        RECT 75.135 183.545 80.645 184.355 ;
        RECT 80.655 183.545 82.485 184.355 ;
        RECT 82.965 183.485 83.395 184.270 ;
        RECT 83.415 183.545 88.925 184.355 ;
        RECT 88.935 183.545 94.445 184.355 ;
        RECT 94.455 183.545 99.965 184.355 ;
        RECT 99.975 183.545 105.485 184.355 ;
        RECT 105.495 183.545 108.245 184.355 ;
        RECT 108.725 183.485 109.155 184.270 ;
        RECT 109.175 183.545 114.685 184.355 ;
        RECT 114.695 183.545 120.205 184.355 ;
        RECT 120.215 183.545 125.725 184.355 ;
        RECT 125.735 183.545 129.405 184.355 ;
        RECT 129.875 183.545 131.245 184.355 ;
      LAYER nwell ;
        RECT 57.000 180.325 131.440 183.155 ;
      LAYER pwell ;
        RECT 57.195 179.125 58.565 179.935 ;
        RECT 58.575 179.125 64.085 179.935 ;
        RECT 64.095 179.125 69.605 179.935 ;
        RECT 70.085 179.210 70.515 179.995 ;
        RECT 70.535 179.125 76.045 179.935 ;
        RECT 76.055 179.125 81.565 179.935 ;
        RECT 81.575 179.125 87.085 179.935 ;
        RECT 87.095 179.125 92.605 179.935 ;
        RECT 92.615 179.125 95.365 179.935 ;
        RECT 95.845 179.210 96.275 179.995 ;
        RECT 96.295 179.125 101.805 179.935 ;
        RECT 101.815 179.125 107.325 179.935 ;
        RECT 107.335 179.125 112.845 179.935 ;
        RECT 112.855 179.125 118.365 179.935 ;
        RECT 118.375 179.125 121.125 179.935 ;
        RECT 121.605 179.210 122.035 179.995 ;
        RECT 122.055 179.125 127.565 179.935 ;
        RECT 127.575 179.125 129.405 179.935 ;
        RECT 129.875 179.125 131.245 179.935 ;
        RECT 57.335 178.915 57.505 179.125 ;
        RECT 58.715 178.915 58.885 179.125 ;
        RECT 64.235 178.915 64.405 179.125 ;
        RECT 69.755 179.075 69.925 179.105 ;
        RECT 69.750 178.965 69.925 179.075 ;
        RECT 69.755 178.915 69.925 178.965 ;
        RECT 70.675 178.935 70.845 179.125 ;
        RECT 75.275 178.915 75.445 179.105 ;
        RECT 76.195 178.935 76.365 179.125 ;
        RECT 80.795 178.915 80.965 179.105 ;
        RECT 81.715 178.935 81.885 179.125 ;
        RECT 82.630 178.965 82.750 179.075 ;
        RECT 83.555 178.915 83.725 179.105 ;
        RECT 87.235 178.935 87.405 179.125 ;
        RECT 89.075 178.915 89.245 179.105 ;
        RECT 92.755 178.935 92.925 179.125 ;
        RECT 94.595 178.915 94.765 179.105 ;
        RECT 95.510 178.965 95.630 179.075 ;
        RECT 96.435 178.935 96.605 179.125 ;
        RECT 100.115 178.915 100.285 179.105 ;
        RECT 101.955 178.935 102.125 179.125 ;
        RECT 105.635 178.915 105.805 179.105 ;
        RECT 107.475 178.935 107.645 179.125 ;
        RECT 108.390 178.965 108.510 179.075 ;
        RECT 109.315 178.915 109.485 179.105 ;
        RECT 112.995 178.935 113.165 179.125 ;
        RECT 114.835 178.915 115.005 179.105 ;
        RECT 118.515 178.935 118.685 179.125 ;
        RECT 120.355 178.915 120.525 179.105 ;
        RECT 121.270 178.965 121.390 179.075 ;
        RECT 122.195 178.935 122.365 179.125 ;
        RECT 125.875 178.915 126.045 179.105 ;
        RECT 127.715 178.935 127.885 179.125 ;
        RECT 129.550 178.965 129.670 179.075 ;
        RECT 130.935 178.915 131.105 179.125 ;
        RECT 57.195 178.105 58.565 178.915 ;
        RECT 58.575 178.105 64.085 178.915 ;
        RECT 64.095 178.105 69.605 178.915 ;
        RECT 69.615 178.105 75.125 178.915 ;
        RECT 75.135 178.105 80.645 178.915 ;
        RECT 80.655 178.105 82.485 178.915 ;
        RECT 82.965 178.045 83.395 178.830 ;
        RECT 83.415 178.105 88.925 178.915 ;
        RECT 88.935 178.105 94.445 178.915 ;
        RECT 94.455 178.105 99.965 178.915 ;
        RECT 99.975 178.105 105.485 178.915 ;
        RECT 105.495 178.105 108.245 178.915 ;
        RECT 108.725 178.045 109.155 178.830 ;
        RECT 109.175 178.105 114.685 178.915 ;
        RECT 114.695 178.105 120.205 178.915 ;
        RECT 120.215 178.105 125.725 178.915 ;
        RECT 125.735 178.105 129.405 178.915 ;
        RECT 129.875 178.105 131.245 178.915 ;
      LAYER nwell ;
        RECT 57.000 174.885 131.440 177.715 ;
      LAYER pwell ;
        RECT 57.195 173.685 58.565 174.495 ;
        RECT 58.575 173.685 64.085 174.495 ;
        RECT 64.095 173.685 69.605 174.495 ;
        RECT 70.085 173.770 70.515 174.555 ;
        RECT 70.535 173.685 76.045 174.495 ;
        RECT 76.055 173.685 81.565 174.495 ;
        RECT 81.575 173.685 87.085 174.495 ;
        RECT 87.095 173.685 92.605 174.495 ;
        RECT 92.615 173.685 95.365 174.495 ;
        RECT 95.845 173.770 96.275 174.555 ;
        RECT 96.295 173.685 101.805 174.495 ;
        RECT 101.815 173.685 107.325 174.495 ;
        RECT 107.335 173.685 112.845 174.495 ;
        RECT 112.855 173.685 118.365 174.495 ;
        RECT 118.375 173.685 121.125 174.495 ;
        RECT 121.605 173.770 122.035 174.555 ;
        RECT 122.055 173.685 127.565 174.495 ;
        RECT 127.575 173.685 129.405 174.495 ;
        RECT 129.875 173.685 131.245 174.495 ;
        RECT 57.335 173.475 57.505 173.685 ;
        RECT 58.715 173.475 58.885 173.685 ;
        RECT 64.235 173.475 64.405 173.685 ;
        RECT 69.755 173.635 69.925 173.665 ;
        RECT 69.750 173.525 69.925 173.635 ;
        RECT 69.755 173.475 69.925 173.525 ;
        RECT 70.675 173.495 70.845 173.685 ;
        RECT 75.275 173.475 75.445 173.665 ;
        RECT 76.195 173.495 76.365 173.685 ;
        RECT 80.795 173.475 80.965 173.665 ;
        RECT 81.715 173.495 81.885 173.685 ;
        RECT 82.630 173.525 82.750 173.635 ;
        RECT 83.555 173.475 83.725 173.665 ;
        RECT 87.235 173.495 87.405 173.685 ;
        RECT 89.075 173.475 89.245 173.665 ;
        RECT 92.755 173.495 92.925 173.685 ;
        RECT 94.595 173.475 94.765 173.665 ;
        RECT 95.510 173.525 95.630 173.635 ;
        RECT 96.435 173.495 96.605 173.685 ;
        RECT 100.115 173.475 100.285 173.665 ;
        RECT 101.955 173.495 102.125 173.685 ;
        RECT 105.635 173.475 105.805 173.665 ;
        RECT 107.475 173.495 107.645 173.685 ;
        RECT 108.390 173.525 108.510 173.635 ;
        RECT 109.315 173.475 109.485 173.665 ;
        RECT 112.995 173.495 113.165 173.685 ;
        RECT 114.835 173.475 115.005 173.665 ;
        RECT 118.515 173.495 118.685 173.685 ;
        RECT 120.355 173.475 120.525 173.665 ;
        RECT 121.270 173.525 121.390 173.635 ;
        RECT 122.195 173.495 122.365 173.685 ;
        RECT 125.875 173.475 126.045 173.665 ;
        RECT 127.715 173.495 127.885 173.685 ;
        RECT 129.550 173.525 129.670 173.635 ;
        RECT 130.935 173.475 131.105 173.685 ;
        RECT 57.195 172.665 58.565 173.475 ;
        RECT 58.575 172.665 64.085 173.475 ;
        RECT 64.095 172.665 69.605 173.475 ;
        RECT 69.615 172.665 75.125 173.475 ;
        RECT 75.135 172.665 80.645 173.475 ;
        RECT 80.655 172.665 82.485 173.475 ;
        RECT 82.965 172.605 83.395 173.390 ;
        RECT 83.415 172.665 88.925 173.475 ;
        RECT 88.935 172.665 94.445 173.475 ;
        RECT 94.455 172.665 99.965 173.475 ;
        RECT 99.975 172.665 105.485 173.475 ;
        RECT 105.495 172.665 108.245 173.475 ;
        RECT 108.725 172.605 109.155 173.390 ;
        RECT 109.175 172.665 114.685 173.475 ;
        RECT 114.695 172.665 120.205 173.475 ;
        RECT 120.215 172.665 125.725 173.475 ;
        RECT 125.735 172.665 129.405 173.475 ;
        RECT 129.875 172.665 131.245 173.475 ;
      LAYER nwell ;
        RECT 57.000 169.445 131.440 172.275 ;
      LAYER pwell ;
        RECT 57.195 168.245 58.565 169.055 ;
        RECT 58.575 168.245 64.085 169.055 ;
        RECT 64.095 168.245 69.605 169.055 ;
        RECT 70.085 168.330 70.515 169.115 ;
        RECT 70.535 168.245 76.045 169.055 ;
        RECT 76.055 168.245 81.565 169.055 ;
        RECT 81.575 168.245 87.085 169.055 ;
        RECT 87.095 168.245 92.605 169.055 ;
        RECT 92.615 168.245 95.365 169.055 ;
        RECT 95.845 168.330 96.275 169.115 ;
        RECT 96.295 168.245 101.805 169.055 ;
        RECT 101.815 168.245 107.325 169.055 ;
        RECT 107.335 168.245 112.845 169.055 ;
        RECT 112.855 168.245 118.365 169.055 ;
        RECT 118.375 168.245 121.125 169.055 ;
        RECT 121.605 168.330 122.035 169.115 ;
        RECT 122.055 168.245 127.565 169.055 ;
        RECT 127.575 168.245 129.405 169.055 ;
        RECT 129.875 168.245 131.245 169.055 ;
        RECT 57.335 168.035 57.505 168.245 ;
        RECT 58.715 168.035 58.885 168.245 ;
        RECT 64.235 168.035 64.405 168.245 ;
        RECT 69.755 168.195 69.925 168.225 ;
        RECT 69.750 168.085 69.925 168.195 ;
        RECT 69.755 168.035 69.925 168.085 ;
        RECT 70.675 168.055 70.845 168.245 ;
        RECT 75.275 168.035 75.445 168.225 ;
        RECT 76.195 168.055 76.365 168.245 ;
        RECT 80.795 168.035 80.965 168.225 ;
        RECT 81.715 168.055 81.885 168.245 ;
        RECT 82.630 168.085 82.750 168.195 ;
        RECT 83.555 168.035 83.725 168.225 ;
        RECT 87.235 168.055 87.405 168.245 ;
        RECT 89.075 168.035 89.245 168.225 ;
        RECT 92.755 168.055 92.925 168.245 ;
        RECT 94.595 168.035 94.765 168.225 ;
        RECT 95.510 168.085 95.630 168.195 ;
        RECT 96.435 168.055 96.605 168.245 ;
        RECT 100.115 168.035 100.285 168.225 ;
        RECT 101.955 168.055 102.125 168.245 ;
        RECT 105.635 168.035 105.805 168.225 ;
        RECT 107.475 168.055 107.645 168.245 ;
        RECT 108.390 168.085 108.510 168.195 ;
        RECT 109.315 168.035 109.485 168.225 ;
        RECT 112.995 168.055 113.165 168.245 ;
        RECT 114.835 168.035 115.005 168.225 ;
        RECT 118.515 168.055 118.685 168.245 ;
        RECT 120.355 168.035 120.525 168.225 ;
        RECT 121.270 168.085 121.390 168.195 ;
        RECT 122.195 168.055 122.365 168.245 ;
        RECT 125.875 168.035 126.045 168.225 ;
        RECT 127.715 168.055 127.885 168.245 ;
        RECT 129.550 168.085 129.670 168.195 ;
        RECT 130.935 168.035 131.105 168.245 ;
        RECT 57.195 167.225 58.565 168.035 ;
        RECT 58.575 167.225 64.085 168.035 ;
        RECT 64.095 167.225 69.605 168.035 ;
        RECT 69.615 167.225 75.125 168.035 ;
        RECT 75.135 167.225 80.645 168.035 ;
        RECT 80.655 167.225 82.485 168.035 ;
        RECT 82.965 167.165 83.395 167.950 ;
        RECT 83.415 167.225 88.925 168.035 ;
        RECT 88.935 167.225 94.445 168.035 ;
        RECT 94.455 167.225 99.965 168.035 ;
        RECT 99.975 167.225 105.485 168.035 ;
        RECT 105.495 167.225 108.245 168.035 ;
        RECT 108.725 167.165 109.155 167.950 ;
        RECT 109.175 167.225 114.685 168.035 ;
        RECT 114.695 167.225 120.205 168.035 ;
        RECT 120.215 167.225 125.725 168.035 ;
        RECT 125.735 167.225 129.405 168.035 ;
        RECT 129.875 167.225 131.245 168.035 ;
      LAYER nwell ;
        RECT 57.000 164.005 131.440 166.835 ;
      LAYER pwell ;
        RECT 57.195 162.805 58.565 163.615 ;
        RECT 58.575 162.805 64.085 163.615 ;
        RECT 64.095 162.805 69.605 163.615 ;
        RECT 70.085 162.890 70.515 163.675 ;
        RECT 70.535 162.805 76.045 163.615 ;
        RECT 76.055 162.805 81.565 163.615 ;
        RECT 81.575 162.805 87.085 163.615 ;
        RECT 87.095 162.805 92.605 163.615 ;
        RECT 92.615 162.805 95.365 163.615 ;
        RECT 95.845 162.890 96.275 163.675 ;
        RECT 96.295 162.805 101.805 163.615 ;
        RECT 101.815 162.805 107.325 163.615 ;
        RECT 107.335 162.805 112.845 163.615 ;
        RECT 112.855 162.805 118.365 163.615 ;
        RECT 118.375 162.805 121.125 163.615 ;
        RECT 121.605 162.890 122.035 163.675 ;
        RECT 122.055 162.805 127.565 163.615 ;
        RECT 127.575 162.805 129.405 163.615 ;
        RECT 129.875 162.805 131.245 163.615 ;
        RECT 57.335 162.595 57.505 162.805 ;
        RECT 58.715 162.595 58.885 162.805 ;
        RECT 64.235 162.595 64.405 162.805 ;
        RECT 69.755 162.755 69.925 162.785 ;
        RECT 69.750 162.645 69.925 162.755 ;
        RECT 69.755 162.595 69.925 162.645 ;
        RECT 70.675 162.615 70.845 162.805 ;
        RECT 75.275 162.595 75.445 162.785 ;
        RECT 76.195 162.615 76.365 162.805 ;
        RECT 80.795 162.595 80.965 162.785 ;
        RECT 81.715 162.615 81.885 162.805 ;
        RECT 82.630 162.645 82.750 162.755 ;
        RECT 83.555 162.595 83.725 162.785 ;
        RECT 87.235 162.615 87.405 162.805 ;
        RECT 89.075 162.595 89.245 162.785 ;
        RECT 92.755 162.615 92.925 162.805 ;
        RECT 94.595 162.595 94.765 162.785 ;
        RECT 95.510 162.645 95.630 162.755 ;
        RECT 96.435 162.615 96.605 162.805 ;
        RECT 100.115 162.595 100.285 162.785 ;
        RECT 101.955 162.615 102.125 162.805 ;
        RECT 105.635 162.595 105.805 162.785 ;
        RECT 107.475 162.615 107.645 162.805 ;
        RECT 108.390 162.645 108.510 162.755 ;
        RECT 109.315 162.595 109.485 162.785 ;
        RECT 112.995 162.615 113.165 162.805 ;
        RECT 114.835 162.595 115.005 162.785 ;
        RECT 118.515 162.615 118.685 162.805 ;
        RECT 120.355 162.595 120.525 162.785 ;
        RECT 121.270 162.645 121.390 162.755 ;
        RECT 122.195 162.615 122.365 162.805 ;
        RECT 125.875 162.595 126.045 162.785 ;
        RECT 127.715 162.615 127.885 162.805 ;
        RECT 129.550 162.645 129.670 162.755 ;
        RECT 130.935 162.595 131.105 162.805 ;
        RECT 57.195 161.785 58.565 162.595 ;
        RECT 58.575 161.785 64.085 162.595 ;
        RECT 64.095 161.785 69.605 162.595 ;
        RECT 69.615 161.785 75.125 162.595 ;
        RECT 75.135 161.785 80.645 162.595 ;
        RECT 80.655 161.785 82.485 162.595 ;
        RECT 82.965 161.725 83.395 162.510 ;
        RECT 83.415 161.785 88.925 162.595 ;
        RECT 88.935 161.785 94.445 162.595 ;
        RECT 94.455 161.785 99.965 162.595 ;
        RECT 99.975 161.785 105.485 162.595 ;
        RECT 105.495 161.785 108.245 162.595 ;
        RECT 108.725 161.725 109.155 162.510 ;
        RECT 109.175 161.785 114.685 162.595 ;
        RECT 114.695 161.785 120.205 162.595 ;
        RECT 120.215 161.785 125.725 162.595 ;
        RECT 125.735 161.785 129.405 162.595 ;
        RECT 129.875 161.785 131.245 162.595 ;
      LAYER nwell ;
        RECT 57.000 158.565 131.440 161.395 ;
      LAYER pwell ;
        RECT 57.195 157.365 58.565 158.175 ;
        RECT 58.575 157.365 64.085 158.175 ;
        RECT 64.095 157.365 69.605 158.175 ;
        RECT 70.085 157.450 70.515 158.235 ;
        RECT 70.535 157.365 76.045 158.175 ;
        RECT 76.055 157.365 81.565 158.175 ;
        RECT 81.575 157.365 87.085 158.175 ;
        RECT 87.095 157.365 92.605 158.175 ;
        RECT 92.615 157.365 95.365 158.175 ;
        RECT 95.845 157.450 96.275 158.235 ;
        RECT 96.295 157.365 101.805 158.175 ;
        RECT 101.815 157.365 107.325 158.175 ;
        RECT 107.335 157.365 112.845 158.175 ;
        RECT 112.855 157.365 118.365 158.175 ;
        RECT 118.375 157.365 121.125 158.175 ;
        RECT 121.605 157.450 122.035 158.235 ;
        RECT 122.055 157.365 127.565 158.175 ;
        RECT 127.575 157.365 129.405 158.175 ;
        RECT 129.875 157.365 131.245 158.175 ;
        RECT 57.335 157.155 57.505 157.365 ;
        RECT 58.715 157.155 58.885 157.365 ;
        RECT 64.235 157.155 64.405 157.365 ;
        RECT 69.755 157.315 69.925 157.345 ;
        RECT 69.750 157.205 69.925 157.315 ;
        RECT 69.755 157.155 69.925 157.205 ;
        RECT 70.675 157.175 70.845 157.365 ;
        RECT 75.275 157.155 75.445 157.345 ;
        RECT 76.195 157.175 76.365 157.365 ;
        RECT 80.795 157.155 80.965 157.345 ;
        RECT 81.715 157.175 81.885 157.365 ;
        RECT 82.630 157.205 82.750 157.315 ;
        RECT 83.555 157.155 83.725 157.345 ;
        RECT 87.235 157.175 87.405 157.365 ;
        RECT 89.075 157.155 89.245 157.345 ;
        RECT 92.755 157.175 92.925 157.365 ;
        RECT 94.595 157.155 94.765 157.345 ;
        RECT 95.510 157.205 95.630 157.315 ;
        RECT 96.435 157.175 96.605 157.365 ;
        RECT 100.115 157.155 100.285 157.345 ;
        RECT 101.955 157.175 102.125 157.365 ;
        RECT 105.635 157.155 105.805 157.345 ;
        RECT 107.475 157.175 107.645 157.365 ;
        RECT 108.390 157.205 108.510 157.315 ;
        RECT 109.315 157.155 109.485 157.345 ;
        RECT 112.995 157.175 113.165 157.365 ;
        RECT 114.835 157.155 115.005 157.345 ;
        RECT 118.515 157.175 118.685 157.365 ;
        RECT 120.355 157.155 120.525 157.345 ;
        RECT 121.270 157.205 121.390 157.315 ;
        RECT 122.195 157.175 122.365 157.365 ;
        RECT 125.875 157.155 126.045 157.345 ;
        RECT 127.715 157.175 127.885 157.365 ;
        RECT 129.550 157.205 129.670 157.315 ;
        RECT 130.935 157.155 131.105 157.365 ;
        RECT 57.195 156.345 58.565 157.155 ;
        RECT 58.575 156.345 64.085 157.155 ;
        RECT 64.095 156.345 69.605 157.155 ;
        RECT 69.615 156.345 75.125 157.155 ;
        RECT 75.135 156.345 80.645 157.155 ;
        RECT 80.655 156.345 82.485 157.155 ;
        RECT 82.965 156.285 83.395 157.070 ;
        RECT 83.415 156.345 88.925 157.155 ;
        RECT 88.935 156.345 94.445 157.155 ;
        RECT 94.455 156.345 99.965 157.155 ;
        RECT 99.975 156.345 105.485 157.155 ;
        RECT 105.495 156.345 108.245 157.155 ;
        RECT 108.725 156.285 109.155 157.070 ;
        RECT 109.175 156.345 114.685 157.155 ;
        RECT 114.695 156.345 120.205 157.155 ;
        RECT 120.215 156.345 125.725 157.155 ;
        RECT 125.735 156.345 129.405 157.155 ;
        RECT 129.875 156.345 131.245 157.155 ;
      LAYER nwell ;
        RECT 57.000 153.125 131.440 155.955 ;
      LAYER pwell ;
        RECT 57.195 151.925 58.565 152.735 ;
        RECT 58.575 151.925 64.085 152.735 ;
        RECT 64.095 151.925 69.605 152.735 ;
        RECT 70.085 152.010 70.515 152.795 ;
        RECT 70.535 151.925 76.045 152.735 ;
        RECT 76.055 151.925 81.565 152.735 ;
        RECT 81.575 151.925 87.085 152.735 ;
        RECT 87.095 151.925 92.605 152.735 ;
        RECT 92.615 151.925 95.365 152.735 ;
        RECT 95.845 152.010 96.275 152.795 ;
        RECT 96.295 151.925 101.805 152.735 ;
        RECT 101.815 151.925 107.325 152.735 ;
        RECT 107.335 151.925 112.845 152.735 ;
        RECT 112.855 151.925 118.365 152.735 ;
        RECT 118.375 151.925 121.125 152.735 ;
        RECT 121.605 152.010 122.035 152.795 ;
        RECT 122.055 151.925 127.565 152.735 ;
        RECT 127.575 151.925 129.405 152.735 ;
        RECT 129.875 151.925 131.245 152.735 ;
        RECT 57.335 151.715 57.505 151.925 ;
        RECT 58.715 151.715 58.885 151.925 ;
        RECT 64.235 151.715 64.405 151.925 ;
        RECT 69.755 151.875 69.925 151.905 ;
        RECT 69.750 151.765 69.925 151.875 ;
        RECT 69.755 151.715 69.925 151.765 ;
        RECT 70.675 151.735 70.845 151.925 ;
        RECT 75.275 151.715 75.445 151.905 ;
        RECT 76.195 151.735 76.365 151.925 ;
        RECT 80.795 151.715 80.965 151.905 ;
        RECT 81.715 151.735 81.885 151.925 ;
        RECT 82.630 151.765 82.750 151.875 ;
        RECT 83.555 151.715 83.725 151.905 ;
        RECT 87.235 151.735 87.405 151.925 ;
        RECT 89.075 151.715 89.245 151.905 ;
        RECT 92.755 151.735 92.925 151.925 ;
        RECT 94.595 151.715 94.765 151.905 ;
        RECT 95.510 151.765 95.630 151.875 ;
        RECT 96.435 151.735 96.605 151.925 ;
        RECT 100.115 151.715 100.285 151.905 ;
        RECT 101.955 151.735 102.125 151.925 ;
        RECT 105.635 151.715 105.805 151.905 ;
        RECT 107.475 151.735 107.645 151.925 ;
        RECT 108.390 151.765 108.510 151.875 ;
        RECT 111.615 151.715 111.785 151.905 ;
        RECT 112.075 151.715 112.245 151.905 ;
        RECT 112.995 151.735 113.165 151.925 ;
        RECT 117.595 151.715 117.765 151.905 ;
        RECT 118.515 151.735 118.685 151.925 ;
        RECT 121.270 151.765 121.390 151.875 ;
        RECT 122.195 151.735 122.365 151.925 ;
        RECT 123.115 151.715 123.285 151.905 ;
        RECT 127.715 151.735 127.885 151.925 ;
        RECT 128.635 151.715 128.805 151.905 ;
        RECT 129.550 151.765 129.670 151.875 ;
        RECT 130.935 151.715 131.105 151.925 ;
        RECT 57.195 150.905 58.565 151.715 ;
        RECT 58.575 150.905 64.085 151.715 ;
        RECT 64.095 150.905 69.605 151.715 ;
        RECT 69.615 150.905 75.125 151.715 ;
        RECT 75.135 150.905 80.645 151.715 ;
        RECT 80.655 150.905 82.485 151.715 ;
        RECT 82.965 150.845 83.395 151.630 ;
        RECT 83.415 150.905 88.925 151.715 ;
        RECT 88.935 150.905 94.445 151.715 ;
        RECT 94.455 150.905 99.965 151.715 ;
        RECT 99.975 150.905 105.485 151.715 ;
        RECT 105.495 150.905 108.245 151.715 ;
        RECT 108.725 150.845 109.155 151.630 ;
        RECT 109.185 151.035 111.925 151.715 ;
        RECT 111.935 150.905 117.445 151.715 ;
        RECT 117.455 150.905 122.965 151.715 ;
        RECT 122.975 150.905 128.485 151.715 ;
        RECT 128.495 150.905 129.865 151.715 ;
        RECT 129.875 150.905 131.245 151.715 ;
      LAYER nwell ;
        RECT 57.000 147.685 131.440 150.515 ;
      LAYER pwell ;
        RECT 57.195 146.485 58.565 147.295 ;
        RECT 58.575 146.485 64.085 147.295 ;
        RECT 64.095 146.485 69.605 147.295 ;
        RECT 70.085 146.570 70.515 147.355 ;
        RECT 70.535 146.485 76.045 147.295 ;
        RECT 76.055 146.485 81.565 147.295 ;
        RECT 81.575 146.485 87.085 147.295 ;
        RECT 87.095 146.485 92.605 147.295 ;
        RECT 92.615 146.485 95.365 147.295 ;
        RECT 95.845 146.570 96.275 147.355 ;
        RECT 96.295 146.485 101.805 147.295 ;
        RECT 101.815 146.485 107.325 147.295 ;
        RECT 107.335 146.485 112.845 147.295 ;
        RECT 112.855 146.485 118.365 147.295 ;
        RECT 118.375 146.485 121.125 147.295 ;
        RECT 121.605 146.570 122.035 147.355 ;
        RECT 122.055 146.485 127.565 147.295 ;
        RECT 127.575 146.485 129.405 147.295 ;
        RECT 129.875 146.485 131.245 147.295 ;
        RECT 57.335 146.275 57.505 146.485 ;
        RECT 58.715 146.275 58.885 146.485 ;
        RECT 64.235 146.275 64.405 146.485 ;
        RECT 69.755 146.435 69.925 146.465 ;
        RECT 69.750 146.325 69.925 146.435 ;
        RECT 69.755 146.275 69.925 146.325 ;
        RECT 70.675 146.295 70.845 146.485 ;
        RECT 75.275 146.275 75.445 146.465 ;
        RECT 76.195 146.295 76.365 146.485 ;
        RECT 80.795 146.275 80.965 146.465 ;
        RECT 81.715 146.295 81.885 146.485 ;
        RECT 82.630 146.325 82.750 146.435 ;
        RECT 83.555 146.275 83.725 146.465 ;
        RECT 87.235 146.295 87.405 146.485 ;
        RECT 89.075 146.275 89.245 146.465 ;
        RECT 92.755 146.295 92.925 146.485 ;
        RECT 94.595 146.275 94.765 146.465 ;
        RECT 95.510 146.325 95.630 146.435 ;
        RECT 96.435 146.295 96.605 146.485 ;
        RECT 100.115 146.275 100.285 146.465 ;
        RECT 101.955 146.295 102.125 146.485 ;
        RECT 105.635 146.275 105.805 146.465 ;
        RECT 107.475 146.295 107.645 146.485 ;
        RECT 108.390 146.325 108.510 146.435 ;
        RECT 109.315 146.275 109.485 146.465 ;
        RECT 112.995 146.295 113.165 146.485 ;
        RECT 114.835 146.275 115.005 146.465 ;
        RECT 118.515 146.295 118.685 146.485 ;
        RECT 120.355 146.275 120.525 146.465 ;
        RECT 121.270 146.325 121.390 146.435 ;
        RECT 122.195 146.295 122.365 146.485 ;
        RECT 125.875 146.275 126.045 146.465 ;
        RECT 127.715 146.295 127.885 146.485 ;
        RECT 129.550 146.325 129.670 146.435 ;
        RECT 130.935 146.275 131.105 146.485 ;
        RECT 57.195 145.465 58.565 146.275 ;
        RECT 58.575 145.465 64.085 146.275 ;
        RECT 64.095 145.465 69.605 146.275 ;
        RECT 69.615 145.465 75.125 146.275 ;
        RECT 75.135 145.465 80.645 146.275 ;
        RECT 80.655 145.465 82.485 146.275 ;
        RECT 82.965 145.405 83.395 146.190 ;
        RECT 83.415 145.465 88.925 146.275 ;
        RECT 88.935 145.465 94.445 146.275 ;
        RECT 94.455 145.465 99.965 146.275 ;
        RECT 99.975 145.465 105.485 146.275 ;
        RECT 105.495 145.465 108.245 146.275 ;
        RECT 108.725 145.405 109.155 146.190 ;
        RECT 109.175 145.465 114.685 146.275 ;
        RECT 114.695 145.465 120.205 146.275 ;
        RECT 120.215 145.465 125.725 146.275 ;
        RECT 125.735 145.465 129.405 146.275 ;
        RECT 129.875 145.465 131.245 146.275 ;
      LAYER nwell ;
        RECT 57.000 142.245 131.440 145.075 ;
      LAYER pwell ;
        RECT 57.195 141.045 58.565 141.855 ;
        RECT 58.575 141.045 64.085 141.855 ;
        RECT 64.095 141.045 69.605 141.855 ;
        RECT 70.085 141.130 70.515 141.915 ;
        RECT 70.535 141.045 76.045 141.855 ;
        RECT 76.055 141.045 81.565 141.855 ;
        RECT 81.575 141.045 87.085 141.855 ;
        RECT 87.095 141.045 92.605 141.855 ;
        RECT 92.615 141.045 95.365 141.855 ;
        RECT 95.845 141.130 96.275 141.915 ;
        RECT 96.295 141.045 101.805 141.855 ;
        RECT 101.815 141.045 107.325 141.855 ;
        RECT 107.335 141.045 112.845 141.855 ;
        RECT 112.855 141.045 118.365 141.855 ;
        RECT 118.375 141.045 121.125 141.855 ;
        RECT 121.605 141.130 122.035 141.915 ;
        RECT 122.055 141.045 127.565 141.855 ;
        RECT 127.575 141.045 129.405 141.855 ;
        RECT 129.875 141.045 131.245 141.855 ;
        RECT 57.335 140.835 57.505 141.045 ;
        RECT 58.715 140.835 58.885 141.045 ;
        RECT 64.235 140.835 64.405 141.045 ;
        RECT 69.755 140.995 69.925 141.025 ;
        RECT 69.750 140.885 69.925 140.995 ;
        RECT 69.755 140.835 69.925 140.885 ;
        RECT 70.675 140.855 70.845 141.045 ;
        RECT 75.275 140.835 75.445 141.025 ;
        RECT 76.195 140.855 76.365 141.045 ;
        RECT 80.795 140.835 80.965 141.025 ;
        RECT 81.715 140.855 81.885 141.045 ;
        RECT 82.630 140.885 82.750 140.995 ;
        RECT 83.555 140.835 83.725 141.025 ;
        RECT 87.235 140.855 87.405 141.045 ;
        RECT 89.075 140.835 89.245 141.025 ;
        RECT 92.755 140.855 92.925 141.045 ;
        RECT 94.595 140.835 94.765 141.025 ;
        RECT 95.510 140.885 95.630 140.995 ;
        RECT 96.435 140.855 96.605 141.045 ;
        RECT 100.115 140.835 100.285 141.025 ;
        RECT 101.955 140.855 102.125 141.045 ;
        RECT 105.635 140.835 105.805 141.025 ;
        RECT 107.475 140.855 107.645 141.045 ;
        RECT 108.390 140.885 108.510 140.995 ;
        RECT 109.315 140.835 109.485 141.025 ;
        RECT 112.995 140.855 113.165 141.045 ;
        RECT 114.835 140.835 115.005 141.025 ;
        RECT 118.515 140.855 118.685 141.045 ;
        RECT 120.355 140.835 120.525 141.025 ;
        RECT 121.270 140.885 121.390 140.995 ;
        RECT 122.195 140.855 122.365 141.045 ;
        RECT 125.875 140.835 126.045 141.025 ;
        RECT 127.715 140.855 127.885 141.045 ;
        RECT 129.550 140.885 129.670 140.995 ;
        RECT 130.935 140.835 131.105 141.045 ;
        RECT 57.195 140.025 58.565 140.835 ;
        RECT 58.575 140.025 64.085 140.835 ;
        RECT 64.095 140.025 69.605 140.835 ;
        RECT 69.615 140.025 75.125 140.835 ;
        RECT 75.135 140.025 80.645 140.835 ;
        RECT 80.655 140.025 82.485 140.835 ;
        RECT 82.965 139.965 83.395 140.750 ;
        RECT 83.415 140.025 88.925 140.835 ;
        RECT 88.935 140.025 94.445 140.835 ;
        RECT 94.455 140.025 99.965 140.835 ;
        RECT 99.975 140.025 105.485 140.835 ;
        RECT 105.495 140.025 108.245 140.835 ;
        RECT 108.725 139.965 109.155 140.750 ;
        RECT 109.175 140.025 114.685 140.835 ;
        RECT 114.695 140.025 120.205 140.835 ;
        RECT 120.215 140.025 125.725 140.835 ;
        RECT 125.735 140.025 129.405 140.835 ;
        RECT 129.875 140.025 131.245 140.835 ;
      LAYER nwell ;
        RECT 57.000 136.805 131.440 139.635 ;
      LAYER pwell ;
        RECT 57.195 135.605 58.565 136.415 ;
        RECT 58.575 135.605 64.085 136.415 ;
        RECT 64.095 135.605 69.605 136.415 ;
        RECT 70.085 135.690 70.515 136.475 ;
        RECT 70.535 135.605 76.045 136.415 ;
        RECT 76.055 135.605 81.565 136.415 ;
        RECT 81.575 135.605 87.085 136.415 ;
        RECT 87.095 135.605 92.605 136.415 ;
        RECT 92.615 135.605 95.365 136.415 ;
        RECT 95.845 135.690 96.275 136.475 ;
        RECT 96.295 135.605 101.805 136.415 ;
        RECT 101.815 135.605 107.325 136.415 ;
        RECT 107.335 135.605 112.845 136.415 ;
        RECT 112.855 135.605 118.365 136.415 ;
        RECT 118.375 135.605 121.125 136.415 ;
        RECT 121.605 135.690 122.035 136.475 ;
        RECT 122.055 135.605 127.565 136.415 ;
        RECT 127.575 135.605 129.405 136.415 ;
        RECT 129.875 135.605 131.245 136.415 ;
        RECT 57.335 135.395 57.505 135.605 ;
        RECT 58.715 135.395 58.885 135.605 ;
        RECT 64.235 135.395 64.405 135.605 ;
        RECT 69.755 135.555 69.925 135.585 ;
        RECT 69.750 135.445 69.925 135.555 ;
        RECT 69.755 135.395 69.925 135.445 ;
        RECT 70.675 135.415 70.845 135.605 ;
        RECT 75.275 135.395 75.445 135.585 ;
        RECT 76.195 135.415 76.365 135.605 ;
        RECT 80.795 135.395 80.965 135.585 ;
        RECT 81.715 135.415 81.885 135.605 ;
        RECT 82.630 135.445 82.750 135.555 ;
        RECT 83.555 135.395 83.725 135.585 ;
        RECT 87.235 135.415 87.405 135.605 ;
        RECT 89.075 135.395 89.245 135.585 ;
        RECT 92.755 135.415 92.925 135.605 ;
        RECT 94.595 135.395 94.765 135.585 ;
        RECT 95.510 135.445 95.630 135.555 ;
        RECT 96.435 135.415 96.605 135.605 ;
        RECT 100.115 135.395 100.285 135.585 ;
        RECT 101.955 135.415 102.125 135.605 ;
        RECT 105.635 135.395 105.805 135.585 ;
        RECT 107.475 135.415 107.645 135.605 ;
        RECT 108.390 135.445 108.510 135.555 ;
        RECT 109.315 135.395 109.485 135.585 ;
        RECT 112.995 135.415 113.165 135.605 ;
        RECT 114.835 135.395 115.005 135.585 ;
        RECT 118.515 135.415 118.685 135.605 ;
        RECT 120.355 135.395 120.525 135.585 ;
        RECT 121.270 135.445 121.390 135.555 ;
        RECT 122.195 135.415 122.365 135.605 ;
        RECT 125.875 135.395 126.045 135.585 ;
        RECT 127.715 135.415 127.885 135.605 ;
        RECT 129.550 135.445 129.670 135.555 ;
        RECT 130.935 135.395 131.105 135.605 ;
        RECT 57.195 134.585 58.565 135.395 ;
        RECT 58.575 134.585 64.085 135.395 ;
        RECT 64.095 134.585 69.605 135.395 ;
        RECT 69.615 134.585 75.125 135.395 ;
        RECT 75.135 134.585 80.645 135.395 ;
        RECT 80.655 134.585 82.485 135.395 ;
        RECT 82.965 134.525 83.395 135.310 ;
        RECT 83.415 134.585 88.925 135.395 ;
        RECT 88.935 134.585 94.445 135.395 ;
        RECT 94.455 134.585 99.965 135.395 ;
        RECT 99.975 134.585 105.485 135.395 ;
        RECT 105.495 134.585 108.245 135.395 ;
        RECT 108.725 134.525 109.155 135.310 ;
        RECT 109.175 134.585 114.685 135.395 ;
        RECT 114.695 134.585 120.205 135.395 ;
        RECT 120.215 134.585 125.725 135.395 ;
        RECT 125.735 134.585 129.405 135.395 ;
        RECT 129.875 134.585 131.245 135.395 ;
      LAYER nwell ;
        RECT 57.000 131.365 131.440 134.195 ;
      LAYER pwell ;
        RECT 57.195 130.165 58.565 130.975 ;
        RECT 58.575 130.165 64.085 130.975 ;
        RECT 64.095 130.165 69.605 130.975 ;
        RECT 70.085 130.250 70.515 131.035 ;
        RECT 70.535 130.165 76.045 130.975 ;
        RECT 76.055 130.165 81.565 130.975 ;
        RECT 81.575 130.165 82.945 130.975 ;
        RECT 82.965 130.250 83.395 131.035 ;
        RECT 83.415 130.165 88.925 130.975 ;
        RECT 88.935 130.165 94.445 130.975 ;
        RECT 94.455 130.165 95.825 130.975 ;
        RECT 95.845 130.250 96.275 131.035 ;
        RECT 96.295 130.165 101.805 130.975 ;
        RECT 101.815 130.165 107.325 130.975 ;
        RECT 107.335 130.165 108.705 130.975 ;
        RECT 108.725 130.250 109.155 131.035 ;
        RECT 109.175 130.165 114.685 130.975 ;
        RECT 114.695 130.165 120.205 130.975 ;
        RECT 120.215 130.165 121.585 130.975 ;
        RECT 121.605 130.250 122.035 131.035 ;
        RECT 122.055 130.165 127.565 130.975 ;
        RECT 127.575 130.165 129.405 130.975 ;
        RECT 129.875 130.165 131.245 130.975 ;
        RECT 57.335 129.975 57.505 130.165 ;
        RECT 58.715 129.975 58.885 130.165 ;
        RECT 64.235 129.975 64.405 130.165 ;
        RECT 69.750 130.005 69.870 130.115 ;
        RECT 70.675 129.975 70.845 130.165 ;
        RECT 76.195 129.975 76.365 130.165 ;
        RECT 81.715 129.975 81.885 130.165 ;
        RECT 83.555 129.975 83.725 130.165 ;
        RECT 89.075 129.975 89.245 130.165 ;
        RECT 94.595 129.975 94.765 130.165 ;
        RECT 96.435 129.975 96.605 130.165 ;
        RECT 101.955 129.975 102.125 130.165 ;
        RECT 107.475 129.975 107.645 130.165 ;
        RECT 109.315 129.975 109.485 130.165 ;
        RECT 114.835 129.975 115.005 130.165 ;
        RECT 120.355 129.975 120.525 130.165 ;
        RECT 122.195 129.975 122.365 130.165 ;
        RECT 127.715 129.975 127.885 130.165 ;
        RECT 129.550 130.005 129.670 130.115 ;
        RECT 130.935 129.975 131.105 130.165 ;
        RECT 137.120 86.570 144.290 88.580 ;
        RECT 147.120 86.570 154.290 88.580 ;
        RECT 138.120 80.570 141.130 84.470 ;
        RECT 142.120 80.570 145.130 84.470 ;
        RECT 147.120 80.570 150.130 84.470 ;
        RECT 151.120 80.570 154.130 84.470 ;
        RECT 140.120 74.570 143.130 78.470 ;
        RECT 149.120 74.570 152.130 78.470 ;
      LAYER li1 ;
        RECT 57.190 203.415 131.250 203.585 ;
        RECT 57.275 202.325 58.485 203.415 ;
        RECT 58.655 202.325 60.325 203.415 ;
        RECT 57.275 201.615 57.795 202.155 ;
        RECT 57.965 201.785 58.485 202.325 ;
        RECT 58.655 201.635 59.405 202.155 ;
        RECT 59.575 201.805 60.325 202.325 ;
        RECT 61.035 202.485 61.215 203.245 ;
        RECT 61.395 202.655 61.725 203.415 ;
        RECT 61.035 202.315 61.710 202.485 ;
        RECT 61.895 202.340 62.165 203.245 ;
        RECT 62.335 202.980 67.680 203.415 ;
        RECT 61.540 202.170 61.710 202.315 ;
        RECT 60.975 201.765 61.315 202.135 ;
        RECT 61.540 201.840 61.815 202.170 ;
        RECT 57.275 200.865 58.485 201.615 ;
        RECT 58.655 200.865 60.325 201.635 ;
        RECT 61.540 201.585 61.710 201.840 ;
        RECT 61.045 201.415 61.710 201.585 ;
        RECT 61.985 201.540 62.165 202.340 ;
        RECT 61.045 201.035 61.215 201.415 ;
        RECT 61.395 200.865 61.725 201.245 ;
        RECT 61.905 201.035 62.165 201.540 ;
        RECT 63.920 201.410 64.260 202.240 ;
        RECT 65.740 201.730 66.090 202.980 ;
        RECT 67.855 202.325 69.525 203.415 ;
        RECT 67.855 201.635 68.605 202.155 ;
        RECT 68.775 201.805 69.525 202.325 ;
        RECT 70.155 202.250 70.445 203.415 ;
        RECT 70.615 202.445 70.885 203.215 ;
        RECT 71.055 202.635 71.385 203.415 ;
        RECT 71.590 202.810 71.775 203.215 ;
        RECT 71.945 202.990 72.280 203.415 ;
        RECT 71.590 202.635 72.255 202.810 ;
        RECT 70.615 202.275 71.745 202.445 ;
        RECT 62.335 200.865 67.680 201.410 ;
        RECT 67.855 200.865 69.525 201.635 ;
        RECT 70.155 200.865 70.445 201.590 ;
        RECT 70.615 201.365 70.785 202.275 ;
        RECT 70.955 201.525 71.315 202.105 ;
        RECT 71.495 201.775 71.745 202.275 ;
        RECT 71.915 201.605 72.255 202.635 ;
        RECT 72.455 202.325 75.045 203.415 ;
        RECT 75.220 202.615 75.535 203.415 ;
        RECT 75.800 203.060 76.880 203.230 ;
        RECT 75.800 202.445 75.970 203.060 ;
        RECT 71.570 201.435 72.255 201.605 ;
        RECT 72.455 201.635 73.665 202.155 ;
        RECT 73.835 201.805 75.045 202.325 ;
        RECT 70.615 201.035 70.875 201.365 ;
        RECT 71.085 200.865 71.360 201.345 ;
        RECT 71.570 201.035 71.775 201.435 ;
        RECT 71.945 200.865 72.280 201.265 ;
        RECT 72.455 200.865 75.045 201.635 ;
        RECT 75.215 201.435 75.485 202.445 ;
        RECT 75.655 202.275 75.970 202.445 ;
        RECT 75.655 201.605 75.825 202.275 ;
        RECT 76.140 202.105 76.375 202.785 ;
        RECT 76.545 202.275 76.880 203.060 ;
        RECT 77.055 202.325 79.645 203.415 ;
        RECT 75.995 201.775 76.375 202.105 ;
        RECT 76.545 201.775 76.880 202.105 ;
        RECT 77.055 201.635 78.265 202.155 ;
        RECT 78.435 201.805 79.645 202.325 ;
        RECT 80.355 202.485 80.535 203.245 ;
        RECT 80.715 202.655 81.045 203.415 ;
        RECT 80.355 202.315 81.030 202.485 ;
        RECT 81.215 202.340 81.485 203.245 ;
        RECT 80.860 202.170 81.030 202.315 ;
        RECT 80.295 201.765 80.635 202.135 ;
        RECT 80.860 201.840 81.135 202.170 ;
        RECT 75.655 201.435 76.880 201.605 ;
        RECT 75.285 200.865 75.615 201.265 ;
        RECT 75.785 201.165 75.955 201.435 ;
        RECT 76.125 200.865 76.455 201.265 ;
        RECT 76.625 201.165 76.880 201.435 ;
        RECT 77.055 200.865 79.645 201.635 ;
        RECT 80.860 201.585 81.030 201.840 ;
        RECT 80.365 201.415 81.030 201.585 ;
        RECT 81.305 201.540 81.485 202.340 ;
        RECT 81.655 202.325 82.865 203.415 ;
        RECT 80.365 201.035 80.535 201.415 ;
        RECT 80.715 200.865 81.045 201.245 ;
        RECT 81.225 201.035 81.485 201.540 ;
        RECT 81.655 201.615 82.175 202.155 ;
        RECT 82.345 201.785 82.865 202.325 ;
        RECT 83.035 202.250 83.325 203.415 ;
        RECT 83.495 202.325 85.165 203.415 ;
        RECT 83.495 201.635 84.245 202.155 ;
        RECT 84.415 201.805 85.165 202.325 ;
        RECT 85.395 202.275 85.605 203.415 ;
        RECT 85.775 202.265 86.105 203.245 ;
        RECT 86.275 202.275 86.505 203.415 ;
        RECT 86.715 202.275 87.100 203.245 ;
        RECT 87.270 202.955 87.595 203.415 ;
        RECT 88.115 202.785 88.395 203.245 ;
        RECT 87.270 202.565 88.395 202.785 ;
        RECT 81.655 200.865 82.865 201.615 ;
        RECT 83.035 200.865 83.325 201.590 ;
        RECT 83.495 200.865 85.165 201.635 ;
        RECT 85.395 200.865 85.605 201.685 ;
        RECT 85.775 201.665 86.025 202.265 ;
        RECT 86.195 201.855 86.525 202.105 ;
        RECT 85.775 201.035 86.105 201.665 ;
        RECT 86.275 200.865 86.505 201.685 ;
        RECT 86.715 201.605 86.995 202.275 ;
        RECT 87.270 202.105 87.720 202.565 ;
        RECT 88.585 202.395 88.985 203.245 ;
        RECT 89.385 202.955 89.655 203.415 ;
        RECT 89.825 202.785 90.110 203.245 ;
        RECT 87.165 201.775 87.720 202.105 ;
        RECT 87.890 201.835 88.985 202.395 ;
        RECT 87.270 201.665 87.720 201.775 ;
        RECT 86.715 201.035 87.100 201.605 ;
        RECT 87.270 201.495 88.395 201.665 ;
        RECT 87.270 200.865 87.595 201.325 ;
        RECT 88.115 201.035 88.395 201.495 ;
        RECT 88.585 201.035 88.985 201.835 ;
        RECT 89.155 202.565 90.110 202.785 ;
        RECT 89.155 201.665 89.365 202.565 ;
        RECT 90.485 202.485 90.655 203.245 ;
        RECT 90.835 202.655 91.165 203.415 ;
        RECT 89.535 201.835 90.225 202.395 ;
        RECT 90.485 202.315 91.150 202.485 ;
        RECT 91.335 202.340 91.605 203.245 ;
        RECT 90.980 202.170 91.150 202.315 ;
        RECT 90.415 201.765 90.745 202.135 ;
        RECT 90.980 201.840 91.265 202.170 ;
        RECT 89.155 201.495 90.110 201.665 ;
        RECT 90.980 201.585 91.150 201.840 ;
        RECT 89.385 200.865 89.655 201.325 ;
        RECT 89.825 201.035 90.110 201.495 ;
        RECT 90.485 201.415 91.150 201.585 ;
        RECT 91.435 201.540 91.605 202.340 ;
        RECT 91.775 202.325 95.285 203.415 ;
        RECT 90.485 201.035 90.655 201.415 ;
        RECT 90.835 200.865 91.165 201.245 ;
        RECT 91.345 201.035 91.605 201.540 ;
        RECT 91.775 201.635 93.425 202.155 ;
        RECT 93.595 201.805 95.285 202.325 ;
        RECT 95.915 202.250 96.205 203.415 ;
        RECT 97.385 202.485 97.555 203.245 ;
        RECT 97.735 202.655 98.065 203.415 ;
        RECT 97.385 202.315 98.050 202.485 ;
        RECT 98.235 202.340 98.505 203.245 ;
        RECT 98.675 202.820 98.935 203.000 ;
        RECT 99.140 202.990 99.500 203.415 ;
        RECT 100.015 202.990 100.345 203.415 ;
        RECT 100.525 202.905 101.725 203.145 ;
        RECT 98.675 202.735 100.310 202.820 ;
        RECT 102.930 202.785 103.215 203.245 ;
        RECT 103.385 202.955 103.655 203.415 ;
        RECT 98.675 202.650 101.250 202.735 ;
        RECT 98.675 202.590 99.355 202.650 ;
        RECT 97.880 202.170 98.050 202.315 ;
        RECT 97.315 201.765 97.645 202.135 ;
        RECT 97.880 201.840 98.165 202.170 ;
        RECT 91.775 200.865 95.285 201.635 ;
        RECT 95.915 200.865 96.205 201.590 ;
        RECT 97.880 201.585 98.050 201.840 ;
        RECT 97.385 201.415 98.050 201.585 ;
        RECT 98.335 201.540 98.505 202.340 ;
        RECT 98.675 201.855 99.015 202.420 ;
        RECT 99.185 201.685 99.355 202.590 ;
        RECT 100.140 202.565 101.250 202.650 ;
        RECT 97.385 201.035 97.555 201.415 ;
        RECT 97.735 200.865 98.065 201.245 ;
        RECT 98.245 201.035 98.505 201.540 ;
        RECT 98.675 201.515 99.355 201.685 ;
        RECT 99.525 202.275 99.920 202.480 ;
        RECT 98.675 201.070 98.935 201.515 ;
        RECT 99.525 201.375 99.695 202.275 ;
        RECT 99.865 201.715 100.035 202.105 ;
        RECT 100.285 201.855 100.820 202.395 ;
        RECT 101.080 202.105 101.250 202.565 ;
        RECT 101.420 202.275 101.725 202.705 ;
        RECT 102.930 202.565 103.885 202.785 ;
        RECT 101.080 201.775 101.380 202.105 ;
        RECT 99.865 201.685 100.185 201.715 ;
        RECT 99.865 201.605 100.750 201.685 ;
        RECT 101.555 201.605 101.725 202.275 ;
        RECT 102.815 201.835 103.505 202.395 ;
        RECT 103.675 201.665 103.885 202.565 ;
        RECT 99.865 201.545 101.725 201.605 ;
        RECT 100.015 201.515 101.725 201.545 ;
        RECT 100.580 201.435 101.725 201.515 ;
        RECT 99.185 200.865 99.355 201.345 ;
        RECT 99.525 201.045 99.875 201.375 ;
        RECT 100.110 200.865 100.280 201.345 ;
        RECT 100.580 201.085 100.750 201.435 ;
        RECT 101.420 201.385 101.725 201.435 ;
        RECT 102.930 201.495 103.885 201.665 ;
        RECT 104.055 202.395 104.455 203.245 ;
        RECT 104.645 202.785 104.925 203.245 ;
        RECT 105.445 202.955 105.770 203.415 ;
        RECT 104.645 202.565 105.770 202.785 ;
        RECT 104.055 201.835 105.150 202.395 ;
        RECT 105.320 202.105 105.770 202.565 ;
        RECT 105.940 202.275 106.325 203.245 ;
        RECT 106.495 202.325 108.165 203.415 ;
        RECT 100.920 200.865 101.250 201.265 ;
        RECT 101.420 201.085 101.675 201.385 ;
        RECT 102.930 201.035 103.215 201.495 ;
        RECT 103.385 200.865 103.655 201.325 ;
        RECT 104.055 201.035 104.455 201.835 ;
        RECT 105.320 201.775 105.875 202.105 ;
        RECT 105.320 201.665 105.770 201.775 ;
        RECT 104.645 201.495 105.770 201.665 ;
        RECT 106.045 201.605 106.325 202.275 ;
        RECT 104.645 201.035 104.925 201.495 ;
        RECT 105.445 200.865 105.770 201.325 ;
        RECT 105.940 201.035 106.325 201.605 ;
        RECT 106.495 201.635 107.245 202.155 ;
        RECT 107.415 201.805 108.165 202.325 ;
        RECT 108.795 202.250 109.085 203.415 ;
        RECT 109.255 202.820 109.690 203.245 ;
        RECT 109.860 202.990 110.245 203.415 ;
        RECT 109.255 202.650 110.245 202.820 ;
        RECT 109.255 201.775 109.740 202.480 ;
        RECT 109.910 202.105 110.245 202.650 ;
        RECT 110.415 202.455 110.840 203.245 ;
        RECT 111.010 202.820 111.285 203.245 ;
        RECT 111.455 202.990 111.840 203.415 ;
        RECT 111.010 202.625 111.840 202.820 ;
        RECT 110.415 202.275 111.320 202.455 ;
        RECT 109.910 201.775 110.320 202.105 ;
        RECT 110.490 201.775 111.320 202.275 ;
        RECT 111.490 202.105 111.840 202.625 ;
        RECT 112.010 202.455 112.255 203.245 ;
        RECT 112.445 202.820 112.700 203.245 ;
        RECT 112.870 202.990 113.255 203.415 ;
        RECT 112.445 202.625 113.255 202.820 ;
        RECT 112.010 202.275 112.735 202.455 ;
        RECT 111.490 201.775 111.915 202.105 ;
        RECT 112.085 201.775 112.735 202.275 ;
        RECT 112.905 202.105 113.255 202.625 ;
        RECT 113.425 202.275 113.685 203.245 ;
        RECT 114.045 202.690 114.375 203.415 ;
        RECT 112.905 201.775 113.330 202.105 ;
        RECT 106.495 200.865 108.165 201.635 ;
        RECT 109.910 201.605 110.245 201.775 ;
        RECT 110.490 201.605 110.840 201.775 ;
        RECT 111.490 201.605 111.840 201.775 ;
        RECT 112.085 201.605 112.255 201.775 ;
        RECT 112.905 201.605 113.255 201.775 ;
        RECT 113.500 201.605 113.685 202.275 ;
        RECT 108.795 200.865 109.085 201.590 ;
        RECT 109.255 201.435 110.245 201.605 ;
        RECT 109.255 201.035 109.690 201.435 ;
        RECT 109.860 200.865 110.245 201.265 ;
        RECT 110.415 201.035 110.840 201.605 ;
        RECT 111.030 201.435 111.840 201.605 ;
        RECT 111.030 201.035 111.285 201.435 ;
        RECT 111.455 200.865 111.840 201.265 ;
        RECT 112.010 201.035 112.255 201.605 ;
        RECT 112.445 201.435 113.255 201.605 ;
        RECT 112.445 201.035 112.700 201.435 ;
        RECT 112.870 200.865 113.255 201.265 ;
        RECT 113.425 201.035 113.685 201.605 ;
        RECT 113.855 201.035 114.375 202.520 ;
        RECT 114.545 201.695 115.065 203.245 ;
        RECT 115.235 202.325 118.745 203.415 ;
        RECT 115.235 201.635 116.885 202.155 ;
        RECT 117.055 201.805 118.745 202.325 ;
        RECT 119.005 202.485 119.175 203.245 ;
        RECT 119.355 202.655 119.685 203.415 ;
        RECT 119.005 202.315 119.670 202.485 ;
        RECT 119.855 202.340 120.125 203.245 ;
        RECT 119.500 202.170 119.670 202.315 ;
        RECT 118.935 201.765 119.265 202.135 ;
        RECT 119.500 201.840 119.785 202.170 ;
        RECT 114.545 200.865 114.885 201.525 ;
        RECT 115.235 200.865 118.745 201.635 ;
        RECT 119.500 201.585 119.670 201.840 ;
        RECT 119.005 201.415 119.670 201.585 ;
        RECT 119.955 201.540 120.125 202.340 ;
        RECT 120.295 202.325 121.505 203.415 ;
        RECT 119.005 201.035 119.175 201.415 ;
        RECT 119.355 200.865 119.685 201.245 ;
        RECT 119.865 201.035 120.125 201.540 ;
        RECT 120.295 201.615 120.815 202.155 ;
        RECT 120.985 201.785 121.505 202.325 ;
        RECT 121.675 202.250 121.965 203.415 ;
        RECT 122.135 202.980 127.480 203.415 ;
        RECT 120.295 200.865 121.505 201.615 ;
        RECT 121.675 200.865 121.965 201.590 ;
        RECT 123.720 201.410 124.060 202.240 ;
        RECT 125.540 201.730 125.890 202.980 ;
        RECT 127.655 202.325 129.325 203.415 ;
        RECT 127.655 201.635 128.405 202.155 ;
        RECT 128.575 201.805 129.325 202.325 ;
        RECT 129.955 202.325 131.165 203.415 ;
        RECT 129.955 201.785 130.475 202.325 ;
        RECT 122.135 200.865 127.480 201.410 ;
        RECT 127.655 200.865 129.325 201.635 ;
        RECT 130.645 201.615 131.165 202.155 ;
        RECT 129.955 200.865 131.165 201.615 ;
        RECT 57.190 200.695 131.250 200.865 ;
        RECT 57.275 199.945 58.485 200.695 ;
        RECT 58.655 200.150 64.000 200.695 ;
        RECT 64.175 200.150 69.520 200.695 ;
        RECT 57.275 199.405 57.795 199.945 ;
        RECT 57.965 199.235 58.485 199.775 ;
        RECT 60.240 199.320 60.580 200.150 ;
        RECT 57.275 198.145 58.485 199.235 ;
        RECT 62.060 198.580 62.410 199.830 ;
        RECT 65.760 199.320 66.100 200.150 ;
        RECT 69.695 199.925 71.365 200.695 ;
        RECT 72.045 200.305 72.375 200.695 ;
        RECT 72.545 200.125 72.715 200.445 ;
        RECT 72.885 200.305 73.215 200.695 ;
        RECT 73.630 200.295 74.585 200.465 ;
        RECT 71.995 199.955 74.245 200.125 ;
        RECT 67.580 198.580 67.930 199.830 ;
        RECT 69.695 199.405 70.445 199.925 ;
        RECT 70.615 199.235 71.365 199.755 ;
        RECT 58.655 198.145 64.000 198.580 ;
        RECT 64.175 198.145 69.520 198.580 ;
        RECT 69.695 198.145 71.365 199.235 ;
        RECT 71.995 198.995 72.165 199.955 ;
        RECT 72.335 199.335 72.580 199.785 ;
        RECT 72.750 199.505 73.300 199.705 ;
        RECT 73.470 199.535 73.845 199.705 ;
        RECT 73.470 199.335 73.640 199.535 ;
        RECT 74.015 199.455 74.245 199.955 ;
        RECT 72.335 199.165 73.640 199.335 ;
        RECT 74.415 199.415 74.585 200.295 ;
        RECT 74.755 199.860 75.045 200.695 ;
        RECT 75.215 200.315 76.600 200.525 ;
        RECT 75.215 200.045 75.505 200.315 ;
        RECT 75.675 199.955 76.100 200.145 ;
        RECT 76.270 200.125 76.600 200.315 ;
        RECT 76.835 200.295 77.165 200.695 ;
        RECT 77.340 200.125 77.670 200.525 ;
        RECT 77.875 200.135 78.045 200.695 ;
        RECT 76.270 199.955 77.670 200.125 ;
        RECT 78.215 199.955 78.725 200.525 ;
        RECT 75.215 199.455 75.490 199.785 ;
        RECT 74.415 199.245 75.045 199.415 ;
        RECT 71.995 198.315 72.375 198.995 ;
        RECT 72.965 198.145 73.135 198.995 ;
        RECT 73.305 198.825 74.545 198.995 ;
        RECT 73.305 198.315 73.635 198.825 ;
        RECT 73.805 198.145 73.975 198.655 ;
        RECT 74.145 198.315 74.545 198.825 ;
        RECT 74.725 198.315 75.045 199.245 ;
        RECT 75.215 198.145 75.505 199.285 ;
        RECT 75.675 198.945 75.845 199.955 ;
        RECT 76.015 199.120 76.370 199.785 ;
        RECT 76.555 199.120 76.830 199.785 ;
        RECT 77.000 199.455 77.345 199.785 ;
        RECT 77.635 199.705 77.805 199.785 ;
        RECT 78.175 199.705 78.365 199.785 ;
        RECT 77.555 199.455 77.805 199.705 ;
        RECT 78.000 199.455 78.365 199.705 ;
        RECT 75.675 198.695 76.630 198.945 ;
        RECT 76.300 198.485 76.630 198.695 ;
        RECT 77.000 198.655 77.325 199.455 ;
        RECT 78.000 199.285 78.170 199.455 ;
        RECT 78.550 199.285 78.725 199.955 ;
        RECT 79.820 199.930 80.275 200.695 ;
        RECT 80.550 200.315 81.850 200.525 ;
        RECT 82.105 200.335 82.435 200.695 ;
        RECT 81.680 200.165 81.850 200.315 ;
        RECT 82.605 200.195 82.865 200.525 ;
        RECT 80.750 199.705 80.970 200.105 ;
        RECT 79.815 199.505 80.305 199.705 ;
        RECT 80.495 199.495 80.970 199.705 ;
        RECT 81.215 199.705 81.425 200.105 ;
        RECT 81.680 200.040 82.435 200.165 ;
        RECT 81.680 199.995 82.525 200.040 ;
        RECT 82.255 199.875 82.525 199.995 ;
        RECT 81.215 199.495 81.545 199.705 ;
        RECT 81.715 199.435 82.125 199.740 ;
        RECT 77.495 199.115 78.170 199.285 ;
        RECT 77.495 198.485 77.665 199.115 ;
        RECT 76.300 198.315 77.665 198.485 ;
        RECT 77.835 198.145 78.125 198.945 ;
        RECT 78.340 198.325 78.725 199.285 ;
        RECT 79.820 199.265 80.995 199.325 ;
        RECT 82.355 199.300 82.525 199.875 ;
        RECT 82.325 199.265 82.525 199.300 ;
        RECT 79.820 199.155 82.525 199.265 ;
        RECT 79.820 198.535 80.075 199.155 ;
        RECT 80.665 199.095 82.465 199.155 ;
        RECT 80.665 199.065 80.995 199.095 ;
        RECT 82.695 198.995 82.865 200.195 ;
        RECT 83.035 199.970 83.325 200.695 ;
        RECT 83.585 200.015 83.755 200.390 ;
        RECT 83.555 199.845 83.755 200.015 ;
        RECT 83.945 200.165 84.175 200.470 ;
        RECT 84.345 200.335 84.675 200.695 ;
        RECT 84.870 200.165 85.160 200.515 ;
        RECT 83.945 199.995 85.160 200.165 ;
        RECT 85.845 200.040 86.175 200.475 ;
        RECT 86.345 200.085 86.515 200.695 ;
        RECT 83.585 199.825 83.755 199.845 ;
        RECT 85.795 199.955 86.175 200.040 ;
        RECT 86.685 199.955 87.015 200.480 ;
        RECT 87.275 200.165 87.485 200.695 ;
        RECT 87.760 200.245 88.545 200.415 ;
        RECT 88.715 200.245 89.120 200.415 ;
        RECT 85.795 199.915 86.020 199.955 ;
        RECT 83.585 199.655 84.105 199.825 ;
        RECT 80.325 198.895 80.510 198.985 ;
        RECT 81.100 198.895 81.935 198.905 ;
        RECT 80.325 198.695 81.935 198.895 ;
        RECT 80.325 198.655 80.555 198.695 ;
        RECT 79.820 198.315 80.155 198.535 ;
        RECT 81.160 198.145 81.515 198.525 ;
        RECT 81.685 198.315 81.935 198.695 ;
        RECT 82.185 198.145 82.435 198.925 ;
        RECT 82.605 198.315 82.865 198.995 ;
        RECT 83.035 198.145 83.325 199.310 ;
        RECT 83.500 199.125 83.745 199.485 ;
        RECT 83.935 199.275 84.105 199.655 ;
        RECT 84.275 199.455 84.660 199.785 ;
        RECT 84.840 199.675 85.100 199.785 ;
        RECT 84.840 199.505 85.105 199.675 ;
        RECT 84.840 199.455 85.100 199.505 ;
        RECT 83.935 198.995 84.285 199.275 ;
        RECT 83.500 198.145 83.755 198.945 ;
        RECT 83.955 198.315 84.285 198.995 ;
        RECT 84.465 198.405 84.660 199.455 ;
        RECT 85.795 199.335 85.965 199.915 ;
        RECT 86.685 199.785 86.885 199.955 ;
        RECT 87.760 199.785 87.930 200.245 ;
        RECT 86.135 199.455 86.885 199.785 ;
        RECT 87.055 199.455 87.930 199.785 ;
        RECT 85.795 199.285 86.010 199.335 ;
        RECT 84.840 198.145 85.160 199.285 ;
        RECT 85.795 199.205 86.185 199.285 ;
        RECT 85.855 198.360 86.185 199.205 ;
        RECT 86.695 199.250 86.885 199.455 ;
        RECT 86.355 198.145 86.525 199.155 ;
        RECT 86.695 198.875 87.590 199.250 ;
        RECT 86.695 198.315 87.035 198.875 ;
        RECT 87.265 198.145 87.580 198.645 ;
        RECT 87.760 198.615 87.930 199.455 ;
        RECT 88.100 199.745 88.565 200.075 ;
        RECT 88.950 200.015 89.120 200.245 ;
        RECT 89.300 200.195 89.670 200.695 ;
        RECT 89.990 200.245 90.665 200.415 ;
        RECT 90.860 200.245 91.195 200.415 ;
        RECT 88.100 198.785 88.420 199.745 ;
        RECT 88.950 199.715 89.780 200.015 ;
        RECT 88.590 198.815 88.780 199.535 ;
        RECT 88.950 198.645 89.120 199.715 ;
        RECT 89.580 199.685 89.780 199.715 ;
        RECT 89.290 199.465 89.460 199.535 ;
        RECT 89.990 199.465 90.160 200.245 ;
        RECT 91.025 200.105 91.195 200.245 ;
        RECT 91.365 200.235 91.615 200.695 ;
        RECT 89.290 199.295 90.160 199.465 ;
        RECT 90.330 199.825 90.855 200.045 ;
        RECT 91.025 199.975 91.250 200.105 ;
        RECT 89.290 199.205 89.800 199.295 ;
        RECT 87.760 198.445 88.645 198.615 ;
        RECT 88.870 198.315 89.120 198.645 ;
        RECT 89.290 198.145 89.460 198.945 ;
        RECT 89.630 198.590 89.800 199.205 ;
        RECT 90.330 199.125 90.500 199.825 ;
        RECT 89.970 198.760 90.500 199.125 ;
        RECT 90.670 199.060 90.910 199.655 ;
        RECT 91.080 198.870 91.250 199.975 ;
        RECT 91.420 199.115 91.700 200.065 ;
        RECT 90.945 198.740 91.250 198.870 ;
        RECT 89.630 198.420 90.735 198.590 ;
        RECT 90.945 198.315 91.195 198.740 ;
        RECT 91.365 198.145 91.630 198.605 ;
        RECT 91.870 198.315 92.055 200.435 ;
        RECT 92.225 200.315 92.555 200.695 ;
        RECT 92.725 200.145 92.895 200.435 ;
        RECT 92.230 199.975 92.895 200.145 ;
        RECT 93.245 200.145 93.415 200.435 ;
        RECT 93.585 200.315 93.915 200.695 ;
        RECT 93.245 199.975 93.910 200.145 ;
        RECT 92.230 198.985 92.460 199.975 ;
        RECT 92.630 199.155 92.980 199.805 ;
        RECT 93.160 199.155 93.510 199.805 ;
        RECT 93.680 198.985 93.910 199.975 ;
        RECT 92.230 198.815 92.895 198.985 ;
        RECT 92.225 198.145 92.555 198.645 ;
        RECT 92.725 198.315 92.895 198.815 ;
        RECT 93.245 198.815 93.910 198.985 ;
        RECT 93.245 198.315 93.415 198.815 ;
        RECT 93.585 198.145 93.915 198.645 ;
        RECT 94.085 198.315 94.270 200.435 ;
        RECT 94.525 200.235 94.775 200.695 ;
        RECT 94.945 200.245 95.280 200.415 ;
        RECT 95.475 200.245 96.150 200.415 ;
        RECT 94.945 200.105 95.115 200.245 ;
        RECT 94.440 199.115 94.720 200.065 ;
        RECT 94.890 199.975 95.115 200.105 ;
        RECT 94.890 198.870 95.060 199.975 ;
        RECT 95.285 199.825 95.810 200.045 ;
        RECT 95.230 199.060 95.470 199.655 ;
        RECT 95.640 199.125 95.810 199.825 ;
        RECT 95.980 199.465 96.150 200.245 ;
        RECT 96.470 200.195 96.840 200.695 ;
        RECT 97.020 200.245 97.425 200.415 ;
        RECT 97.595 200.245 98.380 200.415 ;
        RECT 97.020 200.015 97.190 200.245 ;
        RECT 96.360 199.715 97.190 200.015 ;
        RECT 97.575 199.745 98.040 200.075 ;
        RECT 96.360 199.685 96.560 199.715 ;
        RECT 96.680 199.465 96.850 199.535 ;
        RECT 95.980 199.295 96.850 199.465 ;
        RECT 96.340 199.205 96.850 199.295 ;
        RECT 94.890 198.740 95.195 198.870 ;
        RECT 95.640 198.760 96.170 199.125 ;
        RECT 94.510 198.145 94.775 198.605 ;
        RECT 94.945 198.315 95.195 198.740 ;
        RECT 96.340 198.590 96.510 199.205 ;
        RECT 95.405 198.420 96.510 198.590 ;
        RECT 96.680 198.145 96.850 198.945 ;
        RECT 97.020 198.645 97.190 199.715 ;
        RECT 97.360 198.815 97.550 199.535 ;
        RECT 97.720 198.785 98.040 199.745 ;
        RECT 98.210 199.785 98.380 200.245 ;
        RECT 98.655 200.165 98.865 200.695 ;
        RECT 99.125 199.955 99.455 200.480 ;
        RECT 99.625 200.085 99.795 200.695 ;
        RECT 99.965 200.040 100.295 200.475 ;
        RECT 99.965 199.955 100.345 200.040 ;
        RECT 99.255 199.785 99.455 199.955 ;
        RECT 100.120 199.915 100.345 199.955 ;
        RECT 98.210 199.455 99.085 199.785 ;
        RECT 99.255 199.455 100.005 199.785 ;
        RECT 97.020 198.315 97.270 198.645 ;
        RECT 98.210 198.615 98.380 199.455 ;
        RECT 99.255 199.250 99.445 199.455 ;
        RECT 100.175 199.335 100.345 199.915 ;
        RECT 100.790 199.885 101.035 200.490 ;
        RECT 101.255 200.160 101.765 200.695 ;
        RECT 100.130 199.285 100.345 199.335 ;
        RECT 98.550 198.875 99.445 199.250 ;
        RECT 99.955 199.205 100.345 199.285 ;
        RECT 100.515 199.715 101.745 199.885 ;
        RECT 97.495 198.445 98.380 198.615 ;
        RECT 98.560 198.145 98.875 198.645 ;
        RECT 99.105 198.315 99.445 198.875 ;
        RECT 99.615 198.145 99.785 199.155 ;
        RECT 99.955 198.360 100.285 199.205 ;
        RECT 100.515 198.905 100.855 199.715 ;
        RECT 101.025 199.150 101.775 199.340 ;
        RECT 100.515 198.495 101.030 198.905 ;
        RECT 101.265 198.145 101.435 198.905 ;
        RECT 101.605 198.485 101.775 199.150 ;
        RECT 101.945 199.165 102.135 200.525 ;
        RECT 102.305 200.355 102.580 200.525 ;
        RECT 102.305 200.185 102.585 200.355 ;
        RECT 102.305 199.365 102.580 200.185 ;
        RECT 102.770 200.160 103.300 200.525 ;
        RECT 103.725 200.295 104.055 200.695 ;
        RECT 103.125 200.125 103.300 200.160 ;
        RECT 102.785 199.165 102.955 199.965 ;
        RECT 101.945 198.995 102.955 199.165 ;
        RECT 103.125 199.955 104.055 200.125 ;
        RECT 104.225 199.955 104.480 200.525 ;
        RECT 103.125 198.825 103.295 199.955 ;
        RECT 103.885 199.785 104.055 199.955 ;
        RECT 102.170 198.655 103.295 198.825 ;
        RECT 103.465 199.455 103.660 199.785 ;
        RECT 103.885 199.455 104.140 199.785 ;
        RECT 103.465 198.485 103.635 199.455 ;
        RECT 104.310 199.285 104.480 199.955 ;
        RECT 104.715 199.875 104.925 200.695 ;
        RECT 105.095 199.895 105.425 200.525 ;
        RECT 105.095 199.295 105.345 199.895 ;
        RECT 105.595 199.875 105.825 200.695 ;
        RECT 106.035 199.925 108.625 200.695 ;
        RECT 108.795 199.970 109.085 200.695 ;
        RECT 109.255 199.925 110.925 200.695 ;
        RECT 111.560 200.145 111.815 200.435 ;
        RECT 111.985 200.315 112.315 200.695 ;
        RECT 111.560 199.975 112.310 200.145 ;
        RECT 105.515 199.455 105.845 199.705 ;
        RECT 106.035 199.405 107.245 199.925 ;
        RECT 101.605 198.315 103.635 198.485 ;
        RECT 103.805 198.145 103.975 199.285 ;
        RECT 104.145 198.315 104.480 199.285 ;
        RECT 104.715 198.145 104.925 199.285 ;
        RECT 105.095 198.315 105.425 199.295 ;
        RECT 105.595 198.145 105.825 199.285 ;
        RECT 107.415 199.235 108.625 199.755 ;
        RECT 109.255 199.405 110.005 199.925 ;
        RECT 106.035 198.145 108.625 199.235 ;
        RECT 108.795 198.145 109.085 199.310 ;
        RECT 110.175 199.235 110.925 199.755 ;
        RECT 109.255 198.145 110.925 199.235 ;
        RECT 111.560 199.155 111.910 199.805 ;
        RECT 112.080 198.985 112.310 199.975 ;
        RECT 111.560 198.815 112.310 198.985 ;
        RECT 111.560 198.315 111.815 198.815 ;
        RECT 111.985 198.145 112.315 198.645 ;
        RECT 112.485 198.315 112.655 200.435 ;
        RECT 113.015 200.335 113.345 200.695 ;
        RECT 113.515 200.305 114.010 200.475 ;
        RECT 114.215 200.305 115.070 200.475 ;
        RECT 112.885 199.115 113.345 200.165 ;
        RECT 112.825 198.330 113.150 199.115 ;
        RECT 113.515 198.945 113.685 200.305 ;
        RECT 113.855 199.395 114.205 200.015 ;
        RECT 114.375 199.795 114.730 200.015 ;
        RECT 114.375 199.205 114.545 199.795 ;
        RECT 114.900 199.595 115.070 200.305 ;
        RECT 115.945 200.235 116.275 200.695 ;
        RECT 116.485 200.335 116.835 200.505 ;
        RECT 115.275 199.765 116.065 200.015 ;
        RECT 116.485 199.945 116.745 200.335 ;
        RECT 117.055 200.245 118.005 200.525 ;
        RECT 118.175 200.255 118.365 200.695 ;
        RECT 118.535 200.315 119.605 200.485 ;
        RECT 116.235 199.595 116.405 199.775 ;
        RECT 113.515 198.775 113.910 198.945 ;
        RECT 114.080 198.815 114.545 199.205 ;
        RECT 114.715 199.425 116.405 199.595 ;
        RECT 113.740 198.645 113.910 198.775 ;
        RECT 114.715 198.645 114.885 199.425 ;
        RECT 116.575 199.255 116.745 199.945 ;
        RECT 115.245 199.085 116.745 199.255 ;
        RECT 116.935 199.285 117.145 200.075 ;
        RECT 117.315 199.455 117.665 200.075 ;
        RECT 117.835 199.465 118.005 200.245 ;
        RECT 118.535 200.085 118.705 200.315 ;
        RECT 118.175 199.915 118.705 200.085 ;
        RECT 118.175 199.635 118.395 199.915 ;
        RECT 118.875 199.745 119.115 200.145 ;
        RECT 117.835 199.295 118.240 199.465 ;
        RECT 118.575 199.375 119.115 199.745 ;
        RECT 119.285 199.960 119.605 200.315 ;
        RECT 119.850 200.235 120.155 200.695 ;
        RECT 120.325 199.985 120.580 200.515 ;
        RECT 119.285 199.785 119.610 199.960 ;
        RECT 119.285 199.485 120.200 199.785 ;
        RECT 119.460 199.455 120.200 199.485 ;
        RECT 116.935 199.125 117.610 199.285 ;
        RECT 118.070 199.205 118.240 199.295 ;
        RECT 116.935 199.115 117.900 199.125 ;
        RECT 116.575 198.945 116.745 199.085 ;
        RECT 113.320 198.145 113.570 198.605 ;
        RECT 113.740 198.315 113.990 198.645 ;
        RECT 114.205 198.315 114.885 198.645 ;
        RECT 115.055 198.745 116.130 198.915 ;
        RECT 116.575 198.775 117.135 198.945 ;
        RECT 117.440 198.825 117.900 199.115 ;
        RECT 118.070 199.035 119.290 199.205 ;
        RECT 115.055 198.405 115.225 198.745 ;
        RECT 115.460 198.145 115.790 198.575 ;
        RECT 115.960 198.405 116.130 198.745 ;
        RECT 116.425 198.145 116.795 198.605 ;
        RECT 116.965 198.315 117.135 198.775 ;
        RECT 118.070 198.655 118.240 199.035 ;
        RECT 119.460 198.865 119.630 199.455 ;
        RECT 120.370 199.335 120.580 199.985 ;
        RECT 117.370 198.315 118.240 198.655 ;
        RECT 118.830 198.695 119.630 198.865 ;
        RECT 118.410 198.145 118.660 198.605 ;
        RECT 118.830 198.405 119.000 198.695 ;
        RECT 119.180 198.145 119.510 198.525 ;
        RECT 119.850 198.145 120.155 199.285 ;
        RECT 120.325 198.455 120.580 199.335 ;
        RECT 120.755 199.955 121.140 200.525 ;
        RECT 121.310 200.235 121.635 200.695 ;
        RECT 122.155 200.065 122.435 200.525 ;
        RECT 120.755 199.285 121.035 199.955 ;
        RECT 121.310 199.895 122.435 200.065 ;
        RECT 121.310 199.785 121.760 199.895 ;
        RECT 121.205 199.455 121.760 199.785 ;
        RECT 122.625 199.725 123.025 200.525 ;
        RECT 123.425 200.235 123.695 200.695 ;
        RECT 123.865 200.065 124.150 200.525 ;
        RECT 120.755 198.315 121.140 199.285 ;
        RECT 121.310 198.995 121.760 199.455 ;
        RECT 121.930 199.165 123.025 199.725 ;
        RECT 121.310 198.775 122.435 198.995 ;
        RECT 121.310 198.145 121.635 198.605 ;
        RECT 122.155 198.315 122.435 198.775 ;
        RECT 122.625 198.315 123.025 199.165 ;
        RECT 123.195 199.895 124.150 200.065 ;
        RECT 123.195 198.995 123.405 199.895 ;
        RECT 124.475 199.875 124.705 200.695 ;
        RECT 124.875 199.895 125.205 200.525 ;
        RECT 123.575 199.165 124.265 199.725 ;
        RECT 124.455 199.455 124.785 199.705 ;
        RECT 124.955 199.295 125.205 199.895 ;
        RECT 125.375 199.875 125.585 200.695 ;
        RECT 125.815 199.925 129.325 200.695 ;
        RECT 129.955 199.945 131.165 200.695 ;
        RECT 125.815 199.405 127.465 199.925 ;
        RECT 123.195 198.775 124.150 198.995 ;
        RECT 123.425 198.145 123.695 198.605 ;
        RECT 123.865 198.315 124.150 198.775 ;
        RECT 124.475 198.145 124.705 199.285 ;
        RECT 124.875 198.315 125.205 199.295 ;
        RECT 125.375 198.145 125.585 199.285 ;
        RECT 127.635 199.235 129.325 199.755 ;
        RECT 125.815 198.145 129.325 199.235 ;
        RECT 129.955 199.235 130.475 199.775 ;
        RECT 130.645 199.405 131.165 199.945 ;
        RECT 129.955 198.145 131.165 199.235 ;
        RECT 57.190 197.975 131.250 198.145 ;
        RECT 57.275 196.885 58.485 197.975 ;
        RECT 58.655 197.540 64.000 197.975 ;
        RECT 64.175 197.540 69.520 197.975 ;
        RECT 57.275 196.175 57.795 196.715 ;
        RECT 57.965 196.345 58.485 196.885 ;
        RECT 57.275 195.425 58.485 196.175 ;
        RECT 60.240 195.970 60.580 196.800 ;
        RECT 62.060 196.290 62.410 197.540 ;
        RECT 65.760 195.970 66.100 196.800 ;
        RECT 67.580 196.290 67.930 197.540 ;
        RECT 70.155 196.810 70.445 197.975 ;
        RECT 70.615 196.885 74.125 197.975 ;
        RECT 74.295 196.885 75.505 197.975 ;
        RECT 75.685 197.255 76.015 197.975 ;
        RECT 70.615 196.195 72.265 196.715 ;
        RECT 72.435 196.365 74.125 196.885 ;
        RECT 58.655 195.425 64.000 195.970 ;
        RECT 64.175 195.425 69.520 195.970 ;
        RECT 70.155 195.425 70.445 196.150 ;
        RECT 70.615 195.425 74.125 196.195 ;
        RECT 74.295 196.175 74.815 196.715 ;
        RECT 74.985 196.345 75.505 196.885 ;
        RECT 75.675 196.615 75.905 196.955 ;
        RECT 76.195 196.615 76.410 197.730 ;
        RECT 76.605 197.030 76.935 197.805 ;
        RECT 77.105 197.200 77.815 197.975 ;
        RECT 76.605 196.815 77.755 197.030 ;
        RECT 75.675 196.415 76.005 196.615 ;
        RECT 76.195 196.435 76.645 196.615 ;
        RECT 76.315 196.415 76.645 196.435 ;
        RECT 76.815 196.415 77.285 196.645 ;
        RECT 77.470 196.245 77.755 196.815 ;
        RECT 77.985 196.370 78.265 197.805 ;
        RECT 78.435 196.885 81.945 197.975 ;
        RECT 74.295 195.425 75.505 196.175 ;
        RECT 75.675 196.055 76.855 196.245 ;
        RECT 75.675 195.595 76.015 196.055 ;
        RECT 76.525 195.975 76.855 196.055 ;
        RECT 77.045 196.055 77.755 196.245 ;
        RECT 77.045 195.915 77.345 196.055 ;
        RECT 77.030 195.905 77.345 195.915 ;
        RECT 77.020 195.895 77.345 195.905 ;
        RECT 77.010 195.890 77.345 195.895 ;
        RECT 76.185 195.425 76.355 195.885 ;
        RECT 77.005 195.880 77.345 195.890 ;
        RECT 77.000 195.875 77.345 195.880 ;
        RECT 76.995 195.865 77.345 195.875 ;
        RECT 76.990 195.860 77.345 195.865 ;
        RECT 76.985 195.595 77.345 195.860 ;
        RECT 77.585 195.425 77.755 195.885 ;
        RECT 77.925 195.595 78.265 196.370 ;
        RECT 78.435 196.195 80.085 196.715 ;
        RECT 80.255 196.365 81.945 196.885 ;
        RECT 82.575 197.135 82.835 197.805 ;
        RECT 83.005 197.575 83.335 197.975 ;
        RECT 84.205 197.575 84.605 197.975 ;
        RECT 84.895 197.395 85.225 197.630 ;
        RECT 83.145 197.225 85.225 197.395 ;
        RECT 78.435 195.425 81.945 196.195 ;
        RECT 82.575 196.165 82.750 197.135 ;
        RECT 83.145 196.955 83.315 197.225 ;
        RECT 82.920 196.785 83.315 196.955 ;
        RECT 83.485 196.835 84.500 197.055 ;
        RECT 82.920 196.335 83.090 196.785 ;
        RECT 84.225 196.695 84.500 196.835 ;
        RECT 84.670 196.835 85.225 197.225 ;
        RECT 83.260 196.415 83.710 196.615 ;
        RECT 83.880 196.245 84.055 196.440 ;
        RECT 82.575 195.595 82.915 196.165 ;
        RECT 83.110 195.425 83.280 196.090 ;
        RECT 83.560 196.075 84.055 196.245 ;
        RECT 83.560 195.935 83.780 196.075 ;
        RECT 83.555 195.765 83.780 195.935 ;
        RECT 84.225 195.905 84.395 196.695 ;
        RECT 84.670 196.585 84.840 196.835 ;
        RECT 85.395 196.665 85.570 197.765 ;
        RECT 85.740 197.155 86.085 197.975 ;
        RECT 87.185 197.365 87.515 197.795 ;
        RECT 87.695 197.535 87.890 197.975 ;
        RECT 88.060 197.365 88.390 197.795 ;
        RECT 87.185 197.195 88.390 197.365 ;
        RECT 84.645 196.415 84.840 196.585 ;
        RECT 85.010 196.415 85.570 196.665 ;
        RECT 85.740 196.415 86.085 196.985 ;
        RECT 87.185 196.865 88.080 197.195 ;
        RECT 88.560 197.025 88.835 197.795 ;
        RECT 89.590 197.345 89.875 197.805 ;
        RECT 90.045 197.515 90.315 197.975 ;
        RECT 89.590 197.125 90.545 197.345 ;
        RECT 88.250 196.835 88.835 197.025 ;
        RECT 84.645 196.030 84.815 196.415 ;
        RECT 87.190 196.335 87.485 196.665 ;
        RECT 87.665 196.335 88.080 196.665 ;
        RECT 83.560 195.720 83.780 195.765 ;
        RECT 83.950 195.735 84.395 195.905 ;
        RECT 84.565 195.660 84.815 196.030 ;
        RECT 84.985 196.065 86.085 196.245 ;
        RECT 84.985 195.660 85.235 196.065 ;
        RECT 85.405 195.425 85.575 195.895 ;
        RECT 85.745 195.660 86.085 196.065 ;
        RECT 87.185 195.425 87.485 196.155 ;
        RECT 87.665 195.715 87.895 196.335 ;
        RECT 88.250 196.165 88.425 196.835 ;
        RECT 88.095 195.985 88.425 196.165 ;
        RECT 88.595 196.015 88.835 196.665 ;
        RECT 89.475 196.395 90.165 196.955 ;
        RECT 90.335 196.225 90.545 197.125 ;
        RECT 89.590 196.055 90.545 196.225 ;
        RECT 90.715 196.955 91.115 197.805 ;
        RECT 91.305 197.345 91.585 197.805 ;
        RECT 92.105 197.515 92.430 197.975 ;
        RECT 91.305 197.125 92.430 197.345 ;
        RECT 90.715 196.395 91.810 196.955 ;
        RECT 91.980 196.665 92.430 197.125 ;
        RECT 92.600 196.835 92.985 197.805 ;
        RECT 93.155 196.835 93.435 197.975 ;
        RECT 88.095 195.605 88.320 195.985 ;
        RECT 88.490 195.425 88.820 195.815 ;
        RECT 89.590 195.595 89.875 196.055 ;
        RECT 90.045 195.425 90.315 195.885 ;
        RECT 90.715 195.595 91.115 196.395 ;
        RECT 91.980 196.335 92.535 196.665 ;
        RECT 91.980 196.225 92.430 196.335 ;
        RECT 91.305 196.055 92.430 196.225 ;
        RECT 92.705 196.165 92.985 196.835 ;
        RECT 93.605 196.825 93.935 197.805 ;
        RECT 94.105 196.835 94.365 197.975 ;
        RECT 94.535 196.885 95.745 197.975 ;
        RECT 93.670 196.785 93.845 196.825 ;
        RECT 93.165 196.395 93.500 196.665 ;
        RECT 93.670 196.225 93.840 196.785 ;
        RECT 94.010 196.415 94.345 196.665 ;
        RECT 91.305 195.595 91.585 196.055 ;
        RECT 92.105 195.425 92.430 195.885 ;
        RECT 92.600 195.595 92.985 196.165 ;
        RECT 93.155 195.425 93.465 196.225 ;
        RECT 93.670 195.595 94.365 196.225 ;
        RECT 94.535 196.175 95.055 196.715 ;
        RECT 95.225 196.345 95.745 196.885 ;
        RECT 95.915 196.810 96.205 197.975 ;
        RECT 96.375 196.820 96.715 197.805 ;
        RECT 96.885 197.545 97.295 197.975 ;
        RECT 98.040 197.555 98.370 197.975 ;
        RECT 98.540 197.375 98.865 197.805 ;
        RECT 96.885 197.205 98.865 197.375 ;
        RECT 94.535 195.425 95.745 196.175 ;
        RECT 96.375 196.165 96.630 196.820 ;
        RECT 96.885 196.665 97.150 197.205 ;
        RECT 97.365 196.865 97.990 197.035 ;
        RECT 96.800 196.335 97.150 196.665 ;
        RECT 97.320 196.335 97.650 196.665 ;
        RECT 97.820 196.165 97.990 196.865 ;
        RECT 95.915 195.425 96.205 196.150 ;
        RECT 96.375 195.790 96.735 196.165 ;
        RECT 97.000 195.425 97.170 196.165 ;
        RECT 97.450 195.995 97.990 196.165 ;
        RECT 98.160 196.795 98.865 197.205 ;
        RECT 99.340 196.875 99.670 197.975 ;
        RECT 100.060 197.025 100.325 197.795 ;
        RECT 100.495 197.255 100.825 197.975 ;
        RECT 101.015 197.435 101.275 197.795 ;
        RECT 101.445 197.605 101.775 197.975 ;
        RECT 101.945 197.435 102.205 197.795 ;
        RECT 101.015 197.205 102.205 197.435 ;
        RECT 102.775 197.025 103.065 197.795 ;
        RECT 97.450 195.790 97.620 195.995 ;
        RECT 98.160 195.595 98.330 196.795 ;
        RECT 98.500 196.415 99.070 196.625 ;
        RECT 99.240 196.415 99.885 196.625 ;
        RECT 98.560 196.075 99.730 196.245 ;
        RECT 98.560 195.595 98.890 196.075 ;
        RECT 99.060 195.425 99.230 195.895 ;
        RECT 99.400 195.610 99.730 196.075 ;
        RECT 100.060 195.605 100.395 197.025 ;
        RECT 100.570 196.845 103.065 197.025 ;
        RECT 103.275 196.885 104.485 197.975 ;
        RECT 104.745 197.230 105.015 197.975 ;
        RECT 105.645 197.970 111.920 197.975 ;
        RECT 105.185 197.060 105.475 197.800 ;
        RECT 105.645 197.245 105.900 197.970 ;
        RECT 106.085 197.075 106.345 197.800 ;
        RECT 106.515 197.245 106.760 197.970 ;
        RECT 106.945 197.075 107.205 197.800 ;
        RECT 107.375 197.245 107.620 197.970 ;
        RECT 107.805 197.075 108.065 197.800 ;
        RECT 108.235 197.245 108.480 197.970 ;
        RECT 108.650 197.075 108.910 197.800 ;
        RECT 109.080 197.245 109.340 197.970 ;
        RECT 109.510 197.075 109.770 197.800 ;
        RECT 109.940 197.245 110.200 197.970 ;
        RECT 110.370 197.075 110.630 197.800 ;
        RECT 110.800 197.245 111.060 197.970 ;
        RECT 111.230 197.075 111.490 197.800 ;
        RECT 111.660 197.175 111.920 197.970 ;
        RECT 106.085 197.060 111.490 197.075 ;
        RECT 100.570 196.155 100.795 196.845 ;
        RECT 100.995 196.335 101.275 196.665 ;
        RECT 101.455 196.335 102.030 196.665 ;
        RECT 102.210 196.335 102.645 196.665 ;
        RECT 102.825 196.335 103.095 196.665 ;
        RECT 103.275 196.175 103.795 196.715 ;
        RECT 103.965 196.345 104.485 196.885 ;
        RECT 104.745 196.835 111.490 197.060 ;
        RECT 104.745 196.245 105.910 196.835 ;
        RECT 112.090 196.665 112.340 197.800 ;
        RECT 112.520 197.165 112.780 197.975 ;
        RECT 112.955 196.665 113.200 197.805 ;
        RECT 113.380 197.165 113.675 197.975 ;
        RECT 113.860 196.835 114.195 197.805 ;
        RECT 114.365 196.835 114.535 197.975 ;
        RECT 114.705 197.635 116.735 197.805 ;
        RECT 106.080 196.415 113.200 196.665 ;
        RECT 100.570 195.965 103.055 196.155 ;
        RECT 100.575 195.425 101.320 195.795 ;
        RECT 101.885 195.605 102.140 195.965 ;
        RECT 102.320 195.425 102.650 195.795 ;
        RECT 102.830 195.605 103.055 195.965 ;
        RECT 103.275 195.425 104.485 196.175 ;
        RECT 104.745 196.075 111.490 196.245 ;
        RECT 104.745 195.425 105.045 195.905 ;
        RECT 105.215 195.620 105.475 196.075 ;
        RECT 105.645 195.425 105.905 195.905 ;
        RECT 106.085 195.620 106.345 196.075 ;
        RECT 106.515 195.425 106.765 195.905 ;
        RECT 106.945 195.620 107.205 196.075 ;
        RECT 107.375 195.425 107.625 195.905 ;
        RECT 107.805 195.620 108.065 196.075 ;
        RECT 108.235 195.425 108.480 195.905 ;
        RECT 108.650 195.620 108.925 196.075 ;
        RECT 109.095 195.425 109.340 195.905 ;
        RECT 109.510 195.620 109.770 196.075 ;
        RECT 109.940 195.425 110.200 195.905 ;
        RECT 110.370 195.620 110.630 196.075 ;
        RECT 110.800 195.425 111.060 195.905 ;
        RECT 111.230 195.620 111.490 196.075 ;
        RECT 111.660 195.425 111.920 195.985 ;
        RECT 112.090 195.605 112.340 196.415 ;
        RECT 112.520 195.425 112.780 195.950 ;
        RECT 112.950 195.605 113.200 196.415 ;
        RECT 113.370 196.105 113.685 196.665 ;
        RECT 113.860 196.165 114.030 196.835 ;
        RECT 114.705 196.665 114.875 197.635 ;
        RECT 114.200 196.335 114.455 196.665 ;
        RECT 114.680 196.335 114.875 196.665 ;
        RECT 115.045 197.295 116.170 197.465 ;
        RECT 114.285 196.165 114.455 196.335 ;
        RECT 115.045 196.165 115.215 197.295 ;
        RECT 113.380 195.425 113.685 195.935 ;
        RECT 113.860 195.595 114.115 196.165 ;
        RECT 114.285 195.995 115.215 196.165 ;
        RECT 115.385 196.955 116.395 197.125 ;
        RECT 115.385 196.155 115.555 196.955 ;
        RECT 115.040 195.960 115.215 195.995 ;
        RECT 114.285 195.425 114.615 195.825 ;
        RECT 115.040 195.595 115.570 195.960 ;
        RECT 115.760 195.935 116.035 196.755 ;
        RECT 115.755 195.765 116.035 195.935 ;
        RECT 115.760 195.595 116.035 195.765 ;
        RECT 116.205 195.595 116.395 196.955 ;
        RECT 116.565 196.970 116.735 197.635 ;
        RECT 116.905 197.215 117.075 197.975 ;
        RECT 117.310 197.215 117.825 197.625 ;
        RECT 118.000 197.465 119.655 197.755 ;
        RECT 116.565 196.780 117.315 196.970 ;
        RECT 117.485 196.405 117.825 197.215 ;
        RECT 118.000 197.125 119.590 197.295 ;
        RECT 119.825 197.175 120.105 197.975 ;
        RECT 118.000 196.835 118.320 197.125 ;
        RECT 119.420 197.005 119.590 197.125 ;
        RECT 116.595 196.235 117.825 196.405 ;
        RECT 116.575 195.425 117.085 195.960 ;
        RECT 117.305 195.630 117.550 196.235 ;
        RECT 118.000 196.095 118.350 196.665 ;
        RECT 118.520 196.335 119.230 196.955 ;
        RECT 119.420 196.835 120.145 197.005 ;
        RECT 120.315 196.835 120.585 197.805 ;
        RECT 119.975 196.665 120.145 196.835 ;
        RECT 119.400 196.335 119.805 196.665 ;
        RECT 119.975 196.335 120.245 196.665 ;
        RECT 119.975 196.165 120.145 196.335 ;
        RECT 118.535 195.995 120.145 196.165 ;
        RECT 120.415 196.100 120.585 196.835 ;
        RECT 121.675 196.810 121.965 197.975 ;
        RECT 122.135 196.900 122.405 197.805 ;
        RECT 122.575 197.215 122.905 197.975 ;
        RECT 123.085 197.045 123.255 197.805 ;
        RECT 123.515 197.540 128.860 197.975 ;
        RECT 118.005 195.425 118.335 195.925 ;
        RECT 118.535 195.645 118.705 195.995 ;
        RECT 118.905 195.425 119.235 195.825 ;
        RECT 119.405 195.645 119.575 195.995 ;
        RECT 119.745 195.425 120.125 195.825 ;
        RECT 120.315 195.755 120.585 196.100 ;
        RECT 121.675 195.425 121.965 196.150 ;
        RECT 122.135 196.100 122.305 196.900 ;
        RECT 122.590 196.875 123.255 197.045 ;
        RECT 122.590 196.730 122.760 196.875 ;
        RECT 122.475 196.400 122.760 196.730 ;
        RECT 122.590 196.145 122.760 196.400 ;
        RECT 122.995 196.325 123.325 196.695 ;
        RECT 122.135 195.595 122.395 196.100 ;
        RECT 122.590 195.975 123.255 196.145 ;
        RECT 122.575 195.425 122.905 195.805 ;
        RECT 123.085 195.595 123.255 195.975 ;
        RECT 125.100 195.970 125.440 196.800 ;
        RECT 126.920 196.290 127.270 197.540 ;
        RECT 129.955 196.885 131.165 197.975 ;
        RECT 129.955 196.345 130.475 196.885 ;
        RECT 130.645 196.175 131.165 196.715 ;
        RECT 123.515 195.425 128.860 195.970 ;
        RECT 129.955 195.425 131.165 196.175 ;
        RECT 57.190 195.255 131.250 195.425 ;
        RECT 57.275 194.505 58.485 195.255 ;
        RECT 58.655 194.710 64.000 195.255 ;
        RECT 64.175 194.710 69.520 195.255 ;
        RECT 69.695 194.710 75.040 195.255 ;
        RECT 57.275 193.965 57.795 194.505 ;
        RECT 57.965 193.795 58.485 194.335 ;
        RECT 60.240 193.880 60.580 194.710 ;
        RECT 57.275 192.705 58.485 193.795 ;
        RECT 62.060 193.140 62.410 194.390 ;
        RECT 65.760 193.880 66.100 194.710 ;
        RECT 67.580 193.140 67.930 194.390 ;
        RECT 71.280 193.880 71.620 194.710 ;
        RECT 75.215 194.485 77.805 195.255 ;
        RECT 77.980 194.515 78.235 195.085 ;
        RECT 78.405 194.855 78.735 195.255 ;
        RECT 79.160 194.720 79.690 195.085 ;
        RECT 79.160 194.685 79.335 194.720 ;
        RECT 78.405 194.515 79.335 194.685 ;
        RECT 73.100 193.140 73.450 194.390 ;
        RECT 75.215 193.965 76.425 194.485 ;
        RECT 76.595 193.795 77.805 194.315 ;
        RECT 58.655 192.705 64.000 193.140 ;
        RECT 64.175 192.705 69.520 193.140 ;
        RECT 69.695 192.705 75.040 193.140 ;
        RECT 75.215 192.705 77.805 193.795 ;
        RECT 77.980 193.845 78.150 194.515 ;
        RECT 78.405 194.345 78.575 194.515 ;
        RECT 78.320 194.015 78.575 194.345 ;
        RECT 78.800 194.015 78.995 194.345 ;
        RECT 77.980 192.875 78.315 193.845 ;
        RECT 78.485 192.705 78.655 193.845 ;
        RECT 78.825 193.045 78.995 194.015 ;
        RECT 79.165 193.385 79.335 194.515 ;
        RECT 79.505 193.725 79.675 194.525 ;
        RECT 79.880 194.235 80.155 195.085 ;
        RECT 79.875 194.065 80.155 194.235 ;
        RECT 79.880 193.925 80.155 194.065 ;
        RECT 80.325 193.725 80.515 195.085 ;
        RECT 80.695 194.720 81.205 195.255 ;
        RECT 81.425 194.445 81.670 195.050 ;
        RECT 83.035 194.530 83.325 195.255 ;
        RECT 83.585 194.775 83.885 195.255 ;
        RECT 84.055 194.605 84.315 195.060 ;
        RECT 84.485 194.775 84.745 195.255 ;
        RECT 84.925 194.605 85.185 195.060 ;
        RECT 85.355 194.775 85.605 195.255 ;
        RECT 85.785 194.605 86.045 195.060 ;
        RECT 86.215 194.775 86.465 195.255 ;
        RECT 86.645 194.605 86.905 195.060 ;
        RECT 87.075 194.775 87.320 195.255 ;
        RECT 87.490 194.605 87.765 195.060 ;
        RECT 87.935 194.775 88.180 195.255 ;
        RECT 88.350 194.605 88.610 195.060 ;
        RECT 88.780 194.775 89.040 195.255 ;
        RECT 89.210 194.605 89.470 195.060 ;
        RECT 89.640 194.775 89.900 195.255 ;
        RECT 90.070 194.605 90.330 195.060 ;
        RECT 90.500 194.695 90.760 195.255 ;
        RECT 80.715 194.275 81.945 194.445 ;
        RECT 79.505 193.555 80.515 193.725 ;
        RECT 80.685 193.710 81.435 193.900 ;
        RECT 79.165 193.215 80.290 193.385 ;
        RECT 80.685 193.045 80.855 193.710 ;
        RECT 81.605 193.465 81.945 194.275 ;
        RECT 83.585 194.435 90.330 194.605 ;
        RECT 78.825 192.875 80.855 193.045 ;
        RECT 81.025 192.705 81.195 193.465 ;
        RECT 81.430 193.055 81.945 193.465 ;
        RECT 83.035 192.705 83.325 193.870 ;
        RECT 83.585 193.845 84.750 194.435 ;
        RECT 90.930 194.265 91.180 195.075 ;
        RECT 91.360 194.730 91.620 195.255 ;
        RECT 91.790 194.265 92.040 195.075 ;
        RECT 92.220 194.745 92.525 195.255 ;
        RECT 92.785 194.705 92.955 195.085 ;
        RECT 93.135 194.875 93.465 195.255 ;
        RECT 84.920 194.015 92.040 194.265 ;
        RECT 92.210 194.015 92.525 194.575 ;
        RECT 92.785 194.535 93.450 194.705 ;
        RECT 93.645 194.580 93.905 195.085 ;
        RECT 94.075 194.710 99.420 195.255 ;
        RECT 83.585 193.620 90.330 193.845 ;
        RECT 83.585 192.705 83.855 193.450 ;
        RECT 84.025 192.880 84.315 193.620 ;
        RECT 84.925 193.605 90.330 193.620 ;
        RECT 84.485 192.710 84.740 193.435 ;
        RECT 84.925 192.880 85.185 193.605 ;
        RECT 85.355 192.710 85.600 193.435 ;
        RECT 85.785 192.880 86.045 193.605 ;
        RECT 86.215 192.710 86.460 193.435 ;
        RECT 86.645 192.880 86.905 193.605 ;
        RECT 87.075 192.710 87.320 193.435 ;
        RECT 87.490 192.880 87.750 193.605 ;
        RECT 87.920 192.710 88.180 193.435 ;
        RECT 88.350 192.880 88.610 193.605 ;
        RECT 88.780 192.710 89.040 193.435 ;
        RECT 89.210 192.880 89.470 193.605 ;
        RECT 89.640 192.710 89.900 193.435 ;
        RECT 90.070 192.880 90.330 193.605 ;
        RECT 90.500 192.710 90.760 193.505 ;
        RECT 90.930 192.880 91.180 194.015 ;
        RECT 84.485 192.705 90.760 192.710 ;
        RECT 91.360 192.705 91.620 193.515 ;
        RECT 91.795 192.875 92.040 194.015 ;
        RECT 92.715 193.985 93.045 194.355 ;
        RECT 93.280 194.280 93.450 194.535 ;
        RECT 93.280 193.950 93.565 194.280 ;
        RECT 93.280 193.805 93.450 193.950 ;
        RECT 92.785 193.635 93.450 193.805 ;
        RECT 93.735 193.780 93.905 194.580 ;
        RECT 95.660 193.880 96.000 194.710 ;
        RECT 99.595 194.485 103.105 195.255 ;
        RECT 104.395 194.625 104.725 194.985 ;
        RECT 105.345 194.795 105.595 195.255 ;
        RECT 105.765 194.795 106.325 195.085 ;
        RECT 92.220 192.705 92.515 193.515 ;
        RECT 92.785 192.875 92.955 193.635 ;
        RECT 93.135 192.705 93.465 193.465 ;
        RECT 93.635 192.875 93.905 193.780 ;
        RECT 97.480 193.140 97.830 194.390 ;
        RECT 99.595 193.965 101.245 194.485 ;
        RECT 104.395 194.435 105.785 194.625 ;
        RECT 105.615 194.345 105.785 194.435 ;
        RECT 101.415 193.795 103.105 194.315 ;
        RECT 94.075 192.705 99.420 193.140 ;
        RECT 99.595 192.705 103.105 193.795 ;
        RECT 104.210 194.015 104.885 194.265 ;
        RECT 105.105 194.015 105.445 194.265 ;
        RECT 105.615 194.015 105.905 194.345 ;
        RECT 104.210 193.655 104.475 194.015 ;
        RECT 105.615 193.765 105.785 194.015 ;
        RECT 104.845 193.595 105.785 193.765 ;
        RECT 104.395 192.705 104.675 193.375 ;
        RECT 104.845 193.045 105.145 193.595 ;
        RECT 106.075 193.425 106.325 194.795 ;
        RECT 106.515 194.445 106.755 195.255 ;
        RECT 106.925 194.445 107.255 195.085 ;
        RECT 107.425 194.445 107.695 195.255 ;
        RECT 108.795 194.530 109.085 195.255 ;
        RECT 109.255 194.745 109.560 195.255 ;
        RECT 106.495 194.015 106.845 194.265 ;
        RECT 107.015 193.845 107.185 194.445 ;
        RECT 107.355 194.015 107.705 194.265 ;
        RECT 109.255 194.015 109.570 194.575 ;
        RECT 109.740 194.265 109.990 195.075 ;
        RECT 110.160 194.730 110.420 195.255 ;
        RECT 110.600 194.265 110.850 195.075 ;
        RECT 111.020 194.695 111.280 195.255 ;
        RECT 111.450 194.605 111.710 195.060 ;
        RECT 111.880 194.775 112.140 195.255 ;
        RECT 112.310 194.605 112.570 195.060 ;
        RECT 112.740 194.775 113.000 195.255 ;
        RECT 113.170 194.605 113.430 195.060 ;
        RECT 113.600 194.775 113.845 195.255 ;
        RECT 114.015 194.605 114.290 195.060 ;
        RECT 114.460 194.775 114.705 195.255 ;
        RECT 114.875 194.605 115.135 195.060 ;
        RECT 115.315 194.775 115.565 195.255 ;
        RECT 115.735 194.605 115.995 195.060 ;
        RECT 116.175 194.775 116.425 195.255 ;
        RECT 116.595 194.605 116.855 195.060 ;
        RECT 117.035 194.775 117.295 195.255 ;
        RECT 117.465 194.605 117.725 195.060 ;
        RECT 117.895 194.775 118.195 195.255 ;
        RECT 118.455 194.710 123.800 195.255 ;
        RECT 123.975 194.710 129.320 195.255 ;
        RECT 111.450 194.435 118.195 194.605 ;
        RECT 109.740 194.015 116.860 194.265 ;
        RECT 105.345 192.705 105.675 193.425 ;
        RECT 105.865 192.875 106.325 193.425 ;
        RECT 106.505 193.675 107.185 193.845 ;
        RECT 106.505 192.890 106.835 193.675 ;
        RECT 107.365 192.705 107.695 193.845 ;
        RECT 108.795 192.705 109.085 193.870 ;
        RECT 109.265 192.705 109.560 193.515 ;
        RECT 109.740 192.875 109.985 194.015 ;
        RECT 110.160 192.705 110.420 193.515 ;
        RECT 110.600 192.880 110.850 194.015 ;
        RECT 117.030 193.845 118.195 194.435 ;
        RECT 120.040 193.880 120.380 194.710 ;
        RECT 111.450 193.620 118.195 193.845 ;
        RECT 111.450 193.605 116.855 193.620 ;
        RECT 111.020 192.710 111.280 193.505 ;
        RECT 111.450 192.880 111.710 193.605 ;
        RECT 111.880 192.710 112.140 193.435 ;
        RECT 112.310 192.880 112.570 193.605 ;
        RECT 112.740 192.710 113.000 193.435 ;
        RECT 113.170 192.880 113.430 193.605 ;
        RECT 113.600 192.710 113.860 193.435 ;
        RECT 114.030 192.880 114.290 193.605 ;
        RECT 114.460 192.710 114.705 193.435 ;
        RECT 114.875 192.880 115.135 193.605 ;
        RECT 115.320 192.710 115.565 193.435 ;
        RECT 115.735 192.880 115.995 193.605 ;
        RECT 116.180 192.710 116.425 193.435 ;
        RECT 116.595 192.880 116.855 193.605 ;
        RECT 117.040 192.710 117.295 193.435 ;
        RECT 117.465 192.880 117.755 193.620 ;
        RECT 111.020 192.705 117.295 192.710 ;
        RECT 117.925 192.705 118.195 193.450 ;
        RECT 121.860 193.140 122.210 194.390 ;
        RECT 125.560 193.880 125.900 194.710 ;
        RECT 129.955 194.505 131.165 195.255 ;
        RECT 127.380 193.140 127.730 194.390 ;
        RECT 129.955 193.795 130.475 194.335 ;
        RECT 130.645 193.965 131.165 194.505 ;
        RECT 118.455 192.705 123.800 193.140 ;
        RECT 123.975 192.705 129.320 193.140 ;
        RECT 129.955 192.705 131.165 193.795 ;
        RECT 57.190 192.535 131.250 192.705 ;
        RECT 57.275 191.445 58.485 192.535 ;
        RECT 58.655 192.100 64.000 192.535 ;
        RECT 64.175 192.100 69.520 192.535 ;
        RECT 57.275 190.735 57.795 191.275 ;
        RECT 57.965 190.905 58.485 191.445 ;
        RECT 57.275 189.985 58.485 190.735 ;
        RECT 60.240 190.530 60.580 191.360 ;
        RECT 62.060 190.850 62.410 192.100 ;
        RECT 65.760 190.530 66.100 191.360 ;
        RECT 67.580 190.850 67.930 192.100 ;
        RECT 70.155 191.370 70.445 192.535 ;
        RECT 70.615 192.100 75.960 192.535 ;
        RECT 58.655 189.985 64.000 190.530 ;
        RECT 64.175 189.985 69.520 190.530 ;
        RECT 70.155 189.985 70.445 190.710 ;
        RECT 72.200 190.530 72.540 191.360 ;
        RECT 74.020 190.850 74.370 192.100 ;
        RECT 76.135 191.445 77.805 192.535 ;
        RECT 76.135 190.755 76.885 191.275 ;
        RECT 77.055 190.925 77.805 191.445 ;
        RECT 78.435 191.435 78.755 192.365 ;
        RECT 78.935 191.855 79.335 192.365 ;
        RECT 79.505 192.025 79.675 192.535 ;
        RECT 79.845 191.855 80.175 192.365 ;
        RECT 78.935 191.685 80.175 191.855 ;
        RECT 80.345 191.685 80.515 192.535 ;
        RECT 81.105 191.685 81.485 192.365 ;
        RECT 78.435 191.265 79.065 191.435 ;
        RECT 70.615 189.985 75.960 190.530 ;
        RECT 76.135 189.985 77.805 190.755 ;
        RECT 78.435 189.985 78.725 190.820 ;
        RECT 78.895 190.385 79.065 191.265 ;
        RECT 79.840 191.345 81.145 191.515 ;
        RECT 79.235 190.725 79.465 191.225 ;
        RECT 79.840 191.145 80.010 191.345 ;
        RECT 79.635 190.975 80.010 191.145 ;
        RECT 80.180 190.975 80.730 191.175 ;
        RECT 80.900 190.895 81.145 191.345 ;
        RECT 81.315 190.725 81.485 191.685 ;
        RECT 79.235 190.555 81.485 190.725 ;
        RECT 81.655 191.395 81.925 192.365 ;
        RECT 82.135 191.735 82.415 192.535 ;
        RECT 82.595 191.985 83.790 192.315 ;
        RECT 82.920 191.565 83.340 191.815 ;
        RECT 82.095 191.395 83.340 191.565 ;
        RECT 81.655 190.660 81.825 191.395 ;
        RECT 82.095 191.225 82.265 191.395 ;
        RECT 83.565 191.225 83.735 191.785 ;
        RECT 83.985 191.395 84.240 192.535 ;
        RECT 84.415 191.445 85.625 192.535 ;
        RECT 82.035 190.895 82.265 191.225 ;
        RECT 82.995 190.895 83.735 191.225 ;
        RECT 83.905 190.975 84.240 191.225 ;
        RECT 82.095 190.725 82.265 190.895 ;
        RECT 83.485 190.805 83.735 190.895 ;
        RECT 78.895 190.215 79.850 190.385 ;
        RECT 80.265 189.985 80.595 190.375 ;
        RECT 80.765 190.235 80.935 190.555 ;
        RECT 81.105 189.985 81.435 190.375 ;
        RECT 81.655 190.315 81.925 190.660 ;
        RECT 82.095 190.555 82.835 190.725 ;
        RECT 83.485 190.635 84.220 190.805 ;
        RECT 82.115 189.985 82.495 190.385 ;
        RECT 82.665 190.205 82.835 190.555 ;
        RECT 83.005 189.985 83.740 190.465 ;
        RECT 83.910 190.165 84.220 190.635 ;
        RECT 84.415 190.735 84.935 191.275 ;
        RECT 85.105 190.905 85.625 191.445 ;
        RECT 85.980 191.565 86.370 191.740 ;
        RECT 86.855 191.735 87.185 192.535 ;
        RECT 87.355 191.745 87.890 192.365 ;
        RECT 85.980 191.395 87.405 191.565 ;
        RECT 84.415 189.985 85.625 190.735 ;
        RECT 85.855 190.665 86.210 191.225 ;
        RECT 86.380 190.495 86.550 191.395 ;
        RECT 86.720 190.665 86.985 191.225 ;
        RECT 87.235 190.895 87.405 191.395 ;
        RECT 87.575 190.725 87.890 191.745 ;
        RECT 88.155 191.475 88.485 192.320 ;
        RECT 88.655 191.525 88.825 192.535 ;
        RECT 88.995 191.805 89.335 192.365 ;
        RECT 89.565 192.035 89.880 192.535 ;
        RECT 90.060 192.065 90.945 192.235 ;
        RECT 85.960 189.985 86.200 190.495 ;
        RECT 86.380 190.165 86.660 190.495 ;
        RECT 86.890 189.985 87.105 190.495 ;
        RECT 87.275 190.155 87.890 190.725 ;
        RECT 88.095 191.395 88.485 191.475 ;
        RECT 88.995 191.430 89.890 191.805 ;
        RECT 88.095 191.345 88.310 191.395 ;
        RECT 88.095 190.765 88.265 191.345 ;
        RECT 88.995 191.225 89.185 191.430 ;
        RECT 90.060 191.225 90.230 192.065 ;
        RECT 91.170 192.035 91.420 192.365 ;
        RECT 88.435 190.895 89.185 191.225 ;
        RECT 89.355 190.895 90.230 191.225 ;
        RECT 88.095 190.725 88.320 190.765 ;
        RECT 88.985 190.725 89.185 190.895 ;
        RECT 88.095 190.640 88.475 190.725 ;
        RECT 88.145 190.205 88.475 190.640 ;
        RECT 88.645 189.985 88.815 190.595 ;
        RECT 88.985 190.200 89.315 190.725 ;
        RECT 89.575 189.985 89.785 190.515 ;
        RECT 90.060 190.435 90.230 190.895 ;
        RECT 90.400 190.935 90.720 191.895 ;
        RECT 90.890 191.145 91.080 191.865 ;
        RECT 91.250 190.965 91.420 192.035 ;
        RECT 91.590 191.735 91.760 192.535 ;
        RECT 91.930 192.090 93.035 192.260 ;
        RECT 91.930 191.475 92.100 192.090 ;
        RECT 93.245 191.940 93.495 192.365 ;
        RECT 93.665 192.075 93.930 192.535 ;
        RECT 92.270 191.555 92.800 191.920 ;
        RECT 93.245 191.810 93.550 191.940 ;
        RECT 91.590 191.385 92.100 191.475 ;
        RECT 91.590 191.215 92.460 191.385 ;
        RECT 91.590 191.145 91.760 191.215 ;
        RECT 91.880 190.965 92.080 190.995 ;
        RECT 90.400 190.605 90.865 190.935 ;
        RECT 91.250 190.665 92.080 190.965 ;
        RECT 91.250 190.435 91.420 190.665 ;
        RECT 90.060 190.265 90.845 190.435 ;
        RECT 91.015 190.265 91.420 190.435 ;
        RECT 91.600 189.985 91.970 190.485 ;
        RECT 92.290 190.435 92.460 191.215 ;
        RECT 92.630 190.855 92.800 191.555 ;
        RECT 92.970 191.025 93.210 191.620 ;
        RECT 92.630 190.635 93.155 190.855 ;
        RECT 93.380 190.705 93.550 191.810 ;
        RECT 93.325 190.575 93.550 190.705 ;
        RECT 93.720 190.615 94.000 191.565 ;
        RECT 93.325 190.435 93.495 190.575 ;
        RECT 92.290 190.265 92.965 190.435 ;
        RECT 93.160 190.265 93.495 190.435 ;
        RECT 93.665 189.985 93.915 190.445 ;
        RECT 94.170 190.245 94.355 192.365 ;
        RECT 94.525 192.035 94.855 192.535 ;
        RECT 95.025 191.865 95.195 192.365 ;
        RECT 94.530 191.695 95.195 191.865 ;
        RECT 94.530 190.705 94.760 191.695 ;
        RECT 94.930 190.875 95.280 191.525 ;
        RECT 95.915 191.370 96.205 192.535 ;
        RECT 96.435 191.475 96.765 192.320 ;
        RECT 96.935 191.525 97.105 192.535 ;
        RECT 97.275 191.805 97.615 192.365 ;
        RECT 97.845 192.035 98.160 192.535 ;
        RECT 98.340 192.065 99.225 192.235 ;
        RECT 96.375 191.395 96.765 191.475 ;
        RECT 97.275 191.430 98.170 191.805 ;
        RECT 96.375 191.345 96.590 191.395 ;
        RECT 96.375 190.765 96.545 191.345 ;
        RECT 97.275 191.225 97.465 191.430 ;
        RECT 98.340 191.225 98.510 192.065 ;
        RECT 99.450 192.035 99.700 192.365 ;
        RECT 96.715 190.895 97.465 191.225 ;
        RECT 97.635 190.895 98.510 191.225 ;
        RECT 96.375 190.725 96.600 190.765 ;
        RECT 97.265 190.725 97.465 190.895 ;
        RECT 94.530 190.535 95.195 190.705 ;
        RECT 94.525 189.985 94.855 190.365 ;
        RECT 95.025 190.245 95.195 190.535 ;
        RECT 95.915 189.985 96.205 190.710 ;
        RECT 96.375 190.640 96.755 190.725 ;
        RECT 96.425 190.205 96.755 190.640 ;
        RECT 96.925 189.985 97.095 190.595 ;
        RECT 97.265 190.200 97.595 190.725 ;
        RECT 97.855 189.985 98.065 190.515 ;
        RECT 98.340 190.435 98.510 190.895 ;
        RECT 98.680 190.935 99.000 191.895 ;
        RECT 99.170 191.145 99.360 191.865 ;
        RECT 99.530 190.965 99.700 192.035 ;
        RECT 99.870 191.735 100.040 192.535 ;
        RECT 100.210 192.090 101.315 192.260 ;
        RECT 100.210 191.475 100.380 192.090 ;
        RECT 101.525 191.940 101.775 192.365 ;
        RECT 101.945 192.075 102.210 192.535 ;
        RECT 100.550 191.555 101.080 191.920 ;
        RECT 101.525 191.810 101.830 191.940 ;
        RECT 99.870 191.385 100.380 191.475 ;
        RECT 99.870 191.215 100.740 191.385 ;
        RECT 99.870 191.145 100.040 191.215 ;
        RECT 100.160 190.965 100.360 190.995 ;
        RECT 98.680 190.605 99.145 190.935 ;
        RECT 99.530 190.665 100.360 190.965 ;
        RECT 99.530 190.435 99.700 190.665 ;
        RECT 98.340 190.265 99.125 190.435 ;
        RECT 99.295 190.265 99.700 190.435 ;
        RECT 99.880 189.985 100.250 190.485 ;
        RECT 100.570 190.435 100.740 191.215 ;
        RECT 100.910 190.855 101.080 191.555 ;
        RECT 101.250 191.025 101.490 191.620 ;
        RECT 100.910 190.635 101.435 190.855 ;
        RECT 101.660 190.705 101.830 191.810 ;
        RECT 101.605 190.575 101.830 190.705 ;
        RECT 102.000 190.615 102.280 191.565 ;
        RECT 101.605 190.435 101.775 190.575 ;
        RECT 100.570 190.265 101.245 190.435 ;
        RECT 101.440 190.265 101.775 190.435 ;
        RECT 101.945 189.985 102.195 190.445 ;
        RECT 102.450 190.245 102.635 192.365 ;
        RECT 102.805 192.035 103.135 192.535 ;
        RECT 103.305 191.865 103.475 192.365 ;
        RECT 103.735 192.100 109.080 192.535 ;
        RECT 102.810 191.695 103.475 191.865 ;
        RECT 102.810 190.705 103.040 191.695 ;
        RECT 103.210 190.875 103.560 191.525 ;
        RECT 102.810 190.535 103.475 190.705 ;
        RECT 102.805 189.985 103.135 190.365 ;
        RECT 103.305 190.245 103.475 190.535 ;
        RECT 105.320 190.530 105.660 191.360 ;
        RECT 107.140 190.850 107.490 192.100 ;
        RECT 109.315 191.475 109.645 192.320 ;
        RECT 109.815 191.525 109.985 192.535 ;
        RECT 110.155 191.805 110.495 192.365 ;
        RECT 110.725 192.035 111.040 192.535 ;
        RECT 111.220 192.065 112.105 192.235 ;
        RECT 109.255 191.395 109.645 191.475 ;
        RECT 110.155 191.430 111.050 191.805 ;
        RECT 109.255 191.345 109.470 191.395 ;
        RECT 109.255 190.765 109.425 191.345 ;
        RECT 110.155 191.225 110.345 191.430 ;
        RECT 111.220 191.225 111.390 192.065 ;
        RECT 112.330 192.035 112.580 192.365 ;
        RECT 109.595 190.895 110.345 191.225 ;
        RECT 110.515 190.895 111.390 191.225 ;
        RECT 109.255 190.725 109.480 190.765 ;
        RECT 110.145 190.725 110.345 190.895 ;
        RECT 109.255 190.640 109.635 190.725 ;
        RECT 103.735 189.985 109.080 190.530 ;
        RECT 109.305 190.205 109.635 190.640 ;
        RECT 109.805 189.985 109.975 190.595 ;
        RECT 110.145 190.200 110.475 190.725 ;
        RECT 110.735 189.985 110.945 190.515 ;
        RECT 111.220 190.435 111.390 190.895 ;
        RECT 111.560 190.935 111.880 191.895 ;
        RECT 112.050 191.145 112.240 191.865 ;
        RECT 112.410 190.965 112.580 192.035 ;
        RECT 112.750 191.735 112.920 192.535 ;
        RECT 113.090 192.090 114.195 192.260 ;
        RECT 113.090 191.475 113.260 192.090 ;
        RECT 114.405 191.940 114.655 192.365 ;
        RECT 114.825 192.075 115.090 192.535 ;
        RECT 113.430 191.555 113.960 191.920 ;
        RECT 114.405 191.810 114.710 191.940 ;
        RECT 112.750 191.385 113.260 191.475 ;
        RECT 112.750 191.215 113.620 191.385 ;
        RECT 112.750 191.145 112.920 191.215 ;
        RECT 113.040 190.965 113.240 190.995 ;
        RECT 111.560 190.605 112.025 190.935 ;
        RECT 112.410 190.665 113.240 190.965 ;
        RECT 112.410 190.435 112.580 190.665 ;
        RECT 111.220 190.265 112.005 190.435 ;
        RECT 112.175 190.265 112.580 190.435 ;
        RECT 112.760 189.985 113.130 190.485 ;
        RECT 113.450 190.435 113.620 191.215 ;
        RECT 113.790 190.855 113.960 191.555 ;
        RECT 114.130 191.025 114.370 191.620 ;
        RECT 113.790 190.635 114.315 190.855 ;
        RECT 114.540 190.705 114.710 191.810 ;
        RECT 114.485 190.575 114.710 190.705 ;
        RECT 114.880 190.615 115.160 191.565 ;
        RECT 114.485 190.435 114.655 190.575 ;
        RECT 113.450 190.265 114.125 190.435 ;
        RECT 114.320 190.265 114.655 190.435 ;
        RECT 114.825 189.985 115.075 190.445 ;
        RECT 115.330 190.245 115.515 192.365 ;
        RECT 115.685 192.035 116.015 192.535 ;
        RECT 116.185 191.865 116.355 192.365 ;
        RECT 115.690 191.695 116.355 191.865 ;
        RECT 115.690 190.705 115.920 191.695 ;
        RECT 116.090 190.875 116.440 191.525 ;
        RECT 116.615 191.445 120.125 192.535 ;
        RECT 120.295 191.445 121.505 192.535 ;
        RECT 116.615 190.755 118.265 191.275 ;
        RECT 118.435 190.925 120.125 191.445 ;
        RECT 115.690 190.535 116.355 190.705 ;
        RECT 115.685 189.985 116.015 190.365 ;
        RECT 116.185 190.245 116.355 190.535 ;
        RECT 116.615 189.985 120.125 190.755 ;
        RECT 120.295 190.735 120.815 191.275 ;
        RECT 120.985 190.905 121.505 191.445 ;
        RECT 121.675 191.370 121.965 192.535 ;
        RECT 122.135 192.100 127.480 192.535 ;
        RECT 120.295 189.985 121.505 190.735 ;
        RECT 121.675 189.985 121.965 190.710 ;
        RECT 123.720 190.530 124.060 191.360 ;
        RECT 125.540 190.850 125.890 192.100 ;
        RECT 127.655 191.445 129.325 192.535 ;
        RECT 127.655 190.755 128.405 191.275 ;
        RECT 128.575 190.925 129.325 191.445 ;
        RECT 129.955 191.445 131.165 192.535 ;
        RECT 129.955 190.905 130.475 191.445 ;
        RECT 122.135 189.985 127.480 190.530 ;
        RECT 127.655 189.985 129.325 190.755 ;
        RECT 130.645 190.735 131.165 191.275 ;
        RECT 129.955 189.985 131.165 190.735 ;
        RECT 57.190 189.815 131.250 189.985 ;
        RECT 57.275 189.065 58.485 189.815 ;
        RECT 58.655 189.270 64.000 189.815 ;
        RECT 64.175 189.270 69.520 189.815 ;
        RECT 69.695 189.270 75.040 189.815 ;
        RECT 57.275 188.525 57.795 189.065 ;
        RECT 57.965 188.355 58.485 188.895 ;
        RECT 60.240 188.440 60.580 189.270 ;
        RECT 57.275 187.265 58.485 188.355 ;
        RECT 62.060 187.700 62.410 188.950 ;
        RECT 65.760 188.440 66.100 189.270 ;
        RECT 67.580 187.700 67.930 188.950 ;
        RECT 71.280 188.440 71.620 189.270 ;
        RECT 75.215 189.045 78.725 189.815 ;
        RECT 78.920 189.165 79.230 189.635 ;
        RECT 79.400 189.335 80.135 189.815 ;
        RECT 80.305 189.245 80.475 189.595 ;
        RECT 80.645 189.415 81.025 189.815 ;
        RECT 73.100 187.700 73.450 188.950 ;
        RECT 75.215 188.525 76.865 189.045 ;
        RECT 78.920 188.995 79.655 189.165 ;
        RECT 80.305 189.075 81.045 189.245 ;
        RECT 81.215 189.140 81.485 189.485 ;
        RECT 79.405 188.905 79.655 188.995 ;
        RECT 80.875 188.905 81.045 189.075 ;
        RECT 77.035 188.355 78.725 188.875 ;
        RECT 78.900 188.575 79.235 188.825 ;
        RECT 79.405 188.575 80.145 188.905 ;
        RECT 80.875 188.575 81.105 188.905 ;
        RECT 58.655 187.265 64.000 187.700 ;
        RECT 64.175 187.265 69.520 187.700 ;
        RECT 69.695 187.265 75.040 187.700 ;
        RECT 75.215 187.265 78.725 188.355 ;
        RECT 78.900 187.265 79.155 188.405 ;
        RECT 79.405 188.015 79.575 188.575 ;
        RECT 80.875 188.405 81.045 188.575 ;
        RECT 81.315 188.405 81.485 189.140 ;
        RECT 81.655 189.065 82.865 189.815 ;
        RECT 83.035 189.090 83.325 189.815 ;
        RECT 81.655 188.525 82.175 189.065 ;
        RECT 83.495 189.045 87.005 189.815 ;
        RECT 79.800 188.235 81.045 188.405 ;
        RECT 79.800 187.985 80.220 188.235 ;
        RECT 79.350 187.485 80.545 187.815 ;
        RECT 80.725 187.265 81.005 188.065 ;
        RECT 81.215 187.435 81.485 188.405 ;
        RECT 82.345 188.355 82.865 188.895 ;
        RECT 83.495 188.525 85.145 189.045 ;
        RECT 87.635 188.995 87.895 189.815 ;
        RECT 88.065 188.995 88.395 189.415 ;
        RECT 88.575 189.330 89.365 189.595 ;
        RECT 88.145 188.905 88.395 188.995 ;
        RECT 81.655 187.265 82.865 188.355 ;
        RECT 83.035 187.265 83.325 188.430 ;
        RECT 85.315 188.355 87.005 188.875 ;
        RECT 83.495 187.265 87.005 188.355 ;
        RECT 87.635 187.945 87.975 188.825 ;
        RECT 88.145 188.655 88.940 188.905 ;
        RECT 87.635 187.265 87.895 187.775 ;
        RECT 88.145 187.435 88.315 188.655 ;
        RECT 89.110 188.475 89.365 189.330 ;
        RECT 89.535 189.175 89.735 189.595 ;
        RECT 89.925 189.355 90.255 189.815 ;
        RECT 89.535 188.655 89.945 189.175 ;
        RECT 90.425 189.165 90.685 189.645 ;
        RECT 90.855 189.270 96.200 189.815 ;
        RECT 90.115 188.475 90.345 188.905 ;
        RECT 88.555 188.305 90.345 188.475 ;
        RECT 88.555 187.940 88.805 188.305 ;
        RECT 88.975 187.945 89.305 188.135 ;
        RECT 89.525 188.010 90.240 188.305 ;
        RECT 90.515 188.135 90.685 189.165 ;
        RECT 92.440 188.440 92.780 189.270 ;
        RECT 96.950 189.185 97.235 189.645 ;
        RECT 97.405 189.355 97.675 189.815 ;
        RECT 96.950 189.015 97.905 189.185 ;
        RECT 88.975 187.770 89.170 187.945 ;
        RECT 88.555 187.265 89.170 187.770 ;
        RECT 89.340 187.435 89.815 187.775 ;
        RECT 89.985 187.265 90.200 187.810 ;
        RECT 90.410 187.435 90.685 188.135 ;
        RECT 94.260 187.700 94.610 188.950 ;
        RECT 96.835 188.285 97.525 188.845 ;
        RECT 97.695 188.115 97.905 189.015 ;
        RECT 96.950 187.895 97.905 188.115 ;
        RECT 98.075 188.845 98.475 189.645 ;
        RECT 98.665 189.185 98.945 189.645 ;
        RECT 99.465 189.355 99.790 189.815 ;
        RECT 98.665 189.015 99.790 189.185 ;
        RECT 99.960 189.075 100.345 189.645 ;
        RECT 99.340 188.905 99.790 189.015 ;
        RECT 98.075 188.285 99.170 188.845 ;
        RECT 99.340 188.575 99.895 188.905 ;
        RECT 90.855 187.265 96.200 187.700 ;
        RECT 96.950 187.435 97.235 187.895 ;
        RECT 97.405 187.265 97.675 187.725 ;
        RECT 98.075 187.435 98.475 188.285 ;
        RECT 99.340 188.115 99.790 188.575 ;
        RECT 100.065 188.405 100.345 189.075 ;
        RECT 100.525 189.005 100.795 189.815 ;
        RECT 100.965 189.005 101.295 189.645 ;
        RECT 101.465 189.005 101.705 189.815 ;
        RECT 101.895 189.270 107.240 189.815 ;
        RECT 100.515 188.575 100.865 188.825 ;
        RECT 101.035 188.405 101.205 189.005 ;
        RECT 101.375 188.575 101.725 188.825 ;
        RECT 103.480 188.440 103.820 189.270 ;
        RECT 107.415 189.065 108.625 189.815 ;
        RECT 108.795 189.090 109.085 189.815 ;
        RECT 109.255 189.270 114.600 189.815 ;
        RECT 114.775 189.270 120.120 189.815 ;
        RECT 120.295 189.270 125.640 189.815 ;
        RECT 98.665 187.895 99.790 188.115 ;
        RECT 98.665 187.435 98.945 187.895 ;
        RECT 99.465 187.265 99.790 187.725 ;
        RECT 99.960 187.435 100.345 188.405 ;
        RECT 100.525 187.265 100.855 188.405 ;
        RECT 101.035 188.235 101.715 188.405 ;
        RECT 101.385 187.450 101.715 188.235 ;
        RECT 105.300 187.700 105.650 188.950 ;
        RECT 107.415 188.525 107.935 189.065 ;
        RECT 108.105 188.355 108.625 188.895 ;
        RECT 110.840 188.440 111.180 189.270 ;
        RECT 101.895 187.265 107.240 187.700 ;
        RECT 107.415 187.265 108.625 188.355 ;
        RECT 108.795 187.265 109.085 188.430 ;
        RECT 112.660 187.700 113.010 188.950 ;
        RECT 116.360 188.440 116.700 189.270 ;
        RECT 118.180 187.700 118.530 188.950 ;
        RECT 121.880 188.440 122.220 189.270 ;
        RECT 125.815 189.065 127.025 189.815 ;
        RECT 127.285 189.265 127.455 189.645 ;
        RECT 127.670 189.435 128.000 189.815 ;
        RECT 127.285 189.095 128.000 189.265 ;
        RECT 123.700 187.700 124.050 188.950 ;
        RECT 125.815 188.525 126.335 189.065 ;
        RECT 126.505 188.355 127.025 188.895 ;
        RECT 127.195 188.545 127.550 188.915 ;
        RECT 127.830 188.905 128.000 189.095 ;
        RECT 128.170 189.070 128.425 189.645 ;
        RECT 127.830 188.575 128.085 188.905 ;
        RECT 127.830 188.365 128.000 188.575 ;
        RECT 109.255 187.265 114.600 187.700 ;
        RECT 114.775 187.265 120.120 187.700 ;
        RECT 120.295 187.265 125.640 187.700 ;
        RECT 125.815 187.265 127.025 188.355 ;
        RECT 127.285 188.195 128.000 188.365 ;
        RECT 128.255 188.340 128.425 189.070 ;
        RECT 128.600 188.975 128.860 189.815 ;
        RECT 129.955 189.065 131.165 189.815 ;
        RECT 127.285 187.435 127.455 188.195 ;
        RECT 127.670 187.265 128.000 188.025 ;
        RECT 128.170 187.435 128.425 188.340 ;
        RECT 128.600 187.265 128.860 188.415 ;
        RECT 129.955 188.355 130.475 188.895 ;
        RECT 130.645 188.525 131.165 189.065 ;
        RECT 129.955 187.265 131.165 188.355 ;
        RECT 57.190 187.095 131.250 187.265 ;
        RECT 57.275 186.005 58.485 187.095 ;
        RECT 58.655 186.660 64.000 187.095 ;
        RECT 64.175 186.660 69.520 187.095 ;
        RECT 57.275 185.295 57.795 185.835 ;
        RECT 57.965 185.465 58.485 186.005 ;
        RECT 57.275 184.545 58.485 185.295 ;
        RECT 60.240 185.090 60.580 185.920 ;
        RECT 62.060 185.410 62.410 186.660 ;
        RECT 65.760 185.090 66.100 185.920 ;
        RECT 67.580 185.410 67.930 186.660 ;
        RECT 70.155 185.930 70.445 187.095 ;
        RECT 70.615 186.660 75.960 187.095 ;
        RECT 76.135 186.660 81.480 187.095 ;
        RECT 81.655 186.660 87.000 187.095 ;
        RECT 87.175 186.660 92.520 187.095 ;
        RECT 58.655 184.545 64.000 185.090 ;
        RECT 64.175 184.545 69.520 185.090 ;
        RECT 70.155 184.545 70.445 185.270 ;
        RECT 72.200 185.090 72.540 185.920 ;
        RECT 74.020 185.410 74.370 186.660 ;
        RECT 77.720 185.090 78.060 185.920 ;
        RECT 79.540 185.410 79.890 186.660 ;
        RECT 83.240 185.090 83.580 185.920 ;
        RECT 85.060 185.410 85.410 186.660 ;
        RECT 88.760 185.090 89.100 185.920 ;
        RECT 90.580 185.410 90.930 186.660 ;
        RECT 92.695 186.005 95.285 187.095 ;
        RECT 92.695 185.315 93.905 185.835 ;
        RECT 94.075 185.485 95.285 186.005 ;
        RECT 95.915 185.930 96.205 187.095 ;
        RECT 96.375 186.660 101.720 187.095 ;
        RECT 101.895 186.660 107.240 187.095 ;
        RECT 107.415 186.660 112.760 187.095 ;
        RECT 112.935 186.660 118.280 187.095 ;
        RECT 70.615 184.545 75.960 185.090 ;
        RECT 76.135 184.545 81.480 185.090 ;
        RECT 81.655 184.545 87.000 185.090 ;
        RECT 87.175 184.545 92.520 185.090 ;
        RECT 92.695 184.545 95.285 185.315 ;
        RECT 95.915 184.545 96.205 185.270 ;
        RECT 97.960 185.090 98.300 185.920 ;
        RECT 99.780 185.410 100.130 186.660 ;
        RECT 103.480 185.090 103.820 185.920 ;
        RECT 105.300 185.410 105.650 186.660 ;
        RECT 109.000 185.090 109.340 185.920 ;
        RECT 110.820 185.410 111.170 186.660 ;
        RECT 114.520 185.090 114.860 185.920 ;
        RECT 116.340 185.410 116.690 186.660 ;
        RECT 118.455 186.005 121.045 187.095 ;
        RECT 118.455 185.315 119.665 185.835 ;
        RECT 119.835 185.485 121.045 186.005 ;
        RECT 121.675 185.930 121.965 187.095 ;
        RECT 122.135 186.660 127.480 187.095 ;
        RECT 96.375 184.545 101.720 185.090 ;
        RECT 101.895 184.545 107.240 185.090 ;
        RECT 107.415 184.545 112.760 185.090 ;
        RECT 112.935 184.545 118.280 185.090 ;
        RECT 118.455 184.545 121.045 185.315 ;
        RECT 121.675 184.545 121.965 185.270 ;
        RECT 123.720 185.090 124.060 185.920 ;
        RECT 125.540 185.410 125.890 186.660 ;
        RECT 127.655 186.005 129.325 187.095 ;
        RECT 127.655 185.315 128.405 185.835 ;
        RECT 128.575 185.485 129.325 186.005 ;
        RECT 129.955 186.005 131.165 187.095 ;
        RECT 129.955 185.465 130.475 186.005 ;
        RECT 122.135 184.545 127.480 185.090 ;
        RECT 127.655 184.545 129.325 185.315 ;
        RECT 130.645 185.295 131.165 185.835 ;
        RECT 129.955 184.545 131.165 185.295 ;
        RECT 57.190 184.375 131.250 184.545 ;
        RECT 57.275 183.625 58.485 184.375 ;
        RECT 58.655 183.830 64.000 184.375 ;
        RECT 64.175 183.830 69.520 184.375 ;
        RECT 69.695 183.830 75.040 184.375 ;
        RECT 75.215 183.830 80.560 184.375 ;
        RECT 57.275 183.085 57.795 183.625 ;
        RECT 57.965 182.915 58.485 183.455 ;
        RECT 60.240 183.000 60.580 183.830 ;
        RECT 57.275 181.825 58.485 182.915 ;
        RECT 62.060 182.260 62.410 183.510 ;
        RECT 65.760 183.000 66.100 183.830 ;
        RECT 67.580 182.260 67.930 183.510 ;
        RECT 71.280 183.000 71.620 183.830 ;
        RECT 73.100 182.260 73.450 183.510 ;
        RECT 76.800 183.000 77.140 183.830 ;
        RECT 80.735 183.605 82.405 184.375 ;
        RECT 83.035 183.650 83.325 184.375 ;
        RECT 83.495 183.830 88.840 184.375 ;
        RECT 89.015 183.830 94.360 184.375 ;
        RECT 94.535 183.830 99.880 184.375 ;
        RECT 100.055 183.830 105.400 184.375 ;
        RECT 78.620 182.260 78.970 183.510 ;
        RECT 80.735 183.085 81.485 183.605 ;
        RECT 81.655 182.915 82.405 183.435 ;
        RECT 85.080 183.000 85.420 183.830 ;
        RECT 58.655 181.825 64.000 182.260 ;
        RECT 64.175 181.825 69.520 182.260 ;
        RECT 69.695 181.825 75.040 182.260 ;
        RECT 75.215 181.825 80.560 182.260 ;
        RECT 80.735 181.825 82.405 182.915 ;
        RECT 83.035 181.825 83.325 182.990 ;
        RECT 86.900 182.260 87.250 183.510 ;
        RECT 90.600 183.000 90.940 183.830 ;
        RECT 92.420 182.260 92.770 183.510 ;
        RECT 96.120 183.000 96.460 183.830 ;
        RECT 97.940 182.260 98.290 183.510 ;
        RECT 101.640 183.000 101.980 183.830 ;
        RECT 105.575 183.605 108.165 184.375 ;
        RECT 108.795 183.650 109.085 184.375 ;
        RECT 109.255 183.830 114.600 184.375 ;
        RECT 114.775 183.830 120.120 184.375 ;
        RECT 120.295 183.830 125.640 184.375 ;
        RECT 103.460 182.260 103.810 183.510 ;
        RECT 105.575 183.085 106.785 183.605 ;
        RECT 106.955 182.915 108.165 183.435 ;
        RECT 110.840 183.000 111.180 183.830 ;
        RECT 83.495 181.825 88.840 182.260 ;
        RECT 89.015 181.825 94.360 182.260 ;
        RECT 94.535 181.825 99.880 182.260 ;
        RECT 100.055 181.825 105.400 182.260 ;
        RECT 105.575 181.825 108.165 182.915 ;
        RECT 108.795 181.825 109.085 182.990 ;
        RECT 112.660 182.260 113.010 183.510 ;
        RECT 116.360 183.000 116.700 183.830 ;
        RECT 118.180 182.260 118.530 183.510 ;
        RECT 121.880 183.000 122.220 183.830 ;
        RECT 125.815 183.605 129.325 184.375 ;
        RECT 129.955 183.625 131.165 184.375 ;
        RECT 123.700 182.260 124.050 183.510 ;
        RECT 125.815 183.085 127.465 183.605 ;
        RECT 127.635 182.915 129.325 183.435 ;
        RECT 109.255 181.825 114.600 182.260 ;
        RECT 114.775 181.825 120.120 182.260 ;
        RECT 120.295 181.825 125.640 182.260 ;
        RECT 125.815 181.825 129.325 182.915 ;
        RECT 129.955 182.915 130.475 183.455 ;
        RECT 130.645 183.085 131.165 183.625 ;
        RECT 129.955 181.825 131.165 182.915 ;
        RECT 57.190 181.655 131.250 181.825 ;
        RECT 57.275 180.565 58.485 181.655 ;
        RECT 58.655 181.220 64.000 181.655 ;
        RECT 64.175 181.220 69.520 181.655 ;
        RECT 57.275 179.855 57.795 180.395 ;
        RECT 57.965 180.025 58.485 180.565 ;
        RECT 57.275 179.105 58.485 179.855 ;
        RECT 60.240 179.650 60.580 180.480 ;
        RECT 62.060 179.970 62.410 181.220 ;
        RECT 65.760 179.650 66.100 180.480 ;
        RECT 67.580 179.970 67.930 181.220 ;
        RECT 70.155 180.490 70.445 181.655 ;
        RECT 70.615 181.220 75.960 181.655 ;
        RECT 76.135 181.220 81.480 181.655 ;
        RECT 81.655 181.220 87.000 181.655 ;
        RECT 87.175 181.220 92.520 181.655 ;
        RECT 58.655 179.105 64.000 179.650 ;
        RECT 64.175 179.105 69.520 179.650 ;
        RECT 70.155 179.105 70.445 179.830 ;
        RECT 72.200 179.650 72.540 180.480 ;
        RECT 74.020 179.970 74.370 181.220 ;
        RECT 77.720 179.650 78.060 180.480 ;
        RECT 79.540 179.970 79.890 181.220 ;
        RECT 83.240 179.650 83.580 180.480 ;
        RECT 85.060 179.970 85.410 181.220 ;
        RECT 88.760 179.650 89.100 180.480 ;
        RECT 90.580 179.970 90.930 181.220 ;
        RECT 92.695 180.565 95.285 181.655 ;
        RECT 92.695 179.875 93.905 180.395 ;
        RECT 94.075 180.045 95.285 180.565 ;
        RECT 95.915 180.490 96.205 181.655 ;
        RECT 96.375 181.220 101.720 181.655 ;
        RECT 101.895 181.220 107.240 181.655 ;
        RECT 107.415 181.220 112.760 181.655 ;
        RECT 112.935 181.220 118.280 181.655 ;
        RECT 70.615 179.105 75.960 179.650 ;
        RECT 76.135 179.105 81.480 179.650 ;
        RECT 81.655 179.105 87.000 179.650 ;
        RECT 87.175 179.105 92.520 179.650 ;
        RECT 92.695 179.105 95.285 179.875 ;
        RECT 95.915 179.105 96.205 179.830 ;
        RECT 97.960 179.650 98.300 180.480 ;
        RECT 99.780 179.970 100.130 181.220 ;
        RECT 103.480 179.650 103.820 180.480 ;
        RECT 105.300 179.970 105.650 181.220 ;
        RECT 109.000 179.650 109.340 180.480 ;
        RECT 110.820 179.970 111.170 181.220 ;
        RECT 114.520 179.650 114.860 180.480 ;
        RECT 116.340 179.970 116.690 181.220 ;
        RECT 118.455 180.565 121.045 181.655 ;
        RECT 118.455 179.875 119.665 180.395 ;
        RECT 119.835 180.045 121.045 180.565 ;
        RECT 121.675 180.490 121.965 181.655 ;
        RECT 122.135 181.220 127.480 181.655 ;
        RECT 96.375 179.105 101.720 179.650 ;
        RECT 101.895 179.105 107.240 179.650 ;
        RECT 107.415 179.105 112.760 179.650 ;
        RECT 112.935 179.105 118.280 179.650 ;
        RECT 118.455 179.105 121.045 179.875 ;
        RECT 121.675 179.105 121.965 179.830 ;
        RECT 123.720 179.650 124.060 180.480 ;
        RECT 125.540 179.970 125.890 181.220 ;
        RECT 127.655 180.565 129.325 181.655 ;
        RECT 127.655 179.875 128.405 180.395 ;
        RECT 128.575 180.045 129.325 180.565 ;
        RECT 129.955 180.565 131.165 181.655 ;
        RECT 129.955 180.025 130.475 180.565 ;
        RECT 122.135 179.105 127.480 179.650 ;
        RECT 127.655 179.105 129.325 179.875 ;
        RECT 130.645 179.855 131.165 180.395 ;
        RECT 129.955 179.105 131.165 179.855 ;
        RECT 57.190 178.935 131.250 179.105 ;
        RECT 57.275 178.185 58.485 178.935 ;
        RECT 58.655 178.390 64.000 178.935 ;
        RECT 64.175 178.390 69.520 178.935 ;
        RECT 69.695 178.390 75.040 178.935 ;
        RECT 75.215 178.390 80.560 178.935 ;
        RECT 57.275 177.645 57.795 178.185 ;
        RECT 57.965 177.475 58.485 178.015 ;
        RECT 60.240 177.560 60.580 178.390 ;
        RECT 57.275 176.385 58.485 177.475 ;
        RECT 62.060 176.820 62.410 178.070 ;
        RECT 65.760 177.560 66.100 178.390 ;
        RECT 67.580 176.820 67.930 178.070 ;
        RECT 71.280 177.560 71.620 178.390 ;
        RECT 73.100 176.820 73.450 178.070 ;
        RECT 76.800 177.560 77.140 178.390 ;
        RECT 80.735 178.165 82.405 178.935 ;
        RECT 83.035 178.210 83.325 178.935 ;
        RECT 83.495 178.390 88.840 178.935 ;
        RECT 89.015 178.390 94.360 178.935 ;
        RECT 94.535 178.390 99.880 178.935 ;
        RECT 100.055 178.390 105.400 178.935 ;
        RECT 78.620 176.820 78.970 178.070 ;
        RECT 80.735 177.645 81.485 178.165 ;
        RECT 81.655 177.475 82.405 177.995 ;
        RECT 85.080 177.560 85.420 178.390 ;
        RECT 58.655 176.385 64.000 176.820 ;
        RECT 64.175 176.385 69.520 176.820 ;
        RECT 69.695 176.385 75.040 176.820 ;
        RECT 75.215 176.385 80.560 176.820 ;
        RECT 80.735 176.385 82.405 177.475 ;
        RECT 83.035 176.385 83.325 177.550 ;
        RECT 86.900 176.820 87.250 178.070 ;
        RECT 90.600 177.560 90.940 178.390 ;
        RECT 92.420 176.820 92.770 178.070 ;
        RECT 96.120 177.560 96.460 178.390 ;
        RECT 97.940 176.820 98.290 178.070 ;
        RECT 101.640 177.560 101.980 178.390 ;
        RECT 105.575 178.165 108.165 178.935 ;
        RECT 108.795 178.210 109.085 178.935 ;
        RECT 109.255 178.390 114.600 178.935 ;
        RECT 114.775 178.390 120.120 178.935 ;
        RECT 120.295 178.390 125.640 178.935 ;
        RECT 103.460 176.820 103.810 178.070 ;
        RECT 105.575 177.645 106.785 178.165 ;
        RECT 106.955 177.475 108.165 177.995 ;
        RECT 110.840 177.560 111.180 178.390 ;
        RECT 83.495 176.385 88.840 176.820 ;
        RECT 89.015 176.385 94.360 176.820 ;
        RECT 94.535 176.385 99.880 176.820 ;
        RECT 100.055 176.385 105.400 176.820 ;
        RECT 105.575 176.385 108.165 177.475 ;
        RECT 108.795 176.385 109.085 177.550 ;
        RECT 112.660 176.820 113.010 178.070 ;
        RECT 116.360 177.560 116.700 178.390 ;
        RECT 118.180 176.820 118.530 178.070 ;
        RECT 121.880 177.560 122.220 178.390 ;
        RECT 125.815 178.165 129.325 178.935 ;
        RECT 129.955 178.185 131.165 178.935 ;
        RECT 123.700 176.820 124.050 178.070 ;
        RECT 125.815 177.645 127.465 178.165 ;
        RECT 127.635 177.475 129.325 177.995 ;
        RECT 109.255 176.385 114.600 176.820 ;
        RECT 114.775 176.385 120.120 176.820 ;
        RECT 120.295 176.385 125.640 176.820 ;
        RECT 125.815 176.385 129.325 177.475 ;
        RECT 129.955 177.475 130.475 178.015 ;
        RECT 130.645 177.645 131.165 178.185 ;
        RECT 129.955 176.385 131.165 177.475 ;
        RECT 57.190 176.215 131.250 176.385 ;
        RECT 57.275 175.125 58.485 176.215 ;
        RECT 58.655 175.780 64.000 176.215 ;
        RECT 64.175 175.780 69.520 176.215 ;
        RECT 57.275 174.415 57.795 174.955 ;
        RECT 57.965 174.585 58.485 175.125 ;
        RECT 57.275 173.665 58.485 174.415 ;
        RECT 60.240 174.210 60.580 175.040 ;
        RECT 62.060 174.530 62.410 175.780 ;
        RECT 65.760 174.210 66.100 175.040 ;
        RECT 67.580 174.530 67.930 175.780 ;
        RECT 70.155 175.050 70.445 176.215 ;
        RECT 70.615 175.780 75.960 176.215 ;
        RECT 76.135 175.780 81.480 176.215 ;
        RECT 81.655 175.780 87.000 176.215 ;
        RECT 87.175 175.780 92.520 176.215 ;
        RECT 58.655 173.665 64.000 174.210 ;
        RECT 64.175 173.665 69.520 174.210 ;
        RECT 70.155 173.665 70.445 174.390 ;
        RECT 72.200 174.210 72.540 175.040 ;
        RECT 74.020 174.530 74.370 175.780 ;
        RECT 77.720 174.210 78.060 175.040 ;
        RECT 79.540 174.530 79.890 175.780 ;
        RECT 83.240 174.210 83.580 175.040 ;
        RECT 85.060 174.530 85.410 175.780 ;
        RECT 88.760 174.210 89.100 175.040 ;
        RECT 90.580 174.530 90.930 175.780 ;
        RECT 92.695 175.125 95.285 176.215 ;
        RECT 92.695 174.435 93.905 174.955 ;
        RECT 94.075 174.605 95.285 175.125 ;
        RECT 95.915 175.050 96.205 176.215 ;
        RECT 96.375 175.780 101.720 176.215 ;
        RECT 101.895 175.780 107.240 176.215 ;
        RECT 107.415 175.780 112.760 176.215 ;
        RECT 112.935 175.780 118.280 176.215 ;
        RECT 70.615 173.665 75.960 174.210 ;
        RECT 76.135 173.665 81.480 174.210 ;
        RECT 81.655 173.665 87.000 174.210 ;
        RECT 87.175 173.665 92.520 174.210 ;
        RECT 92.695 173.665 95.285 174.435 ;
        RECT 95.915 173.665 96.205 174.390 ;
        RECT 97.960 174.210 98.300 175.040 ;
        RECT 99.780 174.530 100.130 175.780 ;
        RECT 103.480 174.210 103.820 175.040 ;
        RECT 105.300 174.530 105.650 175.780 ;
        RECT 109.000 174.210 109.340 175.040 ;
        RECT 110.820 174.530 111.170 175.780 ;
        RECT 114.520 174.210 114.860 175.040 ;
        RECT 116.340 174.530 116.690 175.780 ;
        RECT 118.455 175.125 121.045 176.215 ;
        RECT 118.455 174.435 119.665 174.955 ;
        RECT 119.835 174.605 121.045 175.125 ;
        RECT 121.675 175.050 121.965 176.215 ;
        RECT 122.135 175.780 127.480 176.215 ;
        RECT 96.375 173.665 101.720 174.210 ;
        RECT 101.895 173.665 107.240 174.210 ;
        RECT 107.415 173.665 112.760 174.210 ;
        RECT 112.935 173.665 118.280 174.210 ;
        RECT 118.455 173.665 121.045 174.435 ;
        RECT 121.675 173.665 121.965 174.390 ;
        RECT 123.720 174.210 124.060 175.040 ;
        RECT 125.540 174.530 125.890 175.780 ;
        RECT 127.655 175.125 129.325 176.215 ;
        RECT 127.655 174.435 128.405 174.955 ;
        RECT 128.575 174.605 129.325 175.125 ;
        RECT 129.955 175.125 131.165 176.215 ;
        RECT 129.955 174.585 130.475 175.125 ;
        RECT 122.135 173.665 127.480 174.210 ;
        RECT 127.655 173.665 129.325 174.435 ;
        RECT 130.645 174.415 131.165 174.955 ;
        RECT 129.955 173.665 131.165 174.415 ;
        RECT 57.190 173.495 131.250 173.665 ;
        RECT 57.275 172.745 58.485 173.495 ;
        RECT 58.655 172.950 64.000 173.495 ;
        RECT 64.175 172.950 69.520 173.495 ;
        RECT 69.695 172.950 75.040 173.495 ;
        RECT 75.215 172.950 80.560 173.495 ;
        RECT 57.275 172.205 57.795 172.745 ;
        RECT 57.965 172.035 58.485 172.575 ;
        RECT 60.240 172.120 60.580 172.950 ;
        RECT 57.275 170.945 58.485 172.035 ;
        RECT 62.060 171.380 62.410 172.630 ;
        RECT 65.760 172.120 66.100 172.950 ;
        RECT 67.580 171.380 67.930 172.630 ;
        RECT 71.280 172.120 71.620 172.950 ;
        RECT 73.100 171.380 73.450 172.630 ;
        RECT 76.800 172.120 77.140 172.950 ;
        RECT 80.735 172.725 82.405 173.495 ;
        RECT 83.035 172.770 83.325 173.495 ;
        RECT 83.495 172.950 88.840 173.495 ;
        RECT 89.015 172.950 94.360 173.495 ;
        RECT 94.535 172.950 99.880 173.495 ;
        RECT 100.055 172.950 105.400 173.495 ;
        RECT 78.620 171.380 78.970 172.630 ;
        RECT 80.735 172.205 81.485 172.725 ;
        RECT 81.655 172.035 82.405 172.555 ;
        RECT 85.080 172.120 85.420 172.950 ;
        RECT 58.655 170.945 64.000 171.380 ;
        RECT 64.175 170.945 69.520 171.380 ;
        RECT 69.695 170.945 75.040 171.380 ;
        RECT 75.215 170.945 80.560 171.380 ;
        RECT 80.735 170.945 82.405 172.035 ;
        RECT 83.035 170.945 83.325 172.110 ;
        RECT 86.900 171.380 87.250 172.630 ;
        RECT 90.600 172.120 90.940 172.950 ;
        RECT 92.420 171.380 92.770 172.630 ;
        RECT 96.120 172.120 96.460 172.950 ;
        RECT 97.940 171.380 98.290 172.630 ;
        RECT 101.640 172.120 101.980 172.950 ;
        RECT 105.575 172.725 108.165 173.495 ;
        RECT 108.795 172.770 109.085 173.495 ;
        RECT 109.255 172.950 114.600 173.495 ;
        RECT 114.775 172.950 120.120 173.495 ;
        RECT 120.295 172.950 125.640 173.495 ;
        RECT 103.460 171.380 103.810 172.630 ;
        RECT 105.575 172.205 106.785 172.725 ;
        RECT 106.955 172.035 108.165 172.555 ;
        RECT 110.840 172.120 111.180 172.950 ;
        RECT 83.495 170.945 88.840 171.380 ;
        RECT 89.015 170.945 94.360 171.380 ;
        RECT 94.535 170.945 99.880 171.380 ;
        RECT 100.055 170.945 105.400 171.380 ;
        RECT 105.575 170.945 108.165 172.035 ;
        RECT 108.795 170.945 109.085 172.110 ;
        RECT 112.660 171.380 113.010 172.630 ;
        RECT 116.360 172.120 116.700 172.950 ;
        RECT 118.180 171.380 118.530 172.630 ;
        RECT 121.880 172.120 122.220 172.950 ;
        RECT 125.815 172.725 129.325 173.495 ;
        RECT 129.955 172.745 131.165 173.495 ;
        RECT 123.700 171.380 124.050 172.630 ;
        RECT 125.815 172.205 127.465 172.725 ;
        RECT 127.635 172.035 129.325 172.555 ;
        RECT 109.255 170.945 114.600 171.380 ;
        RECT 114.775 170.945 120.120 171.380 ;
        RECT 120.295 170.945 125.640 171.380 ;
        RECT 125.815 170.945 129.325 172.035 ;
        RECT 129.955 172.035 130.475 172.575 ;
        RECT 130.645 172.205 131.165 172.745 ;
        RECT 129.955 170.945 131.165 172.035 ;
        RECT 57.190 170.775 131.250 170.945 ;
        RECT 57.275 169.685 58.485 170.775 ;
        RECT 58.655 170.340 64.000 170.775 ;
        RECT 64.175 170.340 69.520 170.775 ;
        RECT 57.275 168.975 57.795 169.515 ;
        RECT 57.965 169.145 58.485 169.685 ;
        RECT 57.275 168.225 58.485 168.975 ;
        RECT 60.240 168.770 60.580 169.600 ;
        RECT 62.060 169.090 62.410 170.340 ;
        RECT 65.760 168.770 66.100 169.600 ;
        RECT 67.580 169.090 67.930 170.340 ;
        RECT 70.155 169.610 70.445 170.775 ;
        RECT 70.615 170.340 75.960 170.775 ;
        RECT 76.135 170.340 81.480 170.775 ;
        RECT 81.655 170.340 87.000 170.775 ;
        RECT 87.175 170.340 92.520 170.775 ;
        RECT 58.655 168.225 64.000 168.770 ;
        RECT 64.175 168.225 69.520 168.770 ;
        RECT 70.155 168.225 70.445 168.950 ;
        RECT 72.200 168.770 72.540 169.600 ;
        RECT 74.020 169.090 74.370 170.340 ;
        RECT 77.720 168.770 78.060 169.600 ;
        RECT 79.540 169.090 79.890 170.340 ;
        RECT 83.240 168.770 83.580 169.600 ;
        RECT 85.060 169.090 85.410 170.340 ;
        RECT 88.760 168.770 89.100 169.600 ;
        RECT 90.580 169.090 90.930 170.340 ;
        RECT 92.695 169.685 95.285 170.775 ;
        RECT 92.695 168.995 93.905 169.515 ;
        RECT 94.075 169.165 95.285 169.685 ;
        RECT 95.915 169.610 96.205 170.775 ;
        RECT 96.375 170.340 101.720 170.775 ;
        RECT 101.895 170.340 107.240 170.775 ;
        RECT 107.415 170.340 112.760 170.775 ;
        RECT 112.935 170.340 118.280 170.775 ;
        RECT 70.615 168.225 75.960 168.770 ;
        RECT 76.135 168.225 81.480 168.770 ;
        RECT 81.655 168.225 87.000 168.770 ;
        RECT 87.175 168.225 92.520 168.770 ;
        RECT 92.695 168.225 95.285 168.995 ;
        RECT 95.915 168.225 96.205 168.950 ;
        RECT 97.960 168.770 98.300 169.600 ;
        RECT 99.780 169.090 100.130 170.340 ;
        RECT 103.480 168.770 103.820 169.600 ;
        RECT 105.300 169.090 105.650 170.340 ;
        RECT 109.000 168.770 109.340 169.600 ;
        RECT 110.820 169.090 111.170 170.340 ;
        RECT 114.520 168.770 114.860 169.600 ;
        RECT 116.340 169.090 116.690 170.340 ;
        RECT 118.455 169.685 121.045 170.775 ;
        RECT 118.455 168.995 119.665 169.515 ;
        RECT 119.835 169.165 121.045 169.685 ;
        RECT 121.675 169.610 121.965 170.775 ;
        RECT 122.135 170.340 127.480 170.775 ;
        RECT 96.375 168.225 101.720 168.770 ;
        RECT 101.895 168.225 107.240 168.770 ;
        RECT 107.415 168.225 112.760 168.770 ;
        RECT 112.935 168.225 118.280 168.770 ;
        RECT 118.455 168.225 121.045 168.995 ;
        RECT 121.675 168.225 121.965 168.950 ;
        RECT 123.720 168.770 124.060 169.600 ;
        RECT 125.540 169.090 125.890 170.340 ;
        RECT 127.655 169.685 129.325 170.775 ;
        RECT 127.655 168.995 128.405 169.515 ;
        RECT 128.575 169.165 129.325 169.685 ;
        RECT 129.955 169.685 131.165 170.775 ;
        RECT 129.955 169.145 130.475 169.685 ;
        RECT 122.135 168.225 127.480 168.770 ;
        RECT 127.655 168.225 129.325 168.995 ;
        RECT 130.645 168.975 131.165 169.515 ;
        RECT 129.955 168.225 131.165 168.975 ;
        RECT 57.190 168.055 131.250 168.225 ;
        RECT 57.275 167.305 58.485 168.055 ;
        RECT 58.655 167.510 64.000 168.055 ;
        RECT 64.175 167.510 69.520 168.055 ;
        RECT 69.695 167.510 75.040 168.055 ;
        RECT 75.215 167.510 80.560 168.055 ;
        RECT 57.275 166.765 57.795 167.305 ;
        RECT 57.965 166.595 58.485 167.135 ;
        RECT 60.240 166.680 60.580 167.510 ;
        RECT 57.275 165.505 58.485 166.595 ;
        RECT 62.060 165.940 62.410 167.190 ;
        RECT 65.760 166.680 66.100 167.510 ;
        RECT 67.580 165.940 67.930 167.190 ;
        RECT 71.280 166.680 71.620 167.510 ;
        RECT 73.100 165.940 73.450 167.190 ;
        RECT 76.800 166.680 77.140 167.510 ;
        RECT 80.735 167.285 82.405 168.055 ;
        RECT 83.035 167.330 83.325 168.055 ;
        RECT 83.495 167.510 88.840 168.055 ;
        RECT 89.015 167.510 94.360 168.055 ;
        RECT 94.535 167.510 99.880 168.055 ;
        RECT 100.055 167.510 105.400 168.055 ;
        RECT 78.620 165.940 78.970 167.190 ;
        RECT 80.735 166.765 81.485 167.285 ;
        RECT 81.655 166.595 82.405 167.115 ;
        RECT 85.080 166.680 85.420 167.510 ;
        RECT 58.655 165.505 64.000 165.940 ;
        RECT 64.175 165.505 69.520 165.940 ;
        RECT 69.695 165.505 75.040 165.940 ;
        RECT 75.215 165.505 80.560 165.940 ;
        RECT 80.735 165.505 82.405 166.595 ;
        RECT 83.035 165.505 83.325 166.670 ;
        RECT 86.900 165.940 87.250 167.190 ;
        RECT 90.600 166.680 90.940 167.510 ;
        RECT 92.420 165.940 92.770 167.190 ;
        RECT 96.120 166.680 96.460 167.510 ;
        RECT 97.940 165.940 98.290 167.190 ;
        RECT 101.640 166.680 101.980 167.510 ;
        RECT 105.575 167.285 108.165 168.055 ;
        RECT 108.795 167.330 109.085 168.055 ;
        RECT 109.255 167.510 114.600 168.055 ;
        RECT 114.775 167.510 120.120 168.055 ;
        RECT 120.295 167.510 125.640 168.055 ;
        RECT 103.460 165.940 103.810 167.190 ;
        RECT 105.575 166.765 106.785 167.285 ;
        RECT 106.955 166.595 108.165 167.115 ;
        RECT 110.840 166.680 111.180 167.510 ;
        RECT 83.495 165.505 88.840 165.940 ;
        RECT 89.015 165.505 94.360 165.940 ;
        RECT 94.535 165.505 99.880 165.940 ;
        RECT 100.055 165.505 105.400 165.940 ;
        RECT 105.575 165.505 108.165 166.595 ;
        RECT 108.795 165.505 109.085 166.670 ;
        RECT 112.660 165.940 113.010 167.190 ;
        RECT 116.360 166.680 116.700 167.510 ;
        RECT 118.180 165.940 118.530 167.190 ;
        RECT 121.880 166.680 122.220 167.510 ;
        RECT 125.815 167.285 129.325 168.055 ;
        RECT 129.955 167.305 131.165 168.055 ;
        RECT 123.700 165.940 124.050 167.190 ;
        RECT 125.815 166.765 127.465 167.285 ;
        RECT 127.635 166.595 129.325 167.115 ;
        RECT 109.255 165.505 114.600 165.940 ;
        RECT 114.775 165.505 120.120 165.940 ;
        RECT 120.295 165.505 125.640 165.940 ;
        RECT 125.815 165.505 129.325 166.595 ;
        RECT 129.955 166.595 130.475 167.135 ;
        RECT 130.645 166.765 131.165 167.305 ;
        RECT 129.955 165.505 131.165 166.595 ;
        RECT 57.190 165.335 131.250 165.505 ;
        RECT 57.275 164.245 58.485 165.335 ;
        RECT 58.655 164.900 64.000 165.335 ;
        RECT 64.175 164.900 69.520 165.335 ;
        RECT 57.275 163.535 57.795 164.075 ;
        RECT 57.965 163.705 58.485 164.245 ;
        RECT 57.275 162.785 58.485 163.535 ;
        RECT 60.240 163.330 60.580 164.160 ;
        RECT 62.060 163.650 62.410 164.900 ;
        RECT 65.760 163.330 66.100 164.160 ;
        RECT 67.580 163.650 67.930 164.900 ;
        RECT 70.155 164.170 70.445 165.335 ;
        RECT 70.615 164.900 75.960 165.335 ;
        RECT 76.135 164.900 81.480 165.335 ;
        RECT 81.655 164.900 87.000 165.335 ;
        RECT 87.175 164.900 92.520 165.335 ;
        RECT 58.655 162.785 64.000 163.330 ;
        RECT 64.175 162.785 69.520 163.330 ;
        RECT 70.155 162.785 70.445 163.510 ;
        RECT 72.200 163.330 72.540 164.160 ;
        RECT 74.020 163.650 74.370 164.900 ;
        RECT 77.720 163.330 78.060 164.160 ;
        RECT 79.540 163.650 79.890 164.900 ;
        RECT 83.240 163.330 83.580 164.160 ;
        RECT 85.060 163.650 85.410 164.900 ;
        RECT 88.760 163.330 89.100 164.160 ;
        RECT 90.580 163.650 90.930 164.900 ;
        RECT 92.695 164.245 95.285 165.335 ;
        RECT 92.695 163.555 93.905 164.075 ;
        RECT 94.075 163.725 95.285 164.245 ;
        RECT 95.915 164.170 96.205 165.335 ;
        RECT 96.375 164.900 101.720 165.335 ;
        RECT 101.895 164.900 107.240 165.335 ;
        RECT 107.415 164.900 112.760 165.335 ;
        RECT 112.935 164.900 118.280 165.335 ;
        RECT 70.615 162.785 75.960 163.330 ;
        RECT 76.135 162.785 81.480 163.330 ;
        RECT 81.655 162.785 87.000 163.330 ;
        RECT 87.175 162.785 92.520 163.330 ;
        RECT 92.695 162.785 95.285 163.555 ;
        RECT 95.915 162.785 96.205 163.510 ;
        RECT 97.960 163.330 98.300 164.160 ;
        RECT 99.780 163.650 100.130 164.900 ;
        RECT 103.480 163.330 103.820 164.160 ;
        RECT 105.300 163.650 105.650 164.900 ;
        RECT 109.000 163.330 109.340 164.160 ;
        RECT 110.820 163.650 111.170 164.900 ;
        RECT 114.520 163.330 114.860 164.160 ;
        RECT 116.340 163.650 116.690 164.900 ;
        RECT 118.455 164.245 121.045 165.335 ;
        RECT 118.455 163.555 119.665 164.075 ;
        RECT 119.835 163.725 121.045 164.245 ;
        RECT 121.675 164.170 121.965 165.335 ;
        RECT 122.135 164.900 127.480 165.335 ;
        RECT 96.375 162.785 101.720 163.330 ;
        RECT 101.895 162.785 107.240 163.330 ;
        RECT 107.415 162.785 112.760 163.330 ;
        RECT 112.935 162.785 118.280 163.330 ;
        RECT 118.455 162.785 121.045 163.555 ;
        RECT 121.675 162.785 121.965 163.510 ;
        RECT 123.720 163.330 124.060 164.160 ;
        RECT 125.540 163.650 125.890 164.900 ;
        RECT 127.655 164.245 129.325 165.335 ;
        RECT 127.655 163.555 128.405 164.075 ;
        RECT 128.575 163.725 129.325 164.245 ;
        RECT 129.955 164.245 131.165 165.335 ;
        RECT 129.955 163.705 130.475 164.245 ;
        RECT 122.135 162.785 127.480 163.330 ;
        RECT 127.655 162.785 129.325 163.555 ;
        RECT 130.645 163.535 131.165 164.075 ;
        RECT 129.955 162.785 131.165 163.535 ;
        RECT 57.190 162.615 131.250 162.785 ;
        RECT 57.275 161.865 58.485 162.615 ;
        RECT 58.655 162.070 64.000 162.615 ;
        RECT 64.175 162.070 69.520 162.615 ;
        RECT 69.695 162.070 75.040 162.615 ;
        RECT 75.215 162.070 80.560 162.615 ;
        RECT 57.275 161.325 57.795 161.865 ;
        RECT 57.965 161.155 58.485 161.695 ;
        RECT 60.240 161.240 60.580 162.070 ;
        RECT 57.275 160.065 58.485 161.155 ;
        RECT 62.060 160.500 62.410 161.750 ;
        RECT 65.760 161.240 66.100 162.070 ;
        RECT 67.580 160.500 67.930 161.750 ;
        RECT 71.280 161.240 71.620 162.070 ;
        RECT 73.100 160.500 73.450 161.750 ;
        RECT 76.800 161.240 77.140 162.070 ;
        RECT 80.735 161.845 82.405 162.615 ;
        RECT 83.035 161.890 83.325 162.615 ;
        RECT 83.495 162.070 88.840 162.615 ;
        RECT 89.015 162.070 94.360 162.615 ;
        RECT 94.535 162.070 99.880 162.615 ;
        RECT 100.055 162.070 105.400 162.615 ;
        RECT 78.620 160.500 78.970 161.750 ;
        RECT 80.735 161.325 81.485 161.845 ;
        RECT 81.655 161.155 82.405 161.675 ;
        RECT 85.080 161.240 85.420 162.070 ;
        RECT 58.655 160.065 64.000 160.500 ;
        RECT 64.175 160.065 69.520 160.500 ;
        RECT 69.695 160.065 75.040 160.500 ;
        RECT 75.215 160.065 80.560 160.500 ;
        RECT 80.735 160.065 82.405 161.155 ;
        RECT 83.035 160.065 83.325 161.230 ;
        RECT 86.900 160.500 87.250 161.750 ;
        RECT 90.600 161.240 90.940 162.070 ;
        RECT 92.420 160.500 92.770 161.750 ;
        RECT 96.120 161.240 96.460 162.070 ;
        RECT 97.940 160.500 98.290 161.750 ;
        RECT 101.640 161.240 101.980 162.070 ;
        RECT 105.575 161.845 108.165 162.615 ;
        RECT 108.795 161.890 109.085 162.615 ;
        RECT 109.255 162.070 114.600 162.615 ;
        RECT 114.775 162.070 120.120 162.615 ;
        RECT 120.295 162.070 125.640 162.615 ;
        RECT 103.460 160.500 103.810 161.750 ;
        RECT 105.575 161.325 106.785 161.845 ;
        RECT 106.955 161.155 108.165 161.675 ;
        RECT 110.840 161.240 111.180 162.070 ;
        RECT 83.495 160.065 88.840 160.500 ;
        RECT 89.015 160.065 94.360 160.500 ;
        RECT 94.535 160.065 99.880 160.500 ;
        RECT 100.055 160.065 105.400 160.500 ;
        RECT 105.575 160.065 108.165 161.155 ;
        RECT 108.795 160.065 109.085 161.230 ;
        RECT 112.660 160.500 113.010 161.750 ;
        RECT 116.360 161.240 116.700 162.070 ;
        RECT 118.180 160.500 118.530 161.750 ;
        RECT 121.880 161.240 122.220 162.070 ;
        RECT 125.815 161.845 129.325 162.615 ;
        RECT 129.955 161.865 131.165 162.615 ;
        RECT 123.700 160.500 124.050 161.750 ;
        RECT 125.815 161.325 127.465 161.845 ;
        RECT 127.635 161.155 129.325 161.675 ;
        RECT 109.255 160.065 114.600 160.500 ;
        RECT 114.775 160.065 120.120 160.500 ;
        RECT 120.295 160.065 125.640 160.500 ;
        RECT 125.815 160.065 129.325 161.155 ;
        RECT 129.955 161.155 130.475 161.695 ;
        RECT 130.645 161.325 131.165 161.865 ;
        RECT 129.955 160.065 131.165 161.155 ;
        RECT 57.190 159.895 131.250 160.065 ;
        RECT 57.275 158.805 58.485 159.895 ;
        RECT 58.655 159.460 64.000 159.895 ;
        RECT 64.175 159.460 69.520 159.895 ;
        RECT 57.275 158.095 57.795 158.635 ;
        RECT 57.965 158.265 58.485 158.805 ;
        RECT 57.275 157.345 58.485 158.095 ;
        RECT 60.240 157.890 60.580 158.720 ;
        RECT 62.060 158.210 62.410 159.460 ;
        RECT 65.760 157.890 66.100 158.720 ;
        RECT 67.580 158.210 67.930 159.460 ;
        RECT 70.155 158.730 70.445 159.895 ;
        RECT 70.615 159.460 75.960 159.895 ;
        RECT 76.135 159.460 81.480 159.895 ;
        RECT 81.655 159.460 87.000 159.895 ;
        RECT 87.175 159.460 92.520 159.895 ;
        RECT 58.655 157.345 64.000 157.890 ;
        RECT 64.175 157.345 69.520 157.890 ;
        RECT 70.155 157.345 70.445 158.070 ;
        RECT 72.200 157.890 72.540 158.720 ;
        RECT 74.020 158.210 74.370 159.460 ;
        RECT 77.720 157.890 78.060 158.720 ;
        RECT 79.540 158.210 79.890 159.460 ;
        RECT 83.240 157.890 83.580 158.720 ;
        RECT 85.060 158.210 85.410 159.460 ;
        RECT 88.760 157.890 89.100 158.720 ;
        RECT 90.580 158.210 90.930 159.460 ;
        RECT 92.695 158.805 95.285 159.895 ;
        RECT 92.695 158.115 93.905 158.635 ;
        RECT 94.075 158.285 95.285 158.805 ;
        RECT 95.915 158.730 96.205 159.895 ;
        RECT 96.375 159.460 101.720 159.895 ;
        RECT 101.895 159.460 107.240 159.895 ;
        RECT 107.415 159.460 112.760 159.895 ;
        RECT 112.935 159.460 118.280 159.895 ;
        RECT 70.615 157.345 75.960 157.890 ;
        RECT 76.135 157.345 81.480 157.890 ;
        RECT 81.655 157.345 87.000 157.890 ;
        RECT 87.175 157.345 92.520 157.890 ;
        RECT 92.695 157.345 95.285 158.115 ;
        RECT 95.915 157.345 96.205 158.070 ;
        RECT 97.960 157.890 98.300 158.720 ;
        RECT 99.780 158.210 100.130 159.460 ;
        RECT 103.480 157.890 103.820 158.720 ;
        RECT 105.300 158.210 105.650 159.460 ;
        RECT 109.000 157.890 109.340 158.720 ;
        RECT 110.820 158.210 111.170 159.460 ;
        RECT 114.520 157.890 114.860 158.720 ;
        RECT 116.340 158.210 116.690 159.460 ;
        RECT 118.455 158.805 121.045 159.895 ;
        RECT 118.455 158.115 119.665 158.635 ;
        RECT 119.835 158.285 121.045 158.805 ;
        RECT 121.675 158.730 121.965 159.895 ;
        RECT 122.135 159.460 127.480 159.895 ;
        RECT 96.375 157.345 101.720 157.890 ;
        RECT 101.895 157.345 107.240 157.890 ;
        RECT 107.415 157.345 112.760 157.890 ;
        RECT 112.935 157.345 118.280 157.890 ;
        RECT 118.455 157.345 121.045 158.115 ;
        RECT 121.675 157.345 121.965 158.070 ;
        RECT 123.720 157.890 124.060 158.720 ;
        RECT 125.540 158.210 125.890 159.460 ;
        RECT 127.655 158.805 129.325 159.895 ;
        RECT 127.655 158.115 128.405 158.635 ;
        RECT 128.575 158.285 129.325 158.805 ;
        RECT 129.955 158.805 131.165 159.895 ;
        RECT 129.955 158.265 130.475 158.805 ;
        RECT 122.135 157.345 127.480 157.890 ;
        RECT 127.655 157.345 129.325 158.115 ;
        RECT 130.645 158.095 131.165 158.635 ;
        RECT 129.955 157.345 131.165 158.095 ;
        RECT 57.190 157.175 131.250 157.345 ;
        RECT 57.275 156.425 58.485 157.175 ;
        RECT 58.655 156.630 64.000 157.175 ;
        RECT 64.175 156.630 69.520 157.175 ;
        RECT 69.695 156.630 75.040 157.175 ;
        RECT 75.215 156.630 80.560 157.175 ;
        RECT 57.275 155.885 57.795 156.425 ;
        RECT 57.965 155.715 58.485 156.255 ;
        RECT 60.240 155.800 60.580 156.630 ;
        RECT 57.275 154.625 58.485 155.715 ;
        RECT 62.060 155.060 62.410 156.310 ;
        RECT 65.760 155.800 66.100 156.630 ;
        RECT 67.580 155.060 67.930 156.310 ;
        RECT 71.280 155.800 71.620 156.630 ;
        RECT 73.100 155.060 73.450 156.310 ;
        RECT 76.800 155.800 77.140 156.630 ;
        RECT 80.735 156.405 82.405 157.175 ;
        RECT 83.035 156.450 83.325 157.175 ;
        RECT 83.495 156.630 88.840 157.175 ;
        RECT 89.015 156.630 94.360 157.175 ;
        RECT 94.535 156.630 99.880 157.175 ;
        RECT 100.055 156.630 105.400 157.175 ;
        RECT 78.620 155.060 78.970 156.310 ;
        RECT 80.735 155.885 81.485 156.405 ;
        RECT 81.655 155.715 82.405 156.235 ;
        RECT 85.080 155.800 85.420 156.630 ;
        RECT 58.655 154.625 64.000 155.060 ;
        RECT 64.175 154.625 69.520 155.060 ;
        RECT 69.695 154.625 75.040 155.060 ;
        RECT 75.215 154.625 80.560 155.060 ;
        RECT 80.735 154.625 82.405 155.715 ;
        RECT 83.035 154.625 83.325 155.790 ;
        RECT 86.900 155.060 87.250 156.310 ;
        RECT 90.600 155.800 90.940 156.630 ;
        RECT 92.420 155.060 92.770 156.310 ;
        RECT 96.120 155.800 96.460 156.630 ;
        RECT 97.940 155.060 98.290 156.310 ;
        RECT 101.640 155.800 101.980 156.630 ;
        RECT 105.575 156.405 108.165 157.175 ;
        RECT 108.795 156.450 109.085 157.175 ;
        RECT 109.255 156.630 114.600 157.175 ;
        RECT 114.775 156.630 120.120 157.175 ;
        RECT 120.295 156.630 125.640 157.175 ;
        RECT 103.460 155.060 103.810 156.310 ;
        RECT 105.575 155.885 106.785 156.405 ;
        RECT 106.955 155.715 108.165 156.235 ;
        RECT 110.840 155.800 111.180 156.630 ;
        RECT 83.495 154.625 88.840 155.060 ;
        RECT 89.015 154.625 94.360 155.060 ;
        RECT 94.535 154.625 99.880 155.060 ;
        RECT 100.055 154.625 105.400 155.060 ;
        RECT 105.575 154.625 108.165 155.715 ;
        RECT 108.795 154.625 109.085 155.790 ;
        RECT 112.660 155.060 113.010 156.310 ;
        RECT 116.360 155.800 116.700 156.630 ;
        RECT 118.180 155.060 118.530 156.310 ;
        RECT 121.880 155.800 122.220 156.630 ;
        RECT 125.815 156.405 129.325 157.175 ;
        RECT 129.955 156.425 131.165 157.175 ;
        RECT 123.700 155.060 124.050 156.310 ;
        RECT 125.815 155.885 127.465 156.405 ;
        RECT 127.635 155.715 129.325 156.235 ;
        RECT 109.255 154.625 114.600 155.060 ;
        RECT 114.775 154.625 120.120 155.060 ;
        RECT 120.295 154.625 125.640 155.060 ;
        RECT 125.815 154.625 129.325 155.715 ;
        RECT 129.955 155.715 130.475 156.255 ;
        RECT 130.645 155.885 131.165 156.425 ;
        RECT 129.955 154.625 131.165 155.715 ;
        RECT 57.190 154.455 131.250 154.625 ;
        RECT 57.275 153.365 58.485 154.455 ;
        RECT 58.655 154.020 64.000 154.455 ;
        RECT 64.175 154.020 69.520 154.455 ;
        RECT 57.275 152.655 57.795 153.195 ;
        RECT 57.965 152.825 58.485 153.365 ;
        RECT 57.275 151.905 58.485 152.655 ;
        RECT 60.240 152.450 60.580 153.280 ;
        RECT 62.060 152.770 62.410 154.020 ;
        RECT 65.760 152.450 66.100 153.280 ;
        RECT 67.580 152.770 67.930 154.020 ;
        RECT 70.155 153.290 70.445 154.455 ;
        RECT 70.615 154.020 75.960 154.455 ;
        RECT 76.135 154.020 81.480 154.455 ;
        RECT 81.655 154.020 87.000 154.455 ;
        RECT 87.175 154.020 92.520 154.455 ;
        RECT 58.655 151.905 64.000 152.450 ;
        RECT 64.175 151.905 69.520 152.450 ;
        RECT 70.155 151.905 70.445 152.630 ;
        RECT 72.200 152.450 72.540 153.280 ;
        RECT 74.020 152.770 74.370 154.020 ;
        RECT 77.720 152.450 78.060 153.280 ;
        RECT 79.540 152.770 79.890 154.020 ;
        RECT 83.240 152.450 83.580 153.280 ;
        RECT 85.060 152.770 85.410 154.020 ;
        RECT 88.760 152.450 89.100 153.280 ;
        RECT 90.580 152.770 90.930 154.020 ;
        RECT 92.695 153.365 95.285 154.455 ;
        RECT 92.695 152.675 93.905 153.195 ;
        RECT 94.075 152.845 95.285 153.365 ;
        RECT 95.915 153.290 96.205 154.455 ;
        RECT 96.375 154.020 101.720 154.455 ;
        RECT 101.895 154.020 107.240 154.455 ;
        RECT 107.415 154.020 112.760 154.455 ;
        RECT 112.935 154.020 118.280 154.455 ;
        RECT 70.615 151.905 75.960 152.450 ;
        RECT 76.135 151.905 81.480 152.450 ;
        RECT 81.655 151.905 87.000 152.450 ;
        RECT 87.175 151.905 92.520 152.450 ;
        RECT 92.695 151.905 95.285 152.675 ;
        RECT 95.915 151.905 96.205 152.630 ;
        RECT 97.960 152.450 98.300 153.280 ;
        RECT 99.780 152.770 100.130 154.020 ;
        RECT 103.480 152.450 103.820 153.280 ;
        RECT 105.300 152.770 105.650 154.020 ;
        RECT 109.000 152.450 109.340 153.280 ;
        RECT 110.820 152.770 111.170 154.020 ;
        RECT 114.520 152.450 114.860 153.280 ;
        RECT 116.340 152.770 116.690 154.020 ;
        RECT 118.455 153.365 121.045 154.455 ;
        RECT 118.455 152.675 119.665 153.195 ;
        RECT 119.835 152.845 121.045 153.365 ;
        RECT 121.675 153.290 121.965 154.455 ;
        RECT 122.135 154.020 127.480 154.455 ;
        RECT 96.375 151.905 101.720 152.450 ;
        RECT 101.895 151.905 107.240 152.450 ;
        RECT 107.415 151.905 112.760 152.450 ;
        RECT 112.935 151.905 118.280 152.450 ;
        RECT 118.455 151.905 121.045 152.675 ;
        RECT 121.675 151.905 121.965 152.630 ;
        RECT 123.720 152.450 124.060 153.280 ;
        RECT 125.540 152.770 125.890 154.020 ;
        RECT 127.655 153.365 129.325 154.455 ;
        RECT 127.655 152.675 128.405 153.195 ;
        RECT 128.575 152.845 129.325 153.365 ;
        RECT 129.955 153.365 131.165 154.455 ;
        RECT 129.955 152.825 130.475 153.365 ;
        RECT 122.135 151.905 127.480 152.450 ;
        RECT 127.655 151.905 129.325 152.675 ;
        RECT 130.645 152.655 131.165 153.195 ;
        RECT 129.955 151.905 131.165 152.655 ;
        RECT 57.190 151.735 131.250 151.905 ;
        RECT 57.275 150.985 58.485 151.735 ;
        RECT 58.655 151.190 64.000 151.735 ;
        RECT 64.175 151.190 69.520 151.735 ;
        RECT 69.695 151.190 75.040 151.735 ;
        RECT 75.215 151.190 80.560 151.735 ;
        RECT 57.275 150.445 57.795 150.985 ;
        RECT 57.965 150.275 58.485 150.815 ;
        RECT 60.240 150.360 60.580 151.190 ;
        RECT 57.275 149.185 58.485 150.275 ;
        RECT 62.060 149.620 62.410 150.870 ;
        RECT 65.760 150.360 66.100 151.190 ;
        RECT 67.580 149.620 67.930 150.870 ;
        RECT 71.280 150.360 71.620 151.190 ;
        RECT 73.100 149.620 73.450 150.870 ;
        RECT 76.800 150.360 77.140 151.190 ;
        RECT 80.735 150.965 82.405 151.735 ;
        RECT 83.035 151.010 83.325 151.735 ;
        RECT 83.495 151.190 88.840 151.735 ;
        RECT 89.015 151.190 94.360 151.735 ;
        RECT 94.535 151.190 99.880 151.735 ;
        RECT 100.055 151.190 105.400 151.735 ;
        RECT 78.620 149.620 78.970 150.870 ;
        RECT 80.735 150.445 81.485 150.965 ;
        RECT 81.655 150.275 82.405 150.795 ;
        RECT 85.080 150.360 85.420 151.190 ;
        RECT 58.655 149.185 64.000 149.620 ;
        RECT 64.175 149.185 69.520 149.620 ;
        RECT 69.695 149.185 75.040 149.620 ;
        RECT 75.215 149.185 80.560 149.620 ;
        RECT 80.735 149.185 82.405 150.275 ;
        RECT 83.035 149.185 83.325 150.350 ;
        RECT 86.900 149.620 87.250 150.870 ;
        RECT 90.600 150.360 90.940 151.190 ;
        RECT 92.420 149.620 92.770 150.870 ;
        RECT 96.120 150.360 96.460 151.190 ;
        RECT 97.940 149.620 98.290 150.870 ;
        RECT 101.640 150.360 101.980 151.190 ;
        RECT 105.575 150.965 108.165 151.735 ;
        RECT 108.795 151.010 109.085 151.735 ;
        RECT 109.315 151.255 109.595 151.735 ;
        RECT 109.765 151.085 110.025 151.475 ;
        RECT 110.200 151.255 110.455 151.735 ;
        RECT 110.625 151.085 110.920 151.475 ;
        RECT 111.100 151.255 111.375 151.735 ;
        RECT 111.545 151.235 111.845 151.565 ;
        RECT 103.460 149.620 103.810 150.870 ;
        RECT 105.575 150.445 106.785 150.965 ;
        RECT 109.270 150.915 110.920 151.085 ;
        RECT 106.955 150.275 108.165 150.795 ;
        RECT 109.270 150.405 109.675 150.915 ;
        RECT 109.845 150.575 110.985 150.745 ;
        RECT 83.495 149.185 88.840 149.620 ;
        RECT 89.015 149.185 94.360 149.620 ;
        RECT 94.535 149.185 99.880 149.620 ;
        RECT 100.055 149.185 105.400 149.620 ;
        RECT 105.575 149.185 108.165 150.275 ;
        RECT 108.795 149.185 109.085 150.350 ;
        RECT 109.270 150.235 110.025 150.405 ;
        RECT 109.310 149.185 109.595 150.055 ;
        RECT 109.765 149.985 110.025 150.235 ;
        RECT 110.815 150.325 110.985 150.575 ;
        RECT 111.155 150.495 111.505 151.065 ;
        RECT 111.675 150.325 111.845 151.235 ;
        RECT 112.015 151.190 117.360 151.735 ;
        RECT 117.535 151.190 122.880 151.735 ;
        RECT 123.055 151.190 128.400 151.735 ;
        RECT 113.600 150.360 113.940 151.190 ;
        RECT 110.815 150.155 111.845 150.325 ;
        RECT 109.765 149.815 110.885 149.985 ;
        RECT 109.765 149.355 110.025 149.815 ;
        RECT 110.200 149.185 110.455 149.645 ;
        RECT 110.625 149.355 110.885 149.815 ;
        RECT 111.055 149.185 111.365 149.985 ;
        RECT 111.535 149.355 111.845 150.155 ;
        RECT 115.420 149.620 115.770 150.870 ;
        RECT 119.120 150.360 119.460 151.190 ;
        RECT 120.940 149.620 121.290 150.870 ;
        RECT 124.640 150.360 124.980 151.190 ;
        RECT 128.575 150.985 129.785 151.735 ;
        RECT 129.955 150.985 131.165 151.735 ;
        RECT 126.460 149.620 126.810 150.870 ;
        RECT 128.575 150.445 129.095 150.985 ;
        RECT 129.265 150.275 129.785 150.815 ;
        RECT 112.015 149.185 117.360 149.620 ;
        RECT 117.535 149.185 122.880 149.620 ;
        RECT 123.055 149.185 128.400 149.620 ;
        RECT 128.575 149.185 129.785 150.275 ;
        RECT 129.955 150.275 130.475 150.815 ;
        RECT 130.645 150.445 131.165 150.985 ;
        RECT 129.955 149.185 131.165 150.275 ;
        RECT 57.190 149.015 131.250 149.185 ;
        RECT 57.275 147.925 58.485 149.015 ;
        RECT 58.655 148.580 64.000 149.015 ;
        RECT 64.175 148.580 69.520 149.015 ;
        RECT 57.275 147.215 57.795 147.755 ;
        RECT 57.965 147.385 58.485 147.925 ;
        RECT 57.275 146.465 58.485 147.215 ;
        RECT 60.240 147.010 60.580 147.840 ;
        RECT 62.060 147.330 62.410 148.580 ;
        RECT 65.760 147.010 66.100 147.840 ;
        RECT 67.580 147.330 67.930 148.580 ;
        RECT 70.155 147.850 70.445 149.015 ;
        RECT 70.615 148.580 75.960 149.015 ;
        RECT 76.135 148.580 81.480 149.015 ;
        RECT 81.655 148.580 87.000 149.015 ;
        RECT 87.175 148.580 92.520 149.015 ;
        RECT 58.655 146.465 64.000 147.010 ;
        RECT 64.175 146.465 69.520 147.010 ;
        RECT 70.155 146.465 70.445 147.190 ;
        RECT 72.200 147.010 72.540 147.840 ;
        RECT 74.020 147.330 74.370 148.580 ;
        RECT 77.720 147.010 78.060 147.840 ;
        RECT 79.540 147.330 79.890 148.580 ;
        RECT 83.240 147.010 83.580 147.840 ;
        RECT 85.060 147.330 85.410 148.580 ;
        RECT 88.760 147.010 89.100 147.840 ;
        RECT 90.580 147.330 90.930 148.580 ;
        RECT 92.695 147.925 95.285 149.015 ;
        RECT 92.695 147.235 93.905 147.755 ;
        RECT 94.075 147.405 95.285 147.925 ;
        RECT 95.915 147.850 96.205 149.015 ;
        RECT 96.375 148.580 101.720 149.015 ;
        RECT 101.895 148.580 107.240 149.015 ;
        RECT 107.415 148.580 112.760 149.015 ;
        RECT 112.935 148.580 118.280 149.015 ;
        RECT 70.615 146.465 75.960 147.010 ;
        RECT 76.135 146.465 81.480 147.010 ;
        RECT 81.655 146.465 87.000 147.010 ;
        RECT 87.175 146.465 92.520 147.010 ;
        RECT 92.695 146.465 95.285 147.235 ;
        RECT 95.915 146.465 96.205 147.190 ;
        RECT 97.960 147.010 98.300 147.840 ;
        RECT 99.780 147.330 100.130 148.580 ;
        RECT 103.480 147.010 103.820 147.840 ;
        RECT 105.300 147.330 105.650 148.580 ;
        RECT 109.000 147.010 109.340 147.840 ;
        RECT 110.820 147.330 111.170 148.580 ;
        RECT 114.520 147.010 114.860 147.840 ;
        RECT 116.340 147.330 116.690 148.580 ;
        RECT 118.455 147.925 121.045 149.015 ;
        RECT 118.455 147.235 119.665 147.755 ;
        RECT 119.835 147.405 121.045 147.925 ;
        RECT 121.675 147.850 121.965 149.015 ;
        RECT 122.135 148.580 127.480 149.015 ;
        RECT 96.375 146.465 101.720 147.010 ;
        RECT 101.895 146.465 107.240 147.010 ;
        RECT 107.415 146.465 112.760 147.010 ;
        RECT 112.935 146.465 118.280 147.010 ;
        RECT 118.455 146.465 121.045 147.235 ;
        RECT 121.675 146.465 121.965 147.190 ;
        RECT 123.720 147.010 124.060 147.840 ;
        RECT 125.540 147.330 125.890 148.580 ;
        RECT 127.655 147.925 129.325 149.015 ;
        RECT 127.655 147.235 128.405 147.755 ;
        RECT 128.575 147.405 129.325 147.925 ;
        RECT 129.955 147.925 131.165 149.015 ;
        RECT 129.955 147.385 130.475 147.925 ;
        RECT 122.135 146.465 127.480 147.010 ;
        RECT 127.655 146.465 129.325 147.235 ;
        RECT 130.645 147.215 131.165 147.755 ;
        RECT 129.955 146.465 131.165 147.215 ;
        RECT 57.190 146.295 131.250 146.465 ;
        RECT 57.275 145.545 58.485 146.295 ;
        RECT 58.655 145.750 64.000 146.295 ;
        RECT 64.175 145.750 69.520 146.295 ;
        RECT 69.695 145.750 75.040 146.295 ;
        RECT 75.215 145.750 80.560 146.295 ;
        RECT 57.275 145.005 57.795 145.545 ;
        RECT 57.965 144.835 58.485 145.375 ;
        RECT 60.240 144.920 60.580 145.750 ;
        RECT 57.275 143.745 58.485 144.835 ;
        RECT 62.060 144.180 62.410 145.430 ;
        RECT 65.760 144.920 66.100 145.750 ;
        RECT 67.580 144.180 67.930 145.430 ;
        RECT 71.280 144.920 71.620 145.750 ;
        RECT 73.100 144.180 73.450 145.430 ;
        RECT 76.800 144.920 77.140 145.750 ;
        RECT 80.735 145.525 82.405 146.295 ;
        RECT 83.035 145.570 83.325 146.295 ;
        RECT 83.495 145.750 88.840 146.295 ;
        RECT 89.015 145.750 94.360 146.295 ;
        RECT 94.535 145.750 99.880 146.295 ;
        RECT 100.055 145.750 105.400 146.295 ;
        RECT 78.620 144.180 78.970 145.430 ;
        RECT 80.735 145.005 81.485 145.525 ;
        RECT 81.655 144.835 82.405 145.355 ;
        RECT 85.080 144.920 85.420 145.750 ;
        RECT 58.655 143.745 64.000 144.180 ;
        RECT 64.175 143.745 69.520 144.180 ;
        RECT 69.695 143.745 75.040 144.180 ;
        RECT 75.215 143.745 80.560 144.180 ;
        RECT 80.735 143.745 82.405 144.835 ;
        RECT 83.035 143.745 83.325 144.910 ;
        RECT 86.900 144.180 87.250 145.430 ;
        RECT 90.600 144.920 90.940 145.750 ;
        RECT 92.420 144.180 92.770 145.430 ;
        RECT 96.120 144.920 96.460 145.750 ;
        RECT 97.940 144.180 98.290 145.430 ;
        RECT 101.640 144.920 101.980 145.750 ;
        RECT 105.575 145.525 108.165 146.295 ;
        RECT 108.795 145.570 109.085 146.295 ;
        RECT 109.255 145.750 114.600 146.295 ;
        RECT 114.775 145.750 120.120 146.295 ;
        RECT 120.295 145.750 125.640 146.295 ;
        RECT 103.460 144.180 103.810 145.430 ;
        RECT 105.575 145.005 106.785 145.525 ;
        RECT 106.955 144.835 108.165 145.355 ;
        RECT 110.840 144.920 111.180 145.750 ;
        RECT 83.495 143.745 88.840 144.180 ;
        RECT 89.015 143.745 94.360 144.180 ;
        RECT 94.535 143.745 99.880 144.180 ;
        RECT 100.055 143.745 105.400 144.180 ;
        RECT 105.575 143.745 108.165 144.835 ;
        RECT 108.795 143.745 109.085 144.910 ;
        RECT 112.660 144.180 113.010 145.430 ;
        RECT 116.360 144.920 116.700 145.750 ;
        RECT 118.180 144.180 118.530 145.430 ;
        RECT 121.880 144.920 122.220 145.750 ;
        RECT 125.815 145.525 129.325 146.295 ;
        RECT 129.955 145.545 131.165 146.295 ;
        RECT 123.700 144.180 124.050 145.430 ;
        RECT 125.815 145.005 127.465 145.525 ;
        RECT 127.635 144.835 129.325 145.355 ;
        RECT 109.255 143.745 114.600 144.180 ;
        RECT 114.775 143.745 120.120 144.180 ;
        RECT 120.295 143.745 125.640 144.180 ;
        RECT 125.815 143.745 129.325 144.835 ;
        RECT 129.955 144.835 130.475 145.375 ;
        RECT 130.645 145.005 131.165 145.545 ;
        RECT 129.955 143.745 131.165 144.835 ;
        RECT 57.190 143.575 131.250 143.745 ;
        RECT 57.275 142.485 58.485 143.575 ;
        RECT 58.655 143.140 64.000 143.575 ;
        RECT 64.175 143.140 69.520 143.575 ;
        RECT 57.275 141.775 57.795 142.315 ;
        RECT 57.965 141.945 58.485 142.485 ;
        RECT 57.275 141.025 58.485 141.775 ;
        RECT 60.240 141.570 60.580 142.400 ;
        RECT 62.060 141.890 62.410 143.140 ;
        RECT 65.760 141.570 66.100 142.400 ;
        RECT 67.580 141.890 67.930 143.140 ;
        RECT 70.155 142.410 70.445 143.575 ;
        RECT 70.615 143.140 75.960 143.575 ;
        RECT 76.135 143.140 81.480 143.575 ;
        RECT 81.655 143.140 87.000 143.575 ;
        RECT 87.175 143.140 92.520 143.575 ;
        RECT 58.655 141.025 64.000 141.570 ;
        RECT 64.175 141.025 69.520 141.570 ;
        RECT 70.155 141.025 70.445 141.750 ;
        RECT 72.200 141.570 72.540 142.400 ;
        RECT 74.020 141.890 74.370 143.140 ;
        RECT 77.720 141.570 78.060 142.400 ;
        RECT 79.540 141.890 79.890 143.140 ;
        RECT 83.240 141.570 83.580 142.400 ;
        RECT 85.060 141.890 85.410 143.140 ;
        RECT 88.760 141.570 89.100 142.400 ;
        RECT 90.580 141.890 90.930 143.140 ;
        RECT 92.695 142.485 95.285 143.575 ;
        RECT 92.695 141.795 93.905 142.315 ;
        RECT 94.075 141.965 95.285 142.485 ;
        RECT 95.915 142.410 96.205 143.575 ;
        RECT 96.375 143.140 101.720 143.575 ;
        RECT 101.895 143.140 107.240 143.575 ;
        RECT 107.415 143.140 112.760 143.575 ;
        RECT 112.935 143.140 118.280 143.575 ;
        RECT 70.615 141.025 75.960 141.570 ;
        RECT 76.135 141.025 81.480 141.570 ;
        RECT 81.655 141.025 87.000 141.570 ;
        RECT 87.175 141.025 92.520 141.570 ;
        RECT 92.695 141.025 95.285 141.795 ;
        RECT 95.915 141.025 96.205 141.750 ;
        RECT 97.960 141.570 98.300 142.400 ;
        RECT 99.780 141.890 100.130 143.140 ;
        RECT 103.480 141.570 103.820 142.400 ;
        RECT 105.300 141.890 105.650 143.140 ;
        RECT 109.000 141.570 109.340 142.400 ;
        RECT 110.820 141.890 111.170 143.140 ;
        RECT 114.520 141.570 114.860 142.400 ;
        RECT 116.340 141.890 116.690 143.140 ;
        RECT 118.455 142.485 121.045 143.575 ;
        RECT 118.455 141.795 119.665 142.315 ;
        RECT 119.835 141.965 121.045 142.485 ;
        RECT 121.675 142.410 121.965 143.575 ;
        RECT 122.135 143.140 127.480 143.575 ;
        RECT 96.375 141.025 101.720 141.570 ;
        RECT 101.895 141.025 107.240 141.570 ;
        RECT 107.415 141.025 112.760 141.570 ;
        RECT 112.935 141.025 118.280 141.570 ;
        RECT 118.455 141.025 121.045 141.795 ;
        RECT 121.675 141.025 121.965 141.750 ;
        RECT 123.720 141.570 124.060 142.400 ;
        RECT 125.540 141.890 125.890 143.140 ;
        RECT 127.655 142.485 129.325 143.575 ;
        RECT 127.655 141.795 128.405 142.315 ;
        RECT 128.575 141.965 129.325 142.485 ;
        RECT 129.955 142.485 131.165 143.575 ;
        RECT 129.955 141.945 130.475 142.485 ;
        RECT 122.135 141.025 127.480 141.570 ;
        RECT 127.655 141.025 129.325 141.795 ;
        RECT 130.645 141.775 131.165 142.315 ;
        RECT 129.955 141.025 131.165 141.775 ;
        RECT 57.190 140.855 131.250 141.025 ;
        RECT 57.275 140.105 58.485 140.855 ;
        RECT 58.655 140.310 64.000 140.855 ;
        RECT 64.175 140.310 69.520 140.855 ;
        RECT 69.695 140.310 75.040 140.855 ;
        RECT 75.215 140.310 80.560 140.855 ;
        RECT 57.275 139.565 57.795 140.105 ;
        RECT 57.965 139.395 58.485 139.935 ;
        RECT 60.240 139.480 60.580 140.310 ;
        RECT 57.275 138.305 58.485 139.395 ;
        RECT 62.060 138.740 62.410 139.990 ;
        RECT 65.760 139.480 66.100 140.310 ;
        RECT 67.580 138.740 67.930 139.990 ;
        RECT 71.280 139.480 71.620 140.310 ;
        RECT 73.100 138.740 73.450 139.990 ;
        RECT 76.800 139.480 77.140 140.310 ;
        RECT 80.735 140.085 82.405 140.855 ;
        RECT 83.035 140.130 83.325 140.855 ;
        RECT 83.495 140.310 88.840 140.855 ;
        RECT 89.015 140.310 94.360 140.855 ;
        RECT 94.535 140.310 99.880 140.855 ;
        RECT 100.055 140.310 105.400 140.855 ;
        RECT 78.620 138.740 78.970 139.990 ;
        RECT 80.735 139.565 81.485 140.085 ;
        RECT 81.655 139.395 82.405 139.915 ;
        RECT 85.080 139.480 85.420 140.310 ;
        RECT 58.655 138.305 64.000 138.740 ;
        RECT 64.175 138.305 69.520 138.740 ;
        RECT 69.695 138.305 75.040 138.740 ;
        RECT 75.215 138.305 80.560 138.740 ;
        RECT 80.735 138.305 82.405 139.395 ;
        RECT 83.035 138.305 83.325 139.470 ;
        RECT 86.900 138.740 87.250 139.990 ;
        RECT 90.600 139.480 90.940 140.310 ;
        RECT 92.420 138.740 92.770 139.990 ;
        RECT 96.120 139.480 96.460 140.310 ;
        RECT 97.940 138.740 98.290 139.990 ;
        RECT 101.640 139.480 101.980 140.310 ;
        RECT 105.575 140.085 108.165 140.855 ;
        RECT 108.795 140.130 109.085 140.855 ;
        RECT 109.255 140.310 114.600 140.855 ;
        RECT 114.775 140.310 120.120 140.855 ;
        RECT 120.295 140.310 125.640 140.855 ;
        RECT 103.460 138.740 103.810 139.990 ;
        RECT 105.575 139.565 106.785 140.085 ;
        RECT 106.955 139.395 108.165 139.915 ;
        RECT 110.840 139.480 111.180 140.310 ;
        RECT 83.495 138.305 88.840 138.740 ;
        RECT 89.015 138.305 94.360 138.740 ;
        RECT 94.535 138.305 99.880 138.740 ;
        RECT 100.055 138.305 105.400 138.740 ;
        RECT 105.575 138.305 108.165 139.395 ;
        RECT 108.795 138.305 109.085 139.470 ;
        RECT 112.660 138.740 113.010 139.990 ;
        RECT 116.360 139.480 116.700 140.310 ;
        RECT 118.180 138.740 118.530 139.990 ;
        RECT 121.880 139.480 122.220 140.310 ;
        RECT 125.815 140.085 129.325 140.855 ;
        RECT 129.955 140.105 131.165 140.855 ;
        RECT 123.700 138.740 124.050 139.990 ;
        RECT 125.815 139.565 127.465 140.085 ;
        RECT 127.635 139.395 129.325 139.915 ;
        RECT 109.255 138.305 114.600 138.740 ;
        RECT 114.775 138.305 120.120 138.740 ;
        RECT 120.295 138.305 125.640 138.740 ;
        RECT 125.815 138.305 129.325 139.395 ;
        RECT 129.955 139.395 130.475 139.935 ;
        RECT 130.645 139.565 131.165 140.105 ;
        RECT 129.955 138.305 131.165 139.395 ;
        RECT 57.190 138.135 131.250 138.305 ;
        RECT 57.275 137.045 58.485 138.135 ;
        RECT 58.655 137.700 64.000 138.135 ;
        RECT 64.175 137.700 69.520 138.135 ;
        RECT 57.275 136.335 57.795 136.875 ;
        RECT 57.965 136.505 58.485 137.045 ;
        RECT 57.275 135.585 58.485 136.335 ;
        RECT 60.240 136.130 60.580 136.960 ;
        RECT 62.060 136.450 62.410 137.700 ;
        RECT 65.760 136.130 66.100 136.960 ;
        RECT 67.580 136.450 67.930 137.700 ;
        RECT 70.155 136.970 70.445 138.135 ;
        RECT 70.615 137.700 75.960 138.135 ;
        RECT 76.135 137.700 81.480 138.135 ;
        RECT 81.655 137.700 87.000 138.135 ;
        RECT 87.175 137.700 92.520 138.135 ;
        RECT 58.655 135.585 64.000 136.130 ;
        RECT 64.175 135.585 69.520 136.130 ;
        RECT 70.155 135.585 70.445 136.310 ;
        RECT 72.200 136.130 72.540 136.960 ;
        RECT 74.020 136.450 74.370 137.700 ;
        RECT 77.720 136.130 78.060 136.960 ;
        RECT 79.540 136.450 79.890 137.700 ;
        RECT 83.240 136.130 83.580 136.960 ;
        RECT 85.060 136.450 85.410 137.700 ;
        RECT 88.760 136.130 89.100 136.960 ;
        RECT 90.580 136.450 90.930 137.700 ;
        RECT 92.695 137.045 95.285 138.135 ;
        RECT 92.695 136.355 93.905 136.875 ;
        RECT 94.075 136.525 95.285 137.045 ;
        RECT 95.915 136.970 96.205 138.135 ;
        RECT 96.375 137.700 101.720 138.135 ;
        RECT 101.895 137.700 107.240 138.135 ;
        RECT 107.415 137.700 112.760 138.135 ;
        RECT 112.935 137.700 118.280 138.135 ;
        RECT 70.615 135.585 75.960 136.130 ;
        RECT 76.135 135.585 81.480 136.130 ;
        RECT 81.655 135.585 87.000 136.130 ;
        RECT 87.175 135.585 92.520 136.130 ;
        RECT 92.695 135.585 95.285 136.355 ;
        RECT 95.915 135.585 96.205 136.310 ;
        RECT 97.960 136.130 98.300 136.960 ;
        RECT 99.780 136.450 100.130 137.700 ;
        RECT 103.480 136.130 103.820 136.960 ;
        RECT 105.300 136.450 105.650 137.700 ;
        RECT 109.000 136.130 109.340 136.960 ;
        RECT 110.820 136.450 111.170 137.700 ;
        RECT 114.520 136.130 114.860 136.960 ;
        RECT 116.340 136.450 116.690 137.700 ;
        RECT 118.455 137.045 121.045 138.135 ;
        RECT 118.455 136.355 119.665 136.875 ;
        RECT 119.835 136.525 121.045 137.045 ;
        RECT 121.675 136.970 121.965 138.135 ;
        RECT 122.135 137.700 127.480 138.135 ;
        RECT 96.375 135.585 101.720 136.130 ;
        RECT 101.895 135.585 107.240 136.130 ;
        RECT 107.415 135.585 112.760 136.130 ;
        RECT 112.935 135.585 118.280 136.130 ;
        RECT 118.455 135.585 121.045 136.355 ;
        RECT 121.675 135.585 121.965 136.310 ;
        RECT 123.720 136.130 124.060 136.960 ;
        RECT 125.540 136.450 125.890 137.700 ;
        RECT 127.655 137.045 129.325 138.135 ;
        RECT 127.655 136.355 128.405 136.875 ;
        RECT 128.575 136.525 129.325 137.045 ;
        RECT 129.955 137.045 131.165 138.135 ;
        RECT 129.955 136.505 130.475 137.045 ;
        RECT 122.135 135.585 127.480 136.130 ;
        RECT 127.655 135.585 129.325 136.355 ;
        RECT 130.645 136.335 131.165 136.875 ;
        RECT 129.955 135.585 131.165 136.335 ;
        RECT 57.190 135.415 131.250 135.585 ;
        RECT 57.275 134.665 58.485 135.415 ;
        RECT 58.655 134.870 64.000 135.415 ;
        RECT 64.175 134.870 69.520 135.415 ;
        RECT 69.695 134.870 75.040 135.415 ;
        RECT 75.215 134.870 80.560 135.415 ;
        RECT 57.275 134.125 57.795 134.665 ;
        RECT 57.965 133.955 58.485 134.495 ;
        RECT 60.240 134.040 60.580 134.870 ;
        RECT 57.275 132.865 58.485 133.955 ;
        RECT 62.060 133.300 62.410 134.550 ;
        RECT 65.760 134.040 66.100 134.870 ;
        RECT 67.580 133.300 67.930 134.550 ;
        RECT 71.280 134.040 71.620 134.870 ;
        RECT 73.100 133.300 73.450 134.550 ;
        RECT 76.800 134.040 77.140 134.870 ;
        RECT 80.735 134.645 82.405 135.415 ;
        RECT 83.035 134.690 83.325 135.415 ;
        RECT 83.495 134.870 88.840 135.415 ;
        RECT 89.015 134.870 94.360 135.415 ;
        RECT 94.535 134.870 99.880 135.415 ;
        RECT 100.055 134.870 105.400 135.415 ;
        RECT 78.620 133.300 78.970 134.550 ;
        RECT 80.735 134.125 81.485 134.645 ;
        RECT 81.655 133.955 82.405 134.475 ;
        RECT 85.080 134.040 85.420 134.870 ;
        RECT 58.655 132.865 64.000 133.300 ;
        RECT 64.175 132.865 69.520 133.300 ;
        RECT 69.695 132.865 75.040 133.300 ;
        RECT 75.215 132.865 80.560 133.300 ;
        RECT 80.735 132.865 82.405 133.955 ;
        RECT 83.035 132.865 83.325 134.030 ;
        RECT 86.900 133.300 87.250 134.550 ;
        RECT 90.600 134.040 90.940 134.870 ;
        RECT 92.420 133.300 92.770 134.550 ;
        RECT 96.120 134.040 96.460 134.870 ;
        RECT 97.940 133.300 98.290 134.550 ;
        RECT 101.640 134.040 101.980 134.870 ;
        RECT 105.575 134.645 108.165 135.415 ;
        RECT 108.795 134.690 109.085 135.415 ;
        RECT 109.255 134.870 114.600 135.415 ;
        RECT 114.775 134.870 120.120 135.415 ;
        RECT 120.295 134.870 125.640 135.415 ;
        RECT 103.460 133.300 103.810 134.550 ;
        RECT 105.575 134.125 106.785 134.645 ;
        RECT 106.955 133.955 108.165 134.475 ;
        RECT 110.840 134.040 111.180 134.870 ;
        RECT 83.495 132.865 88.840 133.300 ;
        RECT 89.015 132.865 94.360 133.300 ;
        RECT 94.535 132.865 99.880 133.300 ;
        RECT 100.055 132.865 105.400 133.300 ;
        RECT 105.575 132.865 108.165 133.955 ;
        RECT 108.795 132.865 109.085 134.030 ;
        RECT 112.660 133.300 113.010 134.550 ;
        RECT 116.360 134.040 116.700 134.870 ;
        RECT 118.180 133.300 118.530 134.550 ;
        RECT 121.880 134.040 122.220 134.870 ;
        RECT 125.815 134.645 129.325 135.415 ;
        RECT 129.955 134.665 131.165 135.415 ;
        RECT 123.700 133.300 124.050 134.550 ;
        RECT 125.815 134.125 127.465 134.645 ;
        RECT 127.635 133.955 129.325 134.475 ;
        RECT 109.255 132.865 114.600 133.300 ;
        RECT 114.775 132.865 120.120 133.300 ;
        RECT 120.295 132.865 125.640 133.300 ;
        RECT 125.815 132.865 129.325 133.955 ;
        RECT 129.955 133.955 130.475 134.495 ;
        RECT 130.645 134.125 131.165 134.665 ;
        RECT 129.955 132.865 131.165 133.955 ;
        RECT 57.190 132.695 131.250 132.865 ;
        RECT 57.275 131.605 58.485 132.695 ;
        RECT 58.655 132.260 64.000 132.695 ;
        RECT 64.175 132.260 69.520 132.695 ;
        RECT 57.275 130.895 57.795 131.435 ;
        RECT 57.965 131.065 58.485 131.605 ;
        RECT 57.275 130.145 58.485 130.895 ;
        RECT 60.240 130.690 60.580 131.520 ;
        RECT 62.060 131.010 62.410 132.260 ;
        RECT 65.760 130.690 66.100 131.520 ;
        RECT 67.580 131.010 67.930 132.260 ;
        RECT 70.155 131.530 70.445 132.695 ;
        RECT 70.615 132.260 75.960 132.695 ;
        RECT 76.135 132.260 81.480 132.695 ;
        RECT 58.655 130.145 64.000 130.690 ;
        RECT 64.175 130.145 69.520 130.690 ;
        RECT 70.155 130.145 70.445 130.870 ;
        RECT 72.200 130.690 72.540 131.520 ;
        RECT 74.020 131.010 74.370 132.260 ;
        RECT 77.720 130.690 78.060 131.520 ;
        RECT 79.540 131.010 79.890 132.260 ;
        RECT 81.655 131.605 82.865 132.695 ;
        RECT 81.655 130.895 82.175 131.435 ;
        RECT 82.345 131.065 82.865 131.605 ;
        RECT 83.035 131.530 83.325 132.695 ;
        RECT 83.495 132.260 88.840 132.695 ;
        RECT 89.015 132.260 94.360 132.695 ;
        RECT 70.615 130.145 75.960 130.690 ;
        RECT 76.135 130.145 81.480 130.690 ;
        RECT 81.655 130.145 82.865 130.895 ;
        RECT 83.035 130.145 83.325 130.870 ;
        RECT 85.080 130.690 85.420 131.520 ;
        RECT 86.900 131.010 87.250 132.260 ;
        RECT 90.600 130.690 90.940 131.520 ;
        RECT 92.420 131.010 92.770 132.260 ;
        RECT 94.535 131.605 95.745 132.695 ;
        RECT 94.535 130.895 95.055 131.435 ;
        RECT 95.225 131.065 95.745 131.605 ;
        RECT 95.915 131.530 96.205 132.695 ;
        RECT 96.375 132.260 101.720 132.695 ;
        RECT 101.895 132.260 107.240 132.695 ;
        RECT 83.495 130.145 88.840 130.690 ;
        RECT 89.015 130.145 94.360 130.690 ;
        RECT 94.535 130.145 95.745 130.895 ;
        RECT 95.915 130.145 96.205 130.870 ;
        RECT 97.960 130.690 98.300 131.520 ;
        RECT 99.780 131.010 100.130 132.260 ;
        RECT 103.480 130.690 103.820 131.520 ;
        RECT 105.300 131.010 105.650 132.260 ;
        RECT 107.415 131.605 108.625 132.695 ;
        RECT 107.415 130.895 107.935 131.435 ;
        RECT 108.105 131.065 108.625 131.605 ;
        RECT 108.795 131.530 109.085 132.695 ;
        RECT 109.255 132.260 114.600 132.695 ;
        RECT 114.775 132.260 120.120 132.695 ;
        RECT 96.375 130.145 101.720 130.690 ;
        RECT 101.895 130.145 107.240 130.690 ;
        RECT 107.415 130.145 108.625 130.895 ;
        RECT 108.795 130.145 109.085 130.870 ;
        RECT 110.840 130.690 111.180 131.520 ;
        RECT 112.660 131.010 113.010 132.260 ;
        RECT 116.360 130.690 116.700 131.520 ;
        RECT 118.180 131.010 118.530 132.260 ;
        RECT 120.295 131.605 121.505 132.695 ;
        RECT 120.295 130.895 120.815 131.435 ;
        RECT 120.985 131.065 121.505 131.605 ;
        RECT 121.675 131.530 121.965 132.695 ;
        RECT 122.135 132.260 127.480 132.695 ;
        RECT 109.255 130.145 114.600 130.690 ;
        RECT 114.775 130.145 120.120 130.690 ;
        RECT 120.295 130.145 121.505 130.895 ;
        RECT 121.675 130.145 121.965 130.870 ;
        RECT 123.720 130.690 124.060 131.520 ;
        RECT 125.540 131.010 125.890 132.260 ;
        RECT 127.655 131.605 129.325 132.695 ;
        RECT 127.655 130.915 128.405 131.435 ;
        RECT 128.575 131.085 129.325 131.605 ;
        RECT 129.955 131.605 131.165 132.695 ;
        RECT 129.955 131.065 130.475 131.605 ;
        RECT 122.135 130.145 127.480 130.690 ;
        RECT 127.655 130.145 129.325 130.915 ;
        RECT 130.645 130.895 131.165 131.435 ;
        RECT 129.955 130.145 131.165 130.895 ;
        RECT 57.190 129.975 131.250 130.145 ;
        RECT 137.300 88.230 144.110 88.400 ;
        RECT 137.300 86.920 137.470 88.230 ;
        RECT 137.950 87.400 140.110 87.750 ;
        RECT 141.300 87.400 143.460 87.750 ;
        RECT 138.570 86.920 140.120 87.020 ;
        RECT 143.940 86.920 144.110 88.230 ;
        RECT 137.300 86.750 144.110 86.920 ;
        RECT 147.300 88.230 154.110 88.400 ;
        RECT 147.300 86.920 147.470 88.230 ;
        RECT 147.950 87.400 150.110 87.750 ;
        RECT 151.300 87.400 153.460 87.750 ;
        RECT 150.920 86.920 152.520 86.970 ;
        RECT 153.940 86.920 154.110 88.230 ;
        RECT 147.300 86.750 154.110 86.920 ;
        RECT 138.570 86.620 140.120 86.750 ;
        RECT 150.920 86.670 152.520 86.750 ;
        RECT 138.870 84.290 140.420 84.370 ;
        RECT 142.870 84.290 144.420 84.370 ;
        RECT 138.300 84.120 140.950 84.290 ;
        RECT 138.300 80.920 138.470 84.120 ;
        RECT 139.100 83.610 139.480 83.780 ;
        RECT 139.770 83.610 140.150 83.780 ;
        RECT 138.870 81.600 139.040 83.440 ;
        RECT 139.540 81.600 139.710 83.440 ;
        RECT 140.210 81.600 140.380 83.440 ;
        RECT 139.100 81.260 139.480 81.430 ;
        RECT 139.770 81.260 140.150 81.430 ;
        RECT 140.780 80.920 140.950 84.120 ;
        RECT 138.300 80.750 140.950 80.920 ;
        RECT 142.300 84.120 144.950 84.290 ;
        RECT 142.300 80.920 142.470 84.120 ;
        RECT 143.100 83.610 143.480 83.780 ;
        RECT 143.770 83.610 144.150 83.780 ;
        RECT 142.870 81.600 143.040 83.440 ;
        RECT 143.540 81.600 143.710 83.440 ;
        RECT 144.210 81.600 144.380 83.440 ;
        RECT 143.100 81.260 143.480 81.430 ;
        RECT 143.770 81.260 144.150 81.430 ;
        RECT 144.780 80.920 144.950 84.120 ;
        RECT 142.300 80.750 144.950 80.920 ;
        RECT 147.300 84.120 149.950 84.290 ;
        RECT 147.300 80.920 147.470 84.120 ;
        RECT 148.100 83.610 148.480 83.780 ;
        RECT 148.770 83.610 149.150 83.780 ;
        RECT 147.870 81.600 148.040 83.440 ;
        RECT 148.540 81.600 148.710 83.440 ;
        RECT 149.210 81.600 149.380 83.440 ;
        RECT 148.100 81.260 148.480 81.430 ;
        RECT 148.770 81.260 149.150 81.430 ;
        RECT 149.780 80.920 149.950 84.120 ;
        RECT 147.300 80.750 149.950 80.920 ;
        RECT 151.300 84.120 153.950 84.290 ;
        RECT 151.300 80.920 151.470 84.120 ;
        RECT 152.100 83.610 152.480 83.780 ;
        RECT 152.770 83.610 153.150 83.780 ;
        RECT 151.870 81.600 152.040 83.440 ;
        RECT 152.540 81.600 152.710 83.440 ;
        RECT 153.210 81.600 153.380 83.440 ;
        RECT 152.100 81.260 152.480 81.430 ;
        RECT 152.770 81.260 153.150 81.430 ;
        RECT 153.780 80.920 153.950 84.120 ;
        RECT 151.300 80.750 153.950 80.920 ;
        RECT 147.870 80.670 149.370 80.750 ;
        RECT 151.870 80.670 153.370 80.750 ;
        RECT 140.300 78.120 142.950 78.290 ;
        RECT 140.300 74.920 140.470 78.120 ;
        RECT 141.100 77.610 141.480 77.780 ;
        RECT 141.770 77.610 142.150 77.780 ;
        RECT 142.780 77.720 142.950 78.120 ;
        RECT 149.300 78.120 151.950 78.290 ;
        RECT 149.300 77.720 149.470 78.120 ;
        RECT 140.870 75.600 141.040 77.440 ;
        RECT 141.540 75.600 141.710 77.440 ;
        RECT 142.210 75.600 142.380 77.440 ;
        RECT 142.770 76.920 143.070 77.720 ;
        RECT 149.220 76.920 149.470 77.720 ;
        RECT 150.100 77.610 150.480 77.780 ;
        RECT 150.770 77.610 151.150 77.780 ;
        RECT 141.100 75.260 141.480 75.430 ;
        RECT 141.770 75.260 142.150 75.430 ;
        RECT 142.780 74.920 142.950 76.920 ;
        RECT 140.300 74.750 142.950 74.920 ;
        RECT 145.920 74.905 146.320 75.190 ;
        RECT 149.300 74.920 149.470 76.920 ;
        RECT 149.870 75.600 150.040 77.440 ;
        RECT 150.540 75.600 150.710 77.440 ;
        RECT 151.210 75.600 151.380 77.440 ;
        RECT 150.100 75.260 150.480 75.430 ;
        RECT 150.770 75.260 151.150 75.430 ;
        RECT 151.780 74.920 151.950 78.120 ;
        RECT 149.300 74.750 151.950 74.920 ;
        RECT 145.920 73.620 146.320 73.905 ;
      LAYER mcon ;
        RECT 57.335 203.415 57.505 203.585 ;
        RECT 57.795 203.415 57.965 203.585 ;
        RECT 58.255 203.415 58.425 203.585 ;
        RECT 58.715 203.415 58.885 203.585 ;
        RECT 59.175 203.415 59.345 203.585 ;
        RECT 59.635 203.415 59.805 203.585 ;
        RECT 60.095 203.415 60.265 203.585 ;
        RECT 60.555 203.415 60.725 203.585 ;
        RECT 61.015 203.415 61.185 203.585 ;
        RECT 61.475 203.415 61.645 203.585 ;
        RECT 61.935 203.415 62.105 203.585 ;
        RECT 62.395 203.415 62.565 203.585 ;
        RECT 62.855 203.415 63.025 203.585 ;
        RECT 63.315 203.415 63.485 203.585 ;
        RECT 63.775 203.415 63.945 203.585 ;
        RECT 64.235 203.415 64.405 203.585 ;
        RECT 64.695 203.415 64.865 203.585 ;
        RECT 65.155 203.415 65.325 203.585 ;
        RECT 65.615 203.415 65.785 203.585 ;
        RECT 66.075 203.415 66.245 203.585 ;
        RECT 66.535 203.415 66.705 203.585 ;
        RECT 66.995 203.415 67.165 203.585 ;
        RECT 67.455 203.415 67.625 203.585 ;
        RECT 67.915 203.415 68.085 203.585 ;
        RECT 68.375 203.415 68.545 203.585 ;
        RECT 68.835 203.415 69.005 203.585 ;
        RECT 69.295 203.415 69.465 203.585 ;
        RECT 69.755 203.415 69.925 203.585 ;
        RECT 70.215 203.415 70.385 203.585 ;
        RECT 70.675 203.415 70.845 203.585 ;
        RECT 71.135 203.415 71.305 203.585 ;
        RECT 71.595 203.415 71.765 203.585 ;
        RECT 72.055 203.415 72.225 203.585 ;
        RECT 72.515 203.415 72.685 203.585 ;
        RECT 72.975 203.415 73.145 203.585 ;
        RECT 73.435 203.415 73.605 203.585 ;
        RECT 73.895 203.415 74.065 203.585 ;
        RECT 74.355 203.415 74.525 203.585 ;
        RECT 74.815 203.415 74.985 203.585 ;
        RECT 75.275 203.415 75.445 203.585 ;
        RECT 75.735 203.415 75.905 203.585 ;
        RECT 76.195 203.415 76.365 203.585 ;
        RECT 76.655 203.415 76.825 203.585 ;
        RECT 77.115 203.415 77.285 203.585 ;
        RECT 77.575 203.415 77.745 203.585 ;
        RECT 78.035 203.415 78.205 203.585 ;
        RECT 78.495 203.415 78.665 203.585 ;
        RECT 78.955 203.415 79.125 203.585 ;
        RECT 79.415 203.415 79.585 203.585 ;
        RECT 79.875 203.415 80.045 203.585 ;
        RECT 80.335 203.415 80.505 203.585 ;
        RECT 80.795 203.415 80.965 203.585 ;
        RECT 81.255 203.415 81.425 203.585 ;
        RECT 81.715 203.415 81.885 203.585 ;
        RECT 82.175 203.415 82.345 203.585 ;
        RECT 82.635 203.415 82.805 203.585 ;
        RECT 83.095 203.415 83.265 203.585 ;
        RECT 83.555 203.415 83.725 203.585 ;
        RECT 84.015 203.415 84.185 203.585 ;
        RECT 84.475 203.415 84.645 203.585 ;
        RECT 84.935 203.415 85.105 203.585 ;
        RECT 85.395 203.415 85.565 203.585 ;
        RECT 85.855 203.415 86.025 203.585 ;
        RECT 86.315 203.415 86.485 203.585 ;
        RECT 86.775 203.415 86.945 203.585 ;
        RECT 87.235 203.415 87.405 203.585 ;
        RECT 87.695 203.415 87.865 203.585 ;
        RECT 88.155 203.415 88.325 203.585 ;
        RECT 88.615 203.415 88.785 203.585 ;
        RECT 89.075 203.415 89.245 203.585 ;
        RECT 89.535 203.415 89.705 203.585 ;
        RECT 89.995 203.415 90.165 203.585 ;
        RECT 90.455 203.415 90.625 203.585 ;
        RECT 90.915 203.415 91.085 203.585 ;
        RECT 91.375 203.415 91.545 203.585 ;
        RECT 91.835 203.415 92.005 203.585 ;
        RECT 92.295 203.415 92.465 203.585 ;
        RECT 92.755 203.415 92.925 203.585 ;
        RECT 93.215 203.415 93.385 203.585 ;
        RECT 93.675 203.415 93.845 203.585 ;
        RECT 94.135 203.415 94.305 203.585 ;
        RECT 94.595 203.415 94.765 203.585 ;
        RECT 95.055 203.415 95.225 203.585 ;
        RECT 95.515 203.415 95.685 203.585 ;
        RECT 95.975 203.415 96.145 203.585 ;
        RECT 96.435 203.415 96.605 203.585 ;
        RECT 96.895 203.415 97.065 203.585 ;
        RECT 97.355 203.415 97.525 203.585 ;
        RECT 97.815 203.415 97.985 203.585 ;
        RECT 98.275 203.415 98.445 203.585 ;
        RECT 98.735 203.415 98.905 203.585 ;
        RECT 99.195 203.415 99.365 203.585 ;
        RECT 99.655 203.415 99.825 203.585 ;
        RECT 100.115 203.415 100.285 203.585 ;
        RECT 100.575 203.415 100.745 203.585 ;
        RECT 101.035 203.415 101.205 203.585 ;
        RECT 101.495 203.415 101.665 203.585 ;
        RECT 101.955 203.415 102.125 203.585 ;
        RECT 102.415 203.415 102.585 203.585 ;
        RECT 102.875 203.415 103.045 203.585 ;
        RECT 103.335 203.415 103.505 203.585 ;
        RECT 103.795 203.415 103.965 203.585 ;
        RECT 104.255 203.415 104.425 203.585 ;
        RECT 104.715 203.415 104.885 203.585 ;
        RECT 105.175 203.415 105.345 203.585 ;
        RECT 105.635 203.415 105.805 203.585 ;
        RECT 106.095 203.415 106.265 203.585 ;
        RECT 106.555 203.415 106.725 203.585 ;
        RECT 107.015 203.415 107.185 203.585 ;
        RECT 107.475 203.415 107.645 203.585 ;
        RECT 107.935 203.415 108.105 203.585 ;
        RECT 108.395 203.415 108.565 203.585 ;
        RECT 108.855 203.415 109.025 203.585 ;
        RECT 109.315 203.415 109.485 203.585 ;
        RECT 109.775 203.415 109.945 203.585 ;
        RECT 110.235 203.415 110.405 203.585 ;
        RECT 110.695 203.415 110.865 203.585 ;
        RECT 111.155 203.415 111.325 203.585 ;
        RECT 111.615 203.415 111.785 203.585 ;
        RECT 112.075 203.415 112.245 203.585 ;
        RECT 112.535 203.415 112.705 203.585 ;
        RECT 112.995 203.415 113.165 203.585 ;
        RECT 113.455 203.415 113.625 203.585 ;
        RECT 113.915 203.415 114.085 203.585 ;
        RECT 114.375 203.415 114.545 203.585 ;
        RECT 114.835 203.415 115.005 203.585 ;
        RECT 115.295 203.415 115.465 203.585 ;
        RECT 115.755 203.415 115.925 203.585 ;
        RECT 116.215 203.415 116.385 203.585 ;
        RECT 116.675 203.415 116.845 203.585 ;
        RECT 117.135 203.415 117.305 203.585 ;
        RECT 117.595 203.415 117.765 203.585 ;
        RECT 118.055 203.415 118.225 203.585 ;
        RECT 118.515 203.415 118.685 203.585 ;
        RECT 118.975 203.415 119.145 203.585 ;
        RECT 119.435 203.415 119.605 203.585 ;
        RECT 119.895 203.415 120.065 203.585 ;
        RECT 120.355 203.415 120.525 203.585 ;
        RECT 120.815 203.415 120.985 203.585 ;
        RECT 121.275 203.415 121.445 203.585 ;
        RECT 121.735 203.415 121.905 203.585 ;
        RECT 122.195 203.415 122.365 203.585 ;
        RECT 122.655 203.415 122.825 203.585 ;
        RECT 123.115 203.415 123.285 203.585 ;
        RECT 123.575 203.415 123.745 203.585 ;
        RECT 124.035 203.415 124.205 203.585 ;
        RECT 124.495 203.415 124.665 203.585 ;
        RECT 124.955 203.415 125.125 203.585 ;
        RECT 125.415 203.415 125.585 203.585 ;
        RECT 125.875 203.415 126.045 203.585 ;
        RECT 126.335 203.415 126.505 203.585 ;
        RECT 126.795 203.415 126.965 203.585 ;
        RECT 127.255 203.415 127.425 203.585 ;
        RECT 127.715 203.415 127.885 203.585 ;
        RECT 128.175 203.415 128.345 203.585 ;
        RECT 128.635 203.415 128.805 203.585 ;
        RECT 129.095 203.415 129.265 203.585 ;
        RECT 129.555 203.415 129.725 203.585 ;
        RECT 130.015 203.415 130.185 203.585 ;
        RECT 130.475 203.415 130.645 203.585 ;
        RECT 130.935 203.415 131.105 203.585 ;
        RECT 61.015 201.885 61.185 202.055 ;
        RECT 61.935 201.205 62.105 201.375 ;
        RECT 71.135 201.885 71.305 202.055 ;
        RECT 72.055 202.225 72.225 202.395 ;
        RECT 75.275 202.225 75.445 202.395 ;
        RECT 76.195 202.565 76.365 202.735 ;
        RECT 76.655 201.885 76.825 202.055 ;
        RECT 80.335 201.885 80.505 202.055 ;
        RECT 76.655 201.205 76.825 201.375 ;
        RECT 81.255 201.205 81.425 201.375 ;
        RECT 86.315 201.885 86.485 202.055 ;
        RECT 86.775 201.885 86.945 202.055 ;
        RECT 85.855 201.205 86.025 201.375 ;
        RECT 91.375 202.565 91.545 202.735 ;
        RECT 89.535 201.885 89.705 202.055 ;
        RECT 90.455 201.885 90.625 202.055 ;
        RECT 101.495 202.905 101.665 203.075 ;
        RECT 97.355 201.885 97.525 202.055 ;
        RECT 98.735 201.885 98.905 202.055 ;
        RECT 98.275 201.205 98.445 201.375 ;
        RECT 100.575 201.885 100.745 202.055 ;
        RECT 102.875 201.885 103.045 202.055 ;
        RECT 99.655 201.205 99.825 201.375 ;
        RECT 106.095 201.205 106.265 201.375 ;
        RECT 109.315 202.225 109.485 202.395 ;
        RECT 110.695 201.885 110.865 202.055 ;
        RECT 118.975 201.885 119.145 202.055 ;
        RECT 113.915 201.205 114.085 201.375 ;
        RECT 119.895 201.205 120.065 201.375 ;
        RECT 57.335 200.695 57.505 200.865 ;
        RECT 57.795 200.695 57.965 200.865 ;
        RECT 58.255 200.695 58.425 200.865 ;
        RECT 58.715 200.695 58.885 200.865 ;
        RECT 59.175 200.695 59.345 200.865 ;
        RECT 59.635 200.695 59.805 200.865 ;
        RECT 60.095 200.695 60.265 200.865 ;
        RECT 60.555 200.695 60.725 200.865 ;
        RECT 61.015 200.695 61.185 200.865 ;
        RECT 61.475 200.695 61.645 200.865 ;
        RECT 61.935 200.695 62.105 200.865 ;
        RECT 62.395 200.695 62.565 200.865 ;
        RECT 62.855 200.695 63.025 200.865 ;
        RECT 63.315 200.695 63.485 200.865 ;
        RECT 63.775 200.695 63.945 200.865 ;
        RECT 64.235 200.695 64.405 200.865 ;
        RECT 64.695 200.695 64.865 200.865 ;
        RECT 65.155 200.695 65.325 200.865 ;
        RECT 65.615 200.695 65.785 200.865 ;
        RECT 66.075 200.695 66.245 200.865 ;
        RECT 66.535 200.695 66.705 200.865 ;
        RECT 66.995 200.695 67.165 200.865 ;
        RECT 67.455 200.695 67.625 200.865 ;
        RECT 67.915 200.695 68.085 200.865 ;
        RECT 68.375 200.695 68.545 200.865 ;
        RECT 68.835 200.695 69.005 200.865 ;
        RECT 69.295 200.695 69.465 200.865 ;
        RECT 69.755 200.695 69.925 200.865 ;
        RECT 70.215 200.695 70.385 200.865 ;
        RECT 70.675 200.695 70.845 200.865 ;
        RECT 71.135 200.695 71.305 200.865 ;
        RECT 71.595 200.695 71.765 200.865 ;
        RECT 72.055 200.695 72.225 200.865 ;
        RECT 72.515 200.695 72.685 200.865 ;
        RECT 72.975 200.695 73.145 200.865 ;
        RECT 73.435 200.695 73.605 200.865 ;
        RECT 73.895 200.695 74.065 200.865 ;
        RECT 74.355 200.695 74.525 200.865 ;
        RECT 74.815 200.695 74.985 200.865 ;
        RECT 75.275 200.695 75.445 200.865 ;
        RECT 75.735 200.695 75.905 200.865 ;
        RECT 76.195 200.695 76.365 200.865 ;
        RECT 76.655 200.695 76.825 200.865 ;
        RECT 77.115 200.695 77.285 200.865 ;
        RECT 77.575 200.695 77.745 200.865 ;
        RECT 78.035 200.695 78.205 200.865 ;
        RECT 78.495 200.695 78.665 200.865 ;
        RECT 78.955 200.695 79.125 200.865 ;
        RECT 79.415 200.695 79.585 200.865 ;
        RECT 79.875 200.695 80.045 200.865 ;
        RECT 80.335 200.695 80.505 200.865 ;
        RECT 80.795 200.695 80.965 200.865 ;
        RECT 81.255 200.695 81.425 200.865 ;
        RECT 81.715 200.695 81.885 200.865 ;
        RECT 82.175 200.695 82.345 200.865 ;
        RECT 82.635 200.695 82.805 200.865 ;
        RECT 83.095 200.695 83.265 200.865 ;
        RECT 83.555 200.695 83.725 200.865 ;
        RECT 84.015 200.695 84.185 200.865 ;
        RECT 84.475 200.695 84.645 200.865 ;
        RECT 84.935 200.695 85.105 200.865 ;
        RECT 85.395 200.695 85.565 200.865 ;
        RECT 85.855 200.695 86.025 200.865 ;
        RECT 86.315 200.695 86.485 200.865 ;
        RECT 86.775 200.695 86.945 200.865 ;
        RECT 87.235 200.695 87.405 200.865 ;
        RECT 87.695 200.695 87.865 200.865 ;
        RECT 88.155 200.695 88.325 200.865 ;
        RECT 88.615 200.695 88.785 200.865 ;
        RECT 89.075 200.695 89.245 200.865 ;
        RECT 89.535 200.695 89.705 200.865 ;
        RECT 89.995 200.695 90.165 200.865 ;
        RECT 90.455 200.695 90.625 200.865 ;
        RECT 90.915 200.695 91.085 200.865 ;
        RECT 91.375 200.695 91.545 200.865 ;
        RECT 91.835 200.695 92.005 200.865 ;
        RECT 92.295 200.695 92.465 200.865 ;
        RECT 92.755 200.695 92.925 200.865 ;
        RECT 93.215 200.695 93.385 200.865 ;
        RECT 93.675 200.695 93.845 200.865 ;
        RECT 94.135 200.695 94.305 200.865 ;
        RECT 94.595 200.695 94.765 200.865 ;
        RECT 95.055 200.695 95.225 200.865 ;
        RECT 95.515 200.695 95.685 200.865 ;
        RECT 95.975 200.695 96.145 200.865 ;
        RECT 96.435 200.695 96.605 200.865 ;
        RECT 96.895 200.695 97.065 200.865 ;
        RECT 97.355 200.695 97.525 200.865 ;
        RECT 97.815 200.695 97.985 200.865 ;
        RECT 98.275 200.695 98.445 200.865 ;
        RECT 98.735 200.695 98.905 200.865 ;
        RECT 99.195 200.695 99.365 200.865 ;
        RECT 99.655 200.695 99.825 200.865 ;
        RECT 100.115 200.695 100.285 200.865 ;
        RECT 100.575 200.695 100.745 200.865 ;
        RECT 101.035 200.695 101.205 200.865 ;
        RECT 101.495 200.695 101.665 200.865 ;
        RECT 101.955 200.695 102.125 200.865 ;
        RECT 102.415 200.695 102.585 200.865 ;
        RECT 102.875 200.695 103.045 200.865 ;
        RECT 103.335 200.695 103.505 200.865 ;
        RECT 103.795 200.695 103.965 200.865 ;
        RECT 104.255 200.695 104.425 200.865 ;
        RECT 104.715 200.695 104.885 200.865 ;
        RECT 105.175 200.695 105.345 200.865 ;
        RECT 105.635 200.695 105.805 200.865 ;
        RECT 106.095 200.695 106.265 200.865 ;
        RECT 106.555 200.695 106.725 200.865 ;
        RECT 107.015 200.695 107.185 200.865 ;
        RECT 107.475 200.695 107.645 200.865 ;
        RECT 107.935 200.695 108.105 200.865 ;
        RECT 108.395 200.695 108.565 200.865 ;
        RECT 108.855 200.695 109.025 200.865 ;
        RECT 109.315 200.695 109.485 200.865 ;
        RECT 109.775 200.695 109.945 200.865 ;
        RECT 110.235 200.695 110.405 200.865 ;
        RECT 110.695 200.695 110.865 200.865 ;
        RECT 111.155 200.695 111.325 200.865 ;
        RECT 111.615 200.695 111.785 200.865 ;
        RECT 112.075 200.695 112.245 200.865 ;
        RECT 112.535 200.695 112.705 200.865 ;
        RECT 112.995 200.695 113.165 200.865 ;
        RECT 113.455 200.695 113.625 200.865 ;
        RECT 113.915 200.695 114.085 200.865 ;
        RECT 114.375 200.695 114.545 200.865 ;
        RECT 114.835 200.695 115.005 200.865 ;
        RECT 115.295 200.695 115.465 200.865 ;
        RECT 115.755 200.695 115.925 200.865 ;
        RECT 116.215 200.695 116.385 200.865 ;
        RECT 116.675 200.695 116.845 200.865 ;
        RECT 117.135 200.695 117.305 200.865 ;
        RECT 117.595 200.695 117.765 200.865 ;
        RECT 118.055 200.695 118.225 200.865 ;
        RECT 118.515 200.695 118.685 200.865 ;
        RECT 118.975 200.695 119.145 200.865 ;
        RECT 119.435 200.695 119.605 200.865 ;
        RECT 119.895 200.695 120.065 200.865 ;
        RECT 120.355 200.695 120.525 200.865 ;
        RECT 120.815 200.695 120.985 200.865 ;
        RECT 121.275 200.695 121.445 200.865 ;
        RECT 121.735 200.695 121.905 200.865 ;
        RECT 122.195 200.695 122.365 200.865 ;
        RECT 122.655 200.695 122.825 200.865 ;
        RECT 123.115 200.695 123.285 200.865 ;
        RECT 123.575 200.695 123.745 200.865 ;
        RECT 124.035 200.695 124.205 200.865 ;
        RECT 124.495 200.695 124.665 200.865 ;
        RECT 124.955 200.695 125.125 200.865 ;
        RECT 125.415 200.695 125.585 200.865 ;
        RECT 125.875 200.695 126.045 200.865 ;
        RECT 126.335 200.695 126.505 200.865 ;
        RECT 126.795 200.695 126.965 200.865 ;
        RECT 127.255 200.695 127.425 200.865 ;
        RECT 127.715 200.695 127.885 200.865 ;
        RECT 128.175 200.695 128.345 200.865 ;
        RECT 128.635 200.695 128.805 200.865 ;
        RECT 129.095 200.695 129.265 200.865 ;
        RECT 129.555 200.695 129.725 200.865 ;
        RECT 130.015 200.695 130.185 200.865 ;
        RECT 130.475 200.695 130.645 200.865 ;
        RECT 130.935 200.695 131.105 200.865 ;
        RECT 72.975 199.505 73.145 199.675 ;
        RECT 72.515 199.165 72.685 199.335 ;
        RECT 78.495 200.185 78.665 200.355 ;
        RECT 75.275 199.505 75.445 199.675 ;
        RECT 74.815 199.165 74.985 199.335 ;
        RECT 76.195 199.505 76.365 199.675 ;
        RECT 76.655 199.505 76.825 199.675 ;
        RECT 77.575 199.505 77.745 199.675 ;
        RECT 80.795 199.845 80.965 200.015 ;
        RECT 79.875 199.505 80.045 199.675 ;
        RECT 81.255 199.505 81.425 199.675 ;
        RECT 81.715 199.505 81.885 199.675 ;
        RECT 77.115 198.825 77.285 198.995 ;
        RECT 82.635 198.825 82.805 198.995 ;
        RECT 83.555 199.165 83.725 199.335 ;
        RECT 84.935 199.505 85.105 199.675 ;
        RECT 84.475 198.485 84.645 198.655 ;
        RECT 85.855 198.825 86.025 198.995 ;
        RECT 88.165 199.165 88.335 199.335 ;
        RECT 88.600 198.825 88.770 198.995 ;
        RECT 90.685 199.165 90.855 199.335 ;
        RECT 90.170 198.825 90.340 198.995 ;
        RECT 91.475 199.505 91.645 199.675 ;
        RECT 91.875 199.165 92.045 199.335 ;
        RECT 92.755 199.505 92.925 199.675 ;
        RECT 93.215 199.505 93.385 199.675 ;
        RECT 92.270 198.825 92.440 198.995 ;
        RECT 93.700 198.825 93.870 198.995 ;
        RECT 94.095 199.165 94.265 199.335 ;
        RECT 94.550 199.505 94.720 199.675 ;
        RECT 95.285 199.165 95.455 199.335 ;
        RECT 95.800 198.825 95.970 198.995 ;
        RECT 97.370 198.825 97.540 198.995 ;
        RECT 97.805 199.165 97.975 199.335 ;
        RECT 101.955 200.185 102.125 200.355 ;
        RECT 100.115 198.825 100.285 198.995 ;
        RECT 101.495 199.165 101.665 199.335 ;
        RECT 102.415 200.185 102.585 200.355 ;
        RECT 105.635 199.505 105.805 199.675 ;
        RECT 104.255 198.825 104.425 198.995 ;
        RECT 105.175 198.485 105.345 198.655 ;
        RECT 111.615 199.505 111.785 199.675 ;
        RECT 112.080 199.505 112.250 199.675 ;
        RECT 112.995 199.165 113.165 199.335 ;
        RECT 112.485 198.825 112.655 198.995 ;
        RECT 113.915 199.505 114.085 199.675 ;
        RECT 115.275 199.845 115.445 200.015 ;
        RECT 115.635 199.845 115.805 200.015 ;
        RECT 114.375 198.825 114.545 198.995 ;
        RECT 117.495 199.505 117.665 199.675 ;
        RECT 118.875 199.845 119.045 200.015 ;
        RECT 118.575 199.530 118.745 199.700 ;
        RECT 117.495 198.825 117.665 198.995 ;
        RECT 120.355 199.165 120.525 199.335 ;
        RECT 120.815 198.485 120.985 198.655 ;
        RECT 124.955 199.845 125.125 200.015 ;
        RECT 124.495 199.505 124.665 199.675 ;
        RECT 57.335 197.975 57.505 198.145 ;
        RECT 57.795 197.975 57.965 198.145 ;
        RECT 58.255 197.975 58.425 198.145 ;
        RECT 58.715 197.975 58.885 198.145 ;
        RECT 59.175 197.975 59.345 198.145 ;
        RECT 59.635 197.975 59.805 198.145 ;
        RECT 60.095 197.975 60.265 198.145 ;
        RECT 60.555 197.975 60.725 198.145 ;
        RECT 61.015 197.975 61.185 198.145 ;
        RECT 61.475 197.975 61.645 198.145 ;
        RECT 61.935 197.975 62.105 198.145 ;
        RECT 62.395 197.975 62.565 198.145 ;
        RECT 62.855 197.975 63.025 198.145 ;
        RECT 63.315 197.975 63.485 198.145 ;
        RECT 63.775 197.975 63.945 198.145 ;
        RECT 64.235 197.975 64.405 198.145 ;
        RECT 64.695 197.975 64.865 198.145 ;
        RECT 65.155 197.975 65.325 198.145 ;
        RECT 65.615 197.975 65.785 198.145 ;
        RECT 66.075 197.975 66.245 198.145 ;
        RECT 66.535 197.975 66.705 198.145 ;
        RECT 66.995 197.975 67.165 198.145 ;
        RECT 67.455 197.975 67.625 198.145 ;
        RECT 67.915 197.975 68.085 198.145 ;
        RECT 68.375 197.975 68.545 198.145 ;
        RECT 68.835 197.975 69.005 198.145 ;
        RECT 69.295 197.975 69.465 198.145 ;
        RECT 69.755 197.975 69.925 198.145 ;
        RECT 70.215 197.975 70.385 198.145 ;
        RECT 70.675 197.975 70.845 198.145 ;
        RECT 71.135 197.975 71.305 198.145 ;
        RECT 71.595 197.975 71.765 198.145 ;
        RECT 72.055 197.975 72.225 198.145 ;
        RECT 72.515 197.975 72.685 198.145 ;
        RECT 72.975 197.975 73.145 198.145 ;
        RECT 73.435 197.975 73.605 198.145 ;
        RECT 73.895 197.975 74.065 198.145 ;
        RECT 74.355 197.975 74.525 198.145 ;
        RECT 74.815 197.975 74.985 198.145 ;
        RECT 75.275 197.975 75.445 198.145 ;
        RECT 75.735 197.975 75.905 198.145 ;
        RECT 76.195 197.975 76.365 198.145 ;
        RECT 76.655 197.975 76.825 198.145 ;
        RECT 77.115 197.975 77.285 198.145 ;
        RECT 77.575 197.975 77.745 198.145 ;
        RECT 78.035 197.975 78.205 198.145 ;
        RECT 78.495 197.975 78.665 198.145 ;
        RECT 78.955 197.975 79.125 198.145 ;
        RECT 79.415 197.975 79.585 198.145 ;
        RECT 79.875 197.975 80.045 198.145 ;
        RECT 80.335 197.975 80.505 198.145 ;
        RECT 80.795 197.975 80.965 198.145 ;
        RECT 81.255 197.975 81.425 198.145 ;
        RECT 81.715 197.975 81.885 198.145 ;
        RECT 82.175 197.975 82.345 198.145 ;
        RECT 82.635 197.975 82.805 198.145 ;
        RECT 83.095 197.975 83.265 198.145 ;
        RECT 83.555 197.975 83.725 198.145 ;
        RECT 84.015 197.975 84.185 198.145 ;
        RECT 84.475 197.975 84.645 198.145 ;
        RECT 84.935 197.975 85.105 198.145 ;
        RECT 85.395 197.975 85.565 198.145 ;
        RECT 85.855 197.975 86.025 198.145 ;
        RECT 86.315 197.975 86.485 198.145 ;
        RECT 86.775 197.975 86.945 198.145 ;
        RECT 87.235 197.975 87.405 198.145 ;
        RECT 87.695 197.975 87.865 198.145 ;
        RECT 88.155 197.975 88.325 198.145 ;
        RECT 88.615 197.975 88.785 198.145 ;
        RECT 89.075 197.975 89.245 198.145 ;
        RECT 89.535 197.975 89.705 198.145 ;
        RECT 89.995 197.975 90.165 198.145 ;
        RECT 90.455 197.975 90.625 198.145 ;
        RECT 90.915 197.975 91.085 198.145 ;
        RECT 91.375 197.975 91.545 198.145 ;
        RECT 91.835 197.975 92.005 198.145 ;
        RECT 92.295 197.975 92.465 198.145 ;
        RECT 92.755 197.975 92.925 198.145 ;
        RECT 93.215 197.975 93.385 198.145 ;
        RECT 93.675 197.975 93.845 198.145 ;
        RECT 94.135 197.975 94.305 198.145 ;
        RECT 94.595 197.975 94.765 198.145 ;
        RECT 95.055 197.975 95.225 198.145 ;
        RECT 95.515 197.975 95.685 198.145 ;
        RECT 95.975 197.975 96.145 198.145 ;
        RECT 96.435 197.975 96.605 198.145 ;
        RECT 96.895 197.975 97.065 198.145 ;
        RECT 97.355 197.975 97.525 198.145 ;
        RECT 97.815 197.975 97.985 198.145 ;
        RECT 98.275 197.975 98.445 198.145 ;
        RECT 98.735 197.975 98.905 198.145 ;
        RECT 99.195 197.975 99.365 198.145 ;
        RECT 99.655 197.975 99.825 198.145 ;
        RECT 100.115 197.975 100.285 198.145 ;
        RECT 100.575 197.975 100.745 198.145 ;
        RECT 101.035 197.975 101.205 198.145 ;
        RECT 101.495 197.975 101.665 198.145 ;
        RECT 101.955 197.975 102.125 198.145 ;
        RECT 102.415 197.975 102.585 198.145 ;
        RECT 102.875 197.975 103.045 198.145 ;
        RECT 103.335 197.975 103.505 198.145 ;
        RECT 103.795 197.975 103.965 198.145 ;
        RECT 104.255 197.975 104.425 198.145 ;
        RECT 104.715 197.975 104.885 198.145 ;
        RECT 105.175 197.975 105.345 198.145 ;
        RECT 105.635 197.975 105.805 198.145 ;
        RECT 106.095 197.975 106.265 198.145 ;
        RECT 106.555 197.975 106.725 198.145 ;
        RECT 107.015 197.975 107.185 198.145 ;
        RECT 107.475 197.975 107.645 198.145 ;
        RECT 107.935 197.975 108.105 198.145 ;
        RECT 108.395 197.975 108.565 198.145 ;
        RECT 108.855 197.975 109.025 198.145 ;
        RECT 109.315 197.975 109.485 198.145 ;
        RECT 109.775 197.975 109.945 198.145 ;
        RECT 110.235 197.975 110.405 198.145 ;
        RECT 110.695 197.975 110.865 198.145 ;
        RECT 111.155 197.975 111.325 198.145 ;
        RECT 111.615 197.975 111.785 198.145 ;
        RECT 112.075 197.975 112.245 198.145 ;
        RECT 112.535 197.975 112.705 198.145 ;
        RECT 112.995 197.975 113.165 198.145 ;
        RECT 113.455 197.975 113.625 198.145 ;
        RECT 113.915 197.975 114.085 198.145 ;
        RECT 114.375 197.975 114.545 198.145 ;
        RECT 114.835 197.975 115.005 198.145 ;
        RECT 115.295 197.975 115.465 198.145 ;
        RECT 115.755 197.975 115.925 198.145 ;
        RECT 116.215 197.975 116.385 198.145 ;
        RECT 116.675 197.975 116.845 198.145 ;
        RECT 117.135 197.975 117.305 198.145 ;
        RECT 117.595 197.975 117.765 198.145 ;
        RECT 118.055 197.975 118.225 198.145 ;
        RECT 118.515 197.975 118.685 198.145 ;
        RECT 118.975 197.975 119.145 198.145 ;
        RECT 119.435 197.975 119.605 198.145 ;
        RECT 119.895 197.975 120.065 198.145 ;
        RECT 120.355 197.975 120.525 198.145 ;
        RECT 120.815 197.975 120.985 198.145 ;
        RECT 121.275 197.975 121.445 198.145 ;
        RECT 121.735 197.975 121.905 198.145 ;
        RECT 122.195 197.975 122.365 198.145 ;
        RECT 122.655 197.975 122.825 198.145 ;
        RECT 123.115 197.975 123.285 198.145 ;
        RECT 123.575 197.975 123.745 198.145 ;
        RECT 124.035 197.975 124.205 198.145 ;
        RECT 124.495 197.975 124.665 198.145 ;
        RECT 124.955 197.975 125.125 198.145 ;
        RECT 125.415 197.975 125.585 198.145 ;
        RECT 125.875 197.975 126.045 198.145 ;
        RECT 126.335 197.975 126.505 198.145 ;
        RECT 126.795 197.975 126.965 198.145 ;
        RECT 127.255 197.975 127.425 198.145 ;
        RECT 127.715 197.975 127.885 198.145 ;
        RECT 128.175 197.975 128.345 198.145 ;
        RECT 128.635 197.975 128.805 198.145 ;
        RECT 129.095 197.975 129.265 198.145 ;
        RECT 129.555 197.975 129.725 198.145 ;
        RECT 130.015 197.975 130.185 198.145 ;
        RECT 130.475 197.975 130.645 198.145 ;
        RECT 130.935 197.975 131.105 198.145 ;
        RECT 76.195 197.125 76.365 197.295 ;
        RECT 78.035 197.465 78.205 197.635 ;
        RECT 75.735 196.445 75.905 196.615 ;
        RECT 77.115 196.445 77.285 196.615 ;
        RECT 82.635 197.465 82.805 197.635 ;
        RECT 83.540 196.445 83.710 196.615 ;
        RECT 85.395 196.785 85.565 196.955 ;
        RECT 85.855 196.785 86.025 196.955 ;
        RECT 88.615 197.125 88.785 197.295 ;
        RECT 87.235 196.445 87.405 196.615 ;
        RECT 87.695 196.445 87.865 196.615 ;
        RECT 89.535 196.785 89.705 196.955 ;
        RECT 88.615 196.105 88.785 196.275 ;
        RECT 92.755 197.465 92.925 197.635 ;
        RECT 93.675 196.785 93.845 196.955 ;
        RECT 93.215 196.445 93.385 196.615 ;
        RECT 94.135 196.445 94.305 196.615 ;
        RECT 96.435 197.465 96.605 197.635 ;
        RECT 97.355 196.445 97.525 196.615 ;
        RECT 100.115 196.785 100.285 196.955 ;
        RECT 98.735 196.445 98.905 196.615 ;
        RECT 99.655 196.445 99.825 196.615 ;
        RECT 101.035 196.445 101.205 196.615 ;
        RECT 101.495 196.445 101.665 196.615 ;
        RECT 102.415 196.445 102.585 196.615 ;
        RECT 102.875 196.445 103.045 196.615 ;
        RECT 113.915 197.465 114.085 197.635 ;
        RECT 106.095 195.765 106.265 195.935 ;
        RECT 113.455 196.445 113.625 196.615 ;
        RECT 116.215 196.785 116.385 196.955 ;
        RECT 118.055 197.465 118.225 197.635 ;
        RECT 116.675 196.785 116.845 196.955 ;
        RECT 118.055 196.445 118.225 196.615 ;
        RECT 118.975 196.445 119.145 196.615 ;
        RECT 119.435 196.445 119.605 196.615 ;
        RECT 120.355 195.765 120.525 195.935 ;
        RECT 123.115 196.445 123.285 196.615 ;
        RECT 122.195 195.765 122.365 195.935 ;
        RECT 57.335 195.255 57.505 195.425 ;
        RECT 57.795 195.255 57.965 195.425 ;
        RECT 58.255 195.255 58.425 195.425 ;
        RECT 58.715 195.255 58.885 195.425 ;
        RECT 59.175 195.255 59.345 195.425 ;
        RECT 59.635 195.255 59.805 195.425 ;
        RECT 60.095 195.255 60.265 195.425 ;
        RECT 60.555 195.255 60.725 195.425 ;
        RECT 61.015 195.255 61.185 195.425 ;
        RECT 61.475 195.255 61.645 195.425 ;
        RECT 61.935 195.255 62.105 195.425 ;
        RECT 62.395 195.255 62.565 195.425 ;
        RECT 62.855 195.255 63.025 195.425 ;
        RECT 63.315 195.255 63.485 195.425 ;
        RECT 63.775 195.255 63.945 195.425 ;
        RECT 64.235 195.255 64.405 195.425 ;
        RECT 64.695 195.255 64.865 195.425 ;
        RECT 65.155 195.255 65.325 195.425 ;
        RECT 65.615 195.255 65.785 195.425 ;
        RECT 66.075 195.255 66.245 195.425 ;
        RECT 66.535 195.255 66.705 195.425 ;
        RECT 66.995 195.255 67.165 195.425 ;
        RECT 67.455 195.255 67.625 195.425 ;
        RECT 67.915 195.255 68.085 195.425 ;
        RECT 68.375 195.255 68.545 195.425 ;
        RECT 68.835 195.255 69.005 195.425 ;
        RECT 69.295 195.255 69.465 195.425 ;
        RECT 69.755 195.255 69.925 195.425 ;
        RECT 70.215 195.255 70.385 195.425 ;
        RECT 70.675 195.255 70.845 195.425 ;
        RECT 71.135 195.255 71.305 195.425 ;
        RECT 71.595 195.255 71.765 195.425 ;
        RECT 72.055 195.255 72.225 195.425 ;
        RECT 72.515 195.255 72.685 195.425 ;
        RECT 72.975 195.255 73.145 195.425 ;
        RECT 73.435 195.255 73.605 195.425 ;
        RECT 73.895 195.255 74.065 195.425 ;
        RECT 74.355 195.255 74.525 195.425 ;
        RECT 74.815 195.255 74.985 195.425 ;
        RECT 75.275 195.255 75.445 195.425 ;
        RECT 75.735 195.255 75.905 195.425 ;
        RECT 76.195 195.255 76.365 195.425 ;
        RECT 76.655 195.255 76.825 195.425 ;
        RECT 77.115 195.255 77.285 195.425 ;
        RECT 77.575 195.255 77.745 195.425 ;
        RECT 78.035 195.255 78.205 195.425 ;
        RECT 78.495 195.255 78.665 195.425 ;
        RECT 78.955 195.255 79.125 195.425 ;
        RECT 79.415 195.255 79.585 195.425 ;
        RECT 79.875 195.255 80.045 195.425 ;
        RECT 80.335 195.255 80.505 195.425 ;
        RECT 80.795 195.255 80.965 195.425 ;
        RECT 81.255 195.255 81.425 195.425 ;
        RECT 81.715 195.255 81.885 195.425 ;
        RECT 82.175 195.255 82.345 195.425 ;
        RECT 82.635 195.255 82.805 195.425 ;
        RECT 83.095 195.255 83.265 195.425 ;
        RECT 83.555 195.255 83.725 195.425 ;
        RECT 84.015 195.255 84.185 195.425 ;
        RECT 84.475 195.255 84.645 195.425 ;
        RECT 84.935 195.255 85.105 195.425 ;
        RECT 85.395 195.255 85.565 195.425 ;
        RECT 85.855 195.255 86.025 195.425 ;
        RECT 86.315 195.255 86.485 195.425 ;
        RECT 86.775 195.255 86.945 195.425 ;
        RECT 87.235 195.255 87.405 195.425 ;
        RECT 87.695 195.255 87.865 195.425 ;
        RECT 88.155 195.255 88.325 195.425 ;
        RECT 88.615 195.255 88.785 195.425 ;
        RECT 89.075 195.255 89.245 195.425 ;
        RECT 89.535 195.255 89.705 195.425 ;
        RECT 89.995 195.255 90.165 195.425 ;
        RECT 90.455 195.255 90.625 195.425 ;
        RECT 90.915 195.255 91.085 195.425 ;
        RECT 91.375 195.255 91.545 195.425 ;
        RECT 91.835 195.255 92.005 195.425 ;
        RECT 92.295 195.255 92.465 195.425 ;
        RECT 92.755 195.255 92.925 195.425 ;
        RECT 93.215 195.255 93.385 195.425 ;
        RECT 93.675 195.255 93.845 195.425 ;
        RECT 94.135 195.255 94.305 195.425 ;
        RECT 94.595 195.255 94.765 195.425 ;
        RECT 95.055 195.255 95.225 195.425 ;
        RECT 95.515 195.255 95.685 195.425 ;
        RECT 95.975 195.255 96.145 195.425 ;
        RECT 96.435 195.255 96.605 195.425 ;
        RECT 96.895 195.255 97.065 195.425 ;
        RECT 97.355 195.255 97.525 195.425 ;
        RECT 97.815 195.255 97.985 195.425 ;
        RECT 98.275 195.255 98.445 195.425 ;
        RECT 98.735 195.255 98.905 195.425 ;
        RECT 99.195 195.255 99.365 195.425 ;
        RECT 99.655 195.255 99.825 195.425 ;
        RECT 100.115 195.255 100.285 195.425 ;
        RECT 100.575 195.255 100.745 195.425 ;
        RECT 101.035 195.255 101.205 195.425 ;
        RECT 101.495 195.255 101.665 195.425 ;
        RECT 101.955 195.255 102.125 195.425 ;
        RECT 102.415 195.255 102.585 195.425 ;
        RECT 102.875 195.255 103.045 195.425 ;
        RECT 103.335 195.255 103.505 195.425 ;
        RECT 103.795 195.255 103.965 195.425 ;
        RECT 104.255 195.255 104.425 195.425 ;
        RECT 104.715 195.255 104.885 195.425 ;
        RECT 105.175 195.255 105.345 195.425 ;
        RECT 105.635 195.255 105.805 195.425 ;
        RECT 106.095 195.255 106.265 195.425 ;
        RECT 106.555 195.255 106.725 195.425 ;
        RECT 107.015 195.255 107.185 195.425 ;
        RECT 107.475 195.255 107.645 195.425 ;
        RECT 107.935 195.255 108.105 195.425 ;
        RECT 108.395 195.255 108.565 195.425 ;
        RECT 108.855 195.255 109.025 195.425 ;
        RECT 109.315 195.255 109.485 195.425 ;
        RECT 109.775 195.255 109.945 195.425 ;
        RECT 110.235 195.255 110.405 195.425 ;
        RECT 110.695 195.255 110.865 195.425 ;
        RECT 111.155 195.255 111.325 195.425 ;
        RECT 111.615 195.255 111.785 195.425 ;
        RECT 112.075 195.255 112.245 195.425 ;
        RECT 112.535 195.255 112.705 195.425 ;
        RECT 112.995 195.255 113.165 195.425 ;
        RECT 113.455 195.255 113.625 195.425 ;
        RECT 113.915 195.255 114.085 195.425 ;
        RECT 114.375 195.255 114.545 195.425 ;
        RECT 114.835 195.255 115.005 195.425 ;
        RECT 115.295 195.255 115.465 195.425 ;
        RECT 115.755 195.255 115.925 195.425 ;
        RECT 116.215 195.255 116.385 195.425 ;
        RECT 116.675 195.255 116.845 195.425 ;
        RECT 117.135 195.255 117.305 195.425 ;
        RECT 117.595 195.255 117.765 195.425 ;
        RECT 118.055 195.255 118.225 195.425 ;
        RECT 118.515 195.255 118.685 195.425 ;
        RECT 118.975 195.255 119.145 195.425 ;
        RECT 119.435 195.255 119.605 195.425 ;
        RECT 119.895 195.255 120.065 195.425 ;
        RECT 120.355 195.255 120.525 195.425 ;
        RECT 120.815 195.255 120.985 195.425 ;
        RECT 121.275 195.255 121.445 195.425 ;
        RECT 121.735 195.255 121.905 195.425 ;
        RECT 122.195 195.255 122.365 195.425 ;
        RECT 122.655 195.255 122.825 195.425 ;
        RECT 123.115 195.255 123.285 195.425 ;
        RECT 123.575 195.255 123.745 195.425 ;
        RECT 124.035 195.255 124.205 195.425 ;
        RECT 124.495 195.255 124.665 195.425 ;
        RECT 124.955 195.255 125.125 195.425 ;
        RECT 125.415 195.255 125.585 195.425 ;
        RECT 125.875 195.255 126.045 195.425 ;
        RECT 126.335 195.255 126.505 195.425 ;
        RECT 126.795 195.255 126.965 195.425 ;
        RECT 127.255 195.255 127.425 195.425 ;
        RECT 127.715 195.255 127.885 195.425 ;
        RECT 128.175 195.255 128.345 195.425 ;
        RECT 128.635 195.255 128.805 195.425 ;
        RECT 129.095 195.255 129.265 195.425 ;
        RECT 129.555 195.255 129.725 195.425 ;
        RECT 130.015 195.255 130.185 195.425 ;
        RECT 130.475 195.255 130.645 195.425 ;
        RECT 130.935 195.255 131.105 195.425 ;
        RECT 78.035 194.745 78.205 194.915 ;
        RECT 80.335 193.725 80.505 193.895 ;
        RECT 80.795 193.725 80.965 193.895 ;
        RECT 92.295 194.405 92.465 194.575 ;
        RECT 92.755 194.065 92.925 194.235 ;
        RECT 85.855 193.045 86.025 193.215 ;
        RECT 106.095 194.745 106.265 194.915 ;
        RECT 93.675 193.045 93.845 193.215 ;
        RECT 105.175 194.065 105.345 194.235 ;
        RECT 104.255 193.725 104.425 193.895 ;
        RECT 106.555 194.065 106.725 194.235 ;
        RECT 109.315 194.405 109.485 194.575 ;
        RECT 107.475 194.065 107.645 194.235 ;
        RECT 107.015 193.725 107.185 193.895 ;
        RECT 115.755 193.045 115.925 193.215 ;
        RECT 57.335 192.535 57.505 192.705 ;
        RECT 57.795 192.535 57.965 192.705 ;
        RECT 58.255 192.535 58.425 192.705 ;
        RECT 58.715 192.535 58.885 192.705 ;
        RECT 59.175 192.535 59.345 192.705 ;
        RECT 59.635 192.535 59.805 192.705 ;
        RECT 60.095 192.535 60.265 192.705 ;
        RECT 60.555 192.535 60.725 192.705 ;
        RECT 61.015 192.535 61.185 192.705 ;
        RECT 61.475 192.535 61.645 192.705 ;
        RECT 61.935 192.535 62.105 192.705 ;
        RECT 62.395 192.535 62.565 192.705 ;
        RECT 62.855 192.535 63.025 192.705 ;
        RECT 63.315 192.535 63.485 192.705 ;
        RECT 63.775 192.535 63.945 192.705 ;
        RECT 64.235 192.535 64.405 192.705 ;
        RECT 64.695 192.535 64.865 192.705 ;
        RECT 65.155 192.535 65.325 192.705 ;
        RECT 65.615 192.535 65.785 192.705 ;
        RECT 66.075 192.535 66.245 192.705 ;
        RECT 66.535 192.535 66.705 192.705 ;
        RECT 66.995 192.535 67.165 192.705 ;
        RECT 67.455 192.535 67.625 192.705 ;
        RECT 67.915 192.535 68.085 192.705 ;
        RECT 68.375 192.535 68.545 192.705 ;
        RECT 68.835 192.535 69.005 192.705 ;
        RECT 69.295 192.535 69.465 192.705 ;
        RECT 69.755 192.535 69.925 192.705 ;
        RECT 70.215 192.535 70.385 192.705 ;
        RECT 70.675 192.535 70.845 192.705 ;
        RECT 71.135 192.535 71.305 192.705 ;
        RECT 71.595 192.535 71.765 192.705 ;
        RECT 72.055 192.535 72.225 192.705 ;
        RECT 72.515 192.535 72.685 192.705 ;
        RECT 72.975 192.535 73.145 192.705 ;
        RECT 73.435 192.535 73.605 192.705 ;
        RECT 73.895 192.535 74.065 192.705 ;
        RECT 74.355 192.535 74.525 192.705 ;
        RECT 74.815 192.535 74.985 192.705 ;
        RECT 75.275 192.535 75.445 192.705 ;
        RECT 75.735 192.535 75.905 192.705 ;
        RECT 76.195 192.535 76.365 192.705 ;
        RECT 76.655 192.535 76.825 192.705 ;
        RECT 77.115 192.535 77.285 192.705 ;
        RECT 77.575 192.535 77.745 192.705 ;
        RECT 78.035 192.535 78.205 192.705 ;
        RECT 78.495 192.535 78.665 192.705 ;
        RECT 78.955 192.535 79.125 192.705 ;
        RECT 79.415 192.535 79.585 192.705 ;
        RECT 79.875 192.535 80.045 192.705 ;
        RECT 80.335 192.535 80.505 192.705 ;
        RECT 80.795 192.535 80.965 192.705 ;
        RECT 81.255 192.535 81.425 192.705 ;
        RECT 81.715 192.535 81.885 192.705 ;
        RECT 82.175 192.535 82.345 192.705 ;
        RECT 82.635 192.535 82.805 192.705 ;
        RECT 83.095 192.535 83.265 192.705 ;
        RECT 83.555 192.535 83.725 192.705 ;
        RECT 84.015 192.535 84.185 192.705 ;
        RECT 84.475 192.535 84.645 192.705 ;
        RECT 84.935 192.535 85.105 192.705 ;
        RECT 85.395 192.535 85.565 192.705 ;
        RECT 85.855 192.535 86.025 192.705 ;
        RECT 86.315 192.535 86.485 192.705 ;
        RECT 86.775 192.535 86.945 192.705 ;
        RECT 87.235 192.535 87.405 192.705 ;
        RECT 87.695 192.535 87.865 192.705 ;
        RECT 88.155 192.535 88.325 192.705 ;
        RECT 88.615 192.535 88.785 192.705 ;
        RECT 89.075 192.535 89.245 192.705 ;
        RECT 89.535 192.535 89.705 192.705 ;
        RECT 89.995 192.535 90.165 192.705 ;
        RECT 90.455 192.535 90.625 192.705 ;
        RECT 90.915 192.535 91.085 192.705 ;
        RECT 91.375 192.535 91.545 192.705 ;
        RECT 91.835 192.535 92.005 192.705 ;
        RECT 92.295 192.535 92.465 192.705 ;
        RECT 92.755 192.535 92.925 192.705 ;
        RECT 93.215 192.535 93.385 192.705 ;
        RECT 93.675 192.535 93.845 192.705 ;
        RECT 94.135 192.535 94.305 192.705 ;
        RECT 94.595 192.535 94.765 192.705 ;
        RECT 95.055 192.535 95.225 192.705 ;
        RECT 95.515 192.535 95.685 192.705 ;
        RECT 95.975 192.535 96.145 192.705 ;
        RECT 96.435 192.535 96.605 192.705 ;
        RECT 96.895 192.535 97.065 192.705 ;
        RECT 97.355 192.535 97.525 192.705 ;
        RECT 97.815 192.535 97.985 192.705 ;
        RECT 98.275 192.535 98.445 192.705 ;
        RECT 98.735 192.535 98.905 192.705 ;
        RECT 99.195 192.535 99.365 192.705 ;
        RECT 99.655 192.535 99.825 192.705 ;
        RECT 100.115 192.535 100.285 192.705 ;
        RECT 100.575 192.535 100.745 192.705 ;
        RECT 101.035 192.535 101.205 192.705 ;
        RECT 101.495 192.535 101.665 192.705 ;
        RECT 101.955 192.535 102.125 192.705 ;
        RECT 102.415 192.535 102.585 192.705 ;
        RECT 102.875 192.535 103.045 192.705 ;
        RECT 103.335 192.535 103.505 192.705 ;
        RECT 103.795 192.535 103.965 192.705 ;
        RECT 104.255 192.535 104.425 192.705 ;
        RECT 104.715 192.535 104.885 192.705 ;
        RECT 105.175 192.535 105.345 192.705 ;
        RECT 105.635 192.535 105.805 192.705 ;
        RECT 106.095 192.535 106.265 192.705 ;
        RECT 106.555 192.535 106.725 192.705 ;
        RECT 107.015 192.535 107.185 192.705 ;
        RECT 107.475 192.535 107.645 192.705 ;
        RECT 107.935 192.535 108.105 192.705 ;
        RECT 108.395 192.535 108.565 192.705 ;
        RECT 108.855 192.535 109.025 192.705 ;
        RECT 109.315 192.535 109.485 192.705 ;
        RECT 109.775 192.535 109.945 192.705 ;
        RECT 110.235 192.535 110.405 192.705 ;
        RECT 110.695 192.535 110.865 192.705 ;
        RECT 111.155 192.535 111.325 192.705 ;
        RECT 111.615 192.535 111.785 192.705 ;
        RECT 112.075 192.535 112.245 192.705 ;
        RECT 112.535 192.535 112.705 192.705 ;
        RECT 112.995 192.535 113.165 192.705 ;
        RECT 113.455 192.535 113.625 192.705 ;
        RECT 113.915 192.535 114.085 192.705 ;
        RECT 114.375 192.535 114.545 192.705 ;
        RECT 114.835 192.535 115.005 192.705 ;
        RECT 115.295 192.535 115.465 192.705 ;
        RECT 115.755 192.535 115.925 192.705 ;
        RECT 116.215 192.535 116.385 192.705 ;
        RECT 116.675 192.535 116.845 192.705 ;
        RECT 117.135 192.535 117.305 192.705 ;
        RECT 117.595 192.535 117.765 192.705 ;
        RECT 118.055 192.535 118.225 192.705 ;
        RECT 118.515 192.535 118.685 192.705 ;
        RECT 118.975 192.535 119.145 192.705 ;
        RECT 119.435 192.535 119.605 192.705 ;
        RECT 119.895 192.535 120.065 192.705 ;
        RECT 120.355 192.535 120.525 192.705 ;
        RECT 120.815 192.535 120.985 192.705 ;
        RECT 121.275 192.535 121.445 192.705 ;
        RECT 121.735 192.535 121.905 192.705 ;
        RECT 122.195 192.535 122.365 192.705 ;
        RECT 122.655 192.535 122.825 192.705 ;
        RECT 123.115 192.535 123.285 192.705 ;
        RECT 123.575 192.535 123.745 192.705 ;
        RECT 124.035 192.535 124.205 192.705 ;
        RECT 124.495 192.535 124.665 192.705 ;
        RECT 124.955 192.535 125.125 192.705 ;
        RECT 125.415 192.535 125.585 192.705 ;
        RECT 125.875 192.535 126.045 192.705 ;
        RECT 126.335 192.535 126.505 192.705 ;
        RECT 126.795 192.535 126.965 192.705 ;
        RECT 127.255 192.535 127.425 192.705 ;
        RECT 127.715 192.535 127.885 192.705 ;
        RECT 128.175 192.535 128.345 192.705 ;
        RECT 128.635 192.535 128.805 192.705 ;
        RECT 129.095 192.535 129.265 192.705 ;
        RECT 129.555 192.535 129.725 192.705 ;
        RECT 130.015 192.535 130.185 192.705 ;
        RECT 130.475 192.535 130.645 192.705 ;
        RECT 130.935 192.535 131.105 192.705 ;
        RECT 78.495 192.025 78.665 192.195 ;
        RECT 79.875 191.345 80.045 191.515 ;
        RECT 80.335 191.005 80.505 191.175 ;
        RECT 81.715 192.025 81.885 192.195 ;
        RECT 82.635 192.025 82.805 192.195 ;
        RECT 84.015 191.005 84.185 191.175 ;
        RECT 88.155 192.025 88.325 192.195 ;
        RECT 87.695 191.005 87.865 191.175 ;
        RECT 86.775 190.665 86.945 190.835 ;
        RECT 90.465 191.345 90.635 191.515 ;
        RECT 90.900 191.685 91.070 191.855 ;
        RECT 92.470 191.685 92.640 191.855 ;
        RECT 92.985 191.345 93.155 191.515 ;
        RECT 93.720 190.665 93.890 190.835 ;
        RECT 94.175 191.345 94.345 191.515 ;
        RECT 94.570 191.685 94.740 191.855 ;
        RECT 95.055 191.005 95.225 191.175 ;
        RECT 96.435 190.325 96.605 190.495 ;
        RECT 98.745 191.345 98.915 191.515 ;
        RECT 99.180 191.685 99.350 191.855 ;
        RECT 100.750 191.685 100.920 191.855 ;
        RECT 101.265 191.345 101.435 191.515 ;
        RECT 102.000 190.665 102.170 190.835 ;
        RECT 102.455 191.345 102.625 191.515 ;
        RECT 102.850 191.685 103.020 191.855 ;
        RECT 103.335 191.005 103.505 191.175 ;
        RECT 109.315 192.025 109.485 192.195 ;
        RECT 111.625 191.345 111.795 191.515 ;
        RECT 112.060 191.685 112.230 191.855 ;
        RECT 113.630 191.685 113.800 191.855 ;
        RECT 114.145 191.345 114.315 191.515 ;
        RECT 114.990 190.665 115.160 190.835 ;
        RECT 115.335 191.345 115.505 191.515 ;
        RECT 115.730 191.685 115.900 191.855 ;
        RECT 116.215 191.005 116.385 191.175 ;
        RECT 57.335 189.815 57.505 189.985 ;
        RECT 57.795 189.815 57.965 189.985 ;
        RECT 58.255 189.815 58.425 189.985 ;
        RECT 58.715 189.815 58.885 189.985 ;
        RECT 59.175 189.815 59.345 189.985 ;
        RECT 59.635 189.815 59.805 189.985 ;
        RECT 60.095 189.815 60.265 189.985 ;
        RECT 60.555 189.815 60.725 189.985 ;
        RECT 61.015 189.815 61.185 189.985 ;
        RECT 61.475 189.815 61.645 189.985 ;
        RECT 61.935 189.815 62.105 189.985 ;
        RECT 62.395 189.815 62.565 189.985 ;
        RECT 62.855 189.815 63.025 189.985 ;
        RECT 63.315 189.815 63.485 189.985 ;
        RECT 63.775 189.815 63.945 189.985 ;
        RECT 64.235 189.815 64.405 189.985 ;
        RECT 64.695 189.815 64.865 189.985 ;
        RECT 65.155 189.815 65.325 189.985 ;
        RECT 65.615 189.815 65.785 189.985 ;
        RECT 66.075 189.815 66.245 189.985 ;
        RECT 66.535 189.815 66.705 189.985 ;
        RECT 66.995 189.815 67.165 189.985 ;
        RECT 67.455 189.815 67.625 189.985 ;
        RECT 67.915 189.815 68.085 189.985 ;
        RECT 68.375 189.815 68.545 189.985 ;
        RECT 68.835 189.815 69.005 189.985 ;
        RECT 69.295 189.815 69.465 189.985 ;
        RECT 69.755 189.815 69.925 189.985 ;
        RECT 70.215 189.815 70.385 189.985 ;
        RECT 70.675 189.815 70.845 189.985 ;
        RECT 71.135 189.815 71.305 189.985 ;
        RECT 71.595 189.815 71.765 189.985 ;
        RECT 72.055 189.815 72.225 189.985 ;
        RECT 72.515 189.815 72.685 189.985 ;
        RECT 72.975 189.815 73.145 189.985 ;
        RECT 73.435 189.815 73.605 189.985 ;
        RECT 73.895 189.815 74.065 189.985 ;
        RECT 74.355 189.815 74.525 189.985 ;
        RECT 74.815 189.815 74.985 189.985 ;
        RECT 75.275 189.815 75.445 189.985 ;
        RECT 75.735 189.815 75.905 189.985 ;
        RECT 76.195 189.815 76.365 189.985 ;
        RECT 76.655 189.815 76.825 189.985 ;
        RECT 77.115 189.815 77.285 189.985 ;
        RECT 77.575 189.815 77.745 189.985 ;
        RECT 78.035 189.815 78.205 189.985 ;
        RECT 78.495 189.815 78.665 189.985 ;
        RECT 78.955 189.815 79.125 189.985 ;
        RECT 79.415 189.815 79.585 189.985 ;
        RECT 79.875 189.815 80.045 189.985 ;
        RECT 80.335 189.815 80.505 189.985 ;
        RECT 80.795 189.815 80.965 189.985 ;
        RECT 81.255 189.815 81.425 189.985 ;
        RECT 81.715 189.815 81.885 189.985 ;
        RECT 82.175 189.815 82.345 189.985 ;
        RECT 82.635 189.815 82.805 189.985 ;
        RECT 83.095 189.815 83.265 189.985 ;
        RECT 83.555 189.815 83.725 189.985 ;
        RECT 84.015 189.815 84.185 189.985 ;
        RECT 84.475 189.815 84.645 189.985 ;
        RECT 84.935 189.815 85.105 189.985 ;
        RECT 85.395 189.815 85.565 189.985 ;
        RECT 85.855 189.815 86.025 189.985 ;
        RECT 86.315 189.815 86.485 189.985 ;
        RECT 86.775 189.815 86.945 189.985 ;
        RECT 87.235 189.815 87.405 189.985 ;
        RECT 87.695 189.815 87.865 189.985 ;
        RECT 88.155 189.815 88.325 189.985 ;
        RECT 88.615 189.815 88.785 189.985 ;
        RECT 89.075 189.815 89.245 189.985 ;
        RECT 89.535 189.815 89.705 189.985 ;
        RECT 89.995 189.815 90.165 189.985 ;
        RECT 90.455 189.815 90.625 189.985 ;
        RECT 90.915 189.815 91.085 189.985 ;
        RECT 91.375 189.815 91.545 189.985 ;
        RECT 91.835 189.815 92.005 189.985 ;
        RECT 92.295 189.815 92.465 189.985 ;
        RECT 92.755 189.815 92.925 189.985 ;
        RECT 93.215 189.815 93.385 189.985 ;
        RECT 93.675 189.815 93.845 189.985 ;
        RECT 94.135 189.815 94.305 189.985 ;
        RECT 94.595 189.815 94.765 189.985 ;
        RECT 95.055 189.815 95.225 189.985 ;
        RECT 95.515 189.815 95.685 189.985 ;
        RECT 95.975 189.815 96.145 189.985 ;
        RECT 96.435 189.815 96.605 189.985 ;
        RECT 96.895 189.815 97.065 189.985 ;
        RECT 97.355 189.815 97.525 189.985 ;
        RECT 97.815 189.815 97.985 189.985 ;
        RECT 98.275 189.815 98.445 189.985 ;
        RECT 98.735 189.815 98.905 189.985 ;
        RECT 99.195 189.815 99.365 189.985 ;
        RECT 99.655 189.815 99.825 189.985 ;
        RECT 100.115 189.815 100.285 189.985 ;
        RECT 100.575 189.815 100.745 189.985 ;
        RECT 101.035 189.815 101.205 189.985 ;
        RECT 101.495 189.815 101.665 189.985 ;
        RECT 101.955 189.815 102.125 189.985 ;
        RECT 102.415 189.815 102.585 189.985 ;
        RECT 102.875 189.815 103.045 189.985 ;
        RECT 103.335 189.815 103.505 189.985 ;
        RECT 103.795 189.815 103.965 189.985 ;
        RECT 104.255 189.815 104.425 189.985 ;
        RECT 104.715 189.815 104.885 189.985 ;
        RECT 105.175 189.815 105.345 189.985 ;
        RECT 105.635 189.815 105.805 189.985 ;
        RECT 106.095 189.815 106.265 189.985 ;
        RECT 106.555 189.815 106.725 189.985 ;
        RECT 107.015 189.815 107.185 189.985 ;
        RECT 107.475 189.815 107.645 189.985 ;
        RECT 107.935 189.815 108.105 189.985 ;
        RECT 108.395 189.815 108.565 189.985 ;
        RECT 108.855 189.815 109.025 189.985 ;
        RECT 109.315 189.815 109.485 189.985 ;
        RECT 109.775 189.815 109.945 189.985 ;
        RECT 110.235 189.815 110.405 189.985 ;
        RECT 110.695 189.815 110.865 189.985 ;
        RECT 111.155 189.815 111.325 189.985 ;
        RECT 111.615 189.815 111.785 189.985 ;
        RECT 112.075 189.815 112.245 189.985 ;
        RECT 112.535 189.815 112.705 189.985 ;
        RECT 112.995 189.815 113.165 189.985 ;
        RECT 113.455 189.815 113.625 189.985 ;
        RECT 113.915 189.815 114.085 189.985 ;
        RECT 114.375 189.815 114.545 189.985 ;
        RECT 114.835 189.815 115.005 189.985 ;
        RECT 115.295 189.815 115.465 189.985 ;
        RECT 115.755 189.815 115.925 189.985 ;
        RECT 116.215 189.815 116.385 189.985 ;
        RECT 116.675 189.815 116.845 189.985 ;
        RECT 117.135 189.815 117.305 189.985 ;
        RECT 117.595 189.815 117.765 189.985 ;
        RECT 118.055 189.815 118.225 189.985 ;
        RECT 118.515 189.815 118.685 189.985 ;
        RECT 118.975 189.815 119.145 189.985 ;
        RECT 119.435 189.815 119.605 189.985 ;
        RECT 119.895 189.815 120.065 189.985 ;
        RECT 120.355 189.815 120.525 189.985 ;
        RECT 120.815 189.815 120.985 189.985 ;
        RECT 121.275 189.815 121.445 189.985 ;
        RECT 121.735 189.815 121.905 189.985 ;
        RECT 122.195 189.815 122.365 189.985 ;
        RECT 122.655 189.815 122.825 189.985 ;
        RECT 123.115 189.815 123.285 189.985 ;
        RECT 123.575 189.815 123.745 189.985 ;
        RECT 124.035 189.815 124.205 189.985 ;
        RECT 124.495 189.815 124.665 189.985 ;
        RECT 124.955 189.815 125.125 189.985 ;
        RECT 125.415 189.815 125.585 189.985 ;
        RECT 125.875 189.815 126.045 189.985 ;
        RECT 126.335 189.815 126.505 189.985 ;
        RECT 126.795 189.815 126.965 189.985 ;
        RECT 127.255 189.815 127.425 189.985 ;
        RECT 127.715 189.815 127.885 189.985 ;
        RECT 128.175 189.815 128.345 189.985 ;
        RECT 128.635 189.815 128.805 189.985 ;
        RECT 129.095 189.815 129.265 189.985 ;
        RECT 129.555 189.815 129.725 189.985 ;
        RECT 130.015 189.815 130.185 189.985 ;
        RECT 130.475 189.815 130.645 189.985 ;
        RECT 130.935 189.815 131.105 189.985 ;
        RECT 81.255 189.305 81.425 189.475 ;
        RECT 78.955 188.625 79.125 188.795 ;
        RECT 80.335 187.605 80.505 187.775 ;
        RECT 87.695 188.285 87.865 188.455 ;
        RECT 89.535 189.305 89.705 189.475 ;
        RECT 90.455 189.305 90.625 189.475 ;
        RECT 89.535 187.605 89.705 187.775 ;
        RECT 96.895 188.625 97.065 188.795 ;
        RECT 100.115 189.305 100.285 189.475 ;
        RECT 101.035 189.305 101.205 189.475 ;
        RECT 100.575 188.625 100.745 188.795 ;
        RECT 101.495 188.625 101.665 188.795 ;
        RECT 127.255 188.625 127.425 188.795 ;
        RECT 128.175 187.605 128.345 187.775 ;
        RECT 57.335 187.095 57.505 187.265 ;
        RECT 57.795 187.095 57.965 187.265 ;
        RECT 58.255 187.095 58.425 187.265 ;
        RECT 58.715 187.095 58.885 187.265 ;
        RECT 59.175 187.095 59.345 187.265 ;
        RECT 59.635 187.095 59.805 187.265 ;
        RECT 60.095 187.095 60.265 187.265 ;
        RECT 60.555 187.095 60.725 187.265 ;
        RECT 61.015 187.095 61.185 187.265 ;
        RECT 61.475 187.095 61.645 187.265 ;
        RECT 61.935 187.095 62.105 187.265 ;
        RECT 62.395 187.095 62.565 187.265 ;
        RECT 62.855 187.095 63.025 187.265 ;
        RECT 63.315 187.095 63.485 187.265 ;
        RECT 63.775 187.095 63.945 187.265 ;
        RECT 64.235 187.095 64.405 187.265 ;
        RECT 64.695 187.095 64.865 187.265 ;
        RECT 65.155 187.095 65.325 187.265 ;
        RECT 65.615 187.095 65.785 187.265 ;
        RECT 66.075 187.095 66.245 187.265 ;
        RECT 66.535 187.095 66.705 187.265 ;
        RECT 66.995 187.095 67.165 187.265 ;
        RECT 67.455 187.095 67.625 187.265 ;
        RECT 67.915 187.095 68.085 187.265 ;
        RECT 68.375 187.095 68.545 187.265 ;
        RECT 68.835 187.095 69.005 187.265 ;
        RECT 69.295 187.095 69.465 187.265 ;
        RECT 69.755 187.095 69.925 187.265 ;
        RECT 70.215 187.095 70.385 187.265 ;
        RECT 70.675 187.095 70.845 187.265 ;
        RECT 71.135 187.095 71.305 187.265 ;
        RECT 71.595 187.095 71.765 187.265 ;
        RECT 72.055 187.095 72.225 187.265 ;
        RECT 72.515 187.095 72.685 187.265 ;
        RECT 72.975 187.095 73.145 187.265 ;
        RECT 73.435 187.095 73.605 187.265 ;
        RECT 73.895 187.095 74.065 187.265 ;
        RECT 74.355 187.095 74.525 187.265 ;
        RECT 74.815 187.095 74.985 187.265 ;
        RECT 75.275 187.095 75.445 187.265 ;
        RECT 75.735 187.095 75.905 187.265 ;
        RECT 76.195 187.095 76.365 187.265 ;
        RECT 76.655 187.095 76.825 187.265 ;
        RECT 77.115 187.095 77.285 187.265 ;
        RECT 77.575 187.095 77.745 187.265 ;
        RECT 78.035 187.095 78.205 187.265 ;
        RECT 78.495 187.095 78.665 187.265 ;
        RECT 78.955 187.095 79.125 187.265 ;
        RECT 79.415 187.095 79.585 187.265 ;
        RECT 79.875 187.095 80.045 187.265 ;
        RECT 80.335 187.095 80.505 187.265 ;
        RECT 80.795 187.095 80.965 187.265 ;
        RECT 81.255 187.095 81.425 187.265 ;
        RECT 81.715 187.095 81.885 187.265 ;
        RECT 82.175 187.095 82.345 187.265 ;
        RECT 82.635 187.095 82.805 187.265 ;
        RECT 83.095 187.095 83.265 187.265 ;
        RECT 83.555 187.095 83.725 187.265 ;
        RECT 84.015 187.095 84.185 187.265 ;
        RECT 84.475 187.095 84.645 187.265 ;
        RECT 84.935 187.095 85.105 187.265 ;
        RECT 85.395 187.095 85.565 187.265 ;
        RECT 85.855 187.095 86.025 187.265 ;
        RECT 86.315 187.095 86.485 187.265 ;
        RECT 86.775 187.095 86.945 187.265 ;
        RECT 87.235 187.095 87.405 187.265 ;
        RECT 87.695 187.095 87.865 187.265 ;
        RECT 88.155 187.095 88.325 187.265 ;
        RECT 88.615 187.095 88.785 187.265 ;
        RECT 89.075 187.095 89.245 187.265 ;
        RECT 89.535 187.095 89.705 187.265 ;
        RECT 89.995 187.095 90.165 187.265 ;
        RECT 90.455 187.095 90.625 187.265 ;
        RECT 90.915 187.095 91.085 187.265 ;
        RECT 91.375 187.095 91.545 187.265 ;
        RECT 91.835 187.095 92.005 187.265 ;
        RECT 92.295 187.095 92.465 187.265 ;
        RECT 92.755 187.095 92.925 187.265 ;
        RECT 93.215 187.095 93.385 187.265 ;
        RECT 93.675 187.095 93.845 187.265 ;
        RECT 94.135 187.095 94.305 187.265 ;
        RECT 94.595 187.095 94.765 187.265 ;
        RECT 95.055 187.095 95.225 187.265 ;
        RECT 95.515 187.095 95.685 187.265 ;
        RECT 95.975 187.095 96.145 187.265 ;
        RECT 96.435 187.095 96.605 187.265 ;
        RECT 96.895 187.095 97.065 187.265 ;
        RECT 97.355 187.095 97.525 187.265 ;
        RECT 97.815 187.095 97.985 187.265 ;
        RECT 98.275 187.095 98.445 187.265 ;
        RECT 98.735 187.095 98.905 187.265 ;
        RECT 99.195 187.095 99.365 187.265 ;
        RECT 99.655 187.095 99.825 187.265 ;
        RECT 100.115 187.095 100.285 187.265 ;
        RECT 100.575 187.095 100.745 187.265 ;
        RECT 101.035 187.095 101.205 187.265 ;
        RECT 101.495 187.095 101.665 187.265 ;
        RECT 101.955 187.095 102.125 187.265 ;
        RECT 102.415 187.095 102.585 187.265 ;
        RECT 102.875 187.095 103.045 187.265 ;
        RECT 103.335 187.095 103.505 187.265 ;
        RECT 103.795 187.095 103.965 187.265 ;
        RECT 104.255 187.095 104.425 187.265 ;
        RECT 104.715 187.095 104.885 187.265 ;
        RECT 105.175 187.095 105.345 187.265 ;
        RECT 105.635 187.095 105.805 187.265 ;
        RECT 106.095 187.095 106.265 187.265 ;
        RECT 106.555 187.095 106.725 187.265 ;
        RECT 107.015 187.095 107.185 187.265 ;
        RECT 107.475 187.095 107.645 187.265 ;
        RECT 107.935 187.095 108.105 187.265 ;
        RECT 108.395 187.095 108.565 187.265 ;
        RECT 108.855 187.095 109.025 187.265 ;
        RECT 109.315 187.095 109.485 187.265 ;
        RECT 109.775 187.095 109.945 187.265 ;
        RECT 110.235 187.095 110.405 187.265 ;
        RECT 110.695 187.095 110.865 187.265 ;
        RECT 111.155 187.095 111.325 187.265 ;
        RECT 111.615 187.095 111.785 187.265 ;
        RECT 112.075 187.095 112.245 187.265 ;
        RECT 112.535 187.095 112.705 187.265 ;
        RECT 112.995 187.095 113.165 187.265 ;
        RECT 113.455 187.095 113.625 187.265 ;
        RECT 113.915 187.095 114.085 187.265 ;
        RECT 114.375 187.095 114.545 187.265 ;
        RECT 114.835 187.095 115.005 187.265 ;
        RECT 115.295 187.095 115.465 187.265 ;
        RECT 115.755 187.095 115.925 187.265 ;
        RECT 116.215 187.095 116.385 187.265 ;
        RECT 116.675 187.095 116.845 187.265 ;
        RECT 117.135 187.095 117.305 187.265 ;
        RECT 117.595 187.095 117.765 187.265 ;
        RECT 118.055 187.095 118.225 187.265 ;
        RECT 118.515 187.095 118.685 187.265 ;
        RECT 118.975 187.095 119.145 187.265 ;
        RECT 119.435 187.095 119.605 187.265 ;
        RECT 119.895 187.095 120.065 187.265 ;
        RECT 120.355 187.095 120.525 187.265 ;
        RECT 120.815 187.095 120.985 187.265 ;
        RECT 121.275 187.095 121.445 187.265 ;
        RECT 121.735 187.095 121.905 187.265 ;
        RECT 122.195 187.095 122.365 187.265 ;
        RECT 122.655 187.095 122.825 187.265 ;
        RECT 123.115 187.095 123.285 187.265 ;
        RECT 123.575 187.095 123.745 187.265 ;
        RECT 124.035 187.095 124.205 187.265 ;
        RECT 124.495 187.095 124.665 187.265 ;
        RECT 124.955 187.095 125.125 187.265 ;
        RECT 125.415 187.095 125.585 187.265 ;
        RECT 125.875 187.095 126.045 187.265 ;
        RECT 126.335 187.095 126.505 187.265 ;
        RECT 126.795 187.095 126.965 187.265 ;
        RECT 127.255 187.095 127.425 187.265 ;
        RECT 127.715 187.095 127.885 187.265 ;
        RECT 128.175 187.095 128.345 187.265 ;
        RECT 128.635 187.095 128.805 187.265 ;
        RECT 129.095 187.095 129.265 187.265 ;
        RECT 129.555 187.095 129.725 187.265 ;
        RECT 130.015 187.095 130.185 187.265 ;
        RECT 130.475 187.095 130.645 187.265 ;
        RECT 130.935 187.095 131.105 187.265 ;
        RECT 57.335 184.375 57.505 184.545 ;
        RECT 57.795 184.375 57.965 184.545 ;
        RECT 58.255 184.375 58.425 184.545 ;
        RECT 58.715 184.375 58.885 184.545 ;
        RECT 59.175 184.375 59.345 184.545 ;
        RECT 59.635 184.375 59.805 184.545 ;
        RECT 60.095 184.375 60.265 184.545 ;
        RECT 60.555 184.375 60.725 184.545 ;
        RECT 61.015 184.375 61.185 184.545 ;
        RECT 61.475 184.375 61.645 184.545 ;
        RECT 61.935 184.375 62.105 184.545 ;
        RECT 62.395 184.375 62.565 184.545 ;
        RECT 62.855 184.375 63.025 184.545 ;
        RECT 63.315 184.375 63.485 184.545 ;
        RECT 63.775 184.375 63.945 184.545 ;
        RECT 64.235 184.375 64.405 184.545 ;
        RECT 64.695 184.375 64.865 184.545 ;
        RECT 65.155 184.375 65.325 184.545 ;
        RECT 65.615 184.375 65.785 184.545 ;
        RECT 66.075 184.375 66.245 184.545 ;
        RECT 66.535 184.375 66.705 184.545 ;
        RECT 66.995 184.375 67.165 184.545 ;
        RECT 67.455 184.375 67.625 184.545 ;
        RECT 67.915 184.375 68.085 184.545 ;
        RECT 68.375 184.375 68.545 184.545 ;
        RECT 68.835 184.375 69.005 184.545 ;
        RECT 69.295 184.375 69.465 184.545 ;
        RECT 69.755 184.375 69.925 184.545 ;
        RECT 70.215 184.375 70.385 184.545 ;
        RECT 70.675 184.375 70.845 184.545 ;
        RECT 71.135 184.375 71.305 184.545 ;
        RECT 71.595 184.375 71.765 184.545 ;
        RECT 72.055 184.375 72.225 184.545 ;
        RECT 72.515 184.375 72.685 184.545 ;
        RECT 72.975 184.375 73.145 184.545 ;
        RECT 73.435 184.375 73.605 184.545 ;
        RECT 73.895 184.375 74.065 184.545 ;
        RECT 74.355 184.375 74.525 184.545 ;
        RECT 74.815 184.375 74.985 184.545 ;
        RECT 75.275 184.375 75.445 184.545 ;
        RECT 75.735 184.375 75.905 184.545 ;
        RECT 76.195 184.375 76.365 184.545 ;
        RECT 76.655 184.375 76.825 184.545 ;
        RECT 77.115 184.375 77.285 184.545 ;
        RECT 77.575 184.375 77.745 184.545 ;
        RECT 78.035 184.375 78.205 184.545 ;
        RECT 78.495 184.375 78.665 184.545 ;
        RECT 78.955 184.375 79.125 184.545 ;
        RECT 79.415 184.375 79.585 184.545 ;
        RECT 79.875 184.375 80.045 184.545 ;
        RECT 80.335 184.375 80.505 184.545 ;
        RECT 80.795 184.375 80.965 184.545 ;
        RECT 81.255 184.375 81.425 184.545 ;
        RECT 81.715 184.375 81.885 184.545 ;
        RECT 82.175 184.375 82.345 184.545 ;
        RECT 82.635 184.375 82.805 184.545 ;
        RECT 83.095 184.375 83.265 184.545 ;
        RECT 83.555 184.375 83.725 184.545 ;
        RECT 84.015 184.375 84.185 184.545 ;
        RECT 84.475 184.375 84.645 184.545 ;
        RECT 84.935 184.375 85.105 184.545 ;
        RECT 85.395 184.375 85.565 184.545 ;
        RECT 85.855 184.375 86.025 184.545 ;
        RECT 86.315 184.375 86.485 184.545 ;
        RECT 86.775 184.375 86.945 184.545 ;
        RECT 87.235 184.375 87.405 184.545 ;
        RECT 87.695 184.375 87.865 184.545 ;
        RECT 88.155 184.375 88.325 184.545 ;
        RECT 88.615 184.375 88.785 184.545 ;
        RECT 89.075 184.375 89.245 184.545 ;
        RECT 89.535 184.375 89.705 184.545 ;
        RECT 89.995 184.375 90.165 184.545 ;
        RECT 90.455 184.375 90.625 184.545 ;
        RECT 90.915 184.375 91.085 184.545 ;
        RECT 91.375 184.375 91.545 184.545 ;
        RECT 91.835 184.375 92.005 184.545 ;
        RECT 92.295 184.375 92.465 184.545 ;
        RECT 92.755 184.375 92.925 184.545 ;
        RECT 93.215 184.375 93.385 184.545 ;
        RECT 93.675 184.375 93.845 184.545 ;
        RECT 94.135 184.375 94.305 184.545 ;
        RECT 94.595 184.375 94.765 184.545 ;
        RECT 95.055 184.375 95.225 184.545 ;
        RECT 95.515 184.375 95.685 184.545 ;
        RECT 95.975 184.375 96.145 184.545 ;
        RECT 96.435 184.375 96.605 184.545 ;
        RECT 96.895 184.375 97.065 184.545 ;
        RECT 97.355 184.375 97.525 184.545 ;
        RECT 97.815 184.375 97.985 184.545 ;
        RECT 98.275 184.375 98.445 184.545 ;
        RECT 98.735 184.375 98.905 184.545 ;
        RECT 99.195 184.375 99.365 184.545 ;
        RECT 99.655 184.375 99.825 184.545 ;
        RECT 100.115 184.375 100.285 184.545 ;
        RECT 100.575 184.375 100.745 184.545 ;
        RECT 101.035 184.375 101.205 184.545 ;
        RECT 101.495 184.375 101.665 184.545 ;
        RECT 101.955 184.375 102.125 184.545 ;
        RECT 102.415 184.375 102.585 184.545 ;
        RECT 102.875 184.375 103.045 184.545 ;
        RECT 103.335 184.375 103.505 184.545 ;
        RECT 103.795 184.375 103.965 184.545 ;
        RECT 104.255 184.375 104.425 184.545 ;
        RECT 104.715 184.375 104.885 184.545 ;
        RECT 105.175 184.375 105.345 184.545 ;
        RECT 105.635 184.375 105.805 184.545 ;
        RECT 106.095 184.375 106.265 184.545 ;
        RECT 106.555 184.375 106.725 184.545 ;
        RECT 107.015 184.375 107.185 184.545 ;
        RECT 107.475 184.375 107.645 184.545 ;
        RECT 107.935 184.375 108.105 184.545 ;
        RECT 108.395 184.375 108.565 184.545 ;
        RECT 108.855 184.375 109.025 184.545 ;
        RECT 109.315 184.375 109.485 184.545 ;
        RECT 109.775 184.375 109.945 184.545 ;
        RECT 110.235 184.375 110.405 184.545 ;
        RECT 110.695 184.375 110.865 184.545 ;
        RECT 111.155 184.375 111.325 184.545 ;
        RECT 111.615 184.375 111.785 184.545 ;
        RECT 112.075 184.375 112.245 184.545 ;
        RECT 112.535 184.375 112.705 184.545 ;
        RECT 112.995 184.375 113.165 184.545 ;
        RECT 113.455 184.375 113.625 184.545 ;
        RECT 113.915 184.375 114.085 184.545 ;
        RECT 114.375 184.375 114.545 184.545 ;
        RECT 114.835 184.375 115.005 184.545 ;
        RECT 115.295 184.375 115.465 184.545 ;
        RECT 115.755 184.375 115.925 184.545 ;
        RECT 116.215 184.375 116.385 184.545 ;
        RECT 116.675 184.375 116.845 184.545 ;
        RECT 117.135 184.375 117.305 184.545 ;
        RECT 117.595 184.375 117.765 184.545 ;
        RECT 118.055 184.375 118.225 184.545 ;
        RECT 118.515 184.375 118.685 184.545 ;
        RECT 118.975 184.375 119.145 184.545 ;
        RECT 119.435 184.375 119.605 184.545 ;
        RECT 119.895 184.375 120.065 184.545 ;
        RECT 120.355 184.375 120.525 184.545 ;
        RECT 120.815 184.375 120.985 184.545 ;
        RECT 121.275 184.375 121.445 184.545 ;
        RECT 121.735 184.375 121.905 184.545 ;
        RECT 122.195 184.375 122.365 184.545 ;
        RECT 122.655 184.375 122.825 184.545 ;
        RECT 123.115 184.375 123.285 184.545 ;
        RECT 123.575 184.375 123.745 184.545 ;
        RECT 124.035 184.375 124.205 184.545 ;
        RECT 124.495 184.375 124.665 184.545 ;
        RECT 124.955 184.375 125.125 184.545 ;
        RECT 125.415 184.375 125.585 184.545 ;
        RECT 125.875 184.375 126.045 184.545 ;
        RECT 126.335 184.375 126.505 184.545 ;
        RECT 126.795 184.375 126.965 184.545 ;
        RECT 127.255 184.375 127.425 184.545 ;
        RECT 127.715 184.375 127.885 184.545 ;
        RECT 128.175 184.375 128.345 184.545 ;
        RECT 128.635 184.375 128.805 184.545 ;
        RECT 129.095 184.375 129.265 184.545 ;
        RECT 129.555 184.375 129.725 184.545 ;
        RECT 130.015 184.375 130.185 184.545 ;
        RECT 130.475 184.375 130.645 184.545 ;
        RECT 130.935 184.375 131.105 184.545 ;
        RECT 57.335 181.655 57.505 181.825 ;
        RECT 57.795 181.655 57.965 181.825 ;
        RECT 58.255 181.655 58.425 181.825 ;
        RECT 58.715 181.655 58.885 181.825 ;
        RECT 59.175 181.655 59.345 181.825 ;
        RECT 59.635 181.655 59.805 181.825 ;
        RECT 60.095 181.655 60.265 181.825 ;
        RECT 60.555 181.655 60.725 181.825 ;
        RECT 61.015 181.655 61.185 181.825 ;
        RECT 61.475 181.655 61.645 181.825 ;
        RECT 61.935 181.655 62.105 181.825 ;
        RECT 62.395 181.655 62.565 181.825 ;
        RECT 62.855 181.655 63.025 181.825 ;
        RECT 63.315 181.655 63.485 181.825 ;
        RECT 63.775 181.655 63.945 181.825 ;
        RECT 64.235 181.655 64.405 181.825 ;
        RECT 64.695 181.655 64.865 181.825 ;
        RECT 65.155 181.655 65.325 181.825 ;
        RECT 65.615 181.655 65.785 181.825 ;
        RECT 66.075 181.655 66.245 181.825 ;
        RECT 66.535 181.655 66.705 181.825 ;
        RECT 66.995 181.655 67.165 181.825 ;
        RECT 67.455 181.655 67.625 181.825 ;
        RECT 67.915 181.655 68.085 181.825 ;
        RECT 68.375 181.655 68.545 181.825 ;
        RECT 68.835 181.655 69.005 181.825 ;
        RECT 69.295 181.655 69.465 181.825 ;
        RECT 69.755 181.655 69.925 181.825 ;
        RECT 70.215 181.655 70.385 181.825 ;
        RECT 70.675 181.655 70.845 181.825 ;
        RECT 71.135 181.655 71.305 181.825 ;
        RECT 71.595 181.655 71.765 181.825 ;
        RECT 72.055 181.655 72.225 181.825 ;
        RECT 72.515 181.655 72.685 181.825 ;
        RECT 72.975 181.655 73.145 181.825 ;
        RECT 73.435 181.655 73.605 181.825 ;
        RECT 73.895 181.655 74.065 181.825 ;
        RECT 74.355 181.655 74.525 181.825 ;
        RECT 74.815 181.655 74.985 181.825 ;
        RECT 75.275 181.655 75.445 181.825 ;
        RECT 75.735 181.655 75.905 181.825 ;
        RECT 76.195 181.655 76.365 181.825 ;
        RECT 76.655 181.655 76.825 181.825 ;
        RECT 77.115 181.655 77.285 181.825 ;
        RECT 77.575 181.655 77.745 181.825 ;
        RECT 78.035 181.655 78.205 181.825 ;
        RECT 78.495 181.655 78.665 181.825 ;
        RECT 78.955 181.655 79.125 181.825 ;
        RECT 79.415 181.655 79.585 181.825 ;
        RECT 79.875 181.655 80.045 181.825 ;
        RECT 80.335 181.655 80.505 181.825 ;
        RECT 80.795 181.655 80.965 181.825 ;
        RECT 81.255 181.655 81.425 181.825 ;
        RECT 81.715 181.655 81.885 181.825 ;
        RECT 82.175 181.655 82.345 181.825 ;
        RECT 82.635 181.655 82.805 181.825 ;
        RECT 83.095 181.655 83.265 181.825 ;
        RECT 83.555 181.655 83.725 181.825 ;
        RECT 84.015 181.655 84.185 181.825 ;
        RECT 84.475 181.655 84.645 181.825 ;
        RECT 84.935 181.655 85.105 181.825 ;
        RECT 85.395 181.655 85.565 181.825 ;
        RECT 85.855 181.655 86.025 181.825 ;
        RECT 86.315 181.655 86.485 181.825 ;
        RECT 86.775 181.655 86.945 181.825 ;
        RECT 87.235 181.655 87.405 181.825 ;
        RECT 87.695 181.655 87.865 181.825 ;
        RECT 88.155 181.655 88.325 181.825 ;
        RECT 88.615 181.655 88.785 181.825 ;
        RECT 89.075 181.655 89.245 181.825 ;
        RECT 89.535 181.655 89.705 181.825 ;
        RECT 89.995 181.655 90.165 181.825 ;
        RECT 90.455 181.655 90.625 181.825 ;
        RECT 90.915 181.655 91.085 181.825 ;
        RECT 91.375 181.655 91.545 181.825 ;
        RECT 91.835 181.655 92.005 181.825 ;
        RECT 92.295 181.655 92.465 181.825 ;
        RECT 92.755 181.655 92.925 181.825 ;
        RECT 93.215 181.655 93.385 181.825 ;
        RECT 93.675 181.655 93.845 181.825 ;
        RECT 94.135 181.655 94.305 181.825 ;
        RECT 94.595 181.655 94.765 181.825 ;
        RECT 95.055 181.655 95.225 181.825 ;
        RECT 95.515 181.655 95.685 181.825 ;
        RECT 95.975 181.655 96.145 181.825 ;
        RECT 96.435 181.655 96.605 181.825 ;
        RECT 96.895 181.655 97.065 181.825 ;
        RECT 97.355 181.655 97.525 181.825 ;
        RECT 97.815 181.655 97.985 181.825 ;
        RECT 98.275 181.655 98.445 181.825 ;
        RECT 98.735 181.655 98.905 181.825 ;
        RECT 99.195 181.655 99.365 181.825 ;
        RECT 99.655 181.655 99.825 181.825 ;
        RECT 100.115 181.655 100.285 181.825 ;
        RECT 100.575 181.655 100.745 181.825 ;
        RECT 101.035 181.655 101.205 181.825 ;
        RECT 101.495 181.655 101.665 181.825 ;
        RECT 101.955 181.655 102.125 181.825 ;
        RECT 102.415 181.655 102.585 181.825 ;
        RECT 102.875 181.655 103.045 181.825 ;
        RECT 103.335 181.655 103.505 181.825 ;
        RECT 103.795 181.655 103.965 181.825 ;
        RECT 104.255 181.655 104.425 181.825 ;
        RECT 104.715 181.655 104.885 181.825 ;
        RECT 105.175 181.655 105.345 181.825 ;
        RECT 105.635 181.655 105.805 181.825 ;
        RECT 106.095 181.655 106.265 181.825 ;
        RECT 106.555 181.655 106.725 181.825 ;
        RECT 107.015 181.655 107.185 181.825 ;
        RECT 107.475 181.655 107.645 181.825 ;
        RECT 107.935 181.655 108.105 181.825 ;
        RECT 108.395 181.655 108.565 181.825 ;
        RECT 108.855 181.655 109.025 181.825 ;
        RECT 109.315 181.655 109.485 181.825 ;
        RECT 109.775 181.655 109.945 181.825 ;
        RECT 110.235 181.655 110.405 181.825 ;
        RECT 110.695 181.655 110.865 181.825 ;
        RECT 111.155 181.655 111.325 181.825 ;
        RECT 111.615 181.655 111.785 181.825 ;
        RECT 112.075 181.655 112.245 181.825 ;
        RECT 112.535 181.655 112.705 181.825 ;
        RECT 112.995 181.655 113.165 181.825 ;
        RECT 113.455 181.655 113.625 181.825 ;
        RECT 113.915 181.655 114.085 181.825 ;
        RECT 114.375 181.655 114.545 181.825 ;
        RECT 114.835 181.655 115.005 181.825 ;
        RECT 115.295 181.655 115.465 181.825 ;
        RECT 115.755 181.655 115.925 181.825 ;
        RECT 116.215 181.655 116.385 181.825 ;
        RECT 116.675 181.655 116.845 181.825 ;
        RECT 117.135 181.655 117.305 181.825 ;
        RECT 117.595 181.655 117.765 181.825 ;
        RECT 118.055 181.655 118.225 181.825 ;
        RECT 118.515 181.655 118.685 181.825 ;
        RECT 118.975 181.655 119.145 181.825 ;
        RECT 119.435 181.655 119.605 181.825 ;
        RECT 119.895 181.655 120.065 181.825 ;
        RECT 120.355 181.655 120.525 181.825 ;
        RECT 120.815 181.655 120.985 181.825 ;
        RECT 121.275 181.655 121.445 181.825 ;
        RECT 121.735 181.655 121.905 181.825 ;
        RECT 122.195 181.655 122.365 181.825 ;
        RECT 122.655 181.655 122.825 181.825 ;
        RECT 123.115 181.655 123.285 181.825 ;
        RECT 123.575 181.655 123.745 181.825 ;
        RECT 124.035 181.655 124.205 181.825 ;
        RECT 124.495 181.655 124.665 181.825 ;
        RECT 124.955 181.655 125.125 181.825 ;
        RECT 125.415 181.655 125.585 181.825 ;
        RECT 125.875 181.655 126.045 181.825 ;
        RECT 126.335 181.655 126.505 181.825 ;
        RECT 126.795 181.655 126.965 181.825 ;
        RECT 127.255 181.655 127.425 181.825 ;
        RECT 127.715 181.655 127.885 181.825 ;
        RECT 128.175 181.655 128.345 181.825 ;
        RECT 128.635 181.655 128.805 181.825 ;
        RECT 129.095 181.655 129.265 181.825 ;
        RECT 129.555 181.655 129.725 181.825 ;
        RECT 130.015 181.655 130.185 181.825 ;
        RECT 130.475 181.655 130.645 181.825 ;
        RECT 130.935 181.655 131.105 181.825 ;
        RECT 57.335 178.935 57.505 179.105 ;
        RECT 57.795 178.935 57.965 179.105 ;
        RECT 58.255 178.935 58.425 179.105 ;
        RECT 58.715 178.935 58.885 179.105 ;
        RECT 59.175 178.935 59.345 179.105 ;
        RECT 59.635 178.935 59.805 179.105 ;
        RECT 60.095 178.935 60.265 179.105 ;
        RECT 60.555 178.935 60.725 179.105 ;
        RECT 61.015 178.935 61.185 179.105 ;
        RECT 61.475 178.935 61.645 179.105 ;
        RECT 61.935 178.935 62.105 179.105 ;
        RECT 62.395 178.935 62.565 179.105 ;
        RECT 62.855 178.935 63.025 179.105 ;
        RECT 63.315 178.935 63.485 179.105 ;
        RECT 63.775 178.935 63.945 179.105 ;
        RECT 64.235 178.935 64.405 179.105 ;
        RECT 64.695 178.935 64.865 179.105 ;
        RECT 65.155 178.935 65.325 179.105 ;
        RECT 65.615 178.935 65.785 179.105 ;
        RECT 66.075 178.935 66.245 179.105 ;
        RECT 66.535 178.935 66.705 179.105 ;
        RECT 66.995 178.935 67.165 179.105 ;
        RECT 67.455 178.935 67.625 179.105 ;
        RECT 67.915 178.935 68.085 179.105 ;
        RECT 68.375 178.935 68.545 179.105 ;
        RECT 68.835 178.935 69.005 179.105 ;
        RECT 69.295 178.935 69.465 179.105 ;
        RECT 69.755 178.935 69.925 179.105 ;
        RECT 70.215 178.935 70.385 179.105 ;
        RECT 70.675 178.935 70.845 179.105 ;
        RECT 71.135 178.935 71.305 179.105 ;
        RECT 71.595 178.935 71.765 179.105 ;
        RECT 72.055 178.935 72.225 179.105 ;
        RECT 72.515 178.935 72.685 179.105 ;
        RECT 72.975 178.935 73.145 179.105 ;
        RECT 73.435 178.935 73.605 179.105 ;
        RECT 73.895 178.935 74.065 179.105 ;
        RECT 74.355 178.935 74.525 179.105 ;
        RECT 74.815 178.935 74.985 179.105 ;
        RECT 75.275 178.935 75.445 179.105 ;
        RECT 75.735 178.935 75.905 179.105 ;
        RECT 76.195 178.935 76.365 179.105 ;
        RECT 76.655 178.935 76.825 179.105 ;
        RECT 77.115 178.935 77.285 179.105 ;
        RECT 77.575 178.935 77.745 179.105 ;
        RECT 78.035 178.935 78.205 179.105 ;
        RECT 78.495 178.935 78.665 179.105 ;
        RECT 78.955 178.935 79.125 179.105 ;
        RECT 79.415 178.935 79.585 179.105 ;
        RECT 79.875 178.935 80.045 179.105 ;
        RECT 80.335 178.935 80.505 179.105 ;
        RECT 80.795 178.935 80.965 179.105 ;
        RECT 81.255 178.935 81.425 179.105 ;
        RECT 81.715 178.935 81.885 179.105 ;
        RECT 82.175 178.935 82.345 179.105 ;
        RECT 82.635 178.935 82.805 179.105 ;
        RECT 83.095 178.935 83.265 179.105 ;
        RECT 83.555 178.935 83.725 179.105 ;
        RECT 84.015 178.935 84.185 179.105 ;
        RECT 84.475 178.935 84.645 179.105 ;
        RECT 84.935 178.935 85.105 179.105 ;
        RECT 85.395 178.935 85.565 179.105 ;
        RECT 85.855 178.935 86.025 179.105 ;
        RECT 86.315 178.935 86.485 179.105 ;
        RECT 86.775 178.935 86.945 179.105 ;
        RECT 87.235 178.935 87.405 179.105 ;
        RECT 87.695 178.935 87.865 179.105 ;
        RECT 88.155 178.935 88.325 179.105 ;
        RECT 88.615 178.935 88.785 179.105 ;
        RECT 89.075 178.935 89.245 179.105 ;
        RECT 89.535 178.935 89.705 179.105 ;
        RECT 89.995 178.935 90.165 179.105 ;
        RECT 90.455 178.935 90.625 179.105 ;
        RECT 90.915 178.935 91.085 179.105 ;
        RECT 91.375 178.935 91.545 179.105 ;
        RECT 91.835 178.935 92.005 179.105 ;
        RECT 92.295 178.935 92.465 179.105 ;
        RECT 92.755 178.935 92.925 179.105 ;
        RECT 93.215 178.935 93.385 179.105 ;
        RECT 93.675 178.935 93.845 179.105 ;
        RECT 94.135 178.935 94.305 179.105 ;
        RECT 94.595 178.935 94.765 179.105 ;
        RECT 95.055 178.935 95.225 179.105 ;
        RECT 95.515 178.935 95.685 179.105 ;
        RECT 95.975 178.935 96.145 179.105 ;
        RECT 96.435 178.935 96.605 179.105 ;
        RECT 96.895 178.935 97.065 179.105 ;
        RECT 97.355 178.935 97.525 179.105 ;
        RECT 97.815 178.935 97.985 179.105 ;
        RECT 98.275 178.935 98.445 179.105 ;
        RECT 98.735 178.935 98.905 179.105 ;
        RECT 99.195 178.935 99.365 179.105 ;
        RECT 99.655 178.935 99.825 179.105 ;
        RECT 100.115 178.935 100.285 179.105 ;
        RECT 100.575 178.935 100.745 179.105 ;
        RECT 101.035 178.935 101.205 179.105 ;
        RECT 101.495 178.935 101.665 179.105 ;
        RECT 101.955 178.935 102.125 179.105 ;
        RECT 102.415 178.935 102.585 179.105 ;
        RECT 102.875 178.935 103.045 179.105 ;
        RECT 103.335 178.935 103.505 179.105 ;
        RECT 103.795 178.935 103.965 179.105 ;
        RECT 104.255 178.935 104.425 179.105 ;
        RECT 104.715 178.935 104.885 179.105 ;
        RECT 105.175 178.935 105.345 179.105 ;
        RECT 105.635 178.935 105.805 179.105 ;
        RECT 106.095 178.935 106.265 179.105 ;
        RECT 106.555 178.935 106.725 179.105 ;
        RECT 107.015 178.935 107.185 179.105 ;
        RECT 107.475 178.935 107.645 179.105 ;
        RECT 107.935 178.935 108.105 179.105 ;
        RECT 108.395 178.935 108.565 179.105 ;
        RECT 108.855 178.935 109.025 179.105 ;
        RECT 109.315 178.935 109.485 179.105 ;
        RECT 109.775 178.935 109.945 179.105 ;
        RECT 110.235 178.935 110.405 179.105 ;
        RECT 110.695 178.935 110.865 179.105 ;
        RECT 111.155 178.935 111.325 179.105 ;
        RECT 111.615 178.935 111.785 179.105 ;
        RECT 112.075 178.935 112.245 179.105 ;
        RECT 112.535 178.935 112.705 179.105 ;
        RECT 112.995 178.935 113.165 179.105 ;
        RECT 113.455 178.935 113.625 179.105 ;
        RECT 113.915 178.935 114.085 179.105 ;
        RECT 114.375 178.935 114.545 179.105 ;
        RECT 114.835 178.935 115.005 179.105 ;
        RECT 115.295 178.935 115.465 179.105 ;
        RECT 115.755 178.935 115.925 179.105 ;
        RECT 116.215 178.935 116.385 179.105 ;
        RECT 116.675 178.935 116.845 179.105 ;
        RECT 117.135 178.935 117.305 179.105 ;
        RECT 117.595 178.935 117.765 179.105 ;
        RECT 118.055 178.935 118.225 179.105 ;
        RECT 118.515 178.935 118.685 179.105 ;
        RECT 118.975 178.935 119.145 179.105 ;
        RECT 119.435 178.935 119.605 179.105 ;
        RECT 119.895 178.935 120.065 179.105 ;
        RECT 120.355 178.935 120.525 179.105 ;
        RECT 120.815 178.935 120.985 179.105 ;
        RECT 121.275 178.935 121.445 179.105 ;
        RECT 121.735 178.935 121.905 179.105 ;
        RECT 122.195 178.935 122.365 179.105 ;
        RECT 122.655 178.935 122.825 179.105 ;
        RECT 123.115 178.935 123.285 179.105 ;
        RECT 123.575 178.935 123.745 179.105 ;
        RECT 124.035 178.935 124.205 179.105 ;
        RECT 124.495 178.935 124.665 179.105 ;
        RECT 124.955 178.935 125.125 179.105 ;
        RECT 125.415 178.935 125.585 179.105 ;
        RECT 125.875 178.935 126.045 179.105 ;
        RECT 126.335 178.935 126.505 179.105 ;
        RECT 126.795 178.935 126.965 179.105 ;
        RECT 127.255 178.935 127.425 179.105 ;
        RECT 127.715 178.935 127.885 179.105 ;
        RECT 128.175 178.935 128.345 179.105 ;
        RECT 128.635 178.935 128.805 179.105 ;
        RECT 129.095 178.935 129.265 179.105 ;
        RECT 129.555 178.935 129.725 179.105 ;
        RECT 130.015 178.935 130.185 179.105 ;
        RECT 130.475 178.935 130.645 179.105 ;
        RECT 130.935 178.935 131.105 179.105 ;
        RECT 57.335 176.215 57.505 176.385 ;
        RECT 57.795 176.215 57.965 176.385 ;
        RECT 58.255 176.215 58.425 176.385 ;
        RECT 58.715 176.215 58.885 176.385 ;
        RECT 59.175 176.215 59.345 176.385 ;
        RECT 59.635 176.215 59.805 176.385 ;
        RECT 60.095 176.215 60.265 176.385 ;
        RECT 60.555 176.215 60.725 176.385 ;
        RECT 61.015 176.215 61.185 176.385 ;
        RECT 61.475 176.215 61.645 176.385 ;
        RECT 61.935 176.215 62.105 176.385 ;
        RECT 62.395 176.215 62.565 176.385 ;
        RECT 62.855 176.215 63.025 176.385 ;
        RECT 63.315 176.215 63.485 176.385 ;
        RECT 63.775 176.215 63.945 176.385 ;
        RECT 64.235 176.215 64.405 176.385 ;
        RECT 64.695 176.215 64.865 176.385 ;
        RECT 65.155 176.215 65.325 176.385 ;
        RECT 65.615 176.215 65.785 176.385 ;
        RECT 66.075 176.215 66.245 176.385 ;
        RECT 66.535 176.215 66.705 176.385 ;
        RECT 66.995 176.215 67.165 176.385 ;
        RECT 67.455 176.215 67.625 176.385 ;
        RECT 67.915 176.215 68.085 176.385 ;
        RECT 68.375 176.215 68.545 176.385 ;
        RECT 68.835 176.215 69.005 176.385 ;
        RECT 69.295 176.215 69.465 176.385 ;
        RECT 69.755 176.215 69.925 176.385 ;
        RECT 70.215 176.215 70.385 176.385 ;
        RECT 70.675 176.215 70.845 176.385 ;
        RECT 71.135 176.215 71.305 176.385 ;
        RECT 71.595 176.215 71.765 176.385 ;
        RECT 72.055 176.215 72.225 176.385 ;
        RECT 72.515 176.215 72.685 176.385 ;
        RECT 72.975 176.215 73.145 176.385 ;
        RECT 73.435 176.215 73.605 176.385 ;
        RECT 73.895 176.215 74.065 176.385 ;
        RECT 74.355 176.215 74.525 176.385 ;
        RECT 74.815 176.215 74.985 176.385 ;
        RECT 75.275 176.215 75.445 176.385 ;
        RECT 75.735 176.215 75.905 176.385 ;
        RECT 76.195 176.215 76.365 176.385 ;
        RECT 76.655 176.215 76.825 176.385 ;
        RECT 77.115 176.215 77.285 176.385 ;
        RECT 77.575 176.215 77.745 176.385 ;
        RECT 78.035 176.215 78.205 176.385 ;
        RECT 78.495 176.215 78.665 176.385 ;
        RECT 78.955 176.215 79.125 176.385 ;
        RECT 79.415 176.215 79.585 176.385 ;
        RECT 79.875 176.215 80.045 176.385 ;
        RECT 80.335 176.215 80.505 176.385 ;
        RECT 80.795 176.215 80.965 176.385 ;
        RECT 81.255 176.215 81.425 176.385 ;
        RECT 81.715 176.215 81.885 176.385 ;
        RECT 82.175 176.215 82.345 176.385 ;
        RECT 82.635 176.215 82.805 176.385 ;
        RECT 83.095 176.215 83.265 176.385 ;
        RECT 83.555 176.215 83.725 176.385 ;
        RECT 84.015 176.215 84.185 176.385 ;
        RECT 84.475 176.215 84.645 176.385 ;
        RECT 84.935 176.215 85.105 176.385 ;
        RECT 85.395 176.215 85.565 176.385 ;
        RECT 85.855 176.215 86.025 176.385 ;
        RECT 86.315 176.215 86.485 176.385 ;
        RECT 86.775 176.215 86.945 176.385 ;
        RECT 87.235 176.215 87.405 176.385 ;
        RECT 87.695 176.215 87.865 176.385 ;
        RECT 88.155 176.215 88.325 176.385 ;
        RECT 88.615 176.215 88.785 176.385 ;
        RECT 89.075 176.215 89.245 176.385 ;
        RECT 89.535 176.215 89.705 176.385 ;
        RECT 89.995 176.215 90.165 176.385 ;
        RECT 90.455 176.215 90.625 176.385 ;
        RECT 90.915 176.215 91.085 176.385 ;
        RECT 91.375 176.215 91.545 176.385 ;
        RECT 91.835 176.215 92.005 176.385 ;
        RECT 92.295 176.215 92.465 176.385 ;
        RECT 92.755 176.215 92.925 176.385 ;
        RECT 93.215 176.215 93.385 176.385 ;
        RECT 93.675 176.215 93.845 176.385 ;
        RECT 94.135 176.215 94.305 176.385 ;
        RECT 94.595 176.215 94.765 176.385 ;
        RECT 95.055 176.215 95.225 176.385 ;
        RECT 95.515 176.215 95.685 176.385 ;
        RECT 95.975 176.215 96.145 176.385 ;
        RECT 96.435 176.215 96.605 176.385 ;
        RECT 96.895 176.215 97.065 176.385 ;
        RECT 97.355 176.215 97.525 176.385 ;
        RECT 97.815 176.215 97.985 176.385 ;
        RECT 98.275 176.215 98.445 176.385 ;
        RECT 98.735 176.215 98.905 176.385 ;
        RECT 99.195 176.215 99.365 176.385 ;
        RECT 99.655 176.215 99.825 176.385 ;
        RECT 100.115 176.215 100.285 176.385 ;
        RECT 100.575 176.215 100.745 176.385 ;
        RECT 101.035 176.215 101.205 176.385 ;
        RECT 101.495 176.215 101.665 176.385 ;
        RECT 101.955 176.215 102.125 176.385 ;
        RECT 102.415 176.215 102.585 176.385 ;
        RECT 102.875 176.215 103.045 176.385 ;
        RECT 103.335 176.215 103.505 176.385 ;
        RECT 103.795 176.215 103.965 176.385 ;
        RECT 104.255 176.215 104.425 176.385 ;
        RECT 104.715 176.215 104.885 176.385 ;
        RECT 105.175 176.215 105.345 176.385 ;
        RECT 105.635 176.215 105.805 176.385 ;
        RECT 106.095 176.215 106.265 176.385 ;
        RECT 106.555 176.215 106.725 176.385 ;
        RECT 107.015 176.215 107.185 176.385 ;
        RECT 107.475 176.215 107.645 176.385 ;
        RECT 107.935 176.215 108.105 176.385 ;
        RECT 108.395 176.215 108.565 176.385 ;
        RECT 108.855 176.215 109.025 176.385 ;
        RECT 109.315 176.215 109.485 176.385 ;
        RECT 109.775 176.215 109.945 176.385 ;
        RECT 110.235 176.215 110.405 176.385 ;
        RECT 110.695 176.215 110.865 176.385 ;
        RECT 111.155 176.215 111.325 176.385 ;
        RECT 111.615 176.215 111.785 176.385 ;
        RECT 112.075 176.215 112.245 176.385 ;
        RECT 112.535 176.215 112.705 176.385 ;
        RECT 112.995 176.215 113.165 176.385 ;
        RECT 113.455 176.215 113.625 176.385 ;
        RECT 113.915 176.215 114.085 176.385 ;
        RECT 114.375 176.215 114.545 176.385 ;
        RECT 114.835 176.215 115.005 176.385 ;
        RECT 115.295 176.215 115.465 176.385 ;
        RECT 115.755 176.215 115.925 176.385 ;
        RECT 116.215 176.215 116.385 176.385 ;
        RECT 116.675 176.215 116.845 176.385 ;
        RECT 117.135 176.215 117.305 176.385 ;
        RECT 117.595 176.215 117.765 176.385 ;
        RECT 118.055 176.215 118.225 176.385 ;
        RECT 118.515 176.215 118.685 176.385 ;
        RECT 118.975 176.215 119.145 176.385 ;
        RECT 119.435 176.215 119.605 176.385 ;
        RECT 119.895 176.215 120.065 176.385 ;
        RECT 120.355 176.215 120.525 176.385 ;
        RECT 120.815 176.215 120.985 176.385 ;
        RECT 121.275 176.215 121.445 176.385 ;
        RECT 121.735 176.215 121.905 176.385 ;
        RECT 122.195 176.215 122.365 176.385 ;
        RECT 122.655 176.215 122.825 176.385 ;
        RECT 123.115 176.215 123.285 176.385 ;
        RECT 123.575 176.215 123.745 176.385 ;
        RECT 124.035 176.215 124.205 176.385 ;
        RECT 124.495 176.215 124.665 176.385 ;
        RECT 124.955 176.215 125.125 176.385 ;
        RECT 125.415 176.215 125.585 176.385 ;
        RECT 125.875 176.215 126.045 176.385 ;
        RECT 126.335 176.215 126.505 176.385 ;
        RECT 126.795 176.215 126.965 176.385 ;
        RECT 127.255 176.215 127.425 176.385 ;
        RECT 127.715 176.215 127.885 176.385 ;
        RECT 128.175 176.215 128.345 176.385 ;
        RECT 128.635 176.215 128.805 176.385 ;
        RECT 129.095 176.215 129.265 176.385 ;
        RECT 129.555 176.215 129.725 176.385 ;
        RECT 130.015 176.215 130.185 176.385 ;
        RECT 130.475 176.215 130.645 176.385 ;
        RECT 130.935 176.215 131.105 176.385 ;
        RECT 57.335 173.495 57.505 173.665 ;
        RECT 57.795 173.495 57.965 173.665 ;
        RECT 58.255 173.495 58.425 173.665 ;
        RECT 58.715 173.495 58.885 173.665 ;
        RECT 59.175 173.495 59.345 173.665 ;
        RECT 59.635 173.495 59.805 173.665 ;
        RECT 60.095 173.495 60.265 173.665 ;
        RECT 60.555 173.495 60.725 173.665 ;
        RECT 61.015 173.495 61.185 173.665 ;
        RECT 61.475 173.495 61.645 173.665 ;
        RECT 61.935 173.495 62.105 173.665 ;
        RECT 62.395 173.495 62.565 173.665 ;
        RECT 62.855 173.495 63.025 173.665 ;
        RECT 63.315 173.495 63.485 173.665 ;
        RECT 63.775 173.495 63.945 173.665 ;
        RECT 64.235 173.495 64.405 173.665 ;
        RECT 64.695 173.495 64.865 173.665 ;
        RECT 65.155 173.495 65.325 173.665 ;
        RECT 65.615 173.495 65.785 173.665 ;
        RECT 66.075 173.495 66.245 173.665 ;
        RECT 66.535 173.495 66.705 173.665 ;
        RECT 66.995 173.495 67.165 173.665 ;
        RECT 67.455 173.495 67.625 173.665 ;
        RECT 67.915 173.495 68.085 173.665 ;
        RECT 68.375 173.495 68.545 173.665 ;
        RECT 68.835 173.495 69.005 173.665 ;
        RECT 69.295 173.495 69.465 173.665 ;
        RECT 69.755 173.495 69.925 173.665 ;
        RECT 70.215 173.495 70.385 173.665 ;
        RECT 70.675 173.495 70.845 173.665 ;
        RECT 71.135 173.495 71.305 173.665 ;
        RECT 71.595 173.495 71.765 173.665 ;
        RECT 72.055 173.495 72.225 173.665 ;
        RECT 72.515 173.495 72.685 173.665 ;
        RECT 72.975 173.495 73.145 173.665 ;
        RECT 73.435 173.495 73.605 173.665 ;
        RECT 73.895 173.495 74.065 173.665 ;
        RECT 74.355 173.495 74.525 173.665 ;
        RECT 74.815 173.495 74.985 173.665 ;
        RECT 75.275 173.495 75.445 173.665 ;
        RECT 75.735 173.495 75.905 173.665 ;
        RECT 76.195 173.495 76.365 173.665 ;
        RECT 76.655 173.495 76.825 173.665 ;
        RECT 77.115 173.495 77.285 173.665 ;
        RECT 77.575 173.495 77.745 173.665 ;
        RECT 78.035 173.495 78.205 173.665 ;
        RECT 78.495 173.495 78.665 173.665 ;
        RECT 78.955 173.495 79.125 173.665 ;
        RECT 79.415 173.495 79.585 173.665 ;
        RECT 79.875 173.495 80.045 173.665 ;
        RECT 80.335 173.495 80.505 173.665 ;
        RECT 80.795 173.495 80.965 173.665 ;
        RECT 81.255 173.495 81.425 173.665 ;
        RECT 81.715 173.495 81.885 173.665 ;
        RECT 82.175 173.495 82.345 173.665 ;
        RECT 82.635 173.495 82.805 173.665 ;
        RECT 83.095 173.495 83.265 173.665 ;
        RECT 83.555 173.495 83.725 173.665 ;
        RECT 84.015 173.495 84.185 173.665 ;
        RECT 84.475 173.495 84.645 173.665 ;
        RECT 84.935 173.495 85.105 173.665 ;
        RECT 85.395 173.495 85.565 173.665 ;
        RECT 85.855 173.495 86.025 173.665 ;
        RECT 86.315 173.495 86.485 173.665 ;
        RECT 86.775 173.495 86.945 173.665 ;
        RECT 87.235 173.495 87.405 173.665 ;
        RECT 87.695 173.495 87.865 173.665 ;
        RECT 88.155 173.495 88.325 173.665 ;
        RECT 88.615 173.495 88.785 173.665 ;
        RECT 89.075 173.495 89.245 173.665 ;
        RECT 89.535 173.495 89.705 173.665 ;
        RECT 89.995 173.495 90.165 173.665 ;
        RECT 90.455 173.495 90.625 173.665 ;
        RECT 90.915 173.495 91.085 173.665 ;
        RECT 91.375 173.495 91.545 173.665 ;
        RECT 91.835 173.495 92.005 173.665 ;
        RECT 92.295 173.495 92.465 173.665 ;
        RECT 92.755 173.495 92.925 173.665 ;
        RECT 93.215 173.495 93.385 173.665 ;
        RECT 93.675 173.495 93.845 173.665 ;
        RECT 94.135 173.495 94.305 173.665 ;
        RECT 94.595 173.495 94.765 173.665 ;
        RECT 95.055 173.495 95.225 173.665 ;
        RECT 95.515 173.495 95.685 173.665 ;
        RECT 95.975 173.495 96.145 173.665 ;
        RECT 96.435 173.495 96.605 173.665 ;
        RECT 96.895 173.495 97.065 173.665 ;
        RECT 97.355 173.495 97.525 173.665 ;
        RECT 97.815 173.495 97.985 173.665 ;
        RECT 98.275 173.495 98.445 173.665 ;
        RECT 98.735 173.495 98.905 173.665 ;
        RECT 99.195 173.495 99.365 173.665 ;
        RECT 99.655 173.495 99.825 173.665 ;
        RECT 100.115 173.495 100.285 173.665 ;
        RECT 100.575 173.495 100.745 173.665 ;
        RECT 101.035 173.495 101.205 173.665 ;
        RECT 101.495 173.495 101.665 173.665 ;
        RECT 101.955 173.495 102.125 173.665 ;
        RECT 102.415 173.495 102.585 173.665 ;
        RECT 102.875 173.495 103.045 173.665 ;
        RECT 103.335 173.495 103.505 173.665 ;
        RECT 103.795 173.495 103.965 173.665 ;
        RECT 104.255 173.495 104.425 173.665 ;
        RECT 104.715 173.495 104.885 173.665 ;
        RECT 105.175 173.495 105.345 173.665 ;
        RECT 105.635 173.495 105.805 173.665 ;
        RECT 106.095 173.495 106.265 173.665 ;
        RECT 106.555 173.495 106.725 173.665 ;
        RECT 107.015 173.495 107.185 173.665 ;
        RECT 107.475 173.495 107.645 173.665 ;
        RECT 107.935 173.495 108.105 173.665 ;
        RECT 108.395 173.495 108.565 173.665 ;
        RECT 108.855 173.495 109.025 173.665 ;
        RECT 109.315 173.495 109.485 173.665 ;
        RECT 109.775 173.495 109.945 173.665 ;
        RECT 110.235 173.495 110.405 173.665 ;
        RECT 110.695 173.495 110.865 173.665 ;
        RECT 111.155 173.495 111.325 173.665 ;
        RECT 111.615 173.495 111.785 173.665 ;
        RECT 112.075 173.495 112.245 173.665 ;
        RECT 112.535 173.495 112.705 173.665 ;
        RECT 112.995 173.495 113.165 173.665 ;
        RECT 113.455 173.495 113.625 173.665 ;
        RECT 113.915 173.495 114.085 173.665 ;
        RECT 114.375 173.495 114.545 173.665 ;
        RECT 114.835 173.495 115.005 173.665 ;
        RECT 115.295 173.495 115.465 173.665 ;
        RECT 115.755 173.495 115.925 173.665 ;
        RECT 116.215 173.495 116.385 173.665 ;
        RECT 116.675 173.495 116.845 173.665 ;
        RECT 117.135 173.495 117.305 173.665 ;
        RECT 117.595 173.495 117.765 173.665 ;
        RECT 118.055 173.495 118.225 173.665 ;
        RECT 118.515 173.495 118.685 173.665 ;
        RECT 118.975 173.495 119.145 173.665 ;
        RECT 119.435 173.495 119.605 173.665 ;
        RECT 119.895 173.495 120.065 173.665 ;
        RECT 120.355 173.495 120.525 173.665 ;
        RECT 120.815 173.495 120.985 173.665 ;
        RECT 121.275 173.495 121.445 173.665 ;
        RECT 121.735 173.495 121.905 173.665 ;
        RECT 122.195 173.495 122.365 173.665 ;
        RECT 122.655 173.495 122.825 173.665 ;
        RECT 123.115 173.495 123.285 173.665 ;
        RECT 123.575 173.495 123.745 173.665 ;
        RECT 124.035 173.495 124.205 173.665 ;
        RECT 124.495 173.495 124.665 173.665 ;
        RECT 124.955 173.495 125.125 173.665 ;
        RECT 125.415 173.495 125.585 173.665 ;
        RECT 125.875 173.495 126.045 173.665 ;
        RECT 126.335 173.495 126.505 173.665 ;
        RECT 126.795 173.495 126.965 173.665 ;
        RECT 127.255 173.495 127.425 173.665 ;
        RECT 127.715 173.495 127.885 173.665 ;
        RECT 128.175 173.495 128.345 173.665 ;
        RECT 128.635 173.495 128.805 173.665 ;
        RECT 129.095 173.495 129.265 173.665 ;
        RECT 129.555 173.495 129.725 173.665 ;
        RECT 130.015 173.495 130.185 173.665 ;
        RECT 130.475 173.495 130.645 173.665 ;
        RECT 130.935 173.495 131.105 173.665 ;
        RECT 57.335 170.775 57.505 170.945 ;
        RECT 57.795 170.775 57.965 170.945 ;
        RECT 58.255 170.775 58.425 170.945 ;
        RECT 58.715 170.775 58.885 170.945 ;
        RECT 59.175 170.775 59.345 170.945 ;
        RECT 59.635 170.775 59.805 170.945 ;
        RECT 60.095 170.775 60.265 170.945 ;
        RECT 60.555 170.775 60.725 170.945 ;
        RECT 61.015 170.775 61.185 170.945 ;
        RECT 61.475 170.775 61.645 170.945 ;
        RECT 61.935 170.775 62.105 170.945 ;
        RECT 62.395 170.775 62.565 170.945 ;
        RECT 62.855 170.775 63.025 170.945 ;
        RECT 63.315 170.775 63.485 170.945 ;
        RECT 63.775 170.775 63.945 170.945 ;
        RECT 64.235 170.775 64.405 170.945 ;
        RECT 64.695 170.775 64.865 170.945 ;
        RECT 65.155 170.775 65.325 170.945 ;
        RECT 65.615 170.775 65.785 170.945 ;
        RECT 66.075 170.775 66.245 170.945 ;
        RECT 66.535 170.775 66.705 170.945 ;
        RECT 66.995 170.775 67.165 170.945 ;
        RECT 67.455 170.775 67.625 170.945 ;
        RECT 67.915 170.775 68.085 170.945 ;
        RECT 68.375 170.775 68.545 170.945 ;
        RECT 68.835 170.775 69.005 170.945 ;
        RECT 69.295 170.775 69.465 170.945 ;
        RECT 69.755 170.775 69.925 170.945 ;
        RECT 70.215 170.775 70.385 170.945 ;
        RECT 70.675 170.775 70.845 170.945 ;
        RECT 71.135 170.775 71.305 170.945 ;
        RECT 71.595 170.775 71.765 170.945 ;
        RECT 72.055 170.775 72.225 170.945 ;
        RECT 72.515 170.775 72.685 170.945 ;
        RECT 72.975 170.775 73.145 170.945 ;
        RECT 73.435 170.775 73.605 170.945 ;
        RECT 73.895 170.775 74.065 170.945 ;
        RECT 74.355 170.775 74.525 170.945 ;
        RECT 74.815 170.775 74.985 170.945 ;
        RECT 75.275 170.775 75.445 170.945 ;
        RECT 75.735 170.775 75.905 170.945 ;
        RECT 76.195 170.775 76.365 170.945 ;
        RECT 76.655 170.775 76.825 170.945 ;
        RECT 77.115 170.775 77.285 170.945 ;
        RECT 77.575 170.775 77.745 170.945 ;
        RECT 78.035 170.775 78.205 170.945 ;
        RECT 78.495 170.775 78.665 170.945 ;
        RECT 78.955 170.775 79.125 170.945 ;
        RECT 79.415 170.775 79.585 170.945 ;
        RECT 79.875 170.775 80.045 170.945 ;
        RECT 80.335 170.775 80.505 170.945 ;
        RECT 80.795 170.775 80.965 170.945 ;
        RECT 81.255 170.775 81.425 170.945 ;
        RECT 81.715 170.775 81.885 170.945 ;
        RECT 82.175 170.775 82.345 170.945 ;
        RECT 82.635 170.775 82.805 170.945 ;
        RECT 83.095 170.775 83.265 170.945 ;
        RECT 83.555 170.775 83.725 170.945 ;
        RECT 84.015 170.775 84.185 170.945 ;
        RECT 84.475 170.775 84.645 170.945 ;
        RECT 84.935 170.775 85.105 170.945 ;
        RECT 85.395 170.775 85.565 170.945 ;
        RECT 85.855 170.775 86.025 170.945 ;
        RECT 86.315 170.775 86.485 170.945 ;
        RECT 86.775 170.775 86.945 170.945 ;
        RECT 87.235 170.775 87.405 170.945 ;
        RECT 87.695 170.775 87.865 170.945 ;
        RECT 88.155 170.775 88.325 170.945 ;
        RECT 88.615 170.775 88.785 170.945 ;
        RECT 89.075 170.775 89.245 170.945 ;
        RECT 89.535 170.775 89.705 170.945 ;
        RECT 89.995 170.775 90.165 170.945 ;
        RECT 90.455 170.775 90.625 170.945 ;
        RECT 90.915 170.775 91.085 170.945 ;
        RECT 91.375 170.775 91.545 170.945 ;
        RECT 91.835 170.775 92.005 170.945 ;
        RECT 92.295 170.775 92.465 170.945 ;
        RECT 92.755 170.775 92.925 170.945 ;
        RECT 93.215 170.775 93.385 170.945 ;
        RECT 93.675 170.775 93.845 170.945 ;
        RECT 94.135 170.775 94.305 170.945 ;
        RECT 94.595 170.775 94.765 170.945 ;
        RECT 95.055 170.775 95.225 170.945 ;
        RECT 95.515 170.775 95.685 170.945 ;
        RECT 95.975 170.775 96.145 170.945 ;
        RECT 96.435 170.775 96.605 170.945 ;
        RECT 96.895 170.775 97.065 170.945 ;
        RECT 97.355 170.775 97.525 170.945 ;
        RECT 97.815 170.775 97.985 170.945 ;
        RECT 98.275 170.775 98.445 170.945 ;
        RECT 98.735 170.775 98.905 170.945 ;
        RECT 99.195 170.775 99.365 170.945 ;
        RECT 99.655 170.775 99.825 170.945 ;
        RECT 100.115 170.775 100.285 170.945 ;
        RECT 100.575 170.775 100.745 170.945 ;
        RECT 101.035 170.775 101.205 170.945 ;
        RECT 101.495 170.775 101.665 170.945 ;
        RECT 101.955 170.775 102.125 170.945 ;
        RECT 102.415 170.775 102.585 170.945 ;
        RECT 102.875 170.775 103.045 170.945 ;
        RECT 103.335 170.775 103.505 170.945 ;
        RECT 103.795 170.775 103.965 170.945 ;
        RECT 104.255 170.775 104.425 170.945 ;
        RECT 104.715 170.775 104.885 170.945 ;
        RECT 105.175 170.775 105.345 170.945 ;
        RECT 105.635 170.775 105.805 170.945 ;
        RECT 106.095 170.775 106.265 170.945 ;
        RECT 106.555 170.775 106.725 170.945 ;
        RECT 107.015 170.775 107.185 170.945 ;
        RECT 107.475 170.775 107.645 170.945 ;
        RECT 107.935 170.775 108.105 170.945 ;
        RECT 108.395 170.775 108.565 170.945 ;
        RECT 108.855 170.775 109.025 170.945 ;
        RECT 109.315 170.775 109.485 170.945 ;
        RECT 109.775 170.775 109.945 170.945 ;
        RECT 110.235 170.775 110.405 170.945 ;
        RECT 110.695 170.775 110.865 170.945 ;
        RECT 111.155 170.775 111.325 170.945 ;
        RECT 111.615 170.775 111.785 170.945 ;
        RECT 112.075 170.775 112.245 170.945 ;
        RECT 112.535 170.775 112.705 170.945 ;
        RECT 112.995 170.775 113.165 170.945 ;
        RECT 113.455 170.775 113.625 170.945 ;
        RECT 113.915 170.775 114.085 170.945 ;
        RECT 114.375 170.775 114.545 170.945 ;
        RECT 114.835 170.775 115.005 170.945 ;
        RECT 115.295 170.775 115.465 170.945 ;
        RECT 115.755 170.775 115.925 170.945 ;
        RECT 116.215 170.775 116.385 170.945 ;
        RECT 116.675 170.775 116.845 170.945 ;
        RECT 117.135 170.775 117.305 170.945 ;
        RECT 117.595 170.775 117.765 170.945 ;
        RECT 118.055 170.775 118.225 170.945 ;
        RECT 118.515 170.775 118.685 170.945 ;
        RECT 118.975 170.775 119.145 170.945 ;
        RECT 119.435 170.775 119.605 170.945 ;
        RECT 119.895 170.775 120.065 170.945 ;
        RECT 120.355 170.775 120.525 170.945 ;
        RECT 120.815 170.775 120.985 170.945 ;
        RECT 121.275 170.775 121.445 170.945 ;
        RECT 121.735 170.775 121.905 170.945 ;
        RECT 122.195 170.775 122.365 170.945 ;
        RECT 122.655 170.775 122.825 170.945 ;
        RECT 123.115 170.775 123.285 170.945 ;
        RECT 123.575 170.775 123.745 170.945 ;
        RECT 124.035 170.775 124.205 170.945 ;
        RECT 124.495 170.775 124.665 170.945 ;
        RECT 124.955 170.775 125.125 170.945 ;
        RECT 125.415 170.775 125.585 170.945 ;
        RECT 125.875 170.775 126.045 170.945 ;
        RECT 126.335 170.775 126.505 170.945 ;
        RECT 126.795 170.775 126.965 170.945 ;
        RECT 127.255 170.775 127.425 170.945 ;
        RECT 127.715 170.775 127.885 170.945 ;
        RECT 128.175 170.775 128.345 170.945 ;
        RECT 128.635 170.775 128.805 170.945 ;
        RECT 129.095 170.775 129.265 170.945 ;
        RECT 129.555 170.775 129.725 170.945 ;
        RECT 130.015 170.775 130.185 170.945 ;
        RECT 130.475 170.775 130.645 170.945 ;
        RECT 130.935 170.775 131.105 170.945 ;
        RECT 57.335 168.055 57.505 168.225 ;
        RECT 57.795 168.055 57.965 168.225 ;
        RECT 58.255 168.055 58.425 168.225 ;
        RECT 58.715 168.055 58.885 168.225 ;
        RECT 59.175 168.055 59.345 168.225 ;
        RECT 59.635 168.055 59.805 168.225 ;
        RECT 60.095 168.055 60.265 168.225 ;
        RECT 60.555 168.055 60.725 168.225 ;
        RECT 61.015 168.055 61.185 168.225 ;
        RECT 61.475 168.055 61.645 168.225 ;
        RECT 61.935 168.055 62.105 168.225 ;
        RECT 62.395 168.055 62.565 168.225 ;
        RECT 62.855 168.055 63.025 168.225 ;
        RECT 63.315 168.055 63.485 168.225 ;
        RECT 63.775 168.055 63.945 168.225 ;
        RECT 64.235 168.055 64.405 168.225 ;
        RECT 64.695 168.055 64.865 168.225 ;
        RECT 65.155 168.055 65.325 168.225 ;
        RECT 65.615 168.055 65.785 168.225 ;
        RECT 66.075 168.055 66.245 168.225 ;
        RECT 66.535 168.055 66.705 168.225 ;
        RECT 66.995 168.055 67.165 168.225 ;
        RECT 67.455 168.055 67.625 168.225 ;
        RECT 67.915 168.055 68.085 168.225 ;
        RECT 68.375 168.055 68.545 168.225 ;
        RECT 68.835 168.055 69.005 168.225 ;
        RECT 69.295 168.055 69.465 168.225 ;
        RECT 69.755 168.055 69.925 168.225 ;
        RECT 70.215 168.055 70.385 168.225 ;
        RECT 70.675 168.055 70.845 168.225 ;
        RECT 71.135 168.055 71.305 168.225 ;
        RECT 71.595 168.055 71.765 168.225 ;
        RECT 72.055 168.055 72.225 168.225 ;
        RECT 72.515 168.055 72.685 168.225 ;
        RECT 72.975 168.055 73.145 168.225 ;
        RECT 73.435 168.055 73.605 168.225 ;
        RECT 73.895 168.055 74.065 168.225 ;
        RECT 74.355 168.055 74.525 168.225 ;
        RECT 74.815 168.055 74.985 168.225 ;
        RECT 75.275 168.055 75.445 168.225 ;
        RECT 75.735 168.055 75.905 168.225 ;
        RECT 76.195 168.055 76.365 168.225 ;
        RECT 76.655 168.055 76.825 168.225 ;
        RECT 77.115 168.055 77.285 168.225 ;
        RECT 77.575 168.055 77.745 168.225 ;
        RECT 78.035 168.055 78.205 168.225 ;
        RECT 78.495 168.055 78.665 168.225 ;
        RECT 78.955 168.055 79.125 168.225 ;
        RECT 79.415 168.055 79.585 168.225 ;
        RECT 79.875 168.055 80.045 168.225 ;
        RECT 80.335 168.055 80.505 168.225 ;
        RECT 80.795 168.055 80.965 168.225 ;
        RECT 81.255 168.055 81.425 168.225 ;
        RECT 81.715 168.055 81.885 168.225 ;
        RECT 82.175 168.055 82.345 168.225 ;
        RECT 82.635 168.055 82.805 168.225 ;
        RECT 83.095 168.055 83.265 168.225 ;
        RECT 83.555 168.055 83.725 168.225 ;
        RECT 84.015 168.055 84.185 168.225 ;
        RECT 84.475 168.055 84.645 168.225 ;
        RECT 84.935 168.055 85.105 168.225 ;
        RECT 85.395 168.055 85.565 168.225 ;
        RECT 85.855 168.055 86.025 168.225 ;
        RECT 86.315 168.055 86.485 168.225 ;
        RECT 86.775 168.055 86.945 168.225 ;
        RECT 87.235 168.055 87.405 168.225 ;
        RECT 87.695 168.055 87.865 168.225 ;
        RECT 88.155 168.055 88.325 168.225 ;
        RECT 88.615 168.055 88.785 168.225 ;
        RECT 89.075 168.055 89.245 168.225 ;
        RECT 89.535 168.055 89.705 168.225 ;
        RECT 89.995 168.055 90.165 168.225 ;
        RECT 90.455 168.055 90.625 168.225 ;
        RECT 90.915 168.055 91.085 168.225 ;
        RECT 91.375 168.055 91.545 168.225 ;
        RECT 91.835 168.055 92.005 168.225 ;
        RECT 92.295 168.055 92.465 168.225 ;
        RECT 92.755 168.055 92.925 168.225 ;
        RECT 93.215 168.055 93.385 168.225 ;
        RECT 93.675 168.055 93.845 168.225 ;
        RECT 94.135 168.055 94.305 168.225 ;
        RECT 94.595 168.055 94.765 168.225 ;
        RECT 95.055 168.055 95.225 168.225 ;
        RECT 95.515 168.055 95.685 168.225 ;
        RECT 95.975 168.055 96.145 168.225 ;
        RECT 96.435 168.055 96.605 168.225 ;
        RECT 96.895 168.055 97.065 168.225 ;
        RECT 97.355 168.055 97.525 168.225 ;
        RECT 97.815 168.055 97.985 168.225 ;
        RECT 98.275 168.055 98.445 168.225 ;
        RECT 98.735 168.055 98.905 168.225 ;
        RECT 99.195 168.055 99.365 168.225 ;
        RECT 99.655 168.055 99.825 168.225 ;
        RECT 100.115 168.055 100.285 168.225 ;
        RECT 100.575 168.055 100.745 168.225 ;
        RECT 101.035 168.055 101.205 168.225 ;
        RECT 101.495 168.055 101.665 168.225 ;
        RECT 101.955 168.055 102.125 168.225 ;
        RECT 102.415 168.055 102.585 168.225 ;
        RECT 102.875 168.055 103.045 168.225 ;
        RECT 103.335 168.055 103.505 168.225 ;
        RECT 103.795 168.055 103.965 168.225 ;
        RECT 104.255 168.055 104.425 168.225 ;
        RECT 104.715 168.055 104.885 168.225 ;
        RECT 105.175 168.055 105.345 168.225 ;
        RECT 105.635 168.055 105.805 168.225 ;
        RECT 106.095 168.055 106.265 168.225 ;
        RECT 106.555 168.055 106.725 168.225 ;
        RECT 107.015 168.055 107.185 168.225 ;
        RECT 107.475 168.055 107.645 168.225 ;
        RECT 107.935 168.055 108.105 168.225 ;
        RECT 108.395 168.055 108.565 168.225 ;
        RECT 108.855 168.055 109.025 168.225 ;
        RECT 109.315 168.055 109.485 168.225 ;
        RECT 109.775 168.055 109.945 168.225 ;
        RECT 110.235 168.055 110.405 168.225 ;
        RECT 110.695 168.055 110.865 168.225 ;
        RECT 111.155 168.055 111.325 168.225 ;
        RECT 111.615 168.055 111.785 168.225 ;
        RECT 112.075 168.055 112.245 168.225 ;
        RECT 112.535 168.055 112.705 168.225 ;
        RECT 112.995 168.055 113.165 168.225 ;
        RECT 113.455 168.055 113.625 168.225 ;
        RECT 113.915 168.055 114.085 168.225 ;
        RECT 114.375 168.055 114.545 168.225 ;
        RECT 114.835 168.055 115.005 168.225 ;
        RECT 115.295 168.055 115.465 168.225 ;
        RECT 115.755 168.055 115.925 168.225 ;
        RECT 116.215 168.055 116.385 168.225 ;
        RECT 116.675 168.055 116.845 168.225 ;
        RECT 117.135 168.055 117.305 168.225 ;
        RECT 117.595 168.055 117.765 168.225 ;
        RECT 118.055 168.055 118.225 168.225 ;
        RECT 118.515 168.055 118.685 168.225 ;
        RECT 118.975 168.055 119.145 168.225 ;
        RECT 119.435 168.055 119.605 168.225 ;
        RECT 119.895 168.055 120.065 168.225 ;
        RECT 120.355 168.055 120.525 168.225 ;
        RECT 120.815 168.055 120.985 168.225 ;
        RECT 121.275 168.055 121.445 168.225 ;
        RECT 121.735 168.055 121.905 168.225 ;
        RECT 122.195 168.055 122.365 168.225 ;
        RECT 122.655 168.055 122.825 168.225 ;
        RECT 123.115 168.055 123.285 168.225 ;
        RECT 123.575 168.055 123.745 168.225 ;
        RECT 124.035 168.055 124.205 168.225 ;
        RECT 124.495 168.055 124.665 168.225 ;
        RECT 124.955 168.055 125.125 168.225 ;
        RECT 125.415 168.055 125.585 168.225 ;
        RECT 125.875 168.055 126.045 168.225 ;
        RECT 126.335 168.055 126.505 168.225 ;
        RECT 126.795 168.055 126.965 168.225 ;
        RECT 127.255 168.055 127.425 168.225 ;
        RECT 127.715 168.055 127.885 168.225 ;
        RECT 128.175 168.055 128.345 168.225 ;
        RECT 128.635 168.055 128.805 168.225 ;
        RECT 129.095 168.055 129.265 168.225 ;
        RECT 129.555 168.055 129.725 168.225 ;
        RECT 130.015 168.055 130.185 168.225 ;
        RECT 130.475 168.055 130.645 168.225 ;
        RECT 130.935 168.055 131.105 168.225 ;
        RECT 57.335 165.335 57.505 165.505 ;
        RECT 57.795 165.335 57.965 165.505 ;
        RECT 58.255 165.335 58.425 165.505 ;
        RECT 58.715 165.335 58.885 165.505 ;
        RECT 59.175 165.335 59.345 165.505 ;
        RECT 59.635 165.335 59.805 165.505 ;
        RECT 60.095 165.335 60.265 165.505 ;
        RECT 60.555 165.335 60.725 165.505 ;
        RECT 61.015 165.335 61.185 165.505 ;
        RECT 61.475 165.335 61.645 165.505 ;
        RECT 61.935 165.335 62.105 165.505 ;
        RECT 62.395 165.335 62.565 165.505 ;
        RECT 62.855 165.335 63.025 165.505 ;
        RECT 63.315 165.335 63.485 165.505 ;
        RECT 63.775 165.335 63.945 165.505 ;
        RECT 64.235 165.335 64.405 165.505 ;
        RECT 64.695 165.335 64.865 165.505 ;
        RECT 65.155 165.335 65.325 165.505 ;
        RECT 65.615 165.335 65.785 165.505 ;
        RECT 66.075 165.335 66.245 165.505 ;
        RECT 66.535 165.335 66.705 165.505 ;
        RECT 66.995 165.335 67.165 165.505 ;
        RECT 67.455 165.335 67.625 165.505 ;
        RECT 67.915 165.335 68.085 165.505 ;
        RECT 68.375 165.335 68.545 165.505 ;
        RECT 68.835 165.335 69.005 165.505 ;
        RECT 69.295 165.335 69.465 165.505 ;
        RECT 69.755 165.335 69.925 165.505 ;
        RECT 70.215 165.335 70.385 165.505 ;
        RECT 70.675 165.335 70.845 165.505 ;
        RECT 71.135 165.335 71.305 165.505 ;
        RECT 71.595 165.335 71.765 165.505 ;
        RECT 72.055 165.335 72.225 165.505 ;
        RECT 72.515 165.335 72.685 165.505 ;
        RECT 72.975 165.335 73.145 165.505 ;
        RECT 73.435 165.335 73.605 165.505 ;
        RECT 73.895 165.335 74.065 165.505 ;
        RECT 74.355 165.335 74.525 165.505 ;
        RECT 74.815 165.335 74.985 165.505 ;
        RECT 75.275 165.335 75.445 165.505 ;
        RECT 75.735 165.335 75.905 165.505 ;
        RECT 76.195 165.335 76.365 165.505 ;
        RECT 76.655 165.335 76.825 165.505 ;
        RECT 77.115 165.335 77.285 165.505 ;
        RECT 77.575 165.335 77.745 165.505 ;
        RECT 78.035 165.335 78.205 165.505 ;
        RECT 78.495 165.335 78.665 165.505 ;
        RECT 78.955 165.335 79.125 165.505 ;
        RECT 79.415 165.335 79.585 165.505 ;
        RECT 79.875 165.335 80.045 165.505 ;
        RECT 80.335 165.335 80.505 165.505 ;
        RECT 80.795 165.335 80.965 165.505 ;
        RECT 81.255 165.335 81.425 165.505 ;
        RECT 81.715 165.335 81.885 165.505 ;
        RECT 82.175 165.335 82.345 165.505 ;
        RECT 82.635 165.335 82.805 165.505 ;
        RECT 83.095 165.335 83.265 165.505 ;
        RECT 83.555 165.335 83.725 165.505 ;
        RECT 84.015 165.335 84.185 165.505 ;
        RECT 84.475 165.335 84.645 165.505 ;
        RECT 84.935 165.335 85.105 165.505 ;
        RECT 85.395 165.335 85.565 165.505 ;
        RECT 85.855 165.335 86.025 165.505 ;
        RECT 86.315 165.335 86.485 165.505 ;
        RECT 86.775 165.335 86.945 165.505 ;
        RECT 87.235 165.335 87.405 165.505 ;
        RECT 87.695 165.335 87.865 165.505 ;
        RECT 88.155 165.335 88.325 165.505 ;
        RECT 88.615 165.335 88.785 165.505 ;
        RECT 89.075 165.335 89.245 165.505 ;
        RECT 89.535 165.335 89.705 165.505 ;
        RECT 89.995 165.335 90.165 165.505 ;
        RECT 90.455 165.335 90.625 165.505 ;
        RECT 90.915 165.335 91.085 165.505 ;
        RECT 91.375 165.335 91.545 165.505 ;
        RECT 91.835 165.335 92.005 165.505 ;
        RECT 92.295 165.335 92.465 165.505 ;
        RECT 92.755 165.335 92.925 165.505 ;
        RECT 93.215 165.335 93.385 165.505 ;
        RECT 93.675 165.335 93.845 165.505 ;
        RECT 94.135 165.335 94.305 165.505 ;
        RECT 94.595 165.335 94.765 165.505 ;
        RECT 95.055 165.335 95.225 165.505 ;
        RECT 95.515 165.335 95.685 165.505 ;
        RECT 95.975 165.335 96.145 165.505 ;
        RECT 96.435 165.335 96.605 165.505 ;
        RECT 96.895 165.335 97.065 165.505 ;
        RECT 97.355 165.335 97.525 165.505 ;
        RECT 97.815 165.335 97.985 165.505 ;
        RECT 98.275 165.335 98.445 165.505 ;
        RECT 98.735 165.335 98.905 165.505 ;
        RECT 99.195 165.335 99.365 165.505 ;
        RECT 99.655 165.335 99.825 165.505 ;
        RECT 100.115 165.335 100.285 165.505 ;
        RECT 100.575 165.335 100.745 165.505 ;
        RECT 101.035 165.335 101.205 165.505 ;
        RECT 101.495 165.335 101.665 165.505 ;
        RECT 101.955 165.335 102.125 165.505 ;
        RECT 102.415 165.335 102.585 165.505 ;
        RECT 102.875 165.335 103.045 165.505 ;
        RECT 103.335 165.335 103.505 165.505 ;
        RECT 103.795 165.335 103.965 165.505 ;
        RECT 104.255 165.335 104.425 165.505 ;
        RECT 104.715 165.335 104.885 165.505 ;
        RECT 105.175 165.335 105.345 165.505 ;
        RECT 105.635 165.335 105.805 165.505 ;
        RECT 106.095 165.335 106.265 165.505 ;
        RECT 106.555 165.335 106.725 165.505 ;
        RECT 107.015 165.335 107.185 165.505 ;
        RECT 107.475 165.335 107.645 165.505 ;
        RECT 107.935 165.335 108.105 165.505 ;
        RECT 108.395 165.335 108.565 165.505 ;
        RECT 108.855 165.335 109.025 165.505 ;
        RECT 109.315 165.335 109.485 165.505 ;
        RECT 109.775 165.335 109.945 165.505 ;
        RECT 110.235 165.335 110.405 165.505 ;
        RECT 110.695 165.335 110.865 165.505 ;
        RECT 111.155 165.335 111.325 165.505 ;
        RECT 111.615 165.335 111.785 165.505 ;
        RECT 112.075 165.335 112.245 165.505 ;
        RECT 112.535 165.335 112.705 165.505 ;
        RECT 112.995 165.335 113.165 165.505 ;
        RECT 113.455 165.335 113.625 165.505 ;
        RECT 113.915 165.335 114.085 165.505 ;
        RECT 114.375 165.335 114.545 165.505 ;
        RECT 114.835 165.335 115.005 165.505 ;
        RECT 115.295 165.335 115.465 165.505 ;
        RECT 115.755 165.335 115.925 165.505 ;
        RECT 116.215 165.335 116.385 165.505 ;
        RECT 116.675 165.335 116.845 165.505 ;
        RECT 117.135 165.335 117.305 165.505 ;
        RECT 117.595 165.335 117.765 165.505 ;
        RECT 118.055 165.335 118.225 165.505 ;
        RECT 118.515 165.335 118.685 165.505 ;
        RECT 118.975 165.335 119.145 165.505 ;
        RECT 119.435 165.335 119.605 165.505 ;
        RECT 119.895 165.335 120.065 165.505 ;
        RECT 120.355 165.335 120.525 165.505 ;
        RECT 120.815 165.335 120.985 165.505 ;
        RECT 121.275 165.335 121.445 165.505 ;
        RECT 121.735 165.335 121.905 165.505 ;
        RECT 122.195 165.335 122.365 165.505 ;
        RECT 122.655 165.335 122.825 165.505 ;
        RECT 123.115 165.335 123.285 165.505 ;
        RECT 123.575 165.335 123.745 165.505 ;
        RECT 124.035 165.335 124.205 165.505 ;
        RECT 124.495 165.335 124.665 165.505 ;
        RECT 124.955 165.335 125.125 165.505 ;
        RECT 125.415 165.335 125.585 165.505 ;
        RECT 125.875 165.335 126.045 165.505 ;
        RECT 126.335 165.335 126.505 165.505 ;
        RECT 126.795 165.335 126.965 165.505 ;
        RECT 127.255 165.335 127.425 165.505 ;
        RECT 127.715 165.335 127.885 165.505 ;
        RECT 128.175 165.335 128.345 165.505 ;
        RECT 128.635 165.335 128.805 165.505 ;
        RECT 129.095 165.335 129.265 165.505 ;
        RECT 129.555 165.335 129.725 165.505 ;
        RECT 130.015 165.335 130.185 165.505 ;
        RECT 130.475 165.335 130.645 165.505 ;
        RECT 130.935 165.335 131.105 165.505 ;
        RECT 57.335 162.615 57.505 162.785 ;
        RECT 57.795 162.615 57.965 162.785 ;
        RECT 58.255 162.615 58.425 162.785 ;
        RECT 58.715 162.615 58.885 162.785 ;
        RECT 59.175 162.615 59.345 162.785 ;
        RECT 59.635 162.615 59.805 162.785 ;
        RECT 60.095 162.615 60.265 162.785 ;
        RECT 60.555 162.615 60.725 162.785 ;
        RECT 61.015 162.615 61.185 162.785 ;
        RECT 61.475 162.615 61.645 162.785 ;
        RECT 61.935 162.615 62.105 162.785 ;
        RECT 62.395 162.615 62.565 162.785 ;
        RECT 62.855 162.615 63.025 162.785 ;
        RECT 63.315 162.615 63.485 162.785 ;
        RECT 63.775 162.615 63.945 162.785 ;
        RECT 64.235 162.615 64.405 162.785 ;
        RECT 64.695 162.615 64.865 162.785 ;
        RECT 65.155 162.615 65.325 162.785 ;
        RECT 65.615 162.615 65.785 162.785 ;
        RECT 66.075 162.615 66.245 162.785 ;
        RECT 66.535 162.615 66.705 162.785 ;
        RECT 66.995 162.615 67.165 162.785 ;
        RECT 67.455 162.615 67.625 162.785 ;
        RECT 67.915 162.615 68.085 162.785 ;
        RECT 68.375 162.615 68.545 162.785 ;
        RECT 68.835 162.615 69.005 162.785 ;
        RECT 69.295 162.615 69.465 162.785 ;
        RECT 69.755 162.615 69.925 162.785 ;
        RECT 70.215 162.615 70.385 162.785 ;
        RECT 70.675 162.615 70.845 162.785 ;
        RECT 71.135 162.615 71.305 162.785 ;
        RECT 71.595 162.615 71.765 162.785 ;
        RECT 72.055 162.615 72.225 162.785 ;
        RECT 72.515 162.615 72.685 162.785 ;
        RECT 72.975 162.615 73.145 162.785 ;
        RECT 73.435 162.615 73.605 162.785 ;
        RECT 73.895 162.615 74.065 162.785 ;
        RECT 74.355 162.615 74.525 162.785 ;
        RECT 74.815 162.615 74.985 162.785 ;
        RECT 75.275 162.615 75.445 162.785 ;
        RECT 75.735 162.615 75.905 162.785 ;
        RECT 76.195 162.615 76.365 162.785 ;
        RECT 76.655 162.615 76.825 162.785 ;
        RECT 77.115 162.615 77.285 162.785 ;
        RECT 77.575 162.615 77.745 162.785 ;
        RECT 78.035 162.615 78.205 162.785 ;
        RECT 78.495 162.615 78.665 162.785 ;
        RECT 78.955 162.615 79.125 162.785 ;
        RECT 79.415 162.615 79.585 162.785 ;
        RECT 79.875 162.615 80.045 162.785 ;
        RECT 80.335 162.615 80.505 162.785 ;
        RECT 80.795 162.615 80.965 162.785 ;
        RECT 81.255 162.615 81.425 162.785 ;
        RECT 81.715 162.615 81.885 162.785 ;
        RECT 82.175 162.615 82.345 162.785 ;
        RECT 82.635 162.615 82.805 162.785 ;
        RECT 83.095 162.615 83.265 162.785 ;
        RECT 83.555 162.615 83.725 162.785 ;
        RECT 84.015 162.615 84.185 162.785 ;
        RECT 84.475 162.615 84.645 162.785 ;
        RECT 84.935 162.615 85.105 162.785 ;
        RECT 85.395 162.615 85.565 162.785 ;
        RECT 85.855 162.615 86.025 162.785 ;
        RECT 86.315 162.615 86.485 162.785 ;
        RECT 86.775 162.615 86.945 162.785 ;
        RECT 87.235 162.615 87.405 162.785 ;
        RECT 87.695 162.615 87.865 162.785 ;
        RECT 88.155 162.615 88.325 162.785 ;
        RECT 88.615 162.615 88.785 162.785 ;
        RECT 89.075 162.615 89.245 162.785 ;
        RECT 89.535 162.615 89.705 162.785 ;
        RECT 89.995 162.615 90.165 162.785 ;
        RECT 90.455 162.615 90.625 162.785 ;
        RECT 90.915 162.615 91.085 162.785 ;
        RECT 91.375 162.615 91.545 162.785 ;
        RECT 91.835 162.615 92.005 162.785 ;
        RECT 92.295 162.615 92.465 162.785 ;
        RECT 92.755 162.615 92.925 162.785 ;
        RECT 93.215 162.615 93.385 162.785 ;
        RECT 93.675 162.615 93.845 162.785 ;
        RECT 94.135 162.615 94.305 162.785 ;
        RECT 94.595 162.615 94.765 162.785 ;
        RECT 95.055 162.615 95.225 162.785 ;
        RECT 95.515 162.615 95.685 162.785 ;
        RECT 95.975 162.615 96.145 162.785 ;
        RECT 96.435 162.615 96.605 162.785 ;
        RECT 96.895 162.615 97.065 162.785 ;
        RECT 97.355 162.615 97.525 162.785 ;
        RECT 97.815 162.615 97.985 162.785 ;
        RECT 98.275 162.615 98.445 162.785 ;
        RECT 98.735 162.615 98.905 162.785 ;
        RECT 99.195 162.615 99.365 162.785 ;
        RECT 99.655 162.615 99.825 162.785 ;
        RECT 100.115 162.615 100.285 162.785 ;
        RECT 100.575 162.615 100.745 162.785 ;
        RECT 101.035 162.615 101.205 162.785 ;
        RECT 101.495 162.615 101.665 162.785 ;
        RECT 101.955 162.615 102.125 162.785 ;
        RECT 102.415 162.615 102.585 162.785 ;
        RECT 102.875 162.615 103.045 162.785 ;
        RECT 103.335 162.615 103.505 162.785 ;
        RECT 103.795 162.615 103.965 162.785 ;
        RECT 104.255 162.615 104.425 162.785 ;
        RECT 104.715 162.615 104.885 162.785 ;
        RECT 105.175 162.615 105.345 162.785 ;
        RECT 105.635 162.615 105.805 162.785 ;
        RECT 106.095 162.615 106.265 162.785 ;
        RECT 106.555 162.615 106.725 162.785 ;
        RECT 107.015 162.615 107.185 162.785 ;
        RECT 107.475 162.615 107.645 162.785 ;
        RECT 107.935 162.615 108.105 162.785 ;
        RECT 108.395 162.615 108.565 162.785 ;
        RECT 108.855 162.615 109.025 162.785 ;
        RECT 109.315 162.615 109.485 162.785 ;
        RECT 109.775 162.615 109.945 162.785 ;
        RECT 110.235 162.615 110.405 162.785 ;
        RECT 110.695 162.615 110.865 162.785 ;
        RECT 111.155 162.615 111.325 162.785 ;
        RECT 111.615 162.615 111.785 162.785 ;
        RECT 112.075 162.615 112.245 162.785 ;
        RECT 112.535 162.615 112.705 162.785 ;
        RECT 112.995 162.615 113.165 162.785 ;
        RECT 113.455 162.615 113.625 162.785 ;
        RECT 113.915 162.615 114.085 162.785 ;
        RECT 114.375 162.615 114.545 162.785 ;
        RECT 114.835 162.615 115.005 162.785 ;
        RECT 115.295 162.615 115.465 162.785 ;
        RECT 115.755 162.615 115.925 162.785 ;
        RECT 116.215 162.615 116.385 162.785 ;
        RECT 116.675 162.615 116.845 162.785 ;
        RECT 117.135 162.615 117.305 162.785 ;
        RECT 117.595 162.615 117.765 162.785 ;
        RECT 118.055 162.615 118.225 162.785 ;
        RECT 118.515 162.615 118.685 162.785 ;
        RECT 118.975 162.615 119.145 162.785 ;
        RECT 119.435 162.615 119.605 162.785 ;
        RECT 119.895 162.615 120.065 162.785 ;
        RECT 120.355 162.615 120.525 162.785 ;
        RECT 120.815 162.615 120.985 162.785 ;
        RECT 121.275 162.615 121.445 162.785 ;
        RECT 121.735 162.615 121.905 162.785 ;
        RECT 122.195 162.615 122.365 162.785 ;
        RECT 122.655 162.615 122.825 162.785 ;
        RECT 123.115 162.615 123.285 162.785 ;
        RECT 123.575 162.615 123.745 162.785 ;
        RECT 124.035 162.615 124.205 162.785 ;
        RECT 124.495 162.615 124.665 162.785 ;
        RECT 124.955 162.615 125.125 162.785 ;
        RECT 125.415 162.615 125.585 162.785 ;
        RECT 125.875 162.615 126.045 162.785 ;
        RECT 126.335 162.615 126.505 162.785 ;
        RECT 126.795 162.615 126.965 162.785 ;
        RECT 127.255 162.615 127.425 162.785 ;
        RECT 127.715 162.615 127.885 162.785 ;
        RECT 128.175 162.615 128.345 162.785 ;
        RECT 128.635 162.615 128.805 162.785 ;
        RECT 129.095 162.615 129.265 162.785 ;
        RECT 129.555 162.615 129.725 162.785 ;
        RECT 130.015 162.615 130.185 162.785 ;
        RECT 130.475 162.615 130.645 162.785 ;
        RECT 130.935 162.615 131.105 162.785 ;
        RECT 57.335 159.895 57.505 160.065 ;
        RECT 57.795 159.895 57.965 160.065 ;
        RECT 58.255 159.895 58.425 160.065 ;
        RECT 58.715 159.895 58.885 160.065 ;
        RECT 59.175 159.895 59.345 160.065 ;
        RECT 59.635 159.895 59.805 160.065 ;
        RECT 60.095 159.895 60.265 160.065 ;
        RECT 60.555 159.895 60.725 160.065 ;
        RECT 61.015 159.895 61.185 160.065 ;
        RECT 61.475 159.895 61.645 160.065 ;
        RECT 61.935 159.895 62.105 160.065 ;
        RECT 62.395 159.895 62.565 160.065 ;
        RECT 62.855 159.895 63.025 160.065 ;
        RECT 63.315 159.895 63.485 160.065 ;
        RECT 63.775 159.895 63.945 160.065 ;
        RECT 64.235 159.895 64.405 160.065 ;
        RECT 64.695 159.895 64.865 160.065 ;
        RECT 65.155 159.895 65.325 160.065 ;
        RECT 65.615 159.895 65.785 160.065 ;
        RECT 66.075 159.895 66.245 160.065 ;
        RECT 66.535 159.895 66.705 160.065 ;
        RECT 66.995 159.895 67.165 160.065 ;
        RECT 67.455 159.895 67.625 160.065 ;
        RECT 67.915 159.895 68.085 160.065 ;
        RECT 68.375 159.895 68.545 160.065 ;
        RECT 68.835 159.895 69.005 160.065 ;
        RECT 69.295 159.895 69.465 160.065 ;
        RECT 69.755 159.895 69.925 160.065 ;
        RECT 70.215 159.895 70.385 160.065 ;
        RECT 70.675 159.895 70.845 160.065 ;
        RECT 71.135 159.895 71.305 160.065 ;
        RECT 71.595 159.895 71.765 160.065 ;
        RECT 72.055 159.895 72.225 160.065 ;
        RECT 72.515 159.895 72.685 160.065 ;
        RECT 72.975 159.895 73.145 160.065 ;
        RECT 73.435 159.895 73.605 160.065 ;
        RECT 73.895 159.895 74.065 160.065 ;
        RECT 74.355 159.895 74.525 160.065 ;
        RECT 74.815 159.895 74.985 160.065 ;
        RECT 75.275 159.895 75.445 160.065 ;
        RECT 75.735 159.895 75.905 160.065 ;
        RECT 76.195 159.895 76.365 160.065 ;
        RECT 76.655 159.895 76.825 160.065 ;
        RECT 77.115 159.895 77.285 160.065 ;
        RECT 77.575 159.895 77.745 160.065 ;
        RECT 78.035 159.895 78.205 160.065 ;
        RECT 78.495 159.895 78.665 160.065 ;
        RECT 78.955 159.895 79.125 160.065 ;
        RECT 79.415 159.895 79.585 160.065 ;
        RECT 79.875 159.895 80.045 160.065 ;
        RECT 80.335 159.895 80.505 160.065 ;
        RECT 80.795 159.895 80.965 160.065 ;
        RECT 81.255 159.895 81.425 160.065 ;
        RECT 81.715 159.895 81.885 160.065 ;
        RECT 82.175 159.895 82.345 160.065 ;
        RECT 82.635 159.895 82.805 160.065 ;
        RECT 83.095 159.895 83.265 160.065 ;
        RECT 83.555 159.895 83.725 160.065 ;
        RECT 84.015 159.895 84.185 160.065 ;
        RECT 84.475 159.895 84.645 160.065 ;
        RECT 84.935 159.895 85.105 160.065 ;
        RECT 85.395 159.895 85.565 160.065 ;
        RECT 85.855 159.895 86.025 160.065 ;
        RECT 86.315 159.895 86.485 160.065 ;
        RECT 86.775 159.895 86.945 160.065 ;
        RECT 87.235 159.895 87.405 160.065 ;
        RECT 87.695 159.895 87.865 160.065 ;
        RECT 88.155 159.895 88.325 160.065 ;
        RECT 88.615 159.895 88.785 160.065 ;
        RECT 89.075 159.895 89.245 160.065 ;
        RECT 89.535 159.895 89.705 160.065 ;
        RECT 89.995 159.895 90.165 160.065 ;
        RECT 90.455 159.895 90.625 160.065 ;
        RECT 90.915 159.895 91.085 160.065 ;
        RECT 91.375 159.895 91.545 160.065 ;
        RECT 91.835 159.895 92.005 160.065 ;
        RECT 92.295 159.895 92.465 160.065 ;
        RECT 92.755 159.895 92.925 160.065 ;
        RECT 93.215 159.895 93.385 160.065 ;
        RECT 93.675 159.895 93.845 160.065 ;
        RECT 94.135 159.895 94.305 160.065 ;
        RECT 94.595 159.895 94.765 160.065 ;
        RECT 95.055 159.895 95.225 160.065 ;
        RECT 95.515 159.895 95.685 160.065 ;
        RECT 95.975 159.895 96.145 160.065 ;
        RECT 96.435 159.895 96.605 160.065 ;
        RECT 96.895 159.895 97.065 160.065 ;
        RECT 97.355 159.895 97.525 160.065 ;
        RECT 97.815 159.895 97.985 160.065 ;
        RECT 98.275 159.895 98.445 160.065 ;
        RECT 98.735 159.895 98.905 160.065 ;
        RECT 99.195 159.895 99.365 160.065 ;
        RECT 99.655 159.895 99.825 160.065 ;
        RECT 100.115 159.895 100.285 160.065 ;
        RECT 100.575 159.895 100.745 160.065 ;
        RECT 101.035 159.895 101.205 160.065 ;
        RECT 101.495 159.895 101.665 160.065 ;
        RECT 101.955 159.895 102.125 160.065 ;
        RECT 102.415 159.895 102.585 160.065 ;
        RECT 102.875 159.895 103.045 160.065 ;
        RECT 103.335 159.895 103.505 160.065 ;
        RECT 103.795 159.895 103.965 160.065 ;
        RECT 104.255 159.895 104.425 160.065 ;
        RECT 104.715 159.895 104.885 160.065 ;
        RECT 105.175 159.895 105.345 160.065 ;
        RECT 105.635 159.895 105.805 160.065 ;
        RECT 106.095 159.895 106.265 160.065 ;
        RECT 106.555 159.895 106.725 160.065 ;
        RECT 107.015 159.895 107.185 160.065 ;
        RECT 107.475 159.895 107.645 160.065 ;
        RECT 107.935 159.895 108.105 160.065 ;
        RECT 108.395 159.895 108.565 160.065 ;
        RECT 108.855 159.895 109.025 160.065 ;
        RECT 109.315 159.895 109.485 160.065 ;
        RECT 109.775 159.895 109.945 160.065 ;
        RECT 110.235 159.895 110.405 160.065 ;
        RECT 110.695 159.895 110.865 160.065 ;
        RECT 111.155 159.895 111.325 160.065 ;
        RECT 111.615 159.895 111.785 160.065 ;
        RECT 112.075 159.895 112.245 160.065 ;
        RECT 112.535 159.895 112.705 160.065 ;
        RECT 112.995 159.895 113.165 160.065 ;
        RECT 113.455 159.895 113.625 160.065 ;
        RECT 113.915 159.895 114.085 160.065 ;
        RECT 114.375 159.895 114.545 160.065 ;
        RECT 114.835 159.895 115.005 160.065 ;
        RECT 115.295 159.895 115.465 160.065 ;
        RECT 115.755 159.895 115.925 160.065 ;
        RECT 116.215 159.895 116.385 160.065 ;
        RECT 116.675 159.895 116.845 160.065 ;
        RECT 117.135 159.895 117.305 160.065 ;
        RECT 117.595 159.895 117.765 160.065 ;
        RECT 118.055 159.895 118.225 160.065 ;
        RECT 118.515 159.895 118.685 160.065 ;
        RECT 118.975 159.895 119.145 160.065 ;
        RECT 119.435 159.895 119.605 160.065 ;
        RECT 119.895 159.895 120.065 160.065 ;
        RECT 120.355 159.895 120.525 160.065 ;
        RECT 120.815 159.895 120.985 160.065 ;
        RECT 121.275 159.895 121.445 160.065 ;
        RECT 121.735 159.895 121.905 160.065 ;
        RECT 122.195 159.895 122.365 160.065 ;
        RECT 122.655 159.895 122.825 160.065 ;
        RECT 123.115 159.895 123.285 160.065 ;
        RECT 123.575 159.895 123.745 160.065 ;
        RECT 124.035 159.895 124.205 160.065 ;
        RECT 124.495 159.895 124.665 160.065 ;
        RECT 124.955 159.895 125.125 160.065 ;
        RECT 125.415 159.895 125.585 160.065 ;
        RECT 125.875 159.895 126.045 160.065 ;
        RECT 126.335 159.895 126.505 160.065 ;
        RECT 126.795 159.895 126.965 160.065 ;
        RECT 127.255 159.895 127.425 160.065 ;
        RECT 127.715 159.895 127.885 160.065 ;
        RECT 128.175 159.895 128.345 160.065 ;
        RECT 128.635 159.895 128.805 160.065 ;
        RECT 129.095 159.895 129.265 160.065 ;
        RECT 129.555 159.895 129.725 160.065 ;
        RECT 130.015 159.895 130.185 160.065 ;
        RECT 130.475 159.895 130.645 160.065 ;
        RECT 130.935 159.895 131.105 160.065 ;
        RECT 57.335 157.175 57.505 157.345 ;
        RECT 57.795 157.175 57.965 157.345 ;
        RECT 58.255 157.175 58.425 157.345 ;
        RECT 58.715 157.175 58.885 157.345 ;
        RECT 59.175 157.175 59.345 157.345 ;
        RECT 59.635 157.175 59.805 157.345 ;
        RECT 60.095 157.175 60.265 157.345 ;
        RECT 60.555 157.175 60.725 157.345 ;
        RECT 61.015 157.175 61.185 157.345 ;
        RECT 61.475 157.175 61.645 157.345 ;
        RECT 61.935 157.175 62.105 157.345 ;
        RECT 62.395 157.175 62.565 157.345 ;
        RECT 62.855 157.175 63.025 157.345 ;
        RECT 63.315 157.175 63.485 157.345 ;
        RECT 63.775 157.175 63.945 157.345 ;
        RECT 64.235 157.175 64.405 157.345 ;
        RECT 64.695 157.175 64.865 157.345 ;
        RECT 65.155 157.175 65.325 157.345 ;
        RECT 65.615 157.175 65.785 157.345 ;
        RECT 66.075 157.175 66.245 157.345 ;
        RECT 66.535 157.175 66.705 157.345 ;
        RECT 66.995 157.175 67.165 157.345 ;
        RECT 67.455 157.175 67.625 157.345 ;
        RECT 67.915 157.175 68.085 157.345 ;
        RECT 68.375 157.175 68.545 157.345 ;
        RECT 68.835 157.175 69.005 157.345 ;
        RECT 69.295 157.175 69.465 157.345 ;
        RECT 69.755 157.175 69.925 157.345 ;
        RECT 70.215 157.175 70.385 157.345 ;
        RECT 70.675 157.175 70.845 157.345 ;
        RECT 71.135 157.175 71.305 157.345 ;
        RECT 71.595 157.175 71.765 157.345 ;
        RECT 72.055 157.175 72.225 157.345 ;
        RECT 72.515 157.175 72.685 157.345 ;
        RECT 72.975 157.175 73.145 157.345 ;
        RECT 73.435 157.175 73.605 157.345 ;
        RECT 73.895 157.175 74.065 157.345 ;
        RECT 74.355 157.175 74.525 157.345 ;
        RECT 74.815 157.175 74.985 157.345 ;
        RECT 75.275 157.175 75.445 157.345 ;
        RECT 75.735 157.175 75.905 157.345 ;
        RECT 76.195 157.175 76.365 157.345 ;
        RECT 76.655 157.175 76.825 157.345 ;
        RECT 77.115 157.175 77.285 157.345 ;
        RECT 77.575 157.175 77.745 157.345 ;
        RECT 78.035 157.175 78.205 157.345 ;
        RECT 78.495 157.175 78.665 157.345 ;
        RECT 78.955 157.175 79.125 157.345 ;
        RECT 79.415 157.175 79.585 157.345 ;
        RECT 79.875 157.175 80.045 157.345 ;
        RECT 80.335 157.175 80.505 157.345 ;
        RECT 80.795 157.175 80.965 157.345 ;
        RECT 81.255 157.175 81.425 157.345 ;
        RECT 81.715 157.175 81.885 157.345 ;
        RECT 82.175 157.175 82.345 157.345 ;
        RECT 82.635 157.175 82.805 157.345 ;
        RECT 83.095 157.175 83.265 157.345 ;
        RECT 83.555 157.175 83.725 157.345 ;
        RECT 84.015 157.175 84.185 157.345 ;
        RECT 84.475 157.175 84.645 157.345 ;
        RECT 84.935 157.175 85.105 157.345 ;
        RECT 85.395 157.175 85.565 157.345 ;
        RECT 85.855 157.175 86.025 157.345 ;
        RECT 86.315 157.175 86.485 157.345 ;
        RECT 86.775 157.175 86.945 157.345 ;
        RECT 87.235 157.175 87.405 157.345 ;
        RECT 87.695 157.175 87.865 157.345 ;
        RECT 88.155 157.175 88.325 157.345 ;
        RECT 88.615 157.175 88.785 157.345 ;
        RECT 89.075 157.175 89.245 157.345 ;
        RECT 89.535 157.175 89.705 157.345 ;
        RECT 89.995 157.175 90.165 157.345 ;
        RECT 90.455 157.175 90.625 157.345 ;
        RECT 90.915 157.175 91.085 157.345 ;
        RECT 91.375 157.175 91.545 157.345 ;
        RECT 91.835 157.175 92.005 157.345 ;
        RECT 92.295 157.175 92.465 157.345 ;
        RECT 92.755 157.175 92.925 157.345 ;
        RECT 93.215 157.175 93.385 157.345 ;
        RECT 93.675 157.175 93.845 157.345 ;
        RECT 94.135 157.175 94.305 157.345 ;
        RECT 94.595 157.175 94.765 157.345 ;
        RECT 95.055 157.175 95.225 157.345 ;
        RECT 95.515 157.175 95.685 157.345 ;
        RECT 95.975 157.175 96.145 157.345 ;
        RECT 96.435 157.175 96.605 157.345 ;
        RECT 96.895 157.175 97.065 157.345 ;
        RECT 97.355 157.175 97.525 157.345 ;
        RECT 97.815 157.175 97.985 157.345 ;
        RECT 98.275 157.175 98.445 157.345 ;
        RECT 98.735 157.175 98.905 157.345 ;
        RECT 99.195 157.175 99.365 157.345 ;
        RECT 99.655 157.175 99.825 157.345 ;
        RECT 100.115 157.175 100.285 157.345 ;
        RECT 100.575 157.175 100.745 157.345 ;
        RECT 101.035 157.175 101.205 157.345 ;
        RECT 101.495 157.175 101.665 157.345 ;
        RECT 101.955 157.175 102.125 157.345 ;
        RECT 102.415 157.175 102.585 157.345 ;
        RECT 102.875 157.175 103.045 157.345 ;
        RECT 103.335 157.175 103.505 157.345 ;
        RECT 103.795 157.175 103.965 157.345 ;
        RECT 104.255 157.175 104.425 157.345 ;
        RECT 104.715 157.175 104.885 157.345 ;
        RECT 105.175 157.175 105.345 157.345 ;
        RECT 105.635 157.175 105.805 157.345 ;
        RECT 106.095 157.175 106.265 157.345 ;
        RECT 106.555 157.175 106.725 157.345 ;
        RECT 107.015 157.175 107.185 157.345 ;
        RECT 107.475 157.175 107.645 157.345 ;
        RECT 107.935 157.175 108.105 157.345 ;
        RECT 108.395 157.175 108.565 157.345 ;
        RECT 108.855 157.175 109.025 157.345 ;
        RECT 109.315 157.175 109.485 157.345 ;
        RECT 109.775 157.175 109.945 157.345 ;
        RECT 110.235 157.175 110.405 157.345 ;
        RECT 110.695 157.175 110.865 157.345 ;
        RECT 111.155 157.175 111.325 157.345 ;
        RECT 111.615 157.175 111.785 157.345 ;
        RECT 112.075 157.175 112.245 157.345 ;
        RECT 112.535 157.175 112.705 157.345 ;
        RECT 112.995 157.175 113.165 157.345 ;
        RECT 113.455 157.175 113.625 157.345 ;
        RECT 113.915 157.175 114.085 157.345 ;
        RECT 114.375 157.175 114.545 157.345 ;
        RECT 114.835 157.175 115.005 157.345 ;
        RECT 115.295 157.175 115.465 157.345 ;
        RECT 115.755 157.175 115.925 157.345 ;
        RECT 116.215 157.175 116.385 157.345 ;
        RECT 116.675 157.175 116.845 157.345 ;
        RECT 117.135 157.175 117.305 157.345 ;
        RECT 117.595 157.175 117.765 157.345 ;
        RECT 118.055 157.175 118.225 157.345 ;
        RECT 118.515 157.175 118.685 157.345 ;
        RECT 118.975 157.175 119.145 157.345 ;
        RECT 119.435 157.175 119.605 157.345 ;
        RECT 119.895 157.175 120.065 157.345 ;
        RECT 120.355 157.175 120.525 157.345 ;
        RECT 120.815 157.175 120.985 157.345 ;
        RECT 121.275 157.175 121.445 157.345 ;
        RECT 121.735 157.175 121.905 157.345 ;
        RECT 122.195 157.175 122.365 157.345 ;
        RECT 122.655 157.175 122.825 157.345 ;
        RECT 123.115 157.175 123.285 157.345 ;
        RECT 123.575 157.175 123.745 157.345 ;
        RECT 124.035 157.175 124.205 157.345 ;
        RECT 124.495 157.175 124.665 157.345 ;
        RECT 124.955 157.175 125.125 157.345 ;
        RECT 125.415 157.175 125.585 157.345 ;
        RECT 125.875 157.175 126.045 157.345 ;
        RECT 126.335 157.175 126.505 157.345 ;
        RECT 126.795 157.175 126.965 157.345 ;
        RECT 127.255 157.175 127.425 157.345 ;
        RECT 127.715 157.175 127.885 157.345 ;
        RECT 128.175 157.175 128.345 157.345 ;
        RECT 128.635 157.175 128.805 157.345 ;
        RECT 129.095 157.175 129.265 157.345 ;
        RECT 129.555 157.175 129.725 157.345 ;
        RECT 130.015 157.175 130.185 157.345 ;
        RECT 130.475 157.175 130.645 157.345 ;
        RECT 130.935 157.175 131.105 157.345 ;
        RECT 57.335 154.455 57.505 154.625 ;
        RECT 57.795 154.455 57.965 154.625 ;
        RECT 58.255 154.455 58.425 154.625 ;
        RECT 58.715 154.455 58.885 154.625 ;
        RECT 59.175 154.455 59.345 154.625 ;
        RECT 59.635 154.455 59.805 154.625 ;
        RECT 60.095 154.455 60.265 154.625 ;
        RECT 60.555 154.455 60.725 154.625 ;
        RECT 61.015 154.455 61.185 154.625 ;
        RECT 61.475 154.455 61.645 154.625 ;
        RECT 61.935 154.455 62.105 154.625 ;
        RECT 62.395 154.455 62.565 154.625 ;
        RECT 62.855 154.455 63.025 154.625 ;
        RECT 63.315 154.455 63.485 154.625 ;
        RECT 63.775 154.455 63.945 154.625 ;
        RECT 64.235 154.455 64.405 154.625 ;
        RECT 64.695 154.455 64.865 154.625 ;
        RECT 65.155 154.455 65.325 154.625 ;
        RECT 65.615 154.455 65.785 154.625 ;
        RECT 66.075 154.455 66.245 154.625 ;
        RECT 66.535 154.455 66.705 154.625 ;
        RECT 66.995 154.455 67.165 154.625 ;
        RECT 67.455 154.455 67.625 154.625 ;
        RECT 67.915 154.455 68.085 154.625 ;
        RECT 68.375 154.455 68.545 154.625 ;
        RECT 68.835 154.455 69.005 154.625 ;
        RECT 69.295 154.455 69.465 154.625 ;
        RECT 69.755 154.455 69.925 154.625 ;
        RECT 70.215 154.455 70.385 154.625 ;
        RECT 70.675 154.455 70.845 154.625 ;
        RECT 71.135 154.455 71.305 154.625 ;
        RECT 71.595 154.455 71.765 154.625 ;
        RECT 72.055 154.455 72.225 154.625 ;
        RECT 72.515 154.455 72.685 154.625 ;
        RECT 72.975 154.455 73.145 154.625 ;
        RECT 73.435 154.455 73.605 154.625 ;
        RECT 73.895 154.455 74.065 154.625 ;
        RECT 74.355 154.455 74.525 154.625 ;
        RECT 74.815 154.455 74.985 154.625 ;
        RECT 75.275 154.455 75.445 154.625 ;
        RECT 75.735 154.455 75.905 154.625 ;
        RECT 76.195 154.455 76.365 154.625 ;
        RECT 76.655 154.455 76.825 154.625 ;
        RECT 77.115 154.455 77.285 154.625 ;
        RECT 77.575 154.455 77.745 154.625 ;
        RECT 78.035 154.455 78.205 154.625 ;
        RECT 78.495 154.455 78.665 154.625 ;
        RECT 78.955 154.455 79.125 154.625 ;
        RECT 79.415 154.455 79.585 154.625 ;
        RECT 79.875 154.455 80.045 154.625 ;
        RECT 80.335 154.455 80.505 154.625 ;
        RECT 80.795 154.455 80.965 154.625 ;
        RECT 81.255 154.455 81.425 154.625 ;
        RECT 81.715 154.455 81.885 154.625 ;
        RECT 82.175 154.455 82.345 154.625 ;
        RECT 82.635 154.455 82.805 154.625 ;
        RECT 83.095 154.455 83.265 154.625 ;
        RECT 83.555 154.455 83.725 154.625 ;
        RECT 84.015 154.455 84.185 154.625 ;
        RECT 84.475 154.455 84.645 154.625 ;
        RECT 84.935 154.455 85.105 154.625 ;
        RECT 85.395 154.455 85.565 154.625 ;
        RECT 85.855 154.455 86.025 154.625 ;
        RECT 86.315 154.455 86.485 154.625 ;
        RECT 86.775 154.455 86.945 154.625 ;
        RECT 87.235 154.455 87.405 154.625 ;
        RECT 87.695 154.455 87.865 154.625 ;
        RECT 88.155 154.455 88.325 154.625 ;
        RECT 88.615 154.455 88.785 154.625 ;
        RECT 89.075 154.455 89.245 154.625 ;
        RECT 89.535 154.455 89.705 154.625 ;
        RECT 89.995 154.455 90.165 154.625 ;
        RECT 90.455 154.455 90.625 154.625 ;
        RECT 90.915 154.455 91.085 154.625 ;
        RECT 91.375 154.455 91.545 154.625 ;
        RECT 91.835 154.455 92.005 154.625 ;
        RECT 92.295 154.455 92.465 154.625 ;
        RECT 92.755 154.455 92.925 154.625 ;
        RECT 93.215 154.455 93.385 154.625 ;
        RECT 93.675 154.455 93.845 154.625 ;
        RECT 94.135 154.455 94.305 154.625 ;
        RECT 94.595 154.455 94.765 154.625 ;
        RECT 95.055 154.455 95.225 154.625 ;
        RECT 95.515 154.455 95.685 154.625 ;
        RECT 95.975 154.455 96.145 154.625 ;
        RECT 96.435 154.455 96.605 154.625 ;
        RECT 96.895 154.455 97.065 154.625 ;
        RECT 97.355 154.455 97.525 154.625 ;
        RECT 97.815 154.455 97.985 154.625 ;
        RECT 98.275 154.455 98.445 154.625 ;
        RECT 98.735 154.455 98.905 154.625 ;
        RECT 99.195 154.455 99.365 154.625 ;
        RECT 99.655 154.455 99.825 154.625 ;
        RECT 100.115 154.455 100.285 154.625 ;
        RECT 100.575 154.455 100.745 154.625 ;
        RECT 101.035 154.455 101.205 154.625 ;
        RECT 101.495 154.455 101.665 154.625 ;
        RECT 101.955 154.455 102.125 154.625 ;
        RECT 102.415 154.455 102.585 154.625 ;
        RECT 102.875 154.455 103.045 154.625 ;
        RECT 103.335 154.455 103.505 154.625 ;
        RECT 103.795 154.455 103.965 154.625 ;
        RECT 104.255 154.455 104.425 154.625 ;
        RECT 104.715 154.455 104.885 154.625 ;
        RECT 105.175 154.455 105.345 154.625 ;
        RECT 105.635 154.455 105.805 154.625 ;
        RECT 106.095 154.455 106.265 154.625 ;
        RECT 106.555 154.455 106.725 154.625 ;
        RECT 107.015 154.455 107.185 154.625 ;
        RECT 107.475 154.455 107.645 154.625 ;
        RECT 107.935 154.455 108.105 154.625 ;
        RECT 108.395 154.455 108.565 154.625 ;
        RECT 108.855 154.455 109.025 154.625 ;
        RECT 109.315 154.455 109.485 154.625 ;
        RECT 109.775 154.455 109.945 154.625 ;
        RECT 110.235 154.455 110.405 154.625 ;
        RECT 110.695 154.455 110.865 154.625 ;
        RECT 111.155 154.455 111.325 154.625 ;
        RECT 111.615 154.455 111.785 154.625 ;
        RECT 112.075 154.455 112.245 154.625 ;
        RECT 112.535 154.455 112.705 154.625 ;
        RECT 112.995 154.455 113.165 154.625 ;
        RECT 113.455 154.455 113.625 154.625 ;
        RECT 113.915 154.455 114.085 154.625 ;
        RECT 114.375 154.455 114.545 154.625 ;
        RECT 114.835 154.455 115.005 154.625 ;
        RECT 115.295 154.455 115.465 154.625 ;
        RECT 115.755 154.455 115.925 154.625 ;
        RECT 116.215 154.455 116.385 154.625 ;
        RECT 116.675 154.455 116.845 154.625 ;
        RECT 117.135 154.455 117.305 154.625 ;
        RECT 117.595 154.455 117.765 154.625 ;
        RECT 118.055 154.455 118.225 154.625 ;
        RECT 118.515 154.455 118.685 154.625 ;
        RECT 118.975 154.455 119.145 154.625 ;
        RECT 119.435 154.455 119.605 154.625 ;
        RECT 119.895 154.455 120.065 154.625 ;
        RECT 120.355 154.455 120.525 154.625 ;
        RECT 120.815 154.455 120.985 154.625 ;
        RECT 121.275 154.455 121.445 154.625 ;
        RECT 121.735 154.455 121.905 154.625 ;
        RECT 122.195 154.455 122.365 154.625 ;
        RECT 122.655 154.455 122.825 154.625 ;
        RECT 123.115 154.455 123.285 154.625 ;
        RECT 123.575 154.455 123.745 154.625 ;
        RECT 124.035 154.455 124.205 154.625 ;
        RECT 124.495 154.455 124.665 154.625 ;
        RECT 124.955 154.455 125.125 154.625 ;
        RECT 125.415 154.455 125.585 154.625 ;
        RECT 125.875 154.455 126.045 154.625 ;
        RECT 126.335 154.455 126.505 154.625 ;
        RECT 126.795 154.455 126.965 154.625 ;
        RECT 127.255 154.455 127.425 154.625 ;
        RECT 127.715 154.455 127.885 154.625 ;
        RECT 128.175 154.455 128.345 154.625 ;
        RECT 128.635 154.455 128.805 154.625 ;
        RECT 129.095 154.455 129.265 154.625 ;
        RECT 129.555 154.455 129.725 154.625 ;
        RECT 130.015 154.455 130.185 154.625 ;
        RECT 130.475 154.455 130.645 154.625 ;
        RECT 130.935 154.455 131.105 154.625 ;
        RECT 57.335 151.735 57.505 151.905 ;
        RECT 57.795 151.735 57.965 151.905 ;
        RECT 58.255 151.735 58.425 151.905 ;
        RECT 58.715 151.735 58.885 151.905 ;
        RECT 59.175 151.735 59.345 151.905 ;
        RECT 59.635 151.735 59.805 151.905 ;
        RECT 60.095 151.735 60.265 151.905 ;
        RECT 60.555 151.735 60.725 151.905 ;
        RECT 61.015 151.735 61.185 151.905 ;
        RECT 61.475 151.735 61.645 151.905 ;
        RECT 61.935 151.735 62.105 151.905 ;
        RECT 62.395 151.735 62.565 151.905 ;
        RECT 62.855 151.735 63.025 151.905 ;
        RECT 63.315 151.735 63.485 151.905 ;
        RECT 63.775 151.735 63.945 151.905 ;
        RECT 64.235 151.735 64.405 151.905 ;
        RECT 64.695 151.735 64.865 151.905 ;
        RECT 65.155 151.735 65.325 151.905 ;
        RECT 65.615 151.735 65.785 151.905 ;
        RECT 66.075 151.735 66.245 151.905 ;
        RECT 66.535 151.735 66.705 151.905 ;
        RECT 66.995 151.735 67.165 151.905 ;
        RECT 67.455 151.735 67.625 151.905 ;
        RECT 67.915 151.735 68.085 151.905 ;
        RECT 68.375 151.735 68.545 151.905 ;
        RECT 68.835 151.735 69.005 151.905 ;
        RECT 69.295 151.735 69.465 151.905 ;
        RECT 69.755 151.735 69.925 151.905 ;
        RECT 70.215 151.735 70.385 151.905 ;
        RECT 70.675 151.735 70.845 151.905 ;
        RECT 71.135 151.735 71.305 151.905 ;
        RECT 71.595 151.735 71.765 151.905 ;
        RECT 72.055 151.735 72.225 151.905 ;
        RECT 72.515 151.735 72.685 151.905 ;
        RECT 72.975 151.735 73.145 151.905 ;
        RECT 73.435 151.735 73.605 151.905 ;
        RECT 73.895 151.735 74.065 151.905 ;
        RECT 74.355 151.735 74.525 151.905 ;
        RECT 74.815 151.735 74.985 151.905 ;
        RECT 75.275 151.735 75.445 151.905 ;
        RECT 75.735 151.735 75.905 151.905 ;
        RECT 76.195 151.735 76.365 151.905 ;
        RECT 76.655 151.735 76.825 151.905 ;
        RECT 77.115 151.735 77.285 151.905 ;
        RECT 77.575 151.735 77.745 151.905 ;
        RECT 78.035 151.735 78.205 151.905 ;
        RECT 78.495 151.735 78.665 151.905 ;
        RECT 78.955 151.735 79.125 151.905 ;
        RECT 79.415 151.735 79.585 151.905 ;
        RECT 79.875 151.735 80.045 151.905 ;
        RECT 80.335 151.735 80.505 151.905 ;
        RECT 80.795 151.735 80.965 151.905 ;
        RECT 81.255 151.735 81.425 151.905 ;
        RECT 81.715 151.735 81.885 151.905 ;
        RECT 82.175 151.735 82.345 151.905 ;
        RECT 82.635 151.735 82.805 151.905 ;
        RECT 83.095 151.735 83.265 151.905 ;
        RECT 83.555 151.735 83.725 151.905 ;
        RECT 84.015 151.735 84.185 151.905 ;
        RECT 84.475 151.735 84.645 151.905 ;
        RECT 84.935 151.735 85.105 151.905 ;
        RECT 85.395 151.735 85.565 151.905 ;
        RECT 85.855 151.735 86.025 151.905 ;
        RECT 86.315 151.735 86.485 151.905 ;
        RECT 86.775 151.735 86.945 151.905 ;
        RECT 87.235 151.735 87.405 151.905 ;
        RECT 87.695 151.735 87.865 151.905 ;
        RECT 88.155 151.735 88.325 151.905 ;
        RECT 88.615 151.735 88.785 151.905 ;
        RECT 89.075 151.735 89.245 151.905 ;
        RECT 89.535 151.735 89.705 151.905 ;
        RECT 89.995 151.735 90.165 151.905 ;
        RECT 90.455 151.735 90.625 151.905 ;
        RECT 90.915 151.735 91.085 151.905 ;
        RECT 91.375 151.735 91.545 151.905 ;
        RECT 91.835 151.735 92.005 151.905 ;
        RECT 92.295 151.735 92.465 151.905 ;
        RECT 92.755 151.735 92.925 151.905 ;
        RECT 93.215 151.735 93.385 151.905 ;
        RECT 93.675 151.735 93.845 151.905 ;
        RECT 94.135 151.735 94.305 151.905 ;
        RECT 94.595 151.735 94.765 151.905 ;
        RECT 95.055 151.735 95.225 151.905 ;
        RECT 95.515 151.735 95.685 151.905 ;
        RECT 95.975 151.735 96.145 151.905 ;
        RECT 96.435 151.735 96.605 151.905 ;
        RECT 96.895 151.735 97.065 151.905 ;
        RECT 97.355 151.735 97.525 151.905 ;
        RECT 97.815 151.735 97.985 151.905 ;
        RECT 98.275 151.735 98.445 151.905 ;
        RECT 98.735 151.735 98.905 151.905 ;
        RECT 99.195 151.735 99.365 151.905 ;
        RECT 99.655 151.735 99.825 151.905 ;
        RECT 100.115 151.735 100.285 151.905 ;
        RECT 100.575 151.735 100.745 151.905 ;
        RECT 101.035 151.735 101.205 151.905 ;
        RECT 101.495 151.735 101.665 151.905 ;
        RECT 101.955 151.735 102.125 151.905 ;
        RECT 102.415 151.735 102.585 151.905 ;
        RECT 102.875 151.735 103.045 151.905 ;
        RECT 103.335 151.735 103.505 151.905 ;
        RECT 103.795 151.735 103.965 151.905 ;
        RECT 104.255 151.735 104.425 151.905 ;
        RECT 104.715 151.735 104.885 151.905 ;
        RECT 105.175 151.735 105.345 151.905 ;
        RECT 105.635 151.735 105.805 151.905 ;
        RECT 106.095 151.735 106.265 151.905 ;
        RECT 106.555 151.735 106.725 151.905 ;
        RECT 107.015 151.735 107.185 151.905 ;
        RECT 107.475 151.735 107.645 151.905 ;
        RECT 107.935 151.735 108.105 151.905 ;
        RECT 108.395 151.735 108.565 151.905 ;
        RECT 108.855 151.735 109.025 151.905 ;
        RECT 109.315 151.735 109.485 151.905 ;
        RECT 109.775 151.735 109.945 151.905 ;
        RECT 110.235 151.735 110.405 151.905 ;
        RECT 110.695 151.735 110.865 151.905 ;
        RECT 111.155 151.735 111.325 151.905 ;
        RECT 111.615 151.735 111.785 151.905 ;
        RECT 112.075 151.735 112.245 151.905 ;
        RECT 112.535 151.735 112.705 151.905 ;
        RECT 112.995 151.735 113.165 151.905 ;
        RECT 113.455 151.735 113.625 151.905 ;
        RECT 113.915 151.735 114.085 151.905 ;
        RECT 114.375 151.735 114.545 151.905 ;
        RECT 114.835 151.735 115.005 151.905 ;
        RECT 115.295 151.735 115.465 151.905 ;
        RECT 115.755 151.735 115.925 151.905 ;
        RECT 116.215 151.735 116.385 151.905 ;
        RECT 116.675 151.735 116.845 151.905 ;
        RECT 117.135 151.735 117.305 151.905 ;
        RECT 117.595 151.735 117.765 151.905 ;
        RECT 118.055 151.735 118.225 151.905 ;
        RECT 118.515 151.735 118.685 151.905 ;
        RECT 118.975 151.735 119.145 151.905 ;
        RECT 119.435 151.735 119.605 151.905 ;
        RECT 119.895 151.735 120.065 151.905 ;
        RECT 120.355 151.735 120.525 151.905 ;
        RECT 120.815 151.735 120.985 151.905 ;
        RECT 121.275 151.735 121.445 151.905 ;
        RECT 121.735 151.735 121.905 151.905 ;
        RECT 122.195 151.735 122.365 151.905 ;
        RECT 122.655 151.735 122.825 151.905 ;
        RECT 123.115 151.735 123.285 151.905 ;
        RECT 123.575 151.735 123.745 151.905 ;
        RECT 124.035 151.735 124.205 151.905 ;
        RECT 124.495 151.735 124.665 151.905 ;
        RECT 124.955 151.735 125.125 151.905 ;
        RECT 125.415 151.735 125.585 151.905 ;
        RECT 125.875 151.735 126.045 151.905 ;
        RECT 126.335 151.735 126.505 151.905 ;
        RECT 126.795 151.735 126.965 151.905 ;
        RECT 127.255 151.735 127.425 151.905 ;
        RECT 127.715 151.735 127.885 151.905 ;
        RECT 128.175 151.735 128.345 151.905 ;
        RECT 128.635 151.735 128.805 151.905 ;
        RECT 129.095 151.735 129.265 151.905 ;
        RECT 129.555 151.735 129.725 151.905 ;
        RECT 130.015 151.735 130.185 151.905 ;
        RECT 130.475 151.735 130.645 151.905 ;
        RECT 130.935 151.735 131.105 151.905 ;
        RECT 111.155 150.885 111.325 151.055 ;
        RECT 110.695 149.525 110.865 149.695 ;
        RECT 57.335 149.015 57.505 149.185 ;
        RECT 57.795 149.015 57.965 149.185 ;
        RECT 58.255 149.015 58.425 149.185 ;
        RECT 58.715 149.015 58.885 149.185 ;
        RECT 59.175 149.015 59.345 149.185 ;
        RECT 59.635 149.015 59.805 149.185 ;
        RECT 60.095 149.015 60.265 149.185 ;
        RECT 60.555 149.015 60.725 149.185 ;
        RECT 61.015 149.015 61.185 149.185 ;
        RECT 61.475 149.015 61.645 149.185 ;
        RECT 61.935 149.015 62.105 149.185 ;
        RECT 62.395 149.015 62.565 149.185 ;
        RECT 62.855 149.015 63.025 149.185 ;
        RECT 63.315 149.015 63.485 149.185 ;
        RECT 63.775 149.015 63.945 149.185 ;
        RECT 64.235 149.015 64.405 149.185 ;
        RECT 64.695 149.015 64.865 149.185 ;
        RECT 65.155 149.015 65.325 149.185 ;
        RECT 65.615 149.015 65.785 149.185 ;
        RECT 66.075 149.015 66.245 149.185 ;
        RECT 66.535 149.015 66.705 149.185 ;
        RECT 66.995 149.015 67.165 149.185 ;
        RECT 67.455 149.015 67.625 149.185 ;
        RECT 67.915 149.015 68.085 149.185 ;
        RECT 68.375 149.015 68.545 149.185 ;
        RECT 68.835 149.015 69.005 149.185 ;
        RECT 69.295 149.015 69.465 149.185 ;
        RECT 69.755 149.015 69.925 149.185 ;
        RECT 70.215 149.015 70.385 149.185 ;
        RECT 70.675 149.015 70.845 149.185 ;
        RECT 71.135 149.015 71.305 149.185 ;
        RECT 71.595 149.015 71.765 149.185 ;
        RECT 72.055 149.015 72.225 149.185 ;
        RECT 72.515 149.015 72.685 149.185 ;
        RECT 72.975 149.015 73.145 149.185 ;
        RECT 73.435 149.015 73.605 149.185 ;
        RECT 73.895 149.015 74.065 149.185 ;
        RECT 74.355 149.015 74.525 149.185 ;
        RECT 74.815 149.015 74.985 149.185 ;
        RECT 75.275 149.015 75.445 149.185 ;
        RECT 75.735 149.015 75.905 149.185 ;
        RECT 76.195 149.015 76.365 149.185 ;
        RECT 76.655 149.015 76.825 149.185 ;
        RECT 77.115 149.015 77.285 149.185 ;
        RECT 77.575 149.015 77.745 149.185 ;
        RECT 78.035 149.015 78.205 149.185 ;
        RECT 78.495 149.015 78.665 149.185 ;
        RECT 78.955 149.015 79.125 149.185 ;
        RECT 79.415 149.015 79.585 149.185 ;
        RECT 79.875 149.015 80.045 149.185 ;
        RECT 80.335 149.015 80.505 149.185 ;
        RECT 80.795 149.015 80.965 149.185 ;
        RECT 81.255 149.015 81.425 149.185 ;
        RECT 81.715 149.015 81.885 149.185 ;
        RECT 82.175 149.015 82.345 149.185 ;
        RECT 82.635 149.015 82.805 149.185 ;
        RECT 83.095 149.015 83.265 149.185 ;
        RECT 83.555 149.015 83.725 149.185 ;
        RECT 84.015 149.015 84.185 149.185 ;
        RECT 84.475 149.015 84.645 149.185 ;
        RECT 84.935 149.015 85.105 149.185 ;
        RECT 85.395 149.015 85.565 149.185 ;
        RECT 85.855 149.015 86.025 149.185 ;
        RECT 86.315 149.015 86.485 149.185 ;
        RECT 86.775 149.015 86.945 149.185 ;
        RECT 87.235 149.015 87.405 149.185 ;
        RECT 87.695 149.015 87.865 149.185 ;
        RECT 88.155 149.015 88.325 149.185 ;
        RECT 88.615 149.015 88.785 149.185 ;
        RECT 89.075 149.015 89.245 149.185 ;
        RECT 89.535 149.015 89.705 149.185 ;
        RECT 89.995 149.015 90.165 149.185 ;
        RECT 90.455 149.015 90.625 149.185 ;
        RECT 90.915 149.015 91.085 149.185 ;
        RECT 91.375 149.015 91.545 149.185 ;
        RECT 91.835 149.015 92.005 149.185 ;
        RECT 92.295 149.015 92.465 149.185 ;
        RECT 92.755 149.015 92.925 149.185 ;
        RECT 93.215 149.015 93.385 149.185 ;
        RECT 93.675 149.015 93.845 149.185 ;
        RECT 94.135 149.015 94.305 149.185 ;
        RECT 94.595 149.015 94.765 149.185 ;
        RECT 95.055 149.015 95.225 149.185 ;
        RECT 95.515 149.015 95.685 149.185 ;
        RECT 95.975 149.015 96.145 149.185 ;
        RECT 96.435 149.015 96.605 149.185 ;
        RECT 96.895 149.015 97.065 149.185 ;
        RECT 97.355 149.015 97.525 149.185 ;
        RECT 97.815 149.015 97.985 149.185 ;
        RECT 98.275 149.015 98.445 149.185 ;
        RECT 98.735 149.015 98.905 149.185 ;
        RECT 99.195 149.015 99.365 149.185 ;
        RECT 99.655 149.015 99.825 149.185 ;
        RECT 100.115 149.015 100.285 149.185 ;
        RECT 100.575 149.015 100.745 149.185 ;
        RECT 101.035 149.015 101.205 149.185 ;
        RECT 101.495 149.015 101.665 149.185 ;
        RECT 101.955 149.015 102.125 149.185 ;
        RECT 102.415 149.015 102.585 149.185 ;
        RECT 102.875 149.015 103.045 149.185 ;
        RECT 103.335 149.015 103.505 149.185 ;
        RECT 103.795 149.015 103.965 149.185 ;
        RECT 104.255 149.015 104.425 149.185 ;
        RECT 104.715 149.015 104.885 149.185 ;
        RECT 105.175 149.015 105.345 149.185 ;
        RECT 105.635 149.015 105.805 149.185 ;
        RECT 106.095 149.015 106.265 149.185 ;
        RECT 106.555 149.015 106.725 149.185 ;
        RECT 107.015 149.015 107.185 149.185 ;
        RECT 107.475 149.015 107.645 149.185 ;
        RECT 107.935 149.015 108.105 149.185 ;
        RECT 108.395 149.015 108.565 149.185 ;
        RECT 108.855 149.015 109.025 149.185 ;
        RECT 109.315 149.015 109.485 149.185 ;
        RECT 109.775 149.015 109.945 149.185 ;
        RECT 110.235 149.015 110.405 149.185 ;
        RECT 110.695 149.015 110.865 149.185 ;
        RECT 111.155 149.015 111.325 149.185 ;
        RECT 111.615 149.015 111.785 149.185 ;
        RECT 112.075 149.015 112.245 149.185 ;
        RECT 112.535 149.015 112.705 149.185 ;
        RECT 112.995 149.015 113.165 149.185 ;
        RECT 113.455 149.015 113.625 149.185 ;
        RECT 113.915 149.015 114.085 149.185 ;
        RECT 114.375 149.015 114.545 149.185 ;
        RECT 114.835 149.015 115.005 149.185 ;
        RECT 115.295 149.015 115.465 149.185 ;
        RECT 115.755 149.015 115.925 149.185 ;
        RECT 116.215 149.015 116.385 149.185 ;
        RECT 116.675 149.015 116.845 149.185 ;
        RECT 117.135 149.015 117.305 149.185 ;
        RECT 117.595 149.015 117.765 149.185 ;
        RECT 118.055 149.015 118.225 149.185 ;
        RECT 118.515 149.015 118.685 149.185 ;
        RECT 118.975 149.015 119.145 149.185 ;
        RECT 119.435 149.015 119.605 149.185 ;
        RECT 119.895 149.015 120.065 149.185 ;
        RECT 120.355 149.015 120.525 149.185 ;
        RECT 120.815 149.015 120.985 149.185 ;
        RECT 121.275 149.015 121.445 149.185 ;
        RECT 121.735 149.015 121.905 149.185 ;
        RECT 122.195 149.015 122.365 149.185 ;
        RECT 122.655 149.015 122.825 149.185 ;
        RECT 123.115 149.015 123.285 149.185 ;
        RECT 123.575 149.015 123.745 149.185 ;
        RECT 124.035 149.015 124.205 149.185 ;
        RECT 124.495 149.015 124.665 149.185 ;
        RECT 124.955 149.015 125.125 149.185 ;
        RECT 125.415 149.015 125.585 149.185 ;
        RECT 125.875 149.015 126.045 149.185 ;
        RECT 126.335 149.015 126.505 149.185 ;
        RECT 126.795 149.015 126.965 149.185 ;
        RECT 127.255 149.015 127.425 149.185 ;
        RECT 127.715 149.015 127.885 149.185 ;
        RECT 128.175 149.015 128.345 149.185 ;
        RECT 128.635 149.015 128.805 149.185 ;
        RECT 129.095 149.015 129.265 149.185 ;
        RECT 129.555 149.015 129.725 149.185 ;
        RECT 130.015 149.015 130.185 149.185 ;
        RECT 130.475 149.015 130.645 149.185 ;
        RECT 130.935 149.015 131.105 149.185 ;
        RECT 57.335 146.295 57.505 146.465 ;
        RECT 57.795 146.295 57.965 146.465 ;
        RECT 58.255 146.295 58.425 146.465 ;
        RECT 58.715 146.295 58.885 146.465 ;
        RECT 59.175 146.295 59.345 146.465 ;
        RECT 59.635 146.295 59.805 146.465 ;
        RECT 60.095 146.295 60.265 146.465 ;
        RECT 60.555 146.295 60.725 146.465 ;
        RECT 61.015 146.295 61.185 146.465 ;
        RECT 61.475 146.295 61.645 146.465 ;
        RECT 61.935 146.295 62.105 146.465 ;
        RECT 62.395 146.295 62.565 146.465 ;
        RECT 62.855 146.295 63.025 146.465 ;
        RECT 63.315 146.295 63.485 146.465 ;
        RECT 63.775 146.295 63.945 146.465 ;
        RECT 64.235 146.295 64.405 146.465 ;
        RECT 64.695 146.295 64.865 146.465 ;
        RECT 65.155 146.295 65.325 146.465 ;
        RECT 65.615 146.295 65.785 146.465 ;
        RECT 66.075 146.295 66.245 146.465 ;
        RECT 66.535 146.295 66.705 146.465 ;
        RECT 66.995 146.295 67.165 146.465 ;
        RECT 67.455 146.295 67.625 146.465 ;
        RECT 67.915 146.295 68.085 146.465 ;
        RECT 68.375 146.295 68.545 146.465 ;
        RECT 68.835 146.295 69.005 146.465 ;
        RECT 69.295 146.295 69.465 146.465 ;
        RECT 69.755 146.295 69.925 146.465 ;
        RECT 70.215 146.295 70.385 146.465 ;
        RECT 70.675 146.295 70.845 146.465 ;
        RECT 71.135 146.295 71.305 146.465 ;
        RECT 71.595 146.295 71.765 146.465 ;
        RECT 72.055 146.295 72.225 146.465 ;
        RECT 72.515 146.295 72.685 146.465 ;
        RECT 72.975 146.295 73.145 146.465 ;
        RECT 73.435 146.295 73.605 146.465 ;
        RECT 73.895 146.295 74.065 146.465 ;
        RECT 74.355 146.295 74.525 146.465 ;
        RECT 74.815 146.295 74.985 146.465 ;
        RECT 75.275 146.295 75.445 146.465 ;
        RECT 75.735 146.295 75.905 146.465 ;
        RECT 76.195 146.295 76.365 146.465 ;
        RECT 76.655 146.295 76.825 146.465 ;
        RECT 77.115 146.295 77.285 146.465 ;
        RECT 77.575 146.295 77.745 146.465 ;
        RECT 78.035 146.295 78.205 146.465 ;
        RECT 78.495 146.295 78.665 146.465 ;
        RECT 78.955 146.295 79.125 146.465 ;
        RECT 79.415 146.295 79.585 146.465 ;
        RECT 79.875 146.295 80.045 146.465 ;
        RECT 80.335 146.295 80.505 146.465 ;
        RECT 80.795 146.295 80.965 146.465 ;
        RECT 81.255 146.295 81.425 146.465 ;
        RECT 81.715 146.295 81.885 146.465 ;
        RECT 82.175 146.295 82.345 146.465 ;
        RECT 82.635 146.295 82.805 146.465 ;
        RECT 83.095 146.295 83.265 146.465 ;
        RECT 83.555 146.295 83.725 146.465 ;
        RECT 84.015 146.295 84.185 146.465 ;
        RECT 84.475 146.295 84.645 146.465 ;
        RECT 84.935 146.295 85.105 146.465 ;
        RECT 85.395 146.295 85.565 146.465 ;
        RECT 85.855 146.295 86.025 146.465 ;
        RECT 86.315 146.295 86.485 146.465 ;
        RECT 86.775 146.295 86.945 146.465 ;
        RECT 87.235 146.295 87.405 146.465 ;
        RECT 87.695 146.295 87.865 146.465 ;
        RECT 88.155 146.295 88.325 146.465 ;
        RECT 88.615 146.295 88.785 146.465 ;
        RECT 89.075 146.295 89.245 146.465 ;
        RECT 89.535 146.295 89.705 146.465 ;
        RECT 89.995 146.295 90.165 146.465 ;
        RECT 90.455 146.295 90.625 146.465 ;
        RECT 90.915 146.295 91.085 146.465 ;
        RECT 91.375 146.295 91.545 146.465 ;
        RECT 91.835 146.295 92.005 146.465 ;
        RECT 92.295 146.295 92.465 146.465 ;
        RECT 92.755 146.295 92.925 146.465 ;
        RECT 93.215 146.295 93.385 146.465 ;
        RECT 93.675 146.295 93.845 146.465 ;
        RECT 94.135 146.295 94.305 146.465 ;
        RECT 94.595 146.295 94.765 146.465 ;
        RECT 95.055 146.295 95.225 146.465 ;
        RECT 95.515 146.295 95.685 146.465 ;
        RECT 95.975 146.295 96.145 146.465 ;
        RECT 96.435 146.295 96.605 146.465 ;
        RECT 96.895 146.295 97.065 146.465 ;
        RECT 97.355 146.295 97.525 146.465 ;
        RECT 97.815 146.295 97.985 146.465 ;
        RECT 98.275 146.295 98.445 146.465 ;
        RECT 98.735 146.295 98.905 146.465 ;
        RECT 99.195 146.295 99.365 146.465 ;
        RECT 99.655 146.295 99.825 146.465 ;
        RECT 100.115 146.295 100.285 146.465 ;
        RECT 100.575 146.295 100.745 146.465 ;
        RECT 101.035 146.295 101.205 146.465 ;
        RECT 101.495 146.295 101.665 146.465 ;
        RECT 101.955 146.295 102.125 146.465 ;
        RECT 102.415 146.295 102.585 146.465 ;
        RECT 102.875 146.295 103.045 146.465 ;
        RECT 103.335 146.295 103.505 146.465 ;
        RECT 103.795 146.295 103.965 146.465 ;
        RECT 104.255 146.295 104.425 146.465 ;
        RECT 104.715 146.295 104.885 146.465 ;
        RECT 105.175 146.295 105.345 146.465 ;
        RECT 105.635 146.295 105.805 146.465 ;
        RECT 106.095 146.295 106.265 146.465 ;
        RECT 106.555 146.295 106.725 146.465 ;
        RECT 107.015 146.295 107.185 146.465 ;
        RECT 107.475 146.295 107.645 146.465 ;
        RECT 107.935 146.295 108.105 146.465 ;
        RECT 108.395 146.295 108.565 146.465 ;
        RECT 108.855 146.295 109.025 146.465 ;
        RECT 109.315 146.295 109.485 146.465 ;
        RECT 109.775 146.295 109.945 146.465 ;
        RECT 110.235 146.295 110.405 146.465 ;
        RECT 110.695 146.295 110.865 146.465 ;
        RECT 111.155 146.295 111.325 146.465 ;
        RECT 111.615 146.295 111.785 146.465 ;
        RECT 112.075 146.295 112.245 146.465 ;
        RECT 112.535 146.295 112.705 146.465 ;
        RECT 112.995 146.295 113.165 146.465 ;
        RECT 113.455 146.295 113.625 146.465 ;
        RECT 113.915 146.295 114.085 146.465 ;
        RECT 114.375 146.295 114.545 146.465 ;
        RECT 114.835 146.295 115.005 146.465 ;
        RECT 115.295 146.295 115.465 146.465 ;
        RECT 115.755 146.295 115.925 146.465 ;
        RECT 116.215 146.295 116.385 146.465 ;
        RECT 116.675 146.295 116.845 146.465 ;
        RECT 117.135 146.295 117.305 146.465 ;
        RECT 117.595 146.295 117.765 146.465 ;
        RECT 118.055 146.295 118.225 146.465 ;
        RECT 118.515 146.295 118.685 146.465 ;
        RECT 118.975 146.295 119.145 146.465 ;
        RECT 119.435 146.295 119.605 146.465 ;
        RECT 119.895 146.295 120.065 146.465 ;
        RECT 120.355 146.295 120.525 146.465 ;
        RECT 120.815 146.295 120.985 146.465 ;
        RECT 121.275 146.295 121.445 146.465 ;
        RECT 121.735 146.295 121.905 146.465 ;
        RECT 122.195 146.295 122.365 146.465 ;
        RECT 122.655 146.295 122.825 146.465 ;
        RECT 123.115 146.295 123.285 146.465 ;
        RECT 123.575 146.295 123.745 146.465 ;
        RECT 124.035 146.295 124.205 146.465 ;
        RECT 124.495 146.295 124.665 146.465 ;
        RECT 124.955 146.295 125.125 146.465 ;
        RECT 125.415 146.295 125.585 146.465 ;
        RECT 125.875 146.295 126.045 146.465 ;
        RECT 126.335 146.295 126.505 146.465 ;
        RECT 126.795 146.295 126.965 146.465 ;
        RECT 127.255 146.295 127.425 146.465 ;
        RECT 127.715 146.295 127.885 146.465 ;
        RECT 128.175 146.295 128.345 146.465 ;
        RECT 128.635 146.295 128.805 146.465 ;
        RECT 129.095 146.295 129.265 146.465 ;
        RECT 129.555 146.295 129.725 146.465 ;
        RECT 130.015 146.295 130.185 146.465 ;
        RECT 130.475 146.295 130.645 146.465 ;
        RECT 130.935 146.295 131.105 146.465 ;
        RECT 57.335 143.575 57.505 143.745 ;
        RECT 57.795 143.575 57.965 143.745 ;
        RECT 58.255 143.575 58.425 143.745 ;
        RECT 58.715 143.575 58.885 143.745 ;
        RECT 59.175 143.575 59.345 143.745 ;
        RECT 59.635 143.575 59.805 143.745 ;
        RECT 60.095 143.575 60.265 143.745 ;
        RECT 60.555 143.575 60.725 143.745 ;
        RECT 61.015 143.575 61.185 143.745 ;
        RECT 61.475 143.575 61.645 143.745 ;
        RECT 61.935 143.575 62.105 143.745 ;
        RECT 62.395 143.575 62.565 143.745 ;
        RECT 62.855 143.575 63.025 143.745 ;
        RECT 63.315 143.575 63.485 143.745 ;
        RECT 63.775 143.575 63.945 143.745 ;
        RECT 64.235 143.575 64.405 143.745 ;
        RECT 64.695 143.575 64.865 143.745 ;
        RECT 65.155 143.575 65.325 143.745 ;
        RECT 65.615 143.575 65.785 143.745 ;
        RECT 66.075 143.575 66.245 143.745 ;
        RECT 66.535 143.575 66.705 143.745 ;
        RECT 66.995 143.575 67.165 143.745 ;
        RECT 67.455 143.575 67.625 143.745 ;
        RECT 67.915 143.575 68.085 143.745 ;
        RECT 68.375 143.575 68.545 143.745 ;
        RECT 68.835 143.575 69.005 143.745 ;
        RECT 69.295 143.575 69.465 143.745 ;
        RECT 69.755 143.575 69.925 143.745 ;
        RECT 70.215 143.575 70.385 143.745 ;
        RECT 70.675 143.575 70.845 143.745 ;
        RECT 71.135 143.575 71.305 143.745 ;
        RECT 71.595 143.575 71.765 143.745 ;
        RECT 72.055 143.575 72.225 143.745 ;
        RECT 72.515 143.575 72.685 143.745 ;
        RECT 72.975 143.575 73.145 143.745 ;
        RECT 73.435 143.575 73.605 143.745 ;
        RECT 73.895 143.575 74.065 143.745 ;
        RECT 74.355 143.575 74.525 143.745 ;
        RECT 74.815 143.575 74.985 143.745 ;
        RECT 75.275 143.575 75.445 143.745 ;
        RECT 75.735 143.575 75.905 143.745 ;
        RECT 76.195 143.575 76.365 143.745 ;
        RECT 76.655 143.575 76.825 143.745 ;
        RECT 77.115 143.575 77.285 143.745 ;
        RECT 77.575 143.575 77.745 143.745 ;
        RECT 78.035 143.575 78.205 143.745 ;
        RECT 78.495 143.575 78.665 143.745 ;
        RECT 78.955 143.575 79.125 143.745 ;
        RECT 79.415 143.575 79.585 143.745 ;
        RECT 79.875 143.575 80.045 143.745 ;
        RECT 80.335 143.575 80.505 143.745 ;
        RECT 80.795 143.575 80.965 143.745 ;
        RECT 81.255 143.575 81.425 143.745 ;
        RECT 81.715 143.575 81.885 143.745 ;
        RECT 82.175 143.575 82.345 143.745 ;
        RECT 82.635 143.575 82.805 143.745 ;
        RECT 83.095 143.575 83.265 143.745 ;
        RECT 83.555 143.575 83.725 143.745 ;
        RECT 84.015 143.575 84.185 143.745 ;
        RECT 84.475 143.575 84.645 143.745 ;
        RECT 84.935 143.575 85.105 143.745 ;
        RECT 85.395 143.575 85.565 143.745 ;
        RECT 85.855 143.575 86.025 143.745 ;
        RECT 86.315 143.575 86.485 143.745 ;
        RECT 86.775 143.575 86.945 143.745 ;
        RECT 87.235 143.575 87.405 143.745 ;
        RECT 87.695 143.575 87.865 143.745 ;
        RECT 88.155 143.575 88.325 143.745 ;
        RECT 88.615 143.575 88.785 143.745 ;
        RECT 89.075 143.575 89.245 143.745 ;
        RECT 89.535 143.575 89.705 143.745 ;
        RECT 89.995 143.575 90.165 143.745 ;
        RECT 90.455 143.575 90.625 143.745 ;
        RECT 90.915 143.575 91.085 143.745 ;
        RECT 91.375 143.575 91.545 143.745 ;
        RECT 91.835 143.575 92.005 143.745 ;
        RECT 92.295 143.575 92.465 143.745 ;
        RECT 92.755 143.575 92.925 143.745 ;
        RECT 93.215 143.575 93.385 143.745 ;
        RECT 93.675 143.575 93.845 143.745 ;
        RECT 94.135 143.575 94.305 143.745 ;
        RECT 94.595 143.575 94.765 143.745 ;
        RECT 95.055 143.575 95.225 143.745 ;
        RECT 95.515 143.575 95.685 143.745 ;
        RECT 95.975 143.575 96.145 143.745 ;
        RECT 96.435 143.575 96.605 143.745 ;
        RECT 96.895 143.575 97.065 143.745 ;
        RECT 97.355 143.575 97.525 143.745 ;
        RECT 97.815 143.575 97.985 143.745 ;
        RECT 98.275 143.575 98.445 143.745 ;
        RECT 98.735 143.575 98.905 143.745 ;
        RECT 99.195 143.575 99.365 143.745 ;
        RECT 99.655 143.575 99.825 143.745 ;
        RECT 100.115 143.575 100.285 143.745 ;
        RECT 100.575 143.575 100.745 143.745 ;
        RECT 101.035 143.575 101.205 143.745 ;
        RECT 101.495 143.575 101.665 143.745 ;
        RECT 101.955 143.575 102.125 143.745 ;
        RECT 102.415 143.575 102.585 143.745 ;
        RECT 102.875 143.575 103.045 143.745 ;
        RECT 103.335 143.575 103.505 143.745 ;
        RECT 103.795 143.575 103.965 143.745 ;
        RECT 104.255 143.575 104.425 143.745 ;
        RECT 104.715 143.575 104.885 143.745 ;
        RECT 105.175 143.575 105.345 143.745 ;
        RECT 105.635 143.575 105.805 143.745 ;
        RECT 106.095 143.575 106.265 143.745 ;
        RECT 106.555 143.575 106.725 143.745 ;
        RECT 107.015 143.575 107.185 143.745 ;
        RECT 107.475 143.575 107.645 143.745 ;
        RECT 107.935 143.575 108.105 143.745 ;
        RECT 108.395 143.575 108.565 143.745 ;
        RECT 108.855 143.575 109.025 143.745 ;
        RECT 109.315 143.575 109.485 143.745 ;
        RECT 109.775 143.575 109.945 143.745 ;
        RECT 110.235 143.575 110.405 143.745 ;
        RECT 110.695 143.575 110.865 143.745 ;
        RECT 111.155 143.575 111.325 143.745 ;
        RECT 111.615 143.575 111.785 143.745 ;
        RECT 112.075 143.575 112.245 143.745 ;
        RECT 112.535 143.575 112.705 143.745 ;
        RECT 112.995 143.575 113.165 143.745 ;
        RECT 113.455 143.575 113.625 143.745 ;
        RECT 113.915 143.575 114.085 143.745 ;
        RECT 114.375 143.575 114.545 143.745 ;
        RECT 114.835 143.575 115.005 143.745 ;
        RECT 115.295 143.575 115.465 143.745 ;
        RECT 115.755 143.575 115.925 143.745 ;
        RECT 116.215 143.575 116.385 143.745 ;
        RECT 116.675 143.575 116.845 143.745 ;
        RECT 117.135 143.575 117.305 143.745 ;
        RECT 117.595 143.575 117.765 143.745 ;
        RECT 118.055 143.575 118.225 143.745 ;
        RECT 118.515 143.575 118.685 143.745 ;
        RECT 118.975 143.575 119.145 143.745 ;
        RECT 119.435 143.575 119.605 143.745 ;
        RECT 119.895 143.575 120.065 143.745 ;
        RECT 120.355 143.575 120.525 143.745 ;
        RECT 120.815 143.575 120.985 143.745 ;
        RECT 121.275 143.575 121.445 143.745 ;
        RECT 121.735 143.575 121.905 143.745 ;
        RECT 122.195 143.575 122.365 143.745 ;
        RECT 122.655 143.575 122.825 143.745 ;
        RECT 123.115 143.575 123.285 143.745 ;
        RECT 123.575 143.575 123.745 143.745 ;
        RECT 124.035 143.575 124.205 143.745 ;
        RECT 124.495 143.575 124.665 143.745 ;
        RECT 124.955 143.575 125.125 143.745 ;
        RECT 125.415 143.575 125.585 143.745 ;
        RECT 125.875 143.575 126.045 143.745 ;
        RECT 126.335 143.575 126.505 143.745 ;
        RECT 126.795 143.575 126.965 143.745 ;
        RECT 127.255 143.575 127.425 143.745 ;
        RECT 127.715 143.575 127.885 143.745 ;
        RECT 128.175 143.575 128.345 143.745 ;
        RECT 128.635 143.575 128.805 143.745 ;
        RECT 129.095 143.575 129.265 143.745 ;
        RECT 129.555 143.575 129.725 143.745 ;
        RECT 130.015 143.575 130.185 143.745 ;
        RECT 130.475 143.575 130.645 143.745 ;
        RECT 130.935 143.575 131.105 143.745 ;
        RECT 57.335 140.855 57.505 141.025 ;
        RECT 57.795 140.855 57.965 141.025 ;
        RECT 58.255 140.855 58.425 141.025 ;
        RECT 58.715 140.855 58.885 141.025 ;
        RECT 59.175 140.855 59.345 141.025 ;
        RECT 59.635 140.855 59.805 141.025 ;
        RECT 60.095 140.855 60.265 141.025 ;
        RECT 60.555 140.855 60.725 141.025 ;
        RECT 61.015 140.855 61.185 141.025 ;
        RECT 61.475 140.855 61.645 141.025 ;
        RECT 61.935 140.855 62.105 141.025 ;
        RECT 62.395 140.855 62.565 141.025 ;
        RECT 62.855 140.855 63.025 141.025 ;
        RECT 63.315 140.855 63.485 141.025 ;
        RECT 63.775 140.855 63.945 141.025 ;
        RECT 64.235 140.855 64.405 141.025 ;
        RECT 64.695 140.855 64.865 141.025 ;
        RECT 65.155 140.855 65.325 141.025 ;
        RECT 65.615 140.855 65.785 141.025 ;
        RECT 66.075 140.855 66.245 141.025 ;
        RECT 66.535 140.855 66.705 141.025 ;
        RECT 66.995 140.855 67.165 141.025 ;
        RECT 67.455 140.855 67.625 141.025 ;
        RECT 67.915 140.855 68.085 141.025 ;
        RECT 68.375 140.855 68.545 141.025 ;
        RECT 68.835 140.855 69.005 141.025 ;
        RECT 69.295 140.855 69.465 141.025 ;
        RECT 69.755 140.855 69.925 141.025 ;
        RECT 70.215 140.855 70.385 141.025 ;
        RECT 70.675 140.855 70.845 141.025 ;
        RECT 71.135 140.855 71.305 141.025 ;
        RECT 71.595 140.855 71.765 141.025 ;
        RECT 72.055 140.855 72.225 141.025 ;
        RECT 72.515 140.855 72.685 141.025 ;
        RECT 72.975 140.855 73.145 141.025 ;
        RECT 73.435 140.855 73.605 141.025 ;
        RECT 73.895 140.855 74.065 141.025 ;
        RECT 74.355 140.855 74.525 141.025 ;
        RECT 74.815 140.855 74.985 141.025 ;
        RECT 75.275 140.855 75.445 141.025 ;
        RECT 75.735 140.855 75.905 141.025 ;
        RECT 76.195 140.855 76.365 141.025 ;
        RECT 76.655 140.855 76.825 141.025 ;
        RECT 77.115 140.855 77.285 141.025 ;
        RECT 77.575 140.855 77.745 141.025 ;
        RECT 78.035 140.855 78.205 141.025 ;
        RECT 78.495 140.855 78.665 141.025 ;
        RECT 78.955 140.855 79.125 141.025 ;
        RECT 79.415 140.855 79.585 141.025 ;
        RECT 79.875 140.855 80.045 141.025 ;
        RECT 80.335 140.855 80.505 141.025 ;
        RECT 80.795 140.855 80.965 141.025 ;
        RECT 81.255 140.855 81.425 141.025 ;
        RECT 81.715 140.855 81.885 141.025 ;
        RECT 82.175 140.855 82.345 141.025 ;
        RECT 82.635 140.855 82.805 141.025 ;
        RECT 83.095 140.855 83.265 141.025 ;
        RECT 83.555 140.855 83.725 141.025 ;
        RECT 84.015 140.855 84.185 141.025 ;
        RECT 84.475 140.855 84.645 141.025 ;
        RECT 84.935 140.855 85.105 141.025 ;
        RECT 85.395 140.855 85.565 141.025 ;
        RECT 85.855 140.855 86.025 141.025 ;
        RECT 86.315 140.855 86.485 141.025 ;
        RECT 86.775 140.855 86.945 141.025 ;
        RECT 87.235 140.855 87.405 141.025 ;
        RECT 87.695 140.855 87.865 141.025 ;
        RECT 88.155 140.855 88.325 141.025 ;
        RECT 88.615 140.855 88.785 141.025 ;
        RECT 89.075 140.855 89.245 141.025 ;
        RECT 89.535 140.855 89.705 141.025 ;
        RECT 89.995 140.855 90.165 141.025 ;
        RECT 90.455 140.855 90.625 141.025 ;
        RECT 90.915 140.855 91.085 141.025 ;
        RECT 91.375 140.855 91.545 141.025 ;
        RECT 91.835 140.855 92.005 141.025 ;
        RECT 92.295 140.855 92.465 141.025 ;
        RECT 92.755 140.855 92.925 141.025 ;
        RECT 93.215 140.855 93.385 141.025 ;
        RECT 93.675 140.855 93.845 141.025 ;
        RECT 94.135 140.855 94.305 141.025 ;
        RECT 94.595 140.855 94.765 141.025 ;
        RECT 95.055 140.855 95.225 141.025 ;
        RECT 95.515 140.855 95.685 141.025 ;
        RECT 95.975 140.855 96.145 141.025 ;
        RECT 96.435 140.855 96.605 141.025 ;
        RECT 96.895 140.855 97.065 141.025 ;
        RECT 97.355 140.855 97.525 141.025 ;
        RECT 97.815 140.855 97.985 141.025 ;
        RECT 98.275 140.855 98.445 141.025 ;
        RECT 98.735 140.855 98.905 141.025 ;
        RECT 99.195 140.855 99.365 141.025 ;
        RECT 99.655 140.855 99.825 141.025 ;
        RECT 100.115 140.855 100.285 141.025 ;
        RECT 100.575 140.855 100.745 141.025 ;
        RECT 101.035 140.855 101.205 141.025 ;
        RECT 101.495 140.855 101.665 141.025 ;
        RECT 101.955 140.855 102.125 141.025 ;
        RECT 102.415 140.855 102.585 141.025 ;
        RECT 102.875 140.855 103.045 141.025 ;
        RECT 103.335 140.855 103.505 141.025 ;
        RECT 103.795 140.855 103.965 141.025 ;
        RECT 104.255 140.855 104.425 141.025 ;
        RECT 104.715 140.855 104.885 141.025 ;
        RECT 105.175 140.855 105.345 141.025 ;
        RECT 105.635 140.855 105.805 141.025 ;
        RECT 106.095 140.855 106.265 141.025 ;
        RECT 106.555 140.855 106.725 141.025 ;
        RECT 107.015 140.855 107.185 141.025 ;
        RECT 107.475 140.855 107.645 141.025 ;
        RECT 107.935 140.855 108.105 141.025 ;
        RECT 108.395 140.855 108.565 141.025 ;
        RECT 108.855 140.855 109.025 141.025 ;
        RECT 109.315 140.855 109.485 141.025 ;
        RECT 109.775 140.855 109.945 141.025 ;
        RECT 110.235 140.855 110.405 141.025 ;
        RECT 110.695 140.855 110.865 141.025 ;
        RECT 111.155 140.855 111.325 141.025 ;
        RECT 111.615 140.855 111.785 141.025 ;
        RECT 112.075 140.855 112.245 141.025 ;
        RECT 112.535 140.855 112.705 141.025 ;
        RECT 112.995 140.855 113.165 141.025 ;
        RECT 113.455 140.855 113.625 141.025 ;
        RECT 113.915 140.855 114.085 141.025 ;
        RECT 114.375 140.855 114.545 141.025 ;
        RECT 114.835 140.855 115.005 141.025 ;
        RECT 115.295 140.855 115.465 141.025 ;
        RECT 115.755 140.855 115.925 141.025 ;
        RECT 116.215 140.855 116.385 141.025 ;
        RECT 116.675 140.855 116.845 141.025 ;
        RECT 117.135 140.855 117.305 141.025 ;
        RECT 117.595 140.855 117.765 141.025 ;
        RECT 118.055 140.855 118.225 141.025 ;
        RECT 118.515 140.855 118.685 141.025 ;
        RECT 118.975 140.855 119.145 141.025 ;
        RECT 119.435 140.855 119.605 141.025 ;
        RECT 119.895 140.855 120.065 141.025 ;
        RECT 120.355 140.855 120.525 141.025 ;
        RECT 120.815 140.855 120.985 141.025 ;
        RECT 121.275 140.855 121.445 141.025 ;
        RECT 121.735 140.855 121.905 141.025 ;
        RECT 122.195 140.855 122.365 141.025 ;
        RECT 122.655 140.855 122.825 141.025 ;
        RECT 123.115 140.855 123.285 141.025 ;
        RECT 123.575 140.855 123.745 141.025 ;
        RECT 124.035 140.855 124.205 141.025 ;
        RECT 124.495 140.855 124.665 141.025 ;
        RECT 124.955 140.855 125.125 141.025 ;
        RECT 125.415 140.855 125.585 141.025 ;
        RECT 125.875 140.855 126.045 141.025 ;
        RECT 126.335 140.855 126.505 141.025 ;
        RECT 126.795 140.855 126.965 141.025 ;
        RECT 127.255 140.855 127.425 141.025 ;
        RECT 127.715 140.855 127.885 141.025 ;
        RECT 128.175 140.855 128.345 141.025 ;
        RECT 128.635 140.855 128.805 141.025 ;
        RECT 129.095 140.855 129.265 141.025 ;
        RECT 129.555 140.855 129.725 141.025 ;
        RECT 130.015 140.855 130.185 141.025 ;
        RECT 130.475 140.855 130.645 141.025 ;
        RECT 130.935 140.855 131.105 141.025 ;
        RECT 57.335 138.135 57.505 138.305 ;
        RECT 57.795 138.135 57.965 138.305 ;
        RECT 58.255 138.135 58.425 138.305 ;
        RECT 58.715 138.135 58.885 138.305 ;
        RECT 59.175 138.135 59.345 138.305 ;
        RECT 59.635 138.135 59.805 138.305 ;
        RECT 60.095 138.135 60.265 138.305 ;
        RECT 60.555 138.135 60.725 138.305 ;
        RECT 61.015 138.135 61.185 138.305 ;
        RECT 61.475 138.135 61.645 138.305 ;
        RECT 61.935 138.135 62.105 138.305 ;
        RECT 62.395 138.135 62.565 138.305 ;
        RECT 62.855 138.135 63.025 138.305 ;
        RECT 63.315 138.135 63.485 138.305 ;
        RECT 63.775 138.135 63.945 138.305 ;
        RECT 64.235 138.135 64.405 138.305 ;
        RECT 64.695 138.135 64.865 138.305 ;
        RECT 65.155 138.135 65.325 138.305 ;
        RECT 65.615 138.135 65.785 138.305 ;
        RECT 66.075 138.135 66.245 138.305 ;
        RECT 66.535 138.135 66.705 138.305 ;
        RECT 66.995 138.135 67.165 138.305 ;
        RECT 67.455 138.135 67.625 138.305 ;
        RECT 67.915 138.135 68.085 138.305 ;
        RECT 68.375 138.135 68.545 138.305 ;
        RECT 68.835 138.135 69.005 138.305 ;
        RECT 69.295 138.135 69.465 138.305 ;
        RECT 69.755 138.135 69.925 138.305 ;
        RECT 70.215 138.135 70.385 138.305 ;
        RECT 70.675 138.135 70.845 138.305 ;
        RECT 71.135 138.135 71.305 138.305 ;
        RECT 71.595 138.135 71.765 138.305 ;
        RECT 72.055 138.135 72.225 138.305 ;
        RECT 72.515 138.135 72.685 138.305 ;
        RECT 72.975 138.135 73.145 138.305 ;
        RECT 73.435 138.135 73.605 138.305 ;
        RECT 73.895 138.135 74.065 138.305 ;
        RECT 74.355 138.135 74.525 138.305 ;
        RECT 74.815 138.135 74.985 138.305 ;
        RECT 75.275 138.135 75.445 138.305 ;
        RECT 75.735 138.135 75.905 138.305 ;
        RECT 76.195 138.135 76.365 138.305 ;
        RECT 76.655 138.135 76.825 138.305 ;
        RECT 77.115 138.135 77.285 138.305 ;
        RECT 77.575 138.135 77.745 138.305 ;
        RECT 78.035 138.135 78.205 138.305 ;
        RECT 78.495 138.135 78.665 138.305 ;
        RECT 78.955 138.135 79.125 138.305 ;
        RECT 79.415 138.135 79.585 138.305 ;
        RECT 79.875 138.135 80.045 138.305 ;
        RECT 80.335 138.135 80.505 138.305 ;
        RECT 80.795 138.135 80.965 138.305 ;
        RECT 81.255 138.135 81.425 138.305 ;
        RECT 81.715 138.135 81.885 138.305 ;
        RECT 82.175 138.135 82.345 138.305 ;
        RECT 82.635 138.135 82.805 138.305 ;
        RECT 83.095 138.135 83.265 138.305 ;
        RECT 83.555 138.135 83.725 138.305 ;
        RECT 84.015 138.135 84.185 138.305 ;
        RECT 84.475 138.135 84.645 138.305 ;
        RECT 84.935 138.135 85.105 138.305 ;
        RECT 85.395 138.135 85.565 138.305 ;
        RECT 85.855 138.135 86.025 138.305 ;
        RECT 86.315 138.135 86.485 138.305 ;
        RECT 86.775 138.135 86.945 138.305 ;
        RECT 87.235 138.135 87.405 138.305 ;
        RECT 87.695 138.135 87.865 138.305 ;
        RECT 88.155 138.135 88.325 138.305 ;
        RECT 88.615 138.135 88.785 138.305 ;
        RECT 89.075 138.135 89.245 138.305 ;
        RECT 89.535 138.135 89.705 138.305 ;
        RECT 89.995 138.135 90.165 138.305 ;
        RECT 90.455 138.135 90.625 138.305 ;
        RECT 90.915 138.135 91.085 138.305 ;
        RECT 91.375 138.135 91.545 138.305 ;
        RECT 91.835 138.135 92.005 138.305 ;
        RECT 92.295 138.135 92.465 138.305 ;
        RECT 92.755 138.135 92.925 138.305 ;
        RECT 93.215 138.135 93.385 138.305 ;
        RECT 93.675 138.135 93.845 138.305 ;
        RECT 94.135 138.135 94.305 138.305 ;
        RECT 94.595 138.135 94.765 138.305 ;
        RECT 95.055 138.135 95.225 138.305 ;
        RECT 95.515 138.135 95.685 138.305 ;
        RECT 95.975 138.135 96.145 138.305 ;
        RECT 96.435 138.135 96.605 138.305 ;
        RECT 96.895 138.135 97.065 138.305 ;
        RECT 97.355 138.135 97.525 138.305 ;
        RECT 97.815 138.135 97.985 138.305 ;
        RECT 98.275 138.135 98.445 138.305 ;
        RECT 98.735 138.135 98.905 138.305 ;
        RECT 99.195 138.135 99.365 138.305 ;
        RECT 99.655 138.135 99.825 138.305 ;
        RECT 100.115 138.135 100.285 138.305 ;
        RECT 100.575 138.135 100.745 138.305 ;
        RECT 101.035 138.135 101.205 138.305 ;
        RECT 101.495 138.135 101.665 138.305 ;
        RECT 101.955 138.135 102.125 138.305 ;
        RECT 102.415 138.135 102.585 138.305 ;
        RECT 102.875 138.135 103.045 138.305 ;
        RECT 103.335 138.135 103.505 138.305 ;
        RECT 103.795 138.135 103.965 138.305 ;
        RECT 104.255 138.135 104.425 138.305 ;
        RECT 104.715 138.135 104.885 138.305 ;
        RECT 105.175 138.135 105.345 138.305 ;
        RECT 105.635 138.135 105.805 138.305 ;
        RECT 106.095 138.135 106.265 138.305 ;
        RECT 106.555 138.135 106.725 138.305 ;
        RECT 107.015 138.135 107.185 138.305 ;
        RECT 107.475 138.135 107.645 138.305 ;
        RECT 107.935 138.135 108.105 138.305 ;
        RECT 108.395 138.135 108.565 138.305 ;
        RECT 108.855 138.135 109.025 138.305 ;
        RECT 109.315 138.135 109.485 138.305 ;
        RECT 109.775 138.135 109.945 138.305 ;
        RECT 110.235 138.135 110.405 138.305 ;
        RECT 110.695 138.135 110.865 138.305 ;
        RECT 111.155 138.135 111.325 138.305 ;
        RECT 111.615 138.135 111.785 138.305 ;
        RECT 112.075 138.135 112.245 138.305 ;
        RECT 112.535 138.135 112.705 138.305 ;
        RECT 112.995 138.135 113.165 138.305 ;
        RECT 113.455 138.135 113.625 138.305 ;
        RECT 113.915 138.135 114.085 138.305 ;
        RECT 114.375 138.135 114.545 138.305 ;
        RECT 114.835 138.135 115.005 138.305 ;
        RECT 115.295 138.135 115.465 138.305 ;
        RECT 115.755 138.135 115.925 138.305 ;
        RECT 116.215 138.135 116.385 138.305 ;
        RECT 116.675 138.135 116.845 138.305 ;
        RECT 117.135 138.135 117.305 138.305 ;
        RECT 117.595 138.135 117.765 138.305 ;
        RECT 118.055 138.135 118.225 138.305 ;
        RECT 118.515 138.135 118.685 138.305 ;
        RECT 118.975 138.135 119.145 138.305 ;
        RECT 119.435 138.135 119.605 138.305 ;
        RECT 119.895 138.135 120.065 138.305 ;
        RECT 120.355 138.135 120.525 138.305 ;
        RECT 120.815 138.135 120.985 138.305 ;
        RECT 121.275 138.135 121.445 138.305 ;
        RECT 121.735 138.135 121.905 138.305 ;
        RECT 122.195 138.135 122.365 138.305 ;
        RECT 122.655 138.135 122.825 138.305 ;
        RECT 123.115 138.135 123.285 138.305 ;
        RECT 123.575 138.135 123.745 138.305 ;
        RECT 124.035 138.135 124.205 138.305 ;
        RECT 124.495 138.135 124.665 138.305 ;
        RECT 124.955 138.135 125.125 138.305 ;
        RECT 125.415 138.135 125.585 138.305 ;
        RECT 125.875 138.135 126.045 138.305 ;
        RECT 126.335 138.135 126.505 138.305 ;
        RECT 126.795 138.135 126.965 138.305 ;
        RECT 127.255 138.135 127.425 138.305 ;
        RECT 127.715 138.135 127.885 138.305 ;
        RECT 128.175 138.135 128.345 138.305 ;
        RECT 128.635 138.135 128.805 138.305 ;
        RECT 129.095 138.135 129.265 138.305 ;
        RECT 129.555 138.135 129.725 138.305 ;
        RECT 130.015 138.135 130.185 138.305 ;
        RECT 130.475 138.135 130.645 138.305 ;
        RECT 130.935 138.135 131.105 138.305 ;
        RECT 57.335 135.415 57.505 135.585 ;
        RECT 57.795 135.415 57.965 135.585 ;
        RECT 58.255 135.415 58.425 135.585 ;
        RECT 58.715 135.415 58.885 135.585 ;
        RECT 59.175 135.415 59.345 135.585 ;
        RECT 59.635 135.415 59.805 135.585 ;
        RECT 60.095 135.415 60.265 135.585 ;
        RECT 60.555 135.415 60.725 135.585 ;
        RECT 61.015 135.415 61.185 135.585 ;
        RECT 61.475 135.415 61.645 135.585 ;
        RECT 61.935 135.415 62.105 135.585 ;
        RECT 62.395 135.415 62.565 135.585 ;
        RECT 62.855 135.415 63.025 135.585 ;
        RECT 63.315 135.415 63.485 135.585 ;
        RECT 63.775 135.415 63.945 135.585 ;
        RECT 64.235 135.415 64.405 135.585 ;
        RECT 64.695 135.415 64.865 135.585 ;
        RECT 65.155 135.415 65.325 135.585 ;
        RECT 65.615 135.415 65.785 135.585 ;
        RECT 66.075 135.415 66.245 135.585 ;
        RECT 66.535 135.415 66.705 135.585 ;
        RECT 66.995 135.415 67.165 135.585 ;
        RECT 67.455 135.415 67.625 135.585 ;
        RECT 67.915 135.415 68.085 135.585 ;
        RECT 68.375 135.415 68.545 135.585 ;
        RECT 68.835 135.415 69.005 135.585 ;
        RECT 69.295 135.415 69.465 135.585 ;
        RECT 69.755 135.415 69.925 135.585 ;
        RECT 70.215 135.415 70.385 135.585 ;
        RECT 70.675 135.415 70.845 135.585 ;
        RECT 71.135 135.415 71.305 135.585 ;
        RECT 71.595 135.415 71.765 135.585 ;
        RECT 72.055 135.415 72.225 135.585 ;
        RECT 72.515 135.415 72.685 135.585 ;
        RECT 72.975 135.415 73.145 135.585 ;
        RECT 73.435 135.415 73.605 135.585 ;
        RECT 73.895 135.415 74.065 135.585 ;
        RECT 74.355 135.415 74.525 135.585 ;
        RECT 74.815 135.415 74.985 135.585 ;
        RECT 75.275 135.415 75.445 135.585 ;
        RECT 75.735 135.415 75.905 135.585 ;
        RECT 76.195 135.415 76.365 135.585 ;
        RECT 76.655 135.415 76.825 135.585 ;
        RECT 77.115 135.415 77.285 135.585 ;
        RECT 77.575 135.415 77.745 135.585 ;
        RECT 78.035 135.415 78.205 135.585 ;
        RECT 78.495 135.415 78.665 135.585 ;
        RECT 78.955 135.415 79.125 135.585 ;
        RECT 79.415 135.415 79.585 135.585 ;
        RECT 79.875 135.415 80.045 135.585 ;
        RECT 80.335 135.415 80.505 135.585 ;
        RECT 80.795 135.415 80.965 135.585 ;
        RECT 81.255 135.415 81.425 135.585 ;
        RECT 81.715 135.415 81.885 135.585 ;
        RECT 82.175 135.415 82.345 135.585 ;
        RECT 82.635 135.415 82.805 135.585 ;
        RECT 83.095 135.415 83.265 135.585 ;
        RECT 83.555 135.415 83.725 135.585 ;
        RECT 84.015 135.415 84.185 135.585 ;
        RECT 84.475 135.415 84.645 135.585 ;
        RECT 84.935 135.415 85.105 135.585 ;
        RECT 85.395 135.415 85.565 135.585 ;
        RECT 85.855 135.415 86.025 135.585 ;
        RECT 86.315 135.415 86.485 135.585 ;
        RECT 86.775 135.415 86.945 135.585 ;
        RECT 87.235 135.415 87.405 135.585 ;
        RECT 87.695 135.415 87.865 135.585 ;
        RECT 88.155 135.415 88.325 135.585 ;
        RECT 88.615 135.415 88.785 135.585 ;
        RECT 89.075 135.415 89.245 135.585 ;
        RECT 89.535 135.415 89.705 135.585 ;
        RECT 89.995 135.415 90.165 135.585 ;
        RECT 90.455 135.415 90.625 135.585 ;
        RECT 90.915 135.415 91.085 135.585 ;
        RECT 91.375 135.415 91.545 135.585 ;
        RECT 91.835 135.415 92.005 135.585 ;
        RECT 92.295 135.415 92.465 135.585 ;
        RECT 92.755 135.415 92.925 135.585 ;
        RECT 93.215 135.415 93.385 135.585 ;
        RECT 93.675 135.415 93.845 135.585 ;
        RECT 94.135 135.415 94.305 135.585 ;
        RECT 94.595 135.415 94.765 135.585 ;
        RECT 95.055 135.415 95.225 135.585 ;
        RECT 95.515 135.415 95.685 135.585 ;
        RECT 95.975 135.415 96.145 135.585 ;
        RECT 96.435 135.415 96.605 135.585 ;
        RECT 96.895 135.415 97.065 135.585 ;
        RECT 97.355 135.415 97.525 135.585 ;
        RECT 97.815 135.415 97.985 135.585 ;
        RECT 98.275 135.415 98.445 135.585 ;
        RECT 98.735 135.415 98.905 135.585 ;
        RECT 99.195 135.415 99.365 135.585 ;
        RECT 99.655 135.415 99.825 135.585 ;
        RECT 100.115 135.415 100.285 135.585 ;
        RECT 100.575 135.415 100.745 135.585 ;
        RECT 101.035 135.415 101.205 135.585 ;
        RECT 101.495 135.415 101.665 135.585 ;
        RECT 101.955 135.415 102.125 135.585 ;
        RECT 102.415 135.415 102.585 135.585 ;
        RECT 102.875 135.415 103.045 135.585 ;
        RECT 103.335 135.415 103.505 135.585 ;
        RECT 103.795 135.415 103.965 135.585 ;
        RECT 104.255 135.415 104.425 135.585 ;
        RECT 104.715 135.415 104.885 135.585 ;
        RECT 105.175 135.415 105.345 135.585 ;
        RECT 105.635 135.415 105.805 135.585 ;
        RECT 106.095 135.415 106.265 135.585 ;
        RECT 106.555 135.415 106.725 135.585 ;
        RECT 107.015 135.415 107.185 135.585 ;
        RECT 107.475 135.415 107.645 135.585 ;
        RECT 107.935 135.415 108.105 135.585 ;
        RECT 108.395 135.415 108.565 135.585 ;
        RECT 108.855 135.415 109.025 135.585 ;
        RECT 109.315 135.415 109.485 135.585 ;
        RECT 109.775 135.415 109.945 135.585 ;
        RECT 110.235 135.415 110.405 135.585 ;
        RECT 110.695 135.415 110.865 135.585 ;
        RECT 111.155 135.415 111.325 135.585 ;
        RECT 111.615 135.415 111.785 135.585 ;
        RECT 112.075 135.415 112.245 135.585 ;
        RECT 112.535 135.415 112.705 135.585 ;
        RECT 112.995 135.415 113.165 135.585 ;
        RECT 113.455 135.415 113.625 135.585 ;
        RECT 113.915 135.415 114.085 135.585 ;
        RECT 114.375 135.415 114.545 135.585 ;
        RECT 114.835 135.415 115.005 135.585 ;
        RECT 115.295 135.415 115.465 135.585 ;
        RECT 115.755 135.415 115.925 135.585 ;
        RECT 116.215 135.415 116.385 135.585 ;
        RECT 116.675 135.415 116.845 135.585 ;
        RECT 117.135 135.415 117.305 135.585 ;
        RECT 117.595 135.415 117.765 135.585 ;
        RECT 118.055 135.415 118.225 135.585 ;
        RECT 118.515 135.415 118.685 135.585 ;
        RECT 118.975 135.415 119.145 135.585 ;
        RECT 119.435 135.415 119.605 135.585 ;
        RECT 119.895 135.415 120.065 135.585 ;
        RECT 120.355 135.415 120.525 135.585 ;
        RECT 120.815 135.415 120.985 135.585 ;
        RECT 121.275 135.415 121.445 135.585 ;
        RECT 121.735 135.415 121.905 135.585 ;
        RECT 122.195 135.415 122.365 135.585 ;
        RECT 122.655 135.415 122.825 135.585 ;
        RECT 123.115 135.415 123.285 135.585 ;
        RECT 123.575 135.415 123.745 135.585 ;
        RECT 124.035 135.415 124.205 135.585 ;
        RECT 124.495 135.415 124.665 135.585 ;
        RECT 124.955 135.415 125.125 135.585 ;
        RECT 125.415 135.415 125.585 135.585 ;
        RECT 125.875 135.415 126.045 135.585 ;
        RECT 126.335 135.415 126.505 135.585 ;
        RECT 126.795 135.415 126.965 135.585 ;
        RECT 127.255 135.415 127.425 135.585 ;
        RECT 127.715 135.415 127.885 135.585 ;
        RECT 128.175 135.415 128.345 135.585 ;
        RECT 128.635 135.415 128.805 135.585 ;
        RECT 129.095 135.415 129.265 135.585 ;
        RECT 129.555 135.415 129.725 135.585 ;
        RECT 130.015 135.415 130.185 135.585 ;
        RECT 130.475 135.415 130.645 135.585 ;
        RECT 130.935 135.415 131.105 135.585 ;
        RECT 57.335 132.695 57.505 132.865 ;
        RECT 57.795 132.695 57.965 132.865 ;
        RECT 58.255 132.695 58.425 132.865 ;
        RECT 58.715 132.695 58.885 132.865 ;
        RECT 59.175 132.695 59.345 132.865 ;
        RECT 59.635 132.695 59.805 132.865 ;
        RECT 60.095 132.695 60.265 132.865 ;
        RECT 60.555 132.695 60.725 132.865 ;
        RECT 61.015 132.695 61.185 132.865 ;
        RECT 61.475 132.695 61.645 132.865 ;
        RECT 61.935 132.695 62.105 132.865 ;
        RECT 62.395 132.695 62.565 132.865 ;
        RECT 62.855 132.695 63.025 132.865 ;
        RECT 63.315 132.695 63.485 132.865 ;
        RECT 63.775 132.695 63.945 132.865 ;
        RECT 64.235 132.695 64.405 132.865 ;
        RECT 64.695 132.695 64.865 132.865 ;
        RECT 65.155 132.695 65.325 132.865 ;
        RECT 65.615 132.695 65.785 132.865 ;
        RECT 66.075 132.695 66.245 132.865 ;
        RECT 66.535 132.695 66.705 132.865 ;
        RECT 66.995 132.695 67.165 132.865 ;
        RECT 67.455 132.695 67.625 132.865 ;
        RECT 67.915 132.695 68.085 132.865 ;
        RECT 68.375 132.695 68.545 132.865 ;
        RECT 68.835 132.695 69.005 132.865 ;
        RECT 69.295 132.695 69.465 132.865 ;
        RECT 69.755 132.695 69.925 132.865 ;
        RECT 70.215 132.695 70.385 132.865 ;
        RECT 70.675 132.695 70.845 132.865 ;
        RECT 71.135 132.695 71.305 132.865 ;
        RECT 71.595 132.695 71.765 132.865 ;
        RECT 72.055 132.695 72.225 132.865 ;
        RECT 72.515 132.695 72.685 132.865 ;
        RECT 72.975 132.695 73.145 132.865 ;
        RECT 73.435 132.695 73.605 132.865 ;
        RECT 73.895 132.695 74.065 132.865 ;
        RECT 74.355 132.695 74.525 132.865 ;
        RECT 74.815 132.695 74.985 132.865 ;
        RECT 75.275 132.695 75.445 132.865 ;
        RECT 75.735 132.695 75.905 132.865 ;
        RECT 76.195 132.695 76.365 132.865 ;
        RECT 76.655 132.695 76.825 132.865 ;
        RECT 77.115 132.695 77.285 132.865 ;
        RECT 77.575 132.695 77.745 132.865 ;
        RECT 78.035 132.695 78.205 132.865 ;
        RECT 78.495 132.695 78.665 132.865 ;
        RECT 78.955 132.695 79.125 132.865 ;
        RECT 79.415 132.695 79.585 132.865 ;
        RECT 79.875 132.695 80.045 132.865 ;
        RECT 80.335 132.695 80.505 132.865 ;
        RECT 80.795 132.695 80.965 132.865 ;
        RECT 81.255 132.695 81.425 132.865 ;
        RECT 81.715 132.695 81.885 132.865 ;
        RECT 82.175 132.695 82.345 132.865 ;
        RECT 82.635 132.695 82.805 132.865 ;
        RECT 83.095 132.695 83.265 132.865 ;
        RECT 83.555 132.695 83.725 132.865 ;
        RECT 84.015 132.695 84.185 132.865 ;
        RECT 84.475 132.695 84.645 132.865 ;
        RECT 84.935 132.695 85.105 132.865 ;
        RECT 85.395 132.695 85.565 132.865 ;
        RECT 85.855 132.695 86.025 132.865 ;
        RECT 86.315 132.695 86.485 132.865 ;
        RECT 86.775 132.695 86.945 132.865 ;
        RECT 87.235 132.695 87.405 132.865 ;
        RECT 87.695 132.695 87.865 132.865 ;
        RECT 88.155 132.695 88.325 132.865 ;
        RECT 88.615 132.695 88.785 132.865 ;
        RECT 89.075 132.695 89.245 132.865 ;
        RECT 89.535 132.695 89.705 132.865 ;
        RECT 89.995 132.695 90.165 132.865 ;
        RECT 90.455 132.695 90.625 132.865 ;
        RECT 90.915 132.695 91.085 132.865 ;
        RECT 91.375 132.695 91.545 132.865 ;
        RECT 91.835 132.695 92.005 132.865 ;
        RECT 92.295 132.695 92.465 132.865 ;
        RECT 92.755 132.695 92.925 132.865 ;
        RECT 93.215 132.695 93.385 132.865 ;
        RECT 93.675 132.695 93.845 132.865 ;
        RECT 94.135 132.695 94.305 132.865 ;
        RECT 94.595 132.695 94.765 132.865 ;
        RECT 95.055 132.695 95.225 132.865 ;
        RECT 95.515 132.695 95.685 132.865 ;
        RECT 95.975 132.695 96.145 132.865 ;
        RECT 96.435 132.695 96.605 132.865 ;
        RECT 96.895 132.695 97.065 132.865 ;
        RECT 97.355 132.695 97.525 132.865 ;
        RECT 97.815 132.695 97.985 132.865 ;
        RECT 98.275 132.695 98.445 132.865 ;
        RECT 98.735 132.695 98.905 132.865 ;
        RECT 99.195 132.695 99.365 132.865 ;
        RECT 99.655 132.695 99.825 132.865 ;
        RECT 100.115 132.695 100.285 132.865 ;
        RECT 100.575 132.695 100.745 132.865 ;
        RECT 101.035 132.695 101.205 132.865 ;
        RECT 101.495 132.695 101.665 132.865 ;
        RECT 101.955 132.695 102.125 132.865 ;
        RECT 102.415 132.695 102.585 132.865 ;
        RECT 102.875 132.695 103.045 132.865 ;
        RECT 103.335 132.695 103.505 132.865 ;
        RECT 103.795 132.695 103.965 132.865 ;
        RECT 104.255 132.695 104.425 132.865 ;
        RECT 104.715 132.695 104.885 132.865 ;
        RECT 105.175 132.695 105.345 132.865 ;
        RECT 105.635 132.695 105.805 132.865 ;
        RECT 106.095 132.695 106.265 132.865 ;
        RECT 106.555 132.695 106.725 132.865 ;
        RECT 107.015 132.695 107.185 132.865 ;
        RECT 107.475 132.695 107.645 132.865 ;
        RECT 107.935 132.695 108.105 132.865 ;
        RECT 108.395 132.695 108.565 132.865 ;
        RECT 108.855 132.695 109.025 132.865 ;
        RECT 109.315 132.695 109.485 132.865 ;
        RECT 109.775 132.695 109.945 132.865 ;
        RECT 110.235 132.695 110.405 132.865 ;
        RECT 110.695 132.695 110.865 132.865 ;
        RECT 111.155 132.695 111.325 132.865 ;
        RECT 111.615 132.695 111.785 132.865 ;
        RECT 112.075 132.695 112.245 132.865 ;
        RECT 112.535 132.695 112.705 132.865 ;
        RECT 112.995 132.695 113.165 132.865 ;
        RECT 113.455 132.695 113.625 132.865 ;
        RECT 113.915 132.695 114.085 132.865 ;
        RECT 114.375 132.695 114.545 132.865 ;
        RECT 114.835 132.695 115.005 132.865 ;
        RECT 115.295 132.695 115.465 132.865 ;
        RECT 115.755 132.695 115.925 132.865 ;
        RECT 116.215 132.695 116.385 132.865 ;
        RECT 116.675 132.695 116.845 132.865 ;
        RECT 117.135 132.695 117.305 132.865 ;
        RECT 117.595 132.695 117.765 132.865 ;
        RECT 118.055 132.695 118.225 132.865 ;
        RECT 118.515 132.695 118.685 132.865 ;
        RECT 118.975 132.695 119.145 132.865 ;
        RECT 119.435 132.695 119.605 132.865 ;
        RECT 119.895 132.695 120.065 132.865 ;
        RECT 120.355 132.695 120.525 132.865 ;
        RECT 120.815 132.695 120.985 132.865 ;
        RECT 121.275 132.695 121.445 132.865 ;
        RECT 121.735 132.695 121.905 132.865 ;
        RECT 122.195 132.695 122.365 132.865 ;
        RECT 122.655 132.695 122.825 132.865 ;
        RECT 123.115 132.695 123.285 132.865 ;
        RECT 123.575 132.695 123.745 132.865 ;
        RECT 124.035 132.695 124.205 132.865 ;
        RECT 124.495 132.695 124.665 132.865 ;
        RECT 124.955 132.695 125.125 132.865 ;
        RECT 125.415 132.695 125.585 132.865 ;
        RECT 125.875 132.695 126.045 132.865 ;
        RECT 126.335 132.695 126.505 132.865 ;
        RECT 126.795 132.695 126.965 132.865 ;
        RECT 127.255 132.695 127.425 132.865 ;
        RECT 127.715 132.695 127.885 132.865 ;
        RECT 128.175 132.695 128.345 132.865 ;
        RECT 128.635 132.695 128.805 132.865 ;
        RECT 129.095 132.695 129.265 132.865 ;
        RECT 129.555 132.695 129.725 132.865 ;
        RECT 130.015 132.695 130.185 132.865 ;
        RECT 130.475 132.695 130.645 132.865 ;
        RECT 130.935 132.695 131.105 132.865 ;
        RECT 57.335 129.975 57.505 130.145 ;
        RECT 57.795 129.975 57.965 130.145 ;
        RECT 58.255 129.975 58.425 130.145 ;
        RECT 58.715 129.975 58.885 130.145 ;
        RECT 59.175 129.975 59.345 130.145 ;
        RECT 59.635 129.975 59.805 130.145 ;
        RECT 60.095 129.975 60.265 130.145 ;
        RECT 60.555 129.975 60.725 130.145 ;
        RECT 61.015 129.975 61.185 130.145 ;
        RECT 61.475 129.975 61.645 130.145 ;
        RECT 61.935 129.975 62.105 130.145 ;
        RECT 62.395 129.975 62.565 130.145 ;
        RECT 62.855 129.975 63.025 130.145 ;
        RECT 63.315 129.975 63.485 130.145 ;
        RECT 63.775 129.975 63.945 130.145 ;
        RECT 64.235 129.975 64.405 130.145 ;
        RECT 64.695 129.975 64.865 130.145 ;
        RECT 65.155 129.975 65.325 130.145 ;
        RECT 65.615 129.975 65.785 130.145 ;
        RECT 66.075 129.975 66.245 130.145 ;
        RECT 66.535 129.975 66.705 130.145 ;
        RECT 66.995 129.975 67.165 130.145 ;
        RECT 67.455 129.975 67.625 130.145 ;
        RECT 67.915 129.975 68.085 130.145 ;
        RECT 68.375 129.975 68.545 130.145 ;
        RECT 68.835 129.975 69.005 130.145 ;
        RECT 69.295 129.975 69.465 130.145 ;
        RECT 69.755 129.975 69.925 130.145 ;
        RECT 70.215 129.975 70.385 130.145 ;
        RECT 70.675 129.975 70.845 130.145 ;
        RECT 71.135 129.975 71.305 130.145 ;
        RECT 71.595 129.975 71.765 130.145 ;
        RECT 72.055 129.975 72.225 130.145 ;
        RECT 72.515 129.975 72.685 130.145 ;
        RECT 72.975 129.975 73.145 130.145 ;
        RECT 73.435 129.975 73.605 130.145 ;
        RECT 73.895 129.975 74.065 130.145 ;
        RECT 74.355 129.975 74.525 130.145 ;
        RECT 74.815 129.975 74.985 130.145 ;
        RECT 75.275 129.975 75.445 130.145 ;
        RECT 75.735 129.975 75.905 130.145 ;
        RECT 76.195 129.975 76.365 130.145 ;
        RECT 76.655 129.975 76.825 130.145 ;
        RECT 77.115 129.975 77.285 130.145 ;
        RECT 77.575 129.975 77.745 130.145 ;
        RECT 78.035 129.975 78.205 130.145 ;
        RECT 78.495 129.975 78.665 130.145 ;
        RECT 78.955 129.975 79.125 130.145 ;
        RECT 79.415 129.975 79.585 130.145 ;
        RECT 79.875 129.975 80.045 130.145 ;
        RECT 80.335 129.975 80.505 130.145 ;
        RECT 80.795 129.975 80.965 130.145 ;
        RECT 81.255 129.975 81.425 130.145 ;
        RECT 81.715 129.975 81.885 130.145 ;
        RECT 82.175 129.975 82.345 130.145 ;
        RECT 82.635 129.975 82.805 130.145 ;
        RECT 83.095 129.975 83.265 130.145 ;
        RECT 83.555 129.975 83.725 130.145 ;
        RECT 84.015 129.975 84.185 130.145 ;
        RECT 84.475 129.975 84.645 130.145 ;
        RECT 84.935 129.975 85.105 130.145 ;
        RECT 85.395 129.975 85.565 130.145 ;
        RECT 85.855 129.975 86.025 130.145 ;
        RECT 86.315 129.975 86.485 130.145 ;
        RECT 86.775 129.975 86.945 130.145 ;
        RECT 87.235 129.975 87.405 130.145 ;
        RECT 87.695 129.975 87.865 130.145 ;
        RECT 88.155 129.975 88.325 130.145 ;
        RECT 88.615 129.975 88.785 130.145 ;
        RECT 89.075 129.975 89.245 130.145 ;
        RECT 89.535 129.975 89.705 130.145 ;
        RECT 89.995 129.975 90.165 130.145 ;
        RECT 90.455 129.975 90.625 130.145 ;
        RECT 90.915 129.975 91.085 130.145 ;
        RECT 91.375 129.975 91.545 130.145 ;
        RECT 91.835 129.975 92.005 130.145 ;
        RECT 92.295 129.975 92.465 130.145 ;
        RECT 92.755 129.975 92.925 130.145 ;
        RECT 93.215 129.975 93.385 130.145 ;
        RECT 93.675 129.975 93.845 130.145 ;
        RECT 94.135 129.975 94.305 130.145 ;
        RECT 94.595 129.975 94.765 130.145 ;
        RECT 95.055 129.975 95.225 130.145 ;
        RECT 95.515 129.975 95.685 130.145 ;
        RECT 95.975 129.975 96.145 130.145 ;
        RECT 96.435 129.975 96.605 130.145 ;
        RECT 96.895 129.975 97.065 130.145 ;
        RECT 97.355 129.975 97.525 130.145 ;
        RECT 97.815 129.975 97.985 130.145 ;
        RECT 98.275 129.975 98.445 130.145 ;
        RECT 98.735 129.975 98.905 130.145 ;
        RECT 99.195 129.975 99.365 130.145 ;
        RECT 99.655 129.975 99.825 130.145 ;
        RECT 100.115 129.975 100.285 130.145 ;
        RECT 100.575 129.975 100.745 130.145 ;
        RECT 101.035 129.975 101.205 130.145 ;
        RECT 101.495 129.975 101.665 130.145 ;
        RECT 101.955 129.975 102.125 130.145 ;
        RECT 102.415 129.975 102.585 130.145 ;
        RECT 102.875 129.975 103.045 130.145 ;
        RECT 103.335 129.975 103.505 130.145 ;
        RECT 103.795 129.975 103.965 130.145 ;
        RECT 104.255 129.975 104.425 130.145 ;
        RECT 104.715 129.975 104.885 130.145 ;
        RECT 105.175 129.975 105.345 130.145 ;
        RECT 105.635 129.975 105.805 130.145 ;
        RECT 106.095 129.975 106.265 130.145 ;
        RECT 106.555 129.975 106.725 130.145 ;
        RECT 107.015 129.975 107.185 130.145 ;
        RECT 107.475 129.975 107.645 130.145 ;
        RECT 107.935 129.975 108.105 130.145 ;
        RECT 108.395 129.975 108.565 130.145 ;
        RECT 108.855 129.975 109.025 130.145 ;
        RECT 109.315 129.975 109.485 130.145 ;
        RECT 109.775 129.975 109.945 130.145 ;
        RECT 110.235 129.975 110.405 130.145 ;
        RECT 110.695 129.975 110.865 130.145 ;
        RECT 111.155 129.975 111.325 130.145 ;
        RECT 111.615 129.975 111.785 130.145 ;
        RECT 112.075 129.975 112.245 130.145 ;
        RECT 112.535 129.975 112.705 130.145 ;
        RECT 112.995 129.975 113.165 130.145 ;
        RECT 113.455 129.975 113.625 130.145 ;
        RECT 113.915 129.975 114.085 130.145 ;
        RECT 114.375 129.975 114.545 130.145 ;
        RECT 114.835 129.975 115.005 130.145 ;
        RECT 115.295 129.975 115.465 130.145 ;
        RECT 115.755 129.975 115.925 130.145 ;
        RECT 116.215 129.975 116.385 130.145 ;
        RECT 116.675 129.975 116.845 130.145 ;
        RECT 117.135 129.975 117.305 130.145 ;
        RECT 117.595 129.975 117.765 130.145 ;
        RECT 118.055 129.975 118.225 130.145 ;
        RECT 118.515 129.975 118.685 130.145 ;
        RECT 118.975 129.975 119.145 130.145 ;
        RECT 119.435 129.975 119.605 130.145 ;
        RECT 119.895 129.975 120.065 130.145 ;
        RECT 120.355 129.975 120.525 130.145 ;
        RECT 120.815 129.975 120.985 130.145 ;
        RECT 121.275 129.975 121.445 130.145 ;
        RECT 121.735 129.975 121.905 130.145 ;
        RECT 122.195 129.975 122.365 130.145 ;
        RECT 122.655 129.975 122.825 130.145 ;
        RECT 123.115 129.975 123.285 130.145 ;
        RECT 123.575 129.975 123.745 130.145 ;
        RECT 124.035 129.975 124.205 130.145 ;
        RECT 124.495 129.975 124.665 130.145 ;
        RECT 124.955 129.975 125.125 130.145 ;
        RECT 125.415 129.975 125.585 130.145 ;
        RECT 125.875 129.975 126.045 130.145 ;
        RECT 126.335 129.975 126.505 130.145 ;
        RECT 126.795 129.975 126.965 130.145 ;
        RECT 127.255 129.975 127.425 130.145 ;
        RECT 127.715 129.975 127.885 130.145 ;
        RECT 128.175 129.975 128.345 130.145 ;
        RECT 128.635 129.975 128.805 130.145 ;
        RECT 129.095 129.975 129.265 130.145 ;
        RECT 129.555 129.975 129.725 130.145 ;
        RECT 130.015 129.975 130.185 130.145 ;
        RECT 130.475 129.975 130.645 130.145 ;
        RECT 130.935 129.975 131.105 130.145 ;
        RECT 138.040 87.480 140.025 87.670 ;
        RECT 141.385 87.480 143.370 87.670 ;
        RECT 148.040 87.480 150.025 87.670 ;
        RECT 151.385 87.480 153.370 87.670 ;
        RECT 138.870 84.170 140.420 84.370 ;
        RECT 139.180 83.610 139.400 83.780 ;
        RECT 139.850 83.610 140.070 83.780 ;
        RECT 138.870 81.680 139.040 83.360 ;
        RECT 139.540 81.680 139.710 83.360 ;
        RECT 140.210 81.680 140.380 83.360 ;
        RECT 139.180 81.260 139.400 81.430 ;
        RECT 139.850 81.260 140.070 81.430 ;
        RECT 142.870 84.170 144.420 84.370 ;
        RECT 143.180 83.610 143.400 83.780 ;
        RECT 143.850 83.610 144.070 83.780 ;
        RECT 142.870 81.680 143.040 83.360 ;
        RECT 143.540 81.680 143.710 83.360 ;
        RECT 144.210 81.680 144.380 83.360 ;
        RECT 143.180 81.260 143.400 81.430 ;
        RECT 143.850 81.260 144.070 81.430 ;
        RECT 148.180 83.610 148.400 83.780 ;
        RECT 148.850 83.610 149.070 83.780 ;
        RECT 147.870 81.680 148.040 83.360 ;
        RECT 148.540 81.680 148.710 83.360 ;
        RECT 149.210 81.680 149.380 83.360 ;
        RECT 148.180 81.260 148.400 81.430 ;
        RECT 148.850 81.260 149.070 81.430 ;
        RECT 152.180 83.610 152.400 83.780 ;
        RECT 152.850 83.610 153.070 83.780 ;
        RECT 151.870 81.680 152.040 83.360 ;
        RECT 152.540 81.680 152.710 83.360 ;
        RECT 153.210 81.680 153.380 83.360 ;
        RECT 152.180 81.260 152.400 81.430 ;
        RECT 152.850 81.260 153.070 81.430 ;
        RECT 141.180 77.610 141.400 77.780 ;
        RECT 141.850 77.610 142.070 77.780 ;
        RECT 140.870 75.680 141.040 77.360 ;
        RECT 141.540 75.680 141.710 77.360 ;
        RECT 142.210 75.680 142.380 77.360 ;
        RECT 142.770 76.920 143.070 77.720 ;
        RECT 149.220 76.920 149.470 77.720 ;
        RECT 150.180 77.610 150.400 77.780 ;
        RECT 150.850 77.610 151.070 77.780 ;
        RECT 141.180 75.260 141.400 75.430 ;
        RECT 141.850 75.260 142.070 75.430 ;
        RECT 146.020 74.920 146.220 75.120 ;
        RECT 149.870 75.680 150.040 77.360 ;
        RECT 150.540 75.680 150.710 77.360 ;
        RECT 151.210 75.680 151.380 77.360 ;
        RECT 150.180 75.260 150.400 75.430 ;
        RECT 150.850 75.260 151.070 75.430 ;
        RECT 146.020 73.670 146.220 73.870 ;
      LAYER met1 ;
        RECT 57.190 203.260 131.250 203.740 ;
        RECT 101.420 203.060 101.740 203.120 ;
        RECT 101.420 202.920 110.850 203.060 ;
        RECT 101.420 202.860 101.740 202.920 ;
        RECT 76.135 202.720 76.425 202.765 ;
        RECT 91.315 202.720 91.605 202.765 ;
        RECT 76.135 202.580 78.190 202.720 ;
        RECT 76.135 202.535 76.425 202.580 ;
        RECT 71.995 202.380 72.285 202.425 ;
        RECT 75.215 202.380 75.505 202.425 ;
        RECT 71.995 202.240 77.270 202.380 ;
        RECT 71.995 202.195 72.285 202.240 ;
        RECT 75.215 202.195 75.505 202.240 ;
        RECT 60.480 202.040 60.800 202.100 ;
        RECT 60.955 202.040 61.245 202.085 ;
        RECT 60.480 201.900 61.245 202.040 ;
        RECT 60.480 201.840 60.800 201.900 ;
        RECT 60.955 201.855 61.245 201.900 ;
        RECT 70.140 202.040 70.460 202.100 ;
        RECT 71.075 202.040 71.365 202.085 ;
        RECT 70.140 201.900 71.365 202.040 ;
        RECT 70.140 201.840 70.460 201.900 ;
        RECT 71.075 201.855 71.365 201.900 ;
        RECT 76.595 201.855 76.885 202.085 ;
        RECT 76.670 201.700 76.810 201.855 ;
        RECT 77.130 201.760 77.270 202.240 ;
        RECT 75.750 201.560 76.810 201.700 ;
        RECT 61.860 201.160 62.180 201.420 ;
        RECT 74.280 201.360 74.600 201.420 ;
        RECT 75.750 201.360 75.890 201.560 ;
        RECT 77.040 201.500 77.360 201.760 ;
        RECT 78.050 201.420 78.190 202.580 ;
        RECT 91.315 202.580 110.390 202.720 ;
        RECT 91.315 202.535 91.605 202.580 ;
        RECT 109.240 202.180 109.560 202.440 ;
        RECT 79.800 202.040 80.120 202.100 ;
        RECT 80.275 202.040 80.565 202.085 ;
        RECT 79.800 201.900 80.565 202.040 ;
        RECT 79.800 201.840 80.120 201.900 ;
        RECT 80.275 201.855 80.565 201.900 ;
        RECT 86.255 202.040 86.545 202.085 ;
        RECT 86.715 202.040 87.005 202.085 ;
        RECT 86.255 201.900 87.005 202.040 ;
        RECT 86.255 201.855 86.545 201.900 ;
        RECT 86.715 201.855 87.005 201.900 ;
        RECT 87.160 202.040 87.480 202.100 ;
        RECT 89.475 202.040 89.765 202.085 ;
        RECT 87.160 201.900 89.765 202.040 ;
        RECT 87.160 201.840 87.480 201.900 ;
        RECT 89.475 201.855 89.765 201.900 ;
        RECT 89.920 202.040 90.240 202.100 ;
        RECT 90.395 202.040 90.685 202.085 ;
        RECT 89.920 201.900 90.685 202.040 ;
        RECT 89.920 201.840 90.240 201.900 ;
        RECT 90.395 201.855 90.685 201.900 ;
        RECT 97.295 202.040 97.585 202.085 ;
        RECT 98.200 202.040 98.520 202.100 ;
        RECT 97.295 201.900 98.520 202.040 ;
        RECT 97.295 201.855 97.585 201.900 ;
        RECT 98.200 201.840 98.520 201.900 ;
        RECT 98.675 201.855 98.965 202.085 ;
        RECT 100.515 201.855 100.805 202.085 ;
        RECT 82.560 201.700 82.880 201.760 ;
        RECT 98.750 201.700 98.890 201.855 ;
        RECT 82.560 201.560 98.890 201.700 ;
        RECT 100.590 201.700 100.730 201.855 ;
        RECT 102.800 201.840 103.120 202.100 ;
        RECT 110.250 201.700 110.390 202.580 ;
        RECT 110.710 202.085 110.850 202.920 ;
        RECT 110.635 202.040 110.925 202.085 ;
        RECT 116.600 202.040 116.920 202.100 ;
        RECT 110.635 201.900 116.920 202.040 ;
        RECT 110.635 201.855 110.925 201.900 ;
        RECT 116.600 201.840 116.920 201.900 ;
        RECT 118.440 202.040 118.760 202.100 ;
        RECT 118.915 202.040 119.205 202.085 ;
        RECT 118.440 201.900 119.205 202.040 ;
        RECT 118.440 201.840 118.760 201.900 ;
        RECT 118.915 201.855 119.205 201.900 ;
        RECT 114.300 201.700 114.620 201.760 ;
        RECT 100.590 201.560 106.710 201.700 ;
        RECT 110.250 201.560 114.620 201.700 ;
        RECT 82.560 201.500 82.880 201.560 ;
        RECT 106.570 201.420 106.710 201.560 ;
        RECT 114.300 201.500 114.620 201.560 ;
        RECT 74.280 201.220 75.890 201.360 ;
        RECT 74.280 201.160 74.600 201.220 ;
        RECT 76.580 201.160 76.900 201.420 ;
        RECT 77.960 201.360 78.280 201.420 ;
        RECT 81.195 201.360 81.485 201.405 ;
        RECT 77.960 201.220 81.485 201.360 ;
        RECT 77.960 201.160 78.280 201.220 ;
        RECT 81.195 201.175 81.485 201.220 ;
        RECT 85.780 201.160 86.100 201.420 ;
        RECT 98.200 201.160 98.520 201.420 ;
        RECT 99.595 201.360 99.885 201.405 ;
        RECT 100.960 201.360 101.280 201.420 ;
        RECT 99.595 201.220 101.280 201.360 ;
        RECT 99.595 201.175 99.885 201.220 ;
        RECT 100.960 201.160 101.280 201.220 ;
        RECT 106.020 201.160 106.340 201.420 ;
        RECT 106.480 201.160 106.800 201.420 ;
        RECT 113.840 201.160 114.160 201.420 ;
        RECT 119.820 201.160 120.140 201.420 ;
        RECT 57.190 200.540 132.030 201.020 ;
        RECT 61.860 200.140 62.180 200.400 ;
        RECT 74.280 200.340 74.600 200.400 ;
        RECT 78.435 200.340 78.725 200.385 ;
        RECT 97.740 200.340 98.060 200.400 ;
        RECT 74.280 200.200 74.970 200.340 ;
        RECT 74.280 200.140 74.600 200.200 ;
        RECT 61.950 199.660 62.090 200.140 ;
        RECT 72.915 199.660 73.205 199.705 ;
        RECT 61.950 199.520 73.205 199.660 ;
        RECT 72.915 199.475 73.205 199.520 ;
        RECT 72.455 199.135 72.745 199.365 ;
        RECT 72.530 198.640 72.670 199.135 ;
        RECT 72.990 198.980 73.130 199.475 ;
        RECT 74.830 199.365 74.970 200.200 ;
        RECT 78.435 200.200 98.060 200.340 ;
        RECT 78.435 200.155 78.725 200.200 ;
        RECT 97.740 200.140 98.060 200.200 ;
        RECT 98.200 200.340 98.520 200.400 ;
        RECT 101.895 200.340 102.185 200.385 ;
        RECT 98.200 200.200 102.185 200.340 ;
        RECT 98.200 200.140 98.520 200.200 ;
        RECT 101.895 200.155 102.185 200.200 ;
        RECT 102.355 200.340 102.645 200.385 ;
        RECT 102.800 200.340 103.120 200.400 ;
        RECT 102.355 200.200 103.120 200.340 ;
        RECT 102.355 200.155 102.645 200.200 ;
        RECT 77.040 200.000 77.360 200.060 ;
        RECT 80.735 200.000 81.025 200.045 ;
        RECT 83.495 200.000 83.785 200.045 ;
        RECT 76.210 199.860 80.490 200.000 ;
        RECT 76.210 199.705 76.350 199.860 ;
        RECT 77.040 199.800 77.360 199.860 ;
        RECT 75.215 199.475 75.505 199.705 ;
        RECT 76.135 199.475 76.425 199.705 ;
        RECT 74.755 199.135 75.045 199.365 ;
        RECT 75.290 199.320 75.430 199.475 ;
        RECT 76.580 199.460 76.900 199.720 ;
        RECT 77.500 199.460 77.820 199.720 ;
        RECT 79.815 199.660 80.105 199.705 ;
        RECT 79.430 199.520 80.105 199.660 ;
        RECT 80.350 199.660 80.490 199.860 ;
        RECT 80.735 199.860 83.785 200.000 ;
        RECT 80.735 199.815 81.025 199.860 ;
        RECT 83.495 199.815 83.785 199.860 ;
        RECT 90.010 199.860 92.910 200.000 ;
        RECT 90.010 199.720 90.150 199.860 ;
        RECT 81.180 199.660 81.500 199.720 ;
        RECT 80.350 199.520 81.500 199.660 ;
        RECT 75.290 199.180 77.730 199.320 ;
        RECT 75.290 198.980 75.430 199.180 ;
        RECT 72.990 198.840 75.430 198.980 ;
        RECT 77.040 198.780 77.360 199.040 ;
        RECT 77.590 198.980 77.730 199.180 ;
        RECT 79.430 198.980 79.570 199.520 ;
        RECT 79.815 199.475 80.105 199.520 ;
        RECT 81.180 199.460 81.500 199.520 ;
        RECT 81.640 199.460 81.960 199.720 ;
        RECT 84.875 199.475 85.165 199.705 ;
        RECT 83.495 199.320 83.785 199.365 ;
        RECT 83.110 199.180 83.785 199.320 ;
        RECT 84.950 199.320 85.090 199.475 ;
        RECT 89.920 199.460 90.240 199.720 ;
        RECT 91.415 199.660 91.705 199.705 ;
        RECT 92.220 199.660 92.540 199.720 ;
        RECT 92.770 199.705 92.910 199.860 ;
        RECT 101.420 199.800 101.740 200.060 ;
        RECT 91.415 199.520 92.540 199.660 ;
        RECT 91.415 199.475 91.705 199.520 ;
        RECT 92.220 199.460 92.540 199.520 ;
        RECT 92.695 199.660 92.985 199.705 ;
        RECT 93.155 199.660 93.445 199.705 ;
        RECT 92.695 199.520 93.445 199.660 ;
        RECT 92.695 199.475 92.985 199.520 ;
        RECT 93.155 199.475 93.445 199.520 ;
        RECT 94.490 199.660 94.780 199.705 ;
        RECT 96.360 199.660 96.680 199.720 ;
        RECT 94.490 199.520 96.680 199.660 ;
        RECT 94.490 199.475 94.780 199.520 ;
        RECT 96.360 199.460 96.680 199.520 ;
        RECT 86.240 199.320 86.560 199.380 ;
        RECT 101.510 199.365 101.650 199.800 ;
        RECT 84.950 199.180 86.560 199.320 ;
        RECT 80.260 198.980 80.580 199.040 ;
        RECT 77.590 198.840 80.580 198.980 ;
        RECT 80.260 198.780 80.580 198.840 ;
        RECT 82.560 198.780 82.880 199.040 ;
        RECT 83.110 198.980 83.250 199.180 ;
        RECT 83.495 199.135 83.785 199.180 ;
        RECT 86.240 199.120 86.560 199.180 ;
        RECT 88.105 199.320 88.395 199.365 ;
        RECT 90.625 199.320 90.915 199.365 ;
        RECT 91.815 199.320 92.105 199.365 ;
        RECT 88.105 199.180 92.105 199.320 ;
        RECT 88.105 199.135 88.395 199.180 ;
        RECT 90.625 199.135 90.915 199.180 ;
        RECT 91.815 199.135 92.105 199.180 ;
        RECT 94.035 199.320 94.325 199.365 ;
        RECT 95.225 199.320 95.515 199.365 ;
        RECT 97.745 199.320 98.035 199.365 ;
        RECT 94.035 199.180 98.035 199.320 ;
        RECT 94.035 199.135 94.325 199.180 ;
        RECT 95.225 199.135 95.515 199.180 ;
        RECT 97.745 199.135 98.035 199.180 ;
        RECT 101.435 199.135 101.725 199.365 ;
        RECT 85.795 198.980 86.085 199.025 ;
        RECT 87.160 198.980 87.480 199.040 ;
        RECT 83.110 198.840 87.480 198.980 ;
        RECT 83.110 198.640 83.250 198.840 ;
        RECT 85.795 198.795 86.085 198.840 ;
        RECT 87.160 198.780 87.480 198.840 ;
        RECT 88.540 198.980 88.830 199.025 ;
        RECT 90.110 198.980 90.400 199.025 ;
        RECT 92.210 198.980 92.500 199.025 ;
        RECT 88.540 198.840 92.500 198.980 ;
        RECT 88.540 198.795 88.830 198.840 ;
        RECT 90.110 198.795 90.400 198.840 ;
        RECT 92.210 198.795 92.500 198.840 ;
        RECT 93.640 198.980 93.930 199.025 ;
        RECT 95.740 198.980 96.030 199.025 ;
        RECT 97.310 198.980 97.600 199.025 ;
        RECT 93.640 198.840 97.600 198.980 ;
        RECT 93.640 198.795 93.930 198.840 ;
        RECT 95.740 198.795 96.030 198.840 ;
        RECT 97.310 198.795 97.600 198.840 ;
        RECT 100.055 198.980 100.345 199.025 ;
        RECT 102.430 198.980 102.570 200.155 ;
        RECT 102.800 200.140 103.120 200.200 ;
        RECT 106.020 200.140 106.340 200.400 ;
        RECT 123.500 200.340 123.820 200.400 ;
        RECT 114.390 200.200 123.820 200.340 ;
        RECT 105.575 199.660 105.865 199.705 ;
        RECT 106.110 199.660 106.250 200.140 ;
        RECT 114.390 200.000 114.530 200.200 ;
        RECT 123.500 200.140 123.820 200.200 ;
        RECT 105.575 199.520 106.250 199.660 ;
        RECT 110.250 199.860 114.530 200.000 ;
        RECT 115.215 200.000 115.865 200.045 ;
        RECT 118.815 200.000 119.105 200.045 ;
        RECT 124.895 200.000 125.185 200.045 ;
        RECT 115.215 199.860 125.185 200.000 ;
        RECT 105.575 199.475 105.865 199.520 ;
        RECT 100.055 198.840 102.570 198.980 ;
        RECT 104.195 198.980 104.485 199.025 ;
        RECT 110.250 198.980 110.390 199.860 ;
        RECT 115.215 199.815 115.865 199.860 ;
        RECT 118.515 199.815 119.105 199.860 ;
        RECT 124.895 199.815 125.185 199.860 ;
        RECT 111.555 199.660 111.845 199.705 ;
        RECT 111.170 199.520 111.845 199.660 ;
        RECT 111.170 199.380 111.310 199.520 ;
        RECT 111.555 199.475 111.845 199.520 ;
        RECT 112.020 199.660 112.310 199.705 ;
        RECT 113.855 199.660 114.145 199.705 ;
        RECT 117.435 199.660 117.725 199.705 ;
        RECT 112.020 199.520 117.725 199.660 ;
        RECT 112.020 199.475 112.310 199.520 ;
        RECT 113.855 199.475 114.145 199.520 ;
        RECT 117.435 199.475 117.725 199.520 ;
        RECT 118.515 199.500 118.805 199.815 ;
        RECT 119.820 199.660 120.140 199.720 ;
        RECT 124.435 199.660 124.725 199.705 ;
        RECT 119.820 199.520 124.725 199.660 ;
        RECT 119.820 199.460 120.140 199.520 ;
        RECT 124.435 199.475 124.725 199.520 ;
        RECT 111.080 199.120 111.400 199.380 ;
        RECT 112.935 199.320 113.225 199.365 ;
        RECT 113.380 199.320 113.700 199.380 ;
        RECT 112.935 199.180 113.700 199.320 ;
        RECT 112.935 199.135 113.225 199.180 ;
        RECT 113.380 199.120 113.700 199.180 ;
        RECT 120.295 199.320 120.585 199.365 ;
        RECT 123.515 199.320 123.805 199.365 ;
        RECT 120.295 199.180 123.805 199.320 ;
        RECT 120.295 199.135 120.585 199.180 ;
        RECT 123.515 199.135 123.805 199.180 ;
        RECT 104.195 198.840 110.390 198.980 ;
        RECT 112.425 198.980 112.715 199.025 ;
        RECT 114.315 198.980 114.605 199.025 ;
        RECT 117.435 198.980 117.725 199.025 ;
        RECT 112.425 198.840 117.725 198.980 ;
        RECT 100.055 198.795 100.345 198.840 ;
        RECT 104.195 198.795 104.485 198.840 ;
        RECT 112.425 198.795 112.715 198.840 ;
        RECT 114.315 198.795 114.605 198.840 ;
        RECT 117.435 198.795 117.725 198.840 ;
        RECT 72.530 198.500 83.250 198.640 ;
        RECT 83.480 198.640 83.800 198.700 ;
        RECT 84.415 198.640 84.705 198.685 ;
        RECT 83.480 198.500 84.705 198.640 ;
        RECT 83.480 198.440 83.800 198.500 ;
        RECT 84.415 198.455 84.705 198.500 ;
        RECT 91.300 198.640 91.620 198.700 ;
        RECT 100.960 198.640 101.280 198.700 ;
        RECT 91.300 198.500 101.280 198.640 ;
        RECT 91.300 198.440 91.620 198.500 ;
        RECT 100.960 198.440 101.280 198.500 ;
        RECT 101.880 198.640 102.200 198.700 ;
        RECT 105.115 198.640 105.405 198.685 ;
        RECT 101.880 198.500 105.405 198.640 ;
        RECT 101.880 198.440 102.200 198.500 ;
        RECT 105.115 198.455 105.405 198.500 ;
        RECT 106.480 198.640 106.800 198.700 ;
        RECT 120.370 198.640 120.510 199.135 ;
        RECT 106.480 198.500 120.510 198.640 ;
        RECT 106.480 198.440 106.800 198.500 ;
        RECT 120.740 198.440 121.060 198.700 ;
        RECT 57.190 197.820 131.250 198.300 ;
        RECT 74.280 197.420 74.600 197.680 ;
        RECT 77.040 197.620 77.360 197.680 ;
        RECT 77.975 197.620 78.265 197.665 ;
        RECT 77.040 197.480 78.265 197.620 ;
        RECT 77.040 197.420 77.360 197.480 ;
        RECT 77.975 197.435 78.265 197.480 ;
        RECT 81.640 197.620 81.960 197.680 ;
        RECT 82.575 197.620 82.865 197.665 ;
        RECT 81.640 197.480 82.865 197.620 ;
        RECT 81.640 197.420 81.960 197.480 ;
        RECT 82.575 197.435 82.865 197.480 ;
        RECT 85.780 197.420 86.100 197.680 ;
        RECT 90.380 197.620 90.700 197.680 ;
        RECT 92.220 197.620 92.540 197.680 ;
        RECT 92.695 197.620 92.985 197.665 ;
        RECT 87.250 197.480 91.990 197.620 ;
        RECT 74.370 196.940 74.510 197.420 ;
        RECT 76.135 197.280 76.425 197.325 ;
        RECT 76.135 197.140 78.190 197.280 ;
        RECT 76.135 197.095 76.425 197.140 ;
        RECT 74.370 196.800 77.270 196.940 ;
        RECT 77.130 196.645 77.270 196.800 ;
        RECT 78.050 196.660 78.190 197.140 ;
        RECT 80.260 196.940 80.580 197.000 ;
        RECT 85.870 196.985 86.010 197.420 ;
        RECT 85.335 196.940 85.625 196.985 ;
        RECT 80.260 196.800 85.625 196.940 ;
        RECT 80.260 196.740 80.580 196.800 ;
        RECT 85.335 196.755 85.625 196.800 ;
        RECT 85.795 196.940 86.085 196.985 ;
        RECT 85.795 196.800 86.930 196.940 ;
        RECT 85.795 196.755 86.085 196.800 ;
        RECT 75.675 196.415 75.965 196.645 ;
        RECT 77.055 196.415 77.345 196.645 ;
        RECT 75.750 196.260 75.890 196.415 ;
        RECT 77.960 196.400 78.280 196.660 ;
        RECT 80.720 196.400 81.040 196.660 ;
        RECT 83.480 196.600 83.770 196.645 ;
        RECT 86.240 196.600 86.560 196.660 ;
        RECT 83.480 196.460 86.560 196.600 ;
        RECT 83.480 196.415 83.770 196.460 ;
        RECT 80.810 196.260 80.950 196.400 ;
        RECT 75.750 196.120 80.950 196.260 ;
        RECT 81.180 195.920 81.500 195.980 ;
        RECT 83.480 195.920 83.800 195.980 ;
        RECT 81.180 195.780 83.800 195.920 ;
        RECT 85.870 195.920 86.010 196.460 ;
        RECT 86.240 196.400 86.560 196.460 ;
        RECT 86.790 196.260 86.930 196.800 ;
        RECT 87.250 196.645 87.390 197.480 ;
        RECT 90.380 197.420 90.700 197.480 ;
        RECT 88.555 197.095 88.845 197.325 ;
        RECT 91.300 197.280 91.620 197.340 ;
        RECT 90.470 197.140 91.620 197.280 ;
        RECT 88.630 196.940 88.770 197.095 ;
        RECT 89.475 196.940 89.765 196.985 ;
        RECT 88.630 196.800 89.765 196.940 ;
        RECT 89.475 196.755 89.765 196.800 ;
        RECT 87.175 196.415 87.465 196.645 ;
        RECT 87.635 196.415 87.925 196.645 ;
        RECT 90.470 196.600 90.610 197.140 ;
        RECT 91.300 197.080 91.620 197.140 ;
        RECT 91.850 196.940 91.990 197.480 ;
        RECT 92.220 197.480 92.985 197.620 ;
        RECT 92.220 197.420 92.540 197.480 ;
        RECT 92.695 197.435 92.985 197.480 ;
        RECT 96.360 197.420 96.680 197.680 ;
        RECT 101.420 197.420 101.740 197.680 ;
        RECT 106.480 197.420 106.800 197.680 ;
        RECT 111.540 197.620 111.860 197.680 ;
        RECT 113.855 197.620 114.145 197.665 ;
        RECT 111.540 197.480 114.145 197.620 ;
        RECT 111.540 197.420 111.860 197.480 ;
        RECT 113.855 197.435 114.145 197.480 ;
        RECT 116.600 197.620 116.920 197.680 ;
        RECT 117.995 197.620 118.285 197.665 ;
        RECT 116.600 197.480 118.285 197.620 ;
        RECT 116.600 197.420 116.920 197.480 ;
        RECT 117.995 197.435 118.285 197.480 ;
        RECT 101.510 197.280 101.650 197.420 ;
        RECT 101.510 197.140 102.570 197.280 ;
        RECT 93.615 196.940 93.905 196.985 ;
        RECT 100.055 196.940 100.345 196.985 ;
        RECT 101.880 196.940 102.200 197.000 ;
        RECT 91.850 196.800 93.905 196.940 ;
        RECT 93.615 196.755 93.905 196.800 ;
        RECT 97.370 196.800 100.345 196.940 ;
        RECT 93.155 196.600 93.445 196.645 ;
        RECT 88.630 196.460 90.610 196.600 ;
        RECT 91.390 196.460 93.445 196.600 ;
        RECT 87.710 196.260 87.850 196.415 ;
        RECT 88.630 196.305 88.770 196.460 ;
        RECT 86.790 196.120 87.850 196.260 ;
        RECT 88.555 196.075 88.845 196.305 ;
        RECT 88.080 195.920 88.400 195.980 ;
        RECT 91.390 195.920 91.530 196.460 ;
        RECT 93.155 196.415 93.445 196.460 ;
        RECT 94.075 196.600 94.365 196.645 ;
        RECT 95.440 196.600 95.760 196.660 ;
        RECT 97.370 196.645 97.510 196.800 ;
        RECT 100.055 196.755 100.345 196.800 ;
        RECT 100.590 196.800 102.200 196.940 ;
        RECT 94.075 196.460 95.760 196.600 ;
        RECT 94.075 196.415 94.365 196.460 ;
        RECT 95.440 196.400 95.760 196.460 ;
        RECT 97.295 196.415 97.585 196.645 ;
        RECT 97.740 196.600 98.060 196.660 ;
        RECT 98.675 196.600 98.965 196.645 ;
        RECT 99.595 196.600 99.885 196.645 ;
        RECT 100.590 196.600 100.730 196.800 ;
        RECT 101.510 196.645 101.650 196.800 ;
        RECT 101.880 196.740 102.200 196.800 ;
        RECT 102.430 196.645 102.570 197.140 ;
        RECT 97.740 196.460 99.350 196.600 ;
        RECT 97.740 196.400 98.060 196.460 ;
        RECT 98.675 196.415 98.965 196.460 ;
        RECT 99.210 196.260 99.350 196.460 ;
        RECT 99.595 196.460 100.730 196.600 ;
        RECT 99.595 196.415 99.885 196.460 ;
        RECT 100.975 196.415 101.265 196.645 ;
        RECT 101.435 196.415 101.725 196.645 ;
        RECT 102.355 196.415 102.645 196.645 ;
        RECT 102.815 196.600 103.105 196.645 ;
        RECT 106.570 196.600 106.710 197.420 ;
        RECT 128.100 197.280 128.420 197.340 ;
        RECT 113.470 197.140 128.420 197.280 ;
        RECT 113.470 196.645 113.610 197.140 ;
        RECT 128.100 197.080 128.420 197.140 ;
        RECT 114.300 196.940 114.620 197.000 ;
        RECT 116.155 196.940 116.445 196.985 ;
        RECT 114.300 196.800 116.445 196.940 ;
        RECT 114.300 196.740 114.620 196.800 ;
        RECT 116.155 196.755 116.445 196.800 ;
        RECT 116.600 196.740 116.920 197.000 ;
        RECT 120.740 196.940 121.060 197.000 ;
        RECT 119.450 196.800 121.060 196.940 ;
        RECT 102.815 196.460 106.710 196.600 ;
        RECT 102.815 196.415 103.105 196.460 ;
        RECT 113.395 196.415 113.685 196.645 ;
        RECT 113.840 196.600 114.160 196.660 ;
        RECT 119.450 196.645 119.590 196.800 ;
        RECT 120.740 196.740 121.060 196.800 ;
        RECT 117.995 196.600 118.285 196.645 ;
        RECT 113.840 196.460 118.285 196.600 ;
        RECT 101.050 196.260 101.190 196.415 ;
        RECT 113.840 196.400 114.160 196.460 ;
        RECT 117.995 196.415 118.285 196.460 ;
        RECT 118.915 196.415 119.205 196.645 ;
        RECT 119.375 196.415 119.665 196.645 ;
        RECT 123.055 196.600 123.345 196.645 ;
        RECT 120.370 196.460 123.345 196.600 ;
        RECT 103.260 196.260 103.580 196.320 ;
        RECT 99.210 196.120 103.580 196.260 ;
        RECT 103.260 196.060 103.580 196.120 ;
        RECT 110.620 196.260 110.940 196.320 ;
        RECT 118.990 196.260 119.130 196.415 ;
        RECT 110.620 196.120 119.130 196.260 ;
        RECT 110.620 196.060 110.940 196.120 ;
        RECT 85.870 195.780 91.530 195.920 ;
        RECT 104.640 195.920 104.960 195.980 ;
        RECT 106.035 195.920 106.325 195.965 ;
        RECT 104.640 195.780 106.325 195.920 ;
        RECT 81.180 195.720 81.500 195.780 ;
        RECT 83.480 195.720 83.800 195.780 ;
        RECT 88.080 195.720 88.400 195.780 ;
        RECT 104.640 195.720 104.960 195.780 ;
        RECT 106.035 195.735 106.325 195.780 ;
        RECT 115.680 195.720 116.000 195.980 ;
        RECT 120.370 195.965 120.510 196.460 ;
        RECT 123.055 196.415 123.345 196.460 ;
        RECT 120.295 195.735 120.585 195.965 ;
        RECT 120.740 195.920 121.060 195.980 ;
        RECT 122.135 195.920 122.425 195.965 ;
        RECT 120.740 195.780 122.425 195.920 ;
        RECT 120.740 195.720 121.060 195.780 ;
        RECT 122.135 195.735 122.425 195.780 ;
        RECT 57.190 195.100 132.030 195.580 ;
        RECT 77.500 194.900 77.820 194.960 ;
        RECT 77.975 194.900 78.265 194.945 ;
        RECT 77.500 194.760 78.265 194.900 ;
        RECT 77.500 194.700 77.820 194.760 ;
        RECT 77.975 194.715 78.265 194.760 ;
        RECT 106.035 194.900 106.325 194.945 ;
        RECT 110.620 194.900 110.940 194.960 ;
        RECT 106.035 194.760 110.940 194.900 ;
        RECT 106.035 194.715 106.325 194.760 ;
        RECT 110.620 194.700 110.940 194.760 ;
        RECT 115.680 194.700 116.000 194.960 ;
        RECT 92.235 194.560 92.525 194.605 ;
        RECT 104.640 194.560 104.960 194.620 ;
        RECT 109.255 194.560 109.545 194.605 ;
        RECT 92.235 194.420 109.545 194.560 ;
        RECT 92.235 194.375 92.525 194.420 ;
        RECT 104.640 194.360 104.960 194.420 ;
        RECT 109.255 194.375 109.545 194.420 ;
        RECT 79.815 194.220 80.105 194.265 ;
        RECT 81.180 194.220 81.500 194.280 ;
        RECT 79.815 194.080 81.500 194.220 ;
        RECT 79.815 194.035 80.105 194.080 ;
        RECT 81.180 194.020 81.500 194.080 ;
        RECT 91.300 194.220 91.620 194.280 ;
        RECT 92.695 194.220 92.985 194.265 ;
        RECT 91.300 194.080 92.985 194.220 ;
        RECT 91.300 194.020 91.620 194.080 ;
        RECT 92.695 194.035 92.985 194.080 ;
        RECT 103.260 194.220 103.580 194.280 ;
        RECT 105.115 194.220 105.405 194.265 ;
        RECT 106.495 194.220 106.785 194.265 ;
        RECT 103.260 194.080 106.785 194.220 ;
        RECT 103.260 194.020 103.580 194.080 ;
        RECT 105.115 194.035 105.405 194.080 ;
        RECT 106.495 194.035 106.785 194.080 ;
        RECT 107.415 194.220 107.705 194.265 ;
        RECT 108.780 194.220 109.100 194.280 ;
        RECT 115.770 194.220 115.910 194.700 ;
        RECT 107.415 194.080 115.910 194.220 ;
        RECT 107.415 194.035 107.705 194.080 ;
        RECT 108.780 194.020 109.100 194.080 ;
        RECT 80.260 193.680 80.580 193.940 ;
        RECT 80.735 193.695 81.025 193.925 ;
        RECT 104.195 193.695 104.485 193.925 ;
        RECT 106.955 193.880 107.245 193.925 ;
        RECT 113.840 193.880 114.160 193.940 ;
        RECT 106.955 193.740 114.160 193.880 ;
        RECT 106.955 193.695 107.245 193.740 ;
        RECT 78.420 193.540 78.740 193.600 ;
        RECT 80.810 193.540 80.950 193.695 ;
        RECT 78.420 193.400 80.950 193.540 ;
        RECT 104.270 193.540 104.410 193.695 ;
        RECT 113.840 193.680 114.160 193.740 ;
        RECT 108.780 193.540 109.100 193.600 ;
        RECT 104.270 193.400 109.100 193.540 ;
        RECT 78.420 193.340 78.740 193.400 ;
        RECT 108.780 193.340 109.100 193.400 ;
        RECT 85.795 193.200 86.085 193.245 ;
        RECT 89.920 193.200 90.240 193.260 ;
        RECT 85.795 193.060 90.240 193.200 ;
        RECT 85.795 193.015 86.085 193.060 ;
        RECT 89.920 193.000 90.240 193.060 ;
        RECT 93.600 193.000 93.920 193.260 ;
        RECT 115.680 193.000 116.000 193.260 ;
        RECT 57.190 192.380 131.250 192.860 ;
        RECT 77.960 191.980 78.280 192.240 ;
        RECT 78.420 191.980 78.740 192.240 ;
        RECT 80.260 192.180 80.580 192.240 ;
        RECT 81.655 192.180 81.945 192.225 ;
        RECT 80.260 192.040 81.945 192.180 ;
        RECT 80.260 191.980 80.580 192.040 ;
        RECT 81.655 191.995 81.945 192.040 ;
        RECT 82.575 191.995 82.865 192.225 ;
        RECT 78.050 191.840 78.190 191.980 ;
        RECT 82.650 191.840 82.790 191.995 ;
        RECT 88.080 191.980 88.400 192.240 ;
        RECT 108.780 192.180 109.100 192.240 ;
        RECT 109.255 192.180 109.545 192.225 ;
        RECT 108.780 192.040 109.545 192.180 ;
        RECT 108.780 191.980 109.100 192.040 ;
        RECT 109.255 191.995 109.545 192.040 ;
        RECT 78.050 191.700 82.790 191.840 ;
        RECT 90.840 191.840 91.130 191.885 ;
        RECT 92.410 191.840 92.700 191.885 ;
        RECT 94.510 191.840 94.800 191.885 ;
        RECT 90.840 191.700 94.800 191.840 ;
        RECT 90.840 191.655 91.130 191.700 ;
        RECT 92.410 191.655 92.700 191.700 ;
        RECT 94.510 191.655 94.800 191.700 ;
        RECT 99.120 191.840 99.410 191.885 ;
        RECT 100.690 191.840 100.980 191.885 ;
        RECT 102.790 191.840 103.080 191.885 ;
        RECT 99.120 191.700 103.080 191.840 ;
        RECT 99.120 191.655 99.410 191.700 ;
        RECT 100.690 191.655 100.980 191.700 ;
        RECT 102.790 191.655 103.080 191.700 ;
        RECT 112.000 191.840 112.290 191.885 ;
        RECT 113.570 191.840 113.860 191.885 ;
        RECT 115.670 191.840 115.960 191.885 ;
        RECT 112.000 191.700 115.960 191.840 ;
        RECT 112.000 191.655 112.290 191.700 ;
        RECT 113.570 191.655 113.860 191.700 ;
        RECT 115.670 191.655 115.960 191.700 ;
        RECT 79.815 191.315 80.105 191.545 ;
        RECT 79.890 190.820 80.030 191.315 ;
        RECT 89.920 191.300 90.240 191.560 ;
        RECT 90.405 191.500 90.695 191.545 ;
        RECT 92.925 191.500 93.215 191.545 ;
        RECT 94.115 191.500 94.405 191.545 ;
        RECT 90.405 191.360 94.405 191.500 ;
        RECT 90.405 191.315 90.695 191.360 ;
        RECT 92.925 191.315 93.215 191.360 ;
        RECT 94.115 191.315 94.405 191.360 ;
        RECT 98.685 191.500 98.975 191.545 ;
        RECT 101.205 191.500 101.495 191.545 ;
        RECT 102.395 191.500 102.685 191.545 ;
        RECT 98.685 191.360 102.685 191.500 ;
        RECT 98.685 191.315 98.975 191.360 ;
        RECT 101.205 191.315 101.495 191.360 ;
        RECT 102.395 191.315 102.685 191.360 ;
        RECT 111.565 191.500 111.855 191.545 ;
        RECT 114.085 191.500 114.375 191.545 ;
        RECT 115.275 191.500 115.565 191.545 ;
        RECT 111.565 191.360 115.565 191.500 ;
        RECT 111.565 191.315 111.855 191.360 ;
        RECT 114.085 191.315 114.375 191.360 ;
        RECT 115.275 191.315 115.565 191.360 ;
        RECT 80.275 191.160 80.565 191.205 ;
        RECT 80.720 191.160 81.040 191.220 ;
        RECT 80.275 191.020 81.040 191.160 ;
        RECT 80.275 190.975 80.565 191.020 ;
        RECT 80.720 190.960 81.040 191.020 ;
        RECT 83.940 191.160 84.260 191.220 ;
        RECT 87.635 191.160 87.925 191.205 ;
        RECT 89.460 191.160 89.780 191.220 ;
        RECT 83.940 191.020 86.930 191.160 ;
        RECT 83.940 190.960 84.260 191.020 ;
        RECT 86.790 190.865 86.930 191.020 ;
        RECT 87.635 191.020 89.780 191.160 ;
        RECT 90.010 191.160 90.150 191.300 ;
        RECT 94.995 191.160 95.285 191.205 ;
        RECT 90.010 191.020 95.285 191.160 ;
        RECT 87.635 190.975 87.925 191.020 ;
        RECT 89.460 190.960 89.780 191.020 ;
        RECT 94.995 190.975 95.285 191.020 ;
        RECT 103.275 191.160 103.565 191.205 ;
        RECT 111.080 191.160 111.400 191.220 ;
        RECT 115.680 191.160 116.000 191.220 ;
        RECT 116.155 191.160 116.445 191.205 ;
        RECT 103.275 191.020 116.445 191.160 ;
        RECT 103.275 190.975 103.565 191.020 ;
        RECT 111.080 190.960 111.400 191.020 ;
        RECT 115.680 190.960 116.000 191.020 ;
        RECT 116.155 190.975 116.445 191.020 ;
        RECT 93.600 190.865 93.920 190.880 ;
        RECT 85.795 190.820 86.085 190.865 ;
        RECT 79.890 190.680 86.085 190.820 ;
        RECT 85.795 190.635 86.085 190.680 ;
        RECT 86.715 190.820 87.005 190.865 ;
        RECT 93.600 190.820 93.950 190.865 ;
        RECT 101.420 190.820 101.740 190.880 ;
        RECT 101.940 190.820 102.230 190.865 ;
        RECT 86.715 190.680 89.690 190.820 ;
        RECT 86.715 190.635 87.005 190.680 ;
        RECT 85.870 190.480 86.010 190.635 ;
        RECT 88.080 190.480 88.400 190.540 ;
        RECT 85.870 190.340 88.400 190.480 ;
        RECT 89.550 190.480 89.690 190.680 ;
        RECT 93.600 190.680 94.115 190.820 ;
        RECT 101.420 190.680 102.230 190.820 ;
        RECT 93.600 190.635 93.950 190.680 ;
        RECT 93.600 190.620 93.920 190.635 ;
        RECT 101.420 190.620 101.740 190.680 ;
        RECT 101.940 190.635 102.230 190.680 ;
        RECT 114.930 190.820 115.220 190.865 ;
        RECT 120.740 190.820 121.060 190.880 ;
        RECT 114.930 190.680 121.060 190.820 ;
        RECT 114.930 190.635 115.220 190.680 ;
        RECT 120.740 190.620 121.060 190.680 ;
        RECT 96.360 190.480 96.680 190.540 ;
        RECT 89.550 190.340 96.680 190.480 ;
        RECT 88.080 190.280 88.400 190.340 ;
        RECT 96.360 190.280 96.680 190.340 ;
        RECT 57.190 189.660 132.030 190.140 ;
        RECT 77.960 189.260 78.280 189.520 ;
        RECT 81.180 189.260 81.500 189.520 ;
        RECT 89.475 189.460 89.765 189.505 ;
        RECT 89.920 189.460 90.240 189.520 ;
        RECT 89.475 189.320 90.240 189.460 ;
        RECT 89.475 189.275 89.765 189.320 ;
        RECT 89.920 189.260 90.240 189.320 ;
        RECT 90.380 189.260 90.700 189.520 ;
        RECT 95.440 189.460 95.760 189.520 ;
        RECT 100.055 189.460 100.345 189.505 ;
        RECT 95.440 189.320 100.345 189.460 ;
        RECT 95.440 189.260 95.760 189.320 ;
        RECT 100.055 189.275 100.345 189.320 ;
        RECT 100.975 189.460 101.265 189.505 ;
        RECT 101.420 189.460 101.740 189.520 ;
        RECT 100.975 189.320 101.740 189.460 ;
        RECT 100.975 189.275 101.265 189.320 ;
        RECT 78.050 188.780 78.190 189.260 ;
        RECT 78.895 188.780 79.185 188.825 ;
        RECT 78.050 188.640 79.185 188.780 ;
        RECT 78.895 188.595 79.185 188.640 ;
        RECT 96.360 188.780 96.680 188.840 ;
        RECT 96.835 188.780 97.125 188.825 ;
        RECT 96.360 188.640 97.125 188.780 ;
        RECT 100.130 188.780 100.270 189.275 ;
        RECT 101.420 189.260 101.740 189.320 ;
        RECT 100.515 188.780 100.805 188.825 ;
        RECT 100.130 188.640 100.805 188.780 ;
        RECT 96.360 188.580 96.680 188.640 ;
        RECT 96.835 188.595 97.125 188.640 ;
        RECT 100.515 188.595 100.805 188.640 ;
        RECT 100.960 188.780 101.280 188.840 ;
        RECT 101.435 188.780 101.725 188.825 ;
        RECT 100.960 188.640 101.725 188.780 ;
        RECT 100.960 188.580 101.280 188.640 ;
        RECT 101.435 188.595 101.725 188.640 ;
        RECT 123.500 188.780 123.820 188.840 ;
        RECT 127.195 188.780 127.485 188.825 ;
        RECT 123.500 188.640 127.485 188.780 ;
        RECT 123.500 188.580 123.820 188.640 ;
        RECT 127.195 188.595 127.485 188.640 ;
        RECT 87.635 188.440 87.925 188.485 ;
        RECT 101.050 188.440 101.190 188.580 ;
        RECT 87.635 188.300 101.190 188.440 ;
        RECT 87.635 188.255 87.925 188.300 ;
        RECT 80.275 187.760 80.565 187.805 ;
        RECT 83.480 187.760 83.800 187.820 ;
        RECT 80.275 187.620 83.800 187.760 ;
        RECT 80.275 187.575 80.565 187.620 ;
        RECT 83.480 187.560 83.800 187.620 ;
        RECT 89.460 187.560 89.780 187.820 ;
        RECT 128.100 187.560 128.420 187.820 ;
        RECT 57.190 186.940 131.250 187.420 ;
        RECT 57.190 184.220 132.030 184.700 ;
        RECT 57.190 181.500 131.250 181.980 ;
        RECT 57.190 178.780 132.030 179.260 ;
        RECT 57.190 176.060 131.250 176.540 ;
        RECT 57.190 173.340 132.030 173.820 ;
        RECT 57.190 170.620 131.250 171.100 ;
        RECT 57.190 167.900 132.030 168.380 ;
        RECT 57.190 165.180 131.250 165.660 ;
        RECT 57.190 162.460 132.030 162.940 ;
        RECT 57.190 159.740 131.250 160.220 ;
        RECT 57.190 157.020 132.030 157.500 ;
        RECT 57.190 154.300 131.250 154.780 ;
        RECT 57.190 151.580 132.030 152.060 ;
        RECT 111.080 150.840 111.400 151.100 ;
        RECT 110.620 149.480 110.940 149.740 ;
        RECT 57.190 148.860 131.250 149.340 ;
        RECT 57.190 146.140 132.030 146.620 ;
        RECT 57.190 143.420 131.250 143.900 ;
        RECT 57.190 140.700 132.030 141.180 ;
        RECT 57.190 137.980 131.250 138.460 ;
        RECT 57.190 135.260 132.030 135.740 ;
        RECT 57.190 132.540 131.250 133.020 ;
        RECT 57.190 129.820 132.030 130.300 ;
        RECT 140.950 99.000 150.000 101.000 ;
        RECT 140.950 95.000 146.000 97.000 ;
        RECT 144.000 92.000 146.000 95.000 ;
        RECT 148.000 92.000 150.000 99.000 ;
        RECT 144.120 91.570 145.120 92.000 ;
        RECT 148.120 91.570 149.120 92.000 ;
        RECT 123.950 89.610 135.000 90.000 ;
        RECT 123.950 89.590 137.790 89.610 ;
        RECT 123.950 89.570 152.120 89.590 ;
        RECT 123.950 88.550 153.520 89.570 ;
        RECT 123.950 88.000 135.000 88.550 ;
        RECT 137.670 88.520 140.320 88.550 ;
        RECT 137.920 87.270 140.120 88.520 ;
        RECT 148.170 87.820 149.070 87.870 ;
        RECT 138.470 86.420 140.220 87.070 ;
        RECT 141.320 85.470 143.470 87.770 ;
        RECT 144.820 84.470 145.320 84.570 ;
        RECT 147.870 84.520 150.120 87.820 ;
        RECT 151.120 87.270 153.520 88.550 ;
        RECT 150.820 86.570 152.620 87.070 ;
        RECT 138.720 84.070 145.320 84.470 ;
        RECT 134.950 83.570 137.000 84.000 ;
        RECT 137.470 83.570 140.170 83.920 ;
        RECT 142.970 83.570 145.670 83.920 ;
        RECT 134.950 82.570 137.820 83.570 ;
        RECT 138.770 82.570 139.170 83.420 ;
        RECT 134.950 82.000 137.000 82.570 ;
        RECT 137.470 81.470 137.820 82.570 ;
        RECT 138.840 81.620 139.070 82.570 ;
        RECT 139.510 82.270 139.740 83.420 ;
        RECT 140.070 82.570 140.570 83.420 ;
        RECT 142.840 83.370 143.070 83.420 ;
        RECT 142.720 82.620 143.170 83.370 ;
        RECT 139.420 81.720 139.820 82.270 ;
        RECT 139.510 81.620 139.740 81.720 ;
        RECT 140.180 81.620 140.410 82.570 ;
        RECT 142.840 81.620 143.070 82.620 ;
        RECT 143.510 82.270 143.740 83.420 ;
        RECT 144.180 83.370 144.410 83.420 ;
        RECT 144.070 82.620 144.470 83.370 ;
        RECT 143.420 81.720 143.820 82.270 ;
        RECT 143.510 81.620 143.740 81.720 ;
        RECT 144.180 81.620 144.410 82.620 ;
        RECT 145.320 81.720 145.670 83.570 ;
        RECT 145.220 81.470 145.670 81.720 ;
        RECT 137.470 81.460 139.320 81.470 ;
        RECT 137.470 81.420 139.460 81.460 ;
        RECT 139.790 81.420 140.130 81.460 ;
        RECT 137.470 81.120 140.170 81.420 ;
        RECT 142.920 81.120 145.670 81.470 ;
        RECT 146.520 83.570 149.220 83.920 ;
        RECT 152.020 83.570 154.720 83.920 ;
        RECT 155.950 83.570 157.050 84.000 ;
        RECT 146.520 81.470 146.870 83.570 ;
        RECT 147.840 83.370 148.070 83.420 ;
        RECT 147.770 82.620 148.170 83.370 ;
        RECT 147.840 81.620 148.070 82.620 ;
        RECT 148.510 82.320 148.740 83.420 ;
        RECT 149.180 83.370 149.410 83.420 ;
        RECT 151.840 83.370 152.070 83.420 ;
        RECT 149.070 82.620 149.520 83.370 ;
        RECT 151.770 82.620 152.170 83.370 ;
        RECT 148.420 81.670 148.870 82.320 ;
        RECT 148.510 81.620 148.740 81.670 ;
        RECT 149.180 81.620 149.410 82.620 ;
        RECT 151.840 81.620 152.070 82.620 ;
        RECT 152.510 82.320 152.740 83.420 ;
        RECT 153.180 83.370 153.410 83.420 ;
        RECT 153.070 82.620 153.520 83.370 ;
        RECT 152.420 81.670 152.820 82.320 ;
        RECT 152.510 81.620 152.740 81.670 ;
        RECT 153.180 81.620 153.410 82.620 ;
        RECT 154.370 82.570 157.050 83.570 ;
        RECT 154.370 81.470 154.820 82.570 ;
        RECT 155.950 82.000 157.050 82.570 ;
        RECT 146.520 81.120 149.220 81.470 ;
        RECT 151.970 81.120 154.820 81.470 ;
        RECT 137.470 80.395 137.820 81.120 ;
        RECT 146.520 80.395 146.870 81.120 ;
        RECT 137.470 80.020 146.870 80.395 ;
        RECT 147.770 80.170 153.620 80.970 ;
        RECT 154.370 79.870 154.820 81.120 ;
        RECT 145.270 79.470 154.820 79.870 ;
        RECT 129.950 77.570 139.000 78.000 ;
        RECT 139.570 77.570 142.220 77.920 ;
        RECT 129.950 77.000 139.870 77.570 ;
        RECT 140.840 77.370 141.070 77.420 ;
        RECT 130.000 76.570 139.870 77.000 ;
        RECT 140.770 76.670 141.170 77.370 ;
        RECT 130.000 76.000 139.000 76.570 ;
        RECT 139.570 75.470 139.870 76.570 ;
        RECT 140.840 75.620 141.070 76.670 ;
        RECT 141.510 76.370 141.740 77.420 ;
        RECT 142.180 77.370 142.410 77.420 ;
        RECT 142.120 76.670 142.520 77.370 ;
        RECT 142.720 76.820 149.570 77.820 ;
        RECT 150.070 77.570 152.720 77.920 ;
        RECT 154.000 77.570 162.050 78.000 ;
        RECT 149.840 77.320 150.070 77.420 ;
        RECT 149.770 76.670 150.170 77.320 ;
        RECT 141.420 75.670 141.820 76.370 ;
        RECT 141.510 75.620 141.740 75.670 ;
        RECT 142.180 75.620 142.410 76.670 ;
        RECT 139.570 75.120 142.220 75.470 ;
        RECT 145.770 74.820 146.470 76.420 ;
        RECT 149.840 75.620 150.070 76.670 ;
        RECT 150.510 76.370 150.740 77.420 ;
        RECT 151.180 77.320 151.410 77.420 ;
        RECT 151.120 76.670 151.520 77.320 ;
        RECT 152.420 77.000 162.050 77.570 ;
        RECT 150.420 75.720 150.820 76.370 ;
        RECT 150.510 75.620 150.740 75.720 ;
        RECT 151.180 75.620 151.410 76.670 ;
        RECT 152.420 76.570 162.000 77.000 ;
        RECT 152.420 75.470 152.720 76.570 ;
        RECT 154.000 76.000 162.000 76.570 ;
        RECT 150.070 75.120 152.720 75.470 ;
        RECT 145.820 73.570 146.470 74.270 ;
        RECT 145.620 73.000 146.620 73.570 ;
        RECT 123.950 71.000 147.000 73.000 ;
      LAYER via ;
        RECT 65.675 203.370 65.935 203.630 ;
        RECT 65.995 203.370 66.255 203.630 ;
        RECT 66.315 203.370 66.575 203.630 ;
        RECT 66.635 203.370 66.895 203.630 ;
        RECT 66.955 203.370 67.215 203.630 ;
        RECT 84.185 203.370 84.445 203.630 ;
        RECT 84.505 203.370 84.765 203.630 ;
        RECT 84.825 203.370 85.085 203.630 ;
        RECT 85.145 203.370 85.405 203.630 ;
        RECT 85.465 203.370 85.725 203.630 ;
        RECT 102.695 203.370 102.955 203.630 ;
        RECT 103.015 203.370 103.275 203.630 ;
        RECT 103.335 203.370 103.595 203.630 ;
        RECT 103.655 203.370 103.915 203.630 ;
        RECT 103.975 203.370 104.235 203.630 ;
        RECT 121.205 203.370 121.465 203.630 ;
        RECT 121.525 203.370 121.785 203.630 ;
        RECT 121.845 203.370 122.105 203.630 ;
        RECT 122.165 203.370 122.425 203.630 ;
        RECT 122.485 203.370 122.745 203.630 ;
        RECT 101.450 202.860 101.710 203.120 ;
        RECT 60.510 201.840 60.770 202.100 ;
        RECT 70.170 201.840 70.430 202.100 ;
        RECT 61.890 201.160 62.150 201.420 ;
        RECT 74.310 201.160 74.570 201.420 ;
        RECT 77.070 201.500 77.330 201.760 ;
        RECT 109.270 202.180 109.530 202.440 ;
        RECT 79.830 201.840 80.090 202.100 ;
        RECT 87.190 201.840 87.450 202.100 ;
        RECT 89.950 201.840 90.210 202.100 ;
        RECT 98.230 201.840 98.490 202.100 ;
        RECT 82.590 201.500 82.850 201.760 ;
        RECT 102.830 201.840 103.090 202.100 ;
        RECT 116.630 201.840 116.890 202.100 ;
        RECT 118.470 201.840 118.730 202.100 ;
        RECT 114.330 201.500 114.590 201.760 ;
        RECT 76.610 201.160 76.870 201.420 ;
        RECT 77.990 201.160 78.250 201.420 ;
        RECT 85.810 201.160 86.070 201.420 ;
        RECT 98.230 201.160 98.490 201.420 ;
        RECT 100.990 201.160 101.250 201.420 ;
        RECT 106.050 201.160 106.310 201.420 ;
        RECT 106.510 201.160 106.770 201.420 ;
        RECT 113.870 201.160 114.130 201.420 ;
        RECT 119.850 201.160 120.110 201.420 ;
        RECT 74.930 200.650 75.190 200.910 ;
        RECT 75.250 200.650 75.510 200.910 ;
        RECT 75.570 200.650 75.830 200.910 ;
        RECT 75.890 200.650 76.150 200.910 ;
        RECT 76.210 200.650 76.470 200.910 ;
        RECT 93.440 200.650 93.700 200.910 ;
        RECT 93.760 200.650 94.020 200.910 ;
        RECT 94.080 200.650 94.340 200.910 ;
        RECT 94.400 200.650 94.660 200.910 ;
        RECT 94.720 200.650 94.980 200.910 ;
        RECT 111.950 200.650 112.210 200.910 ;
        RECT 112.270 200.650 112.530 200.910 ;
        RECT 112.590 200.650 112.850 200.910 ;
        RECT 112.910 200.650 113.170 200.910 ;
        RECT 113.230 200.650 113.490 200.910 ;
        RECT 130.460 200.650 130.720 200.910 ;
        RECT 130.780 200.650 131.040 200.910 ;
        RECT 131.100 200.650 131.360 200.910 ;
        RECT 131.420 200.650 131.680 200.910 ;
        RECT 131.740 200.650 132.000 200.910 ;
        RECT 61.890 200.140 62.150 200.400 ;
        RECT 74.310 200.140 74.570 200.400 ;
        RECT 97.770 200.140 98.030 200.400 ;
        RECT 98.230 200.140 98.490 200.400 ;
        RECT 77.070 199.800 77.330 200.060 ;
        RECT 76.610 199.460 76.870 199.720 ;
        RECT 77.530 199.460 77.790 199.720 ;
        RECT 77.070 198.780 77.330 199.040 ;
        RECT 81.210 199.460 81.470 199.720 ;
        RECT 81.670 199.460 81.930 199.720 ;
        RECT 89.950 199.460 90.210 199.720 ;
        RECT 92.250 199.460 92.510 199.720 ;
        RECT 101.450 199.800 101.710 200.060 ;
        RECT 96.390 199.460 96.650 199.720 ;
        RECT 80.290 198.780 80.550 199.040 ;
        RECT 82.590 198.780 82.850 199.040 ;
        RECT 86.270 199.120 86.530 199.380 ;
        RECT 87.190 198.780 87.450 199.040 ;
        RECT 102.830 200.140 103.090 200.400 ;
        RECT 106.050 200.140 106.310 200.400 ;
        RECT 123.530 200.140 123.790 200.400 ;
        RECT 119.850 199.460 120.110 199.720 ;
        RECT 111.110 199.120 111.370 199.380 ;
        RECT 113.410 199.120 113.670 199.380 ;
        RECT 83.510 198.440 83.770 198.700 ;
        RECT 91.330 198.440 91.590 198.700 ;
        RECT 100.990 198.440 101.250 198.700 ;
        RECT 101.910 198.440 102.170 198.700 ;
        RECT 106.510 198.440 106.770 198.700 ;
        RECT 120.770 198.440 121.030 198.700 ;
        RECT 65.675 197.930 65.935 198.190 ;
        RECT 65.995 197.930 66.255 198.190 ;
        RECT 66.315 197.930 66.575 198.190 ;
        RECT 66.635 197.930 66.895 198.190 ;
        RECT 66.955 197.930 67.215 198.190 ;
        RECT 84.185 197.930 84.445 198.190 ;
        RECT 84.505 197.930 84.765 198.190 ;
        RECT 84.825 197.930 85.085 198.190 ;
        RECT 85.145 197.930 85.405 198.190 ;
        RECT 85.465 197.930 85.725 198.190 ;
        RECT 102.695 197.930 102.955 198.190 ;
        RECT 103.015 197.930 103.275 198.190 ;
        RECT 103.335 197.930 103.595 198.190 ;
        RECT 103.655 197.930 103.915 198.190 ;
        RECT 103.975 197.930 104.235 198.190 ;
        RECT 121.205 197.930 121.465 198.190 ;
        RECT 121.525 197.930 121.785 198.190 ;
        RECT 121.845 197.930 122.105 198.190 ;
        RECT 122.165 197.930 122.425 198.190 ;
        RECT 122.485 197.930 122.745 198.190 ;
        RECT 74.310 197.420 74.570 197.680 ;
        RECT 77.070 197.420 77.330 197.680 ;
        RECT 81.670 197.420 81.930 197.680 ;
        RECT 85.810 197.420 86.070 197.680 ;
        RECT 80.290 196.740 80.550 197.000 ;
        RECT 77.990 196.400 78.250 196.660 ;
        RECT 80.750 196.400 81.010 196.660 ;
        RECT 81.210 195.720 81.470 195.980 ;
        RECT 83.510 195.720 83.770 195.980 ;
        RECT 86.270 196.400 86.530 196.660 ;
        RECT 90.410 197.420 90.670 197.680 ;
        RECT 91.330 197.080 91.590 197.340 ;
        RECT 92.250 197.420 92.510 197.680 ;
        RECT 96.390 197.420 96.650 197.680 ;
        RECT 101.450 197.420 101.710 197.680 ;
        RECT 106.510 197.420 106.770 197.680 ;
        RECT 111.570 197.420 111.830 197.680 ;
        RECT 116.630 197.420 116.890 197.680 ;
        RECT 88.110 195.720 88.370 195.980 ;
        RECT 95.470 196.400 95.730 196.660 ;
        RECT 97.770 196.400 98.030 196.660 ;
        RECT 101.910 196.740 102.170 197.000 ;
        RECT 128.130 197.080 128.390 197.340 ;
        RECT 114.330 196.740 114.590 197.000 ;
        RECT 116.630 196.740 116.890 197.000 ;
        RECT 113.870 196.400 114.130 196.660 ;
        RECT 120.770 196.740 121.030 197.000 ;
        RECT 103.290 196.060 103.550 196.320 ;
        RECT 110.650 196.060 110.910 196.320 ;
        RECT 104.670 195.720 104.930 195.980 ;
        RECT 115.710 195.720 115.970 195.980 ;
        RECT 120.770 195.720 121.030 195.980 ;
        RECT 74.930 195.210 75.190 195.470 ;
        RECT 75.250 195.210 75.510 195.470 ;
        RECT 75.570 195.210 75.830 195.470 ;
        RECT 75.890 195.210 76.150 195.470 ;
        RECT 76.210 195.210 76.470 195.470 ;
        RECT 93.440 195.210 93.700 195.470 ;
        RECT 93.760 195.210 94.020 195.470 ;
        RECT 94.080 195.210 94.340 195.470 ;
        RECT 94.400 195.210 94.660 195.470 ;
        RECT 94.720 195.210 94.980 195.470 ;
        RECT 111.950 195.210 112.210 195.470 ;
        RECT 112.270 195.210 112.530 195.470 ;
        RECT 112.590 195.210 112.850 195.470 ;
        RECT 112.910 195.210 113.170 195.470 ;
        RECT 113.230 195.210 113.490 195.470 ;
        RECT 130.460 195.210 130.720 195.470 ;
        RECT 130.780 195.210 131.040 195.470 ;
        RECT 131.100 195.210 131.360 195.470 ;
        RECT 131.420 195.210 131.680 195.470 ;
        RECT 131.740 195.210 132.000 195.470 ;
        RECT 77.530 194.700 77.790 194.960 ;
        RECT 110.650 194.700 110.910 194.960 ;
        RECT 115.710 194.700 115.970 194.960 ;
        RECT 104.670 194.360 104.930 194.620 ;
        RECT 81.210 194.020 81.470 194.280 ;
        RECT 91.330 194.020 91.590 194.280 ;
        RECT 103.290 194.020 103.550 194.280 ;
        RECT 108.810 194.020 109.070 194.280 ;
        RECT 80.290 193.680 80.550 193.940 ;
        RECT 78.450 193.340 78.710 193.600 ;
        RECT 113.870 193.680 114.130 193.940 ;
        RECT 108.810 193.340 109.070 193.600 ;
        RECT 89.950 193.000 90.210 193.260 ;
        RECT 93.630 193.000 93.890 193.260 ;
        RECT 115.710 193.000 115.970 193.260 ;
        RECT 65.675 192.490 65.935 192.750 ;
        RECT 65.995 192.490 66.255 192.750 ;
        RECT 66.315 192.490 66.575 192.750 ;
        RECT 66.635 192.490 66.895 192.750 ;
        RECT 66.955 192.490 67.215 192.750 ;
        RECT 84.185 192.490 84.445 192.750 ;
        RECT 84.505 192.490 84.765 192.750 ;
        RECT 84.825 192.490 85.085 192.750 ;
        RECT 85.145 192.490 85.405 192.750 ;
        RECT 85.465 192.490 85.725 192.750 ;
        RECT 102.695 192.490 102.955 192.750 ;
        RECT 103.015 192.490 103.275 192.750 ;
        RECT 103.335 192.490 103.595 192.750 ;
        RECT 103.655 192.490 103.915 192.750 ;
        RECT 103.975 192.490 104.235 192.750 ;
        RECT 121.205 192.490 121.465 192.750 ;
        RECT 121.525 192.490 121.785 192.750 ;
        RECT 121.845 192.490 122.105 192.750 ;
        RECT 122.165 192.490 122.425 192.750 ;
        RECT 122.485 192.490 122.745 192.750 ;
        RECT 77.990 191.980 78.250 192.240 ;
        RECT 78.450 191.980 78.710 192.240 ;
        RECT 80.290 191.980 80.550 192.240 ;
        RECT 88.110 191.980 88.370 192.240 ;
        RECT 108.810 191.980 109.070 192.240 ;
        RECT 89.950 191.300 90.210 191.560 ;
        RECT 80.750 190.960 81.010 191.220 ;
        RECT 83.970 190.960 84.230 191.220 ;
        RECT 89.490 190.960 89.750 191.220 ;
        RECT 111.110 190.960 111.370 191.220 ;
        RECT 115.710 190.960 115.970 191.220 ;
        RECT 88.110 190.280 88.370 190.540 ;
        RECT 93.630 190.620 93.890 190.880 ;
        RECT 101.450 190.620 101.710 190.880 ;
        RECT 120.770 190.620 121.030 190.880 ;
        RECT 96.390 190.280 96.650 190.540 ;
        RECT 74.930 189.770 75.190 190.030 ;
        RECT 75.250 189.770 75.510 190.030 ;
        RECT 75.570 189.770 75.830 190.030 ;
        RECT 75.890 189.770 76.150 190.030 ;
        RECT 76.210 189.770 76.470 190.030 ;
        RECT 93.440 189.770 93.700 190.030 ;
        RECT 93.760 189.770 94.020 190.030 ;
        RECT 94.080 189.770 94.340 190.030 ;
        RECT 94.400 189.770 94.660 190.030 ;
        RECT 94.720 189.770 94.980 190.030 ;
        RECT 111.950 189.770 112.210 190.030 ;
        RECT 112.270 189.770 112.530 190.030 ;
        RECT 112.590 189.770 112.850 190.030 ;
        RECT 112.910 189.770 113.170 190.030 ;
        RECT 113.230 189.770 113.490 190.030 ;
        RECT 130.460 189.770 130.720 190.030 ;
        RECT 130.780 189.770 131.040 190.030 ;
        RECT 131.100 189.770 131.360 190.030 ;
        RECT 131.420 189.770 131.680 190.030 ;
        RECT 131.740 189.770 132.000 190.030 ;
        RECT 77.990 189.260 78.250 189.520 ;
        RECT 81.210 189.260 81.470 189.520 ;
        RECT 89.950 189.260 90.210 189.520 ;
        RECT 90.410 189.260 90.670 189.520 ;
        RECT 95.470 189.260 95.730 189.520 ;
        RECT 96.390 188.580 96.650 188.840 ;
        RECT 101.450 189.260 101.710 189.520 ;
        RECT 100.990 188.580 101.250 188.840 ;
        RECT 123.530 188.580 123.790 188.840 ;
        RECT 83.510 187.560 83.770 187.820 ;
        RECT 89.490 187.560 89.750 187.820 ;
        RECT 128.130 187.560 128.390 187.820 ;
        RECT 65.675 187.050 65.935 187.310 ;
        RECT 65.995 187.050 66.255 187.310 ;
        RECT 66.315 187.050 66.575 187.310 ;
        RECT 66.635 187.050 66.895 187.310 ;
        RECT 66.955 187.050 67.215 187.310 ;
        RECT 84.185 187.050 84.445 187.310 ;
        RECT 84.505 187.050 84.765 187.310 ;
        RECT 84.825 187.050 85.085 187.310 ;
        RECT 85.145 187.050 85.405 187.310 ;
        RECT 85.465 187.050 85.725 187.310 ;
        RECT 102.695 187.050 102.955 187.310 ;
        RECT 103.015 187.050 103.275 187.310 ;
        RECT 103.335 187.050 103.595 187.310 ;
        RECT 103.655 187.050 103.915 187.310 ;
        RECT 103.975 187.050 104.235 187.310 ;
        RECT 121.205 187.050 121.465 187.310 ;
        RECT 121.525 187.050 121.785 187.310 ;
        RECT 121.845 187.050 122.105 187.310 ;
        RECT 122.165 187.050 122.425 187.310 ;
        RECT 122.485 187.050 122.745 187.310 ;
        RECT 74.930 184.330 75.190 184.590 ;
        RECT 75.250 184.330 75.510 184.590 ;
        RECT 75.570 184.330 75.830 184.590 ;
        RECT 75.890 184.330 76.150 184.590 ;
        RECT 76.210 184.330 76.470 184.590 ;
        RECT 93.440 184.330 93.700 184.590 ;
        RECT 93.760 184.330 94.020 184.590 ;
        RECT 94.080 184.330 94.340 184.590 ;
        RECT 94.400 184.330 94.660 184.590 ;
        RECT 94.720 184.330 94.980 184.590 ;
        RECT 111.950 184.330 112.210 184.590 ;
        RECT 112.270 184.330 112.530 184.590 ;
        RECT 112.590 184.330 112.850 184.590 ;
        RECT 112.910 184.330 113.170 184.590 ;
        RECT 113.230 184.330 113.490 184.590 ;
        RECT 130.460 184.330 130.720 184.590 ;
        RECT 130.780 184.330 131.040 184.590 ;
        RECT 131.100 184.330 131.360 184.590 ;
        RECT 131.420 184.330 131.680 184.590 ;
        RECT 131.740 184.330 132.000 184.590 ;
        RECT 65.675 181.610 65.935 181.870 ;
        RECT 65.995 181.610 66.255 181.870 ;
        RECT 66.315 181.610 66.575 181.870 ;
        RECT 66.635 181.610 66.895 181.870 ;
        RECT 66.955 181.610 67.215 181.870 ;
        RECT 84.185 181.610 84.445 181.870 ;
        RECT 84.505 181.610 84.765 181.870 ;
        RECT 84.825 181.610 85.085 181.870 ;
        RECT 85.145 181.610 85.405 181.870 ;
        RECT 85.465 181.610 85.725 181.870 ;
        RECT 102.695 181.610 102.955 181.870 ;
        RECT 103.015 181.610 103.275 181.870 ;
        RECT 103.335 181.610 103.595 181.870 ;
        RECT 103.655 181.610 103.915 181.870 ;
        RECT 103.975 181.610 104.235 181.870 ;
        RECT 121.205 181.610 121.465 181.870 ;
        RECT 121.525 181.610 121.785 181.870 ;
        RECT 121.845 181.610 122.105 181.870 ;
        RECT 122.165 181.610 122.425 181.870 ;
        RECT 122.485 181.610 122.745 181.870 ;
        RECT 74.930 178.890 75.190 179.150 ;
        RECT 75.250 178.890 75.510 179.150 ;
        RECT 75.570 178.890 75.830 179.150 ;
        RECT 75.890 178.890 76.150 179.150 ;
        RECT 76.210 178.890 76.470 179.150 ;
        RECT 93.440 178.890 93.700 179.150 ;
        RECT 93.760 178.890 94.020 179.150 ;
        RECT 94.080 178.890 94.340 179.150 ;
        RECT 94.400 178.890 94.660 179.150 ;
        RECT 94.720 178.890 94.980 179.150 ;
        RECT 111.950 178.890 112.210 179.150 ;
        RECT 112.270 178.890 112.530 179.150 ;
        RECT 112.590 178.890 112.850 179.150 ;
        RECT 112.910 178.890 113.170 179.150 ;
        RECT 113.230 178.890 113.490 179.150 ;
        RECT 130.460 178.890 130.720 179.150 ;
        RECT 130.780 178.890 131.040 179.150 ;
        RECT 131.100 178.890 131.360 179.150 ;
        RECT 131.420 178.890 131.680 179.150 ;
        RECT 131.740 178.890 132.000 179.150 ;
        RECT 65.675 176.170 65.935 176.430 ;
        RECT 65.995 176.170 66.255 176.430 ;
        RECT 66.315 176.170 66.575 176.430 ;
        RECT 66.635 176.170 66.895 176.430 ;
        RECT 66.955 176.170 67.215 176.430 ;
        RECT 84.185 176.170 84.445 176.430 ;
        RECT 84.505 176.170 84.765 176.430 ;
        RECT 84.825 176.170 85.085 176.430 ;
        RECT 85.145 176.170 85.405 176.430 ;
        RECT 85.465 176.170 85.725 176.430 ;
        RECT 102.695 176.170 102.955 176.430 ;
        RECT 103.015 176.170 103.275 176.430 ;
        RECT 103.335 176.170 103.595 176.430 ;
        RECT 103.655 176.170 103.915 176.430 ;
        RECT 103.975 176.170 104.235 176.430 ;
        RECT 121.205 176.170 121.465 176.430 ;
        RECT 121.525 176.170 121.785 176.430 ;
        RECT 121.845 176.170 122.105 176.430 ;
        RECT 122.165 176.170 122.425 176.430 ;
        RECT 122.485 176.170 122.745 176.430 ;
        RECT 74.930 173.450 75.190 173.710 ;
        RECT 75.250 173.450 75.510 173.710 ;
        RECT 75.570 173.450 75.830 173.710 ;
        RECT 75.890 173.450 76.150 173.710 ;
        RECT 76.210 173.450 76.470 173.710 ;
        RECT 93.440 173.450 93.700 173.710 ;
        RECT 93.760 173.450 94.020 173.710 ;
        RECT 94.080 173.450 94.340 173.710 ;
        RECT 94.400 173.450 94.660 173.710 ;
        RECT 94.720 173.450 94.980 173.710 ;
        RECT 111.950 173.450 112.210 173.710 ;
        RECT 112.270 173.450 112.530 173.710 ;
        RECT 112.590 173.450 112.850 173.710 ;
        RECT 112.910 173.450 113.170 173.710 ;
        RECT 113.230 173.450 113.490 173.710 ;
        RECT 130.460 173.450 130.720 173.710 ;
        RECT 130.780 173.450 131.040 173.710 ;
        RECT 131.100 173.450 131.360 173.710 ;
        RECT 131.420 173.450 131.680 173.710 ;
        RECT 131.740 173.450 132.000 173.710 ;
        RECT 65.675 170.730 65.935 170.990 ;
        RECT 65.995 170.730 66.255 170.990 ;
        RECT 66.315 170.730 66.575 170.990 ;
        RECT 66.635 170.730 66.895 170.990 ;
        RECT 66.955 170.730 67.215 170.990 ;
        RECT 84.185 170.730 84.445 170.990 ;
        RECT 84.505 170.730 84.765 170.990 ;
        RECT 84.825 170.730 85.085 170.990 ;
        RECT 85.145 170.730 85.405 170.990 ;
        RECT 85.465 170.730 85.725 170.990 ;
        RECT 102.695 170.730 102.955 170.990 ;
        RECT 103.015 170.730 103.275 170.990 ;
        RECT 103.335 170.730 103.595 170.990 ;
        RECT 103.655 170.730 103.915 170.990 ;
        RECT 103.975 170.730 104.235 170.990 ;
        RECT 121.205 170.730 121.465 170.990 ;
        RECT 121.525 170.730 121.785 170.990 ;
        RECT 121.845 170.730 122.105 170.990 ;
        RECT 122.165 170.730 122.425 170.990 ;
        RECT 122.485 170.730 122.745 170.990 ;
        RECT 74.930 168.010 75.190 168.270 ;
        RECT 75.250 168.010 75.510 168.270 ;
        RECT 75.570 168.010 75.830 168.270 ;
        RECT 75.890 168.010 76.150 168.270 ;
        RECT 76.210 168.010 76.470 168.270 ;
        RECT 93.440 168.010 93.700 168.270 ;
        RECT 93.760 168.010 94.020 168.270 ;
        RECT 94.080 168.010 94.340 168.270 ;
        RECT 94.400 168.010 94.660 168.270 ;
        RECT 94.720 168.010 94.980 168.270 ;
        RECT 111.950 168.010 112.210 168.270 ;
        RECT 112.270 168.010 112.530 168.270 ;
        RECT 112.590 168.010 112.850 168.270 ;
        RECT 112.910 168.010 113.170 168.270 ;
        RECT 113.230 168.010 113.490 168.270 ;
        RECT 130.460 168.010 130.720 168.270 ;
        RECT 130.780 168.010 131.040 168.270 ;
        RECT 131.100 168.010 131.360 168.270 ;
        RECT 131.420 168.010 131.680 168.270 ;
        RECT 131.740 168.010 132.000 168.270 ;
        RECT 65.675 165.290 65.935 165.550 ;
        RECT 65.995 165.290 66.255 165.550 ;
        RECT 66.315 165.290 66.575 165.550 ;
        RECT 66.635 165.290 66.895 165.550 ;
        RECT 66.955 165.290 67.215 165.550 ;
        RECT 84.185 165.290 84.445 165.550 ;
        RECT 84.505 165.290 84.765 165.550 ;
        RECT 84.825 165.290 85.085 165.550 ;
        RECT 85.145 165.290 85.405 165.550 ;
        RECT 85.465 165.290 85.725 165.550 ;
        RECT 102.695 165.290 102.955 165.550 ;
        RECT 103.015 165.290 103.275 165.550 ;
        RECT 103.335 165.290 103.595 165.550 ;
        RECT 103.655 165.290 103.915 165.550 ;
        RECT 103.975 165.290 104.235 165.550 ;
        RECT 121.205 165.290 121.465 165.550 ;
        RECT 121.525 165.290 121.785 165.550 ;
        RECT 121.845 165.290 122.105 165.550 ;
        RECT 122.165 165.290 122.425 165.550 ;
        RECT 122.485 165.290 122.745 165.550 ;
        RECT 74.930 162.570 75.190 162.830 ;
        RECT 75.250 162.570 75.510 162.830 ;
        RECT 75.570 162.570 75.830 162.830 ;
        RECT 75.890 162.570 76.150 162.830 ;
        RECT 76.210 162.570 76.470 162.830 ;
        RECT 93.440 162.570 93.700 162.830 ;
        RECT 93.760 162.570 94.020 162.830 ;
        RECT 94.080 162.570 94.340 162.830 ;
        RECT 94.400 162.570 94.660 162.830 ;
        RECT 94.720 162.570 94.980 162.830 ;
        RECT 111.950 162.570 112.210 162.830 ;
        RECT 112.270 162.570 112.530 162.830 ;
        RECT 112.590 162.570 112.850 162.830 ;
        RECT 112.910 162.570 113.170 162.830 ;
        RECT 113.230 162.570 113.490 162.830 ;
        RECT 130.460 162.570 130.720 162.830 ;
        RECT 130.780 162.570 131.040 162.830 ;
        RECT 131.100 162.570 131.360 162.830 ;
        RECT 131.420 162.570 131.680 162.830 ;
        RECT 131.740 162.570 132.000 162.830 ;
        RECT 65.675 159.850 65.935 160.110 ;
        RECT 65.995 159.850 66.255 160.110 ;
        RECT 66.315 159.850 66.575 160.110 ;
        RECT 66.635 159.850 66.895 160.110 ;
        RECT 66.955 159.850 67.215 160.110 ;
        RECT 84.185 159.850 84.445 160.110 ;
        RECT 84.505 159.850 84.765 160.110 ;
        RECT 84.825 159.850 85.085 160.110 ;
        RECT 85.145 159.850 85.405 160.110 ;
        RECT 85.465 159.850 85.725 160.110 ;
        RECT 102.695 159.850 102.955 160.110 ;
        RECT 103.015 159.850 103.275 160.110 ;
        RECT 103.335 159.850 103.595 160.110 ;
        RECT 103.655 159.850 103.915 160.110 ;
        RECT 103.975 159.850 104.235 160.110 ;
        RECT 121.205 159.850 121.465 160.110 ;
        RECT 121.525 159.850 121.785 160.110 ;
        RECT 121.845 159.850 122.105 160.110 ;
        RECT 122.165 159.850 122.425 160.110 ;
        RECT 122.485 159.850 122.745 160.110 ;
        RECT 74.930 157.130 75.190 157.390 ;
        RECT 75.250 157.130 75.510 157.390 ;
        RECT 75.570 157.130 75.830 157.390 ;
        RECT 75.890 157.130 76.150 157.390 ;
        RECT 76.210 157.130 76.470 157.390 ;
        RECT 93.440 157.130 93.700 157.390 ;
        RECT 93.760 157.130 94.020 157.390 ;
        RECT 94.080 157.130 94.340 157.390 ;
        RECT 94.400 157.130 94.660 157.390 ;
        RECT 94.720 157.130 94.980 157.390 ;
        RECT 111.950 157.130 112.210 157.390 ;
        RECT 112.270 157.130 112.530 157.390 ;
        RECT 112.590 157.130 112.850 157.390 ;
        RECT 112.910 157.130 113.170 157.390 ;
        RECT 113.230 157.130 113.490 157.390 ;
        RECT 130.460 157.130 130.720 157.390 ;
        RECT 130.780 157.130 131.040 157.390 ;
        RECT 131.100 157.130 131.360 157.390 ;
        RECT 131.420 157.130 131.680 157.390 ;
        RECT 131.740 157.130 132.000 157.390 ;
        RECT 65.675 154.410 65.935 154.670 ;
        RECT 65.995 154.410 66.255 154.670 ;
        RECT 66.315 154.410 66.575 154.670 ;
        RECT 66.635 154.410 66.895 154.670 ;
        RECT 66.955 154.410 67.215 154.670 ;
        RECT 84.185 154.410 84.445 154.670 ;
        RECT 84.505 154.410 84.765 154.670 ;
        RECT 84.825 154.410 85.085 154.670 ;
        RECT 85.145 154.410 85.405 154.670 ;
        RECT 85.465 154.410 85.725 154.670 ;
        RECT 102.695 154.410 102.955 154.670 ;
        RECT 103.015 154.410 103.275 154.670 ;
        RECT 103.335 154.410 103.595 154.670 ;
        RECT 103.655 154.410 103.915 154.670 ;
        RECT 103.975 154.410 104.235 154.670 ;
        RECT 121.205 154.410 121.465 154.670 ;
        RECT 121.525 154.410 121.785 154.670 ;
        RECT 121.845 154.410 122.105 154.670 ;
        RECT 122.165 154.410 122.425 154.670 ;
        RECT 122.485 154.410 122.745 154.670 ;
        RECT 74.930 151.690 75.190 151.950 ;
        RECT 75.250 151.690 75.510 151.950 ;
        RECT 75.570 151.690 75.830 151.950 ;
        RECT 75.890 151.690 76.150 151.950 ;
        RECT 76.210 151.690 76.470 151.950 ;
        RECT 93.440 151.690 93.700 151.950 ;
        RECT 93.760 151.690 94.020 151.950 ;
        RECT 94.080 151.690 94.340 151.950 ;
        RECT 94.400 151.690 94.660 151.950 ;
        RECT 94.720 151.690 94.980 151.950 ;
        RECT 111.950 151.690 112.210 151.950 ;
        RECT 112.270 151.690 112.530 151.950 ;
        RECT 112.590 151.690 112.850 151.950 ;
        RECT 112.910 151.690 113.170 151.950 ;
        RECT 113.230 151.690 113.490 151.950 ;
        RECT 130.460 151.690 130.720 151.950 ;
        RECT 130.780 151.690 131.040 151.950 ;
        RECT 131.100 151.690 131.360 151.950 ;
        RECT 131.420 151.690 131.680 151.950 ;
        RECT 131.740 151.690 132.000 151.950 ;
        RECT 111.110 150.840 111.370 151.100 ;
        RECT 110.650 149.480 110.910 149.740 ;
        RECT 65.675 148.970 65.935 149.230 ;
        RECT 65.995 148.970 66.255 149.230 ;
        RECT 66.315 148.970 66.575 149.230 ;
        RECT 66.635 148.970 66.895 149.230 ;
        RECT 66.955 148.970 67.215 149.230 ;
        RECT 84.185 148.970 84.445 149.230 ;
        RECT 84.505 148.970 84.765 149.230 ;
        RECT 84.825 148.970 85.085 149.230 ;
        RECT 85.145 148.970 85.405 149.230 ;
        RECT 85.465 148.970 85.725 149.230 ;
        RECT 102.695 148.970 102.955 149.230 ;
        RECT 103.015 148.970 103.275 149.230 ;
        RECT 103.335 148.970 103.595 149.230 ;
        RECT 103.655 148.970 103.915 149.230 ;
        RECT 103.975 148.970 104.235 149.230 ;
        RECT 121.205 148.970 121.465 149.230 ;
        RECT 121.525 148.970 121.785 149.230 ;
        RECT 121.845 148.970 122.105 149.230 ;
        RECT 122.165 148.970 122.425 149.230 ;
        RECT 122.485 148.970 122.745 149.230 ;
        RECT 74.930 146.250 75.190 146.510 ;
        RECT 75.250 146.250 75.510 146.510 ;
        RECT 75.570 146.250 75.830 146.510 ;
        RECT 75.890 146.250 76.150 146.510 ;
        RECT 76.210 146.250 76.470 146.510 ;
        RECT 93.440 146.250 93.700 146.510 ;
        RECT 93.760 146.250 94.020 146.510 ;
        RECT 94.080 146.250 94.340 146.510 ;
        RECT 94.400 146.250 94.660 146.510 ;
        RECT 94.720 146.250 94.980 146.510 ;
        RECT 111.950 146.250 112.210 146.510 ;
        RECT 112.270 146.250 112.530 146.510 ;
        RECT 112.590 146.250 112.850 146.510 ;
        RECT 112.910 146.250 113.170 146.510 ;
        RECT 113.230 146.250 113.490 146.510 ;
        RECT 130.460 146.250 130.720 146.510 ;
        RECT 130.780 146.250 131.040 146.510 ;
        RECT 131.100 146.250 131.360 146.510 ;
        RECT 131.420 146.250 131.680 146.510 ;
        RECT 131.740 146.250 132.000 146.510 ;
        RECT 65.675 143.530 65.935 143.790 ;
        RECT 65.995 143.530 66.255 143.790 ;
        RECT 66.315 143.530 66.575 143.790 ;
        RECT 66.635 143.530 66.895 143.790 ;
        RECT 66.955 143.530 67.215 143.790 ;
        RECT 84.185 143.530 84.445 143.790 ;
        RECT 84.505 143.530 84.765 143.790 ;
        RECT 84.825 143.530 85.085 143.790 ;
        RECT 85.145 143.530 85.405 143.790 ;
        RECT 85.465 143.530 85.725 143.790 ;
        RECT 102.695 143.530 102.955 143.790 ;
        RECT 103.015 143.530 103.275 143.790 ;
        RECT 103.335 143.530 103.595 143.790 ;
        RECT 103.655 143.530 103.915 143.790 ;
        RECT 103.975 143.530 104.235 143.790 ;
        RECT 121.205 143.530 121.465 143.790 ;
        RECT 121.525 143.530 121.785 143.790 ;
        RECT 121.845 143.530 122.105 143.790 ;
        RECT 122.165 143.530 122.425 143.790 ;
        RECT 122.485 143.530 122.745 143.790 ;
        RECT 74.930 140.810 75.190 141.070 ;
        RECT 75.250 140.810 75.510 141.070 ;
        RECT 75.570 140.810 75.830 141.070 ;
        RECT 75.890 140.810 76.150 141.070 ;
        RECT 76.210 140.810 76.470 141.070 ;
        RECT 93.440 140.810 93.700 141.070 ;
        RECT 93.760 140.810 94.020 141.070 ;
        RECT 94.080 140.810 94.340 141.070 ;
        RECT 94.400 140.810 94.660 141.070 ;
        RECT 94.720 140.810 94.980 141.070 ;
        RECT 111.950 140.810 112.210 141.070 ;
        RECT 112.270 140.810 112.530 141.070 ;
        RECT 112.590 140.810 112.850 141.070 ;
        RECT 112.910 140.810 113.170 141.070 ;
        RECT 113.230 140.810 113.490 141.070 ;
        RECT 130.460 140.810 130.720 141.070 ;
        RECT 130.780 140.810 131.040 141.070 ;
        RECT 131.100 140.810 131.360 141.070 ;
        RECT 131.420 140.810 131.680 141.070 ;
        RECT 131.740 140.810 132.000 141.070 ;
        RECT 65.675 138.090 65.935 138.350 ;
        RECT 65.995 138.090 66.255 138.350 ;
        RECT 66.315 138.090 66.575 138.350 ;
        RECT 66.635 138.090 66.895 138.350 ;
        RECT 66.955 138.090 67.215 138.350 ;
        RECT 84.185 138.090 84.445 138.350 ;
        RECT 84.505 138.090 84.765 138.350 ;
        RECT 84.825 138.090 85.085 138.350 ;
        RECT 85.145 138.090 85.405 138.350 ;
        RECT 85.465 138.090 85.725 138.350 ;
        RECT 102.695 138.090 102.955 138.350 ;
        RECT 103.015 138.090 103.275 138.350 ;
        RECT 103.335 138.090 103.595 138.350 ;
        RECT 103.655 138.090 103.915 138.350 ;
        RECT 103.975 138.090 104.235 138.350 ;
        RECT 121.205 138.090 121.465 138.350 ;
        RECT 121.525 138.090 121.785 138.350 ;
        RECT 121.845 138.090 122.105 138.350 ;
        RECT 122.165 138.090 122.425 138.350 ;
        RECT 122.485 138.090 122.745 138.350 ;
        RECT 74.930 135.370 75.190 135.630 ;
        RECT 75.250 135.370 75.510 135.630 ;
        RECT 75.570 135.370 75.830 135.630 ;
        RECT 75.890 135.370 76.150 135.630 ;
        RECT 76.210 135.370 76.470 135.630 ;
        RECT 93.440 135.370 93.700 135.630 ;
        RECT 93.760 135.370 94.020 135.630 ;
        RECT 94.080 135.370 94.340 135.630 ;
        RECT 94.400 135.370 94.660 135.630 ;
        RECT 94.720 135.370 94.980 135.630 ;
        RECT 111.950 135.370 112.210 135.630 ;
        RECT 112.270 135.370 112.530 135.630 ;
        RECT 112.590 135.370 112.850 135.630 ;
        RECT 112.910 135.370 113.170 135.630 ;
        RECT 113.230 135.370 113.490 135.630 ;
        RECT 130.460 135.370 130.720 135.630 ;
        RECT 130.780 135.370 131.040 135.630 ;
        RECT 131.100 135.370 131.360 135.630 ;
        RECT 131.420 135.370 131.680 135.630 ;
        RECT 131.740 135.370 132.000 135.630 ;
        RECT 65.675 132.650 65.935 132.910 ;
        RECT 65.995 132.650 66.255 132.910 ;
        RECT 66.315 132.650 66.575 132.910 ;
        RECT 66.635 132.650 66.895 132.910 ;
        RECT 66.955 132.650 67.215 132.910 ;
        RECT 84.185 132.650 84.445 132.910 ;
        RECT 84.505 132.650 84.765 132.910 ;
        RECT 84.825 132.650 85.085 132.910 ;
        RECT 85.145 132.650 85.405 132.910 ;
        RECT 85.465 132.650 85.725 132.910 ;
        RECT 102.695 132.650 102.955 132.910 ;
        RECT 103.015 132.650 103.275 132.910 ;
        RECT 103.335 132.650 103.595 132.910 ;
        RECT 103.655 132.650 103.915 132.910 ;
        RECT 103.975 132.650 104.235 132.910 ;
        RECT 121.205 132.650 121.465 132.910 ;
        RECT 121.525 132.650 121.785 132.910 ;
        RECT 121.845 132.650 122.105 132.910 ;
        RECT 122.165 132.650 122.425 132.910 ;
        RECT 122.485 132.650 122.745 132.910 ;
        RECT 74.930 129.930 75.190 130.190 ;
        RECT 75.250 129.930 75.510 130.190 ;
        RECT 75.570 129.930 75.830 130.190 ;
        RECT 75.890 129.930 76.150 130.190 ;
        RECT 76.210 129.930 76.470 130.190 ;
        RECT 93.440 129.930 93.700 130.190 ;
        RECT 93.760 129.930 94.020 130.190 ;
        RECT 94.080 129.930 94.340 130.190 ;
        RECT 94.400 129.930 94.660 130.190 ;
        RECT 94.720 129.930 94.980 130.190 ;
        RECT 111.950 129.930 112.210 130.190 ;
        RECT 112.270 129.930 112.530 130.190 ;
        RECT 112.590 129.930 112.850 130.190 ;
        RECT 112.910 129.930 113.170 130.190 ;
        RECT 113.230 129.930 113.490 130.190 ;
        RECT 130.460 129.930 130.720 130.190 ;
        RECT 130.780 129.930 131.040 130.190 ;
        RECT 131.100 129.930 131.360 130.190 ;
        RECT 131.420 129.930 131.680 130.190 ;
        RECT 131.740 129.930 132.000 130.190 ;
        RECT 141.000 99.000 142.000 101.000 ;
        RECT 141.000 95.000 142.000 97.000 ;
        RECT 144.270 91.670 144.920 92.420 ;
        RECT 148.220 91.640 148.960 92.460 ;
        RECT 124.000 88.000 125.000 90.000 ;
        RECT 138.570 86.620 140.120 87.020 ;
        RECT 141.420 85.520 143.420 85.970 ;
        RECT 148.220 87.220 149.020 87.870 ;
        RECT 150.920 86.670 152.520 86.970 ;
        RECT 147.920 84.620 150.020 85.020 ;
        RECT 144.920 84.170 145.220 84.470 ;
        RECT 135.000 82.000 136.000 84.000 ;
        RECT 138.820 82.570 139.120 83.420 ;
        RECT 140.120 82.570 140.520 83.420 ;
        RECT 142.770 82.620 143.120 83.370 ;
        RECT 139.470 81.720 139.770 82.270 ;
        RECT 144.120 82.620 144.420 83.370 ;
        RECT 143.470 81.720 143.770 82.270 ;
        RECT 145.320 81.170 145.620 81.520 ;
        RECT 147.820 82.620 148.120 83.370 ;
        RECT 149.120 82.620 149.470 83.370 ;
        RECT 151.820 82.620 152.120 83.370 ;
        RECT 148.470 81.670 148.820 82.320 ;
        RECT 153.120 82.620 153.470 83.370 ;
        RECT 152.470 81.670 152.770 82.320 ;
        RECT 156.000 82.000 157.000 84.000 ;
        RECT 147.920 80.220 148.470 80.570 ;
        RECT 145.270 79.520 145.620 79.820 ;
        RECT 130.000 77.000 132.000 78.000 ;
        RECT 140.820 76.670 141.120 77.370 ;
        RECT 142.170 76.670 142.470 77.370 ;
        RECT 145.770 77.020 146.470 77.620 ;
        RECT 149.820 76.670 150.120 77.320 ;
        RECT 141.470 75.670 141.770 76.370 ;
        RECT 145.820 75.720 146.420 76.370 ;
        RECT 151.170 76.670 151.470 77.320 ;
        RECT 160.000 77.000 162.000 78.000 ;
        RECT 150.470 75.720 150.770 76.370 ;
        RECT 124.000 71.000 125.000 73.000 ;
        RECT 145.770 72.670 146.470 73.420 ;
      LAYER met2 ;
        RECT 129.000 215.500 129.500 215.550 ;
        RECT 60.500 215.000 129.500 215.500 ;
        RECT 60.500 207.000 61.000 215.000 ;
        RECT 129.000 214.950 129.500 215.000 ;
        RECT 133.000 214.500 133.500 214.550 ;
        RECT 70.000 214.000 133.500 214.500 ;
        RECT 70.000 207.000 70.500 214.000 ;
        RECT 133.000 213.950 133.500 214.000 ;
        RECT 136.500 213.500 137.000 213.550 ;
        RECT 79.500 213.000 137.000 213.500 ;
        RECT 79.500 207.000 80.500 213.000 ;
        RECT 136.500 212.950 137.000 213.000 ;
        RECT 140.000 212.500 140.500 212.550 ;
        RECT 89.500 212.000 140.500 212.500 ;
        RECT 89.500 207.340 90.000 212.000 ;
        RECT 140.000 211.950 140.500 212.000 ;
        RECT 144.000 211.500 144.500 211.550 ;
        RECT 89.480 207.000 90.000 207.340 ;
        RECT 99.000 211.000 144.500 211.500 ;
        RECT 99.000 207.000 99.500 211.000 ;
        RECT 144.000 210.950 144.500 211.000 ;
        RECT 147.500 210.500 148.000 210.550 ;
        RECT 108.500 210.000 148.000 210.500 ;
        RECT 108.500 207.000 109.500 210.000 ;
        RECT 147.500 209.950 148.000 210.000 ;
        RECT 151.000 209.500 151.500 209.550 ;
        RECT 118.500 209.000 151.500 209.500 ;
        RECT 118.500 207.340 119.000 209.000 ;
        RECT 151.000 208.950 151.500 209.000 ;
        RECT 154.745 208.335 155.280 208.355 ;
        RECT 118.460 207.000 119.000 207.340 ;
        RECT 128.120 207.750 155.305 208.335 ;
        RECT 60.500 205.340 60.780 207.000 ;
        RECT 70.160 205.340 70.440 207.000 ;
        RECT 79.820 205.340 80.100 207.000 ;
        RECT 89.480 205.950 89.760 207.000 ;
        RECT 99.140 205.950 99.420 207.000 ;
        RECT 89.480 205.810 90.150 205.950 ;
        RECT 89.480 205.340 89.760 205.810 ;
        RECT 60.570 202.130 60.710 205.340 ;
        RECT 65.675 203.315 67.215 203.685 ;
        RECT 70.230 202.130 70.370 205.340 ;
        RECT 79.890 202.130 80.030 205.340 ;
        RECT 84.185 203.315 85.725 203.685 ;
        RECT 90.010 202.130 90.150 205.810 ;
        RECT 98.290 205.810 99.420 205.950 ;
        RECT 98.290 202.130 98.430 205.810 ;
        RECT 99.140 205.340 99.420 205.810 ;
        RECT 108.800 205.950 109.080 207.000 ;
        RECT 108.800 205.810 109.470 205.950 ;
        RECT 108.800 205.340 109.080 205.810 ;
        RECT 102.695 203.315 104.235 203.685 ;
        RECT 101.450 202.830 101.710 203.150 ;
        RECT 60.510 201.810 60.770 202.130 ;
        RECT 70.170 201.810 70.430 202.130 ;
        RECT 79.830 201.810 80.090 202.130 ;
        RECT 87.190 201.810 87.450 202.130 ;
        RECT 89.950 201.810 90.210 202.130 ;
        RECT 98.230 201.810 98.490 202.130 ;
        RECT 77.070 201.470 77.330 201.790 ;
        RECT 82.590 201.470 82.850 201.790 ;
        RECT 61.890 201.130 62.150 201.450 ;
        RECT 74.310 201.130 74.570 201.450 ;
        RECT 76.610 201.130 76.870 201.450 ;
        RECT 61.950 200.430 62.090 201.130 ;
        RECT 74.370 200.430 74.510 201.130 ;
        RECT 74.930 200.595 76.470 200.965 ;
        RECT 61.890 200.110 62.150 200.430 ;
        RECT 74.310 200.110 74.570 200.430 ;
        RECT 65.675 197.875 67.215 198.245 ;
        RECT 74.370 197.710 74.510 200.110 ;
        RECT 76.670 199.750 76.810 201.130 ;
        RECT 77.130 200.090 77.270 201.470 ;
        RECT 77.990 201.130 78.250 201.450 ;
        RECT 77.070 199.770 77.330 200.090 ;
        RECT 76.610 199.430 76.870 199.750 ;
        RECT 77.530 199.430 77.790 199.750 ;
        RECT 77.070 198.750 77.330 199.070 ;
        RECT 77.130 197.710 77.270 198.750 ;
        RECT 74.310 197.390 74.570 197.710 ;
        RECT 77.070 197.390 77.330 197.710 ;
        RECT 74.930 195.155 76.470 195.525 ;
        RECT 77.590 194.990 77.730 199.430 ;
        RECT 78.050 196.690 78.190 201.130 ;
        RECT 81.210 199.430 81.470 199.750 ;
        RECT 81.670 199.430 81.930 199.750 ;
        RECT 80.290 198.750 80.550 199.070 ;
        RECT 80.350 197.030 80.490 198.750 ;
        RECT 81.270 198.470 81.410 199.430 ;
        RECT 80.810 198.330 81.410 198.470 ;
        RECT 80.290 196.710 80.550 197.030 ;
        RECT 80.810 196.690 80.950 198.330 ;
        RECT 81.730 197.710 81.870 199.430 ;
        RECT 82.650 199.070 82.790 201.470 ;
        RECT 85.810 201.130 86.070 201.450 ;
        RECT 82.590 198.750 82.850 199.070 ;
        RECT 83.510 198.410 83.770 198.730 ;
        RECT 81.670 197.390 81.930 197.710 ;
        RECT 77.990 196.370 78.250 196.690 ;
        RECT 80.750 196.370 81.010 196.690 ;
        RECT 77.530 194.670 77.790 194.990 ;
        RECT 65.675 192.435 67.215 192.805 ;
        RECT 78.050 192.270 78.190 196.370 ;
        RECT 80.290 193.650 80.550 193.970 ;
        RECT 78.450 193.310 78.710 193.630 ;
        RECT 78.510 192.270 78.650 193.310 ;
        RECT 80.350 192.270 80.490 193.650 ;
        RECT 77.990 191.950 78.250 192.270 ;
        RECT 78.450 191.950 78.710 192.270 ;
        RECT 80.290 191.950 80.550 192.270 ;
        RECT 74.930 189.715 76.470 190.085 ;
        RECT 78.050 189.550 78.190 191.950 ;
        RECT 80.810 191.250 80.950 196.370 ;
        RECT 83.570 196.010 83.710 198.410 ;
        RECT 84.185 197.875 85.725 198.245 ;
        RECT 85.870 197.710 86.010 201.130 ;
        RECT 86.270 199.090 86.530 199.410 ;
        RECT 85.810 197.390 86.070 197.710 ;
        RECT 86.330 196.690 86.470 199.090 ;
        RECT 87.250 199.070 87.390 201.810 ;
        RECT 98.230 201.130 98.490 201.450 ;
        RECT 100.990 201.130 101.250 201.450 ;
        RECT 93.440 200.595 94.980 200.965 ;
        RECT 98.290 200.430 98.430 201.130 ;
        RECT 97.770 200.110 98.030 200.430 ;
        RECT 98.230 200.110 98.490 200.430 ;
        RECT 89.950 199.430 90.210 199.750 ;
        RECT 92.250 199.430 92.510 199.750 ;
        RECT 96.390 199.430 96.650 199.750 ;
        RECT 87.190 198.750 87.450 199.070 ;
        RECT 86.270 196.370 86.530 196.690 ;
        RECT 81.210 195.690 81.470 196.010 ;
        RECT 83.510 195.690 83.770 196.010 ;
        RECT 88.110 195.690 88.370 196.010 ;
        RECT 81.270 194.310 81.410 195.690 ;
        RECT 81.210 193.990 81.470 194.310 ;
        RECT 80.750 190.930 81.010 191.250 ;
        RECT 81.270 189.550 81.410 193.990 ;
        RECT 84.185 192.435 85.725 192.805 ;
        RECT 88.170 192.270 88.310 195.690 ;
        RECT 90.010 193.290 90.150 199.430 ;
        RECT 91.330 198.410 91.590 198.730 ;
        RECT 90.410 197.390 90.670 197.710 ;
        RECT 89.950 192.970 90.210 193.290 ;
        RECT 88.110 191.950 88.370 192.270 ;
        RECT 83.970 190.930 84.230 191.250 ;
        RECT 77.990 189.230 78.250 189.550 ;
        RECT 81.210 189.230 81.470 189.550 ;
        RECT 84.030 189.510 84.170 190.930 ;
        RECT 88.170 190.570 88.310 191.950 ;
        RECT 90.010 191.590 90.150 192.970 ;
        RECT 89.950 191.270 90.210 191.590 ;
        RECT 89.490 190.930 89.750 191.250 ;
        RECT 90.470 190.990 90.610 197.390 ;
        RECT 91.390 197.370 91.530 198.410 ;
        RECT 92.310 197.710 92.450 199.430 ;
        RECT 96.450 197.710 96.590 199.430 ;
        RECT 92.250 197.390 92.510 197.710 ;
        RECT 96.390 197.390 96.650 197.710 ;
        RECT 91.330 197.050 91.590 197.370 ;
        RECT 97.830 196.690 97.970 200.110 ;
        RECT 101.050 198.730 101.190 201.130 ;
        RECT 101.510 200.090 101.650 202.830 ;
        RECT 109.330 202.470 109.470 205.810 ;
        RECT 118.460 205.340 118.740 207.000 ;
        RECT 128.120 205.340 128.400 207.750 ;
        RECT 154.745 207.730 155.280 207.750 ;
        RECT 109.270 202.150 109.530 202.470 ;
        RECT 118.530 202.130 118.670 205.340 ;
        RECT 121.205 203.315 122.745 203.685 ;
        RECT 102.830 201.810 103.090 202.130 ;
        RECT 116.630 201.810 116.890 202.130 ;
        RECT 118.470 201.810 118.730 202.130 ;
        RECT 102.890 200.430 103.030 201.810 ;
        RECT 114.330 201.470 114.590 201.790 ;
        RECT 106.050 201.130 106.310 201.450 ;
        RECT 106.510 201.130 106.770 201.450 ;
        RECT 113.870 201.130 114.130 201.450 ;
        RECT 106.110 200.430 106.250 201.130 ;
        RECT 102.830 200.110 103.090 200.430 ;
        RECT 106.050 200.110 106.310 200.430 ;
        RECT 101.450 199.770 101.710 200.090 ;
        RECT 100.990 198.410 101.250 198.730 ;
        RECT 95.470 196.370 95.730 196.690 ;
        RECT 97.770 196.370 98.030 196.690 ;
        RECT 93.440 195.155 94.980 195.525 ;
        RECT 91.330 193.990 91.590 194.310 ;
        RECT 88.110 190.250 88.370 190.570 ;
        RECT 83.570 189.370 84.170 189.510 ;
        RECT 83.570 187.850 83.710 189.370 ;
        RECT 89.550 187.850 89.690 190.930 ;
        RECT 90.010 190.850 90.610 190.990 ;
        RECT 90.010 189.550 90.150 190.850 ;
        RECT 91.390 189.630 91.530 193.990 ;
        RECT 93.630 192.970 93.890 193.290 ;
        RECT 93.690 190.910 93.830 192.970 ;
        RECT 93.630 190.590 93.890 190.910 ;
        RECT 93.440 189.715 94.980 190.085 ;
        RECT 90.470 189.550 91.530 189.630 ;
        RECT 95.530 189.550 95.670 196.370 ;
        RECT 96.390 190.250 96.650 190.570 ;
        RECT 89.950 189.230 90.210 189.550 ;
        RECT 90.410 189.490 91.530 189.550 ;
        RECT 90.410 189.230 90.670 189.490 ;
        RECT 95.470 189.230 95.730 189.550 ;
        RECT 96.450 188.870 96.590 190.250 ;
        RECT 101.050 188.870 101.190 198.410 ;
        RECT 101.510 197.710 101.650 199.770 ;
        RECT 106.570 198.730 106.710 201.130 ;
        RECT 111.950 200.595 113.490 200.965 ;
        RECT 113.930 199.830 114.070 201.130 ;
        RECT 113.470 199.690 114.070 199.830 ;
        RECT 113.470 199.410 113.610 199.690 ;
        RECT 111.110 199.090 111.370 199.410 ;
        RECT 113.410 199.090 113.670 199.410 ;
        RECT 101.910 198.410 102.170 198.730 ;
        RECT 106.510 198.410 106.770 198.730 ;
        RECT 101.450 197.390 101.710 197.710 ;
        RECT 101.970 197.030 102.110 198.410 ;
        RECT 102.695 197.875 104.235 198.245 ;
        RECT 106.570 197.710 106.710 198.410 ;
        RECT 106.510 197.390 106.770 197.710 ;
        RECT 101.910 196.710 102.170 197.030 ;
        RECT 103.290 196.030 103.550 196.350 ;
        RECT 110.650 196.030 110.910 196.350 ;
        RECT 103.350 194.310 103.490 196.030 ;
        RECT 104.670 195.690 104.930 196.010 ;
        RECT 104.730 194.650 104.870 195.690 ;
        RECT 110.710 194.990 110.850 196.030 ;
        RECT 110.650 194.670 110.910 194.990 ;
        RECT 104.670 194.330 104.930 194.650 ;
        RECT 103.290 193.990 103.550 194.310 ;
        RECT 108.810 193.990 109.070 194.310 ;
        RECT 108.870 193.630 109.010 193.990 ;
        RECT 108.810 193.310 109.070 193.630 ;
        RECT 102.695 192.435 104.235 192.805 ;
        RECT 108.870 192.270 109.010 193.310 ;
        RECT 108.810 191.950 109.070 192.270 ;
        RECT 111.170 191.250 111.310 199.090 ;
        RECT 111.570 197.390 111.830 197.710 ;
        RECT 111.110 190.930 111.370 191.250 ;
        RECT 101.450 190.590 101.710 190.910 ;
        RECT 101.510 189.550 101.650 190.590 ;
        RECT 101.450 189.230 101.710 189.550 ;
        RECT 96.390 188.550 96.650 188.870 ;
        RECT 100.990 188.550 101.250 188.870 ;
        RECT 83.510 187.530 83.770 187.850 ;
        RECT 89.490 187.530 89.750 187.850 ;
        RECT 65.675 186.995 67.215 187.365 ;
        RECT 84.185 186.995 85.725 187.365 ;
        RECT 102.695 186.995 104.235 187.365 ;
        RECT 74.930 184.275 76.470 184.645 ;
        RECT 93.440 184.275 94.980 184.645 ;
        RECT 65.675 181.555 67.215 181.925 ;
        RECT 84.185 181.555 85.725 181.925 ;
        RECT 102.695 181.555 104.235 181.925 ;
        RECT 74.930 178.835 76.470 179.205 ;
        RECT 93.440 178.835 94.980 179.205 ;
        RECT 65.675 176.115 67.215 176.485 ;
        RECT 84.185 176.115 85.725 176.485 ;
        RECT 102.695 176.115 104.235 176.485 ;
        RECT 74.930 173.395 76.470 173.765 ;
        RECT 93.440 173.395 94.980 173.765 ;
        RECT 65.675 170.675 67.215 171.045 ;
        RECT 84.185 170.675 85.725 171.045 ;
        RECT 102.695 170.675 104.235 171.045 ;
        RECT 74.930 167.955 76.470 168.325 ;
        RECT 93.440 167.955 94.980 168.325 ;
        RECT 65.675 165.235 67.215 165.605 ;
        RECT 84.185 165.235 85.725 165.605 ;
        RECT 102.695 165.235 104.235 165.605 ;
        RECT 74.930 162.515 76.470 162.885 ;
        RECT 93.440 162.515 94.980 162.885 ;
        RECT 111.630 161.910 111.770 197.390 ;
        RECT 114.390 197.030 114.530 201.470 ;
        RECT 116.690 197.710 116.830 201.810 ;
        RECT 119.850 201.130 120.110 201.450 ;
        RECT 119.910 199.750 120.050 201.130 ;
        RECT 123.530 200.110 123.790 200.430 ;
        RECT 119.850 199.430 120.110 199.750 ;
        RECT 120.770 198.410 121.030 198.730 ;
        RECT 116.630 197.390 116.890 197.710 ;
        RECT 116.690 197.030 116.830 197.390 ;
        RECT 120.830 197.030 120.970 198.410 ;
        RECT 121.205 197.875 122.745 198.245 ;
        RECT 114.330 196.710 114.590 197.030 ;
        RECT 116.630 196.710 116.890 197.030 ;
        RECT 120.770 196.710 121.030 197.030 ;
        RECT 113.870 196.370 114.130 196.690 ;
        RECT 111.950 195.155 113.490 195.525 ;
        RECT 113.930 193.970 114.070 196.370 ;
        RECT 115.710 195.690 115.970 196.010 ;
        RECT 120.770 195.690 121.030 196.010 ;
        RECT 115.770 194.990 115.910 195.690 ;
        RECT 115.710 194.670 115.970 194.990 ;
        RECT 113.870 193.650 114.130 193.970 ;
        RECT 115.710 192.970 115.970 193.290 ;
        RECT 115.770 191.250 115.910 192.970 ;
        RECT 115.710 190.930 115.970 191.250 ;
        RECT 120.830 190.910 120.970 195.690 ;
        RECT 121.205 192.435 122.745 192.805 ;
        RECT 120.770 190.590 121.030 190.910 ;
        RECT 111.950 189.715 113.490 190.085 ;
        RECT 123.590 188.870 123.730 200.110 ;
        RECT 128.190 197.370 128.330 205.340 ;
        RECT 130.460 200.595 132.000 200.965 ;
        RECT 128.130 197.050 128.390 197.370 ;
        RECT 130.460 195.155 132.000 195.525 ;
        RECT 130.460 189.715 132.000 190.085 ;
        RECT 123.530 188.550 123.790 188.870 ;
        RECT 128.130 187.530 128.390 187.850 ;
        RECT 121.205 186.995 122.745 187.365 ;
        RECT 128.190 186.345 128.330 187.530 ;
        RECT 138.000 187.000 139.000 187.050 ;
        RECT 128.120 185.975 128.400 186.345 ;
        RECT 138.000 185.000 150.000 187.000 ;
        RECT 138.000 184.950 139.000 185.000 ;
        RECT 111.950 184.275 113.490 184.645 ;
        RECT 130.460 184.275 132.000 184.645 ;
        RECT 121.205 181.555 122.745 181.925 ;
        RECT 111.950 178.835 113.490 179.205 ;
        RECT 130.460 178.835 132.000 179.205 ;
        RECT 121.205 176.115 122.745 176.485 ;
        RECT 111.950 173.395 113.490 173.765 ;
        RECT 130.460 173.395 132.000 173.765 ;
        RECT 121.205 170.675 122.745 171.045 ;
        RECT 111.950 167.955 113.490 168.325 ;
        RECT 130.460 167.955 132.000 168.325 ;
        RECT 121.205 165.235 122.745 165.605 ;
        RECT 111.950 162.515 113.490 162.885 ;
        RECT 130.460 162.515 132.000 162.885 ;
        RECT 111.170 161.770 111.770 161.910 ;
        RECT 65.675 159.795 67.215 160.165 ;
        RECT 84.185 159.795 85.725 160.165 ;
        RECT 102.695 159.795 104.235 160.165 ;
        RECT 74.930 157.075 76.470 157.445 ;
        RECT 93.440 157.075 94.980 157.445 ;
        RECT 65.675 154.355 67.215 154.725 ;
        RECT 84.185 154.355 85.725 154.725 ;
        RECT 102.695 154.355 104.235 154.725 ;
        RECT 74.930 151.635 76.470 152.005 ;
        RECT 93.440 151.635 94.980 152.005 ;
        RECT 111.170 151.130 111.310 161.770 ;
        RECT 121.205 159.795 122.745 160.165 ;
        RECT 111.950 157.075 113.490 157.445 ;
        RECT 130.460 157.075 132.000 157.445 ;
        RECT 121.205 154.355 122.745 154.725 ;
        RECT 111.950 151.635 113.490 152.005 ;
        RECT 130.460 151.635 132.000 152.005 ;
        RECT 111.110 150.810 111.370 151.130 ;
        RECT 110.650 149.450 110.910 149.770 ;
        RECT 65.675 148.915 67.215 149.285 ;
        RECT 84.185 148.915 85.725 149.285 ;
        RECT 102.695 148.915 104.235 149.285 ;
        RECT 110.710 148.265 110.850 149.450 ;
        RECT 121.205 148.915 122.745 149.285 ;
        RECT 110.640 147.895 110.920 148.265 ;
        RECT 137.000 147.000 138.000 147.050 ;
        RECT 74.930 146.195 76.470 146.565 ;
        RECT 93.440 146.195 94.980 146.565 ;
        RECT 111.950 146.195 113.490 146.565 ;
        RECT 130.460 146.195 132.000 146.565 ;
        RECT 137.000 145.000 146.000 147.000 ;
        RECT 137.000 144.950 138.000 145.000 ;
        RECT 65.675 143.475 67.215 143.845 ;
        RECT 84.185 143.475 85.725 143.845 ;
        RECT 102.695 143.475 104.235 143.845 ;
        RECT 121.205 143.475 122.745 143.845 ;
        RECT 74.930 140.755 76.470 141.125 ;
        RECT 93.440 140.755 94.980 141.125 ;
        RECT 111.950 140.755 113.490 141.125 ;
        RECT 130.460 140.755 132.000 141.125 ;
        RECT 65.675 138.035 67.215 138.405 ;
        RECT 84.185 138.035 85.725 138.405 ;
        RECT 102.695 138.035 104.235 138.405 ;
        RECT 121.205 138.035 122.745 138.405 ;
        RECT 74.930 135.315 76.470 135.685 ;
        RECT 93.440 135.315 94.980 135.685 ;
        RECT 111.950 135.315 113.490 135.685 ;
        RECT 130.460 135.315 132.000 135.685 ;
        RECT 65.675 132.595 67.215 132.965 ;
        RECT 84.185 132.595 85.725 132.965 ;
        RECT 102.695 132.595 104.235 132.965 ;
        RECT 121.205 132.595 122.745 132.965 ;
        RECT 74.930 129.875 76.470 130.245 ;
        RECT 93.440 129.875 94.980 130.245 ;
        RECT 111.950 129.875 113.490 130.245 ;
        RECT 130.460 129.875 132.000 130.245 ;
        RECT 144.000 106.000 146.000 145.000 ;
        RECT 130.000 104.000 146.000 106.000 ;
        RECT 148.000 106.000 150.000 185.000 ;
        RECT 148.000 104.000 162.000 106.000 ;
        RECT 120.000 92.000 121.000 92.050 ;
        RECT 120.000 88.000 125.000 92.000 ;
        RECT 120.000 87.950 121.000 88.000 ;
        RECT 124.000 87.950 125.000 88.000 ;
        RECT 130.000 76.950 132.000 104.000 ;
        RECT 138.000 101.000 139.000 101.050 ;
        RECT 141.000 101.000 142.000 101.050 ;
        RECT 138.000 99.000 142.000 101.000 ;
        RECT 138.000 98.950 139.000 99.000 ;
        RECT 141.000 98.950 142.000 99.000 ;
        RECT 138.000 97.000 139.000 97.050 ;
        RECT 141.000 97.000 142.000 97.050 ;
        RECT 138.000 95.000 142.000 97.000 ;
        RECT 138.000 94.950 139.000 95.000 ;
        RECT 141.000 94.950 142.000 95.000 ;
        RECT 138.470 86.420 140.220 87.070 ;
        RECT 144.220 86.270 144.970 92.470 ;
        RECT 148.170 87.170 149.020 92.520 ;
        RECT 150.820 86.570 152.620 87.070 ;
        RECT 138.770 85.470 153.520 86.270 ;
        RECT 135.000 84.000 136.000 84.050 ;
        RECT 134.000 78.950 136.000 84.000 ;
        RECT 138.770 82.570 140.520 85.470 ;
        RECT 144.820 84.070 145.320 84.570 ;
        RECT 145.470 84.520 150.120 85.120 ;
        RECT 145.470 83.420 146.770 84.520 ;
        RECT 142.770 82.570 149.470 83.420 ;
        RECT 151.820 82.570 153.520 85.470 ;
        RECT 156.000 84.000 157.000 84.050 ;
        RECT 138.820 82.520 139.120 82.570 ;
        RECT 140.120 82.520 140.520 82.570 ;
        RECT 148.470 82.320 148.820 82.370 ;
        RECT 152.470 82.320 152.770 82.370 ;
        RECT 139.420 81.670 143.820 82.320 ;
        RECT 148.470 81.670 152.870 82.320 ;
        RECT 141.270 77.370 142.120 81.670 ;
        RECT 148.470 81.620 148.820 81.670 ;
        RECT 145.270 79.470 145.620 81.570 ;
        RECT 147.720 80.170 148.620 80.620 ;
        RECT 140.720 76.620 142.570 77.370 ;
        RECT 145.670 76.920 146.570 77.720 ;
        RECT 150.170 77.370 151.020 81.670 ;
        RECT 152.470 81.620 152.770 81.670 ;
        RECT 156.000 78.950 158.000 84.000 ;
        RECT 149.720 76.620 151.570 77.370 ;
        RECT 160.000 76.950 162.000 104.000 ;
        RECT 141.420 75.670 150.820 76.420 ;
        RECT 141.470 75.620 141.770 75.670 ;
        RECT 120.000 74.000 121.000 74.050 ;
        RECT 120.000 70.000 125.000 74.000 ;
        RECT 145.620 72.570 146.620 73.570 ;
        RECT 120.000 69.950 121.000 70.000 ;
      LAYER via2 ;
        RECT 129.000 215.000 129.500 215.500 ;
        RECT 133.000 214.000 133.500 214.500 ;
        RECT 136.500 213.000 137.000 213.500 ;
        RECT 140.000 212.000 140.500 212.500 ;
        RECT 144.000 211.000 144.500 211.500 ;
        RECT 147.500 210.000 148.000 210.500 ;
        RECT 151.000 209.000 151.500 209.500 ;
        RECT 154.745 207.775 155.280 208.310 ;
        RECT 65.705 203.360 65.985 203.640 ;
        RECT 66.105 203.360 66.385 203.640 ;
        RECT 66.505 203.360 66.785 203.640 ;
        RECT 66.905 203.360 67.185 203.640 ;
        RECT 84.215 203.360 84.495 203.640 ;
        RECT 84.615 203.360 84.895 203.640 ;
        RECT 85.015 203.360 85.295 203.640 ;
        RECT 85.415 203.360 85.695 203.640 ;
        RECT 102.725 203.360 103.005 203.640 ;
        RECT 103.125 203.360 103.405 203.640 ;
        RECT 103.525 203.360 103.805 203.640 ;
        RECT 103.925 203.360 104.205 203.640 ;
        RECT 74.960 200.640 75.240 200.920 ;
        RECT 75.360 200.640 75.640 200.920 ;
        RECT 75.760 200.640 76.040 200.920 ;
        RECT 76.160 200.640 76.440 200.920 ;
        RECT 65.705 197.920 65.985 198.200 ;
        RECT 66.105 197.920 66.385 198.200 ;
        RECT 66.505 197.920 66.785 198.200 ;
        RECT 66.905 197.920 67.185 198.200 ;
        RECT 74.960 195.200 75.240 195.480 ;
        RECT 75.360 195.200 75.640 195.480 ;
        RECT 75.760 195.200 76.040 195.480 ;
        RECT 76.160 195.200 76.440 195.480 ;
        RECT 65.705 192.480 65.985 192.760 ;
        RECT 66.105 192.480 66.385 192.760 ;
        RECT 66.505 192.480 66.785 192.760 ;
        RECT 66.905 192.480 67.185 192.760 ;
        RECT 74.960 189.760 75.240 190.040 ;
        RECT 75.360 189.760 75.640 190.040 ;
        RECT 75.760 189.760 76.040 190.040 ;
        RECT 76.160 189.760 76.440 190.040 ;
        RECT 84.215 197.920 84.495 198.200 ;
        RECT 84.615 197.920 84.895 198.200 ;
        RECT 85.015 197.920 85.295 198.200 ;
        RECT 85.415 197.920 85.695 198.200 ;
        RECT 93.470 200.640 93.750 200.920 ;
        RECT 93.870 200.640 94.150 200.920 ;
        RECT 94.270 200.640 94.550 200.920 ;
        RECT 94.670 200.640 94.950 200.920 ;
        RECT 84.215 192.480 84.495 192.760 ;
        RECT 84.615 192.480 84.895 192.760 ;
        RECT 85.015 192.480 85.295 192.760 ;
        RECT 85.415 192.480 85.695 192.760 ;
        RECT 121.235 203.360 121.515 203.640 ;
        RECT 121.635 203.360 121.915 203.640 ;
        RECT 122.035 203.360 122.315 203.640 ;
        RECT 122.435 203.360 122.715 203.640 ;
        RECT 93.470 195.200 93.750 195.480 ;
        RECT 93.870 195.200 94.150 195.480 ;
        RECT 94.270 195.200 94.550 195.480 ;
        RECT 94.670 195.200 94.950 195.480 ;
        RECT 93.470 189.760 93.750 190.040 ;
        RECT 93.870 189.760 94.150 190.040 ;
        RECT 94.270 189.760 94.550 190.040 ;
        RECT 94.670 189.760 94.950 190.040 ;
        RECT 111.980 200.640 112.260 200.920 ;
        RECT 112.380 200.640 112.660 200.920 ;
        RECT 112.780 200.640 113.060 200.920 ;
        RECT 113.180 200.640 113.460 200.920 ;
        RECT 102.725 197.920 103.005 198.200 ;
        RECT 103.125 197.920 103.405 198.200 ;
        RECT 103.525 197.920 103.805 198.200 ;
        RECT 103.925 197.920 104.205 198.200 ;
        RECT 102.725 192.480 103.005 192.760 ;
        RECT 103.125 192.480 103.405 192.760 ;
        RECT 103.525 192.480 103.805 192.760 ;
        RECT 103.925 192.480 104.205 192.760 ;
        RECT 65.705 187.040 65.985 187.320 ;
        RECT 66.105 187.040 66.385 187.320 ;
        RECT 66.505 187.040 66.785 187.320 ;
        RECT 66.905 187.040 67.185 187.320 ;
        RECT 84.215 187.040 84.495 187.320 ;
        RECT 84.615 187.040 84.895 187.320 ;
        RECT 85.015 187.040 85.295 187.320 ;
        RECT 85.415 187.040 85.695 187.320 ;
        RECT 102.725 187.040 103.005 187.320 ;
        RECT 103.125 187.040 103.405 187.320 ;
        RECT 103.525 187.040 103.805 187.320 ;
        RECT 103.925 187.040 104.205 187.320 ;
        RECT 74.960 184.320 75.240 184.600 ;
        RECT 75.360 184.320 75.640 184.600 ;
        RECT 75.760 184.320 76.040 184.600 ;
        RECT 76.160 184.320 76.440 184.600 ;
        RECT 93.470 184.320 93.750 184.600 ;
        RECT 93.870 184.320 94.150 184.600 ;
        RECT 94.270 184.320 94.550 184.600 ;
        RECT 94.670 184.320 94.950 184.600 ;
        RECT 65.705 181.600 65.985 181.880 ;
        RECT 66.105 181.600 66.385 181.880 ;
        RECT 66.505 181.600 66.785 181.880 ;
        RECT 66.905 181.600 67.185 181.880 ;
        RECT 84.215 181.600 84.495 181.880 ;
        RECT 84.615 181.600 84.895 181.880 ;
        RECT 85.015 181.600 85.295 181.880 ;
        RECT 85.415 181.600 85.695 181.880 ;
        RECT 102.725 181.600 103.005 181.880 ;
        RECT 103.125 181.600 103.405 181.880 ;
        RECT 103.525 181.600 103.805 181.880 ;
        RECT 103.925 181.600 104.205 181.880 ;
        RECT 74.960 178.880 75.240 179.160 ;
        RECT 75.360 178.880 75.640 179.160 ;
        RECT 75.760 178.880 76.040 179.160 ;
        RECT 76.160 178.880 76.440 179.160 ;
        RECT 93.470 178.880 93.750 179.160 ;
        RECT 93.870 178.880 94.150 179.160 ;
        RECT 94.270 178.880 94.550 179.160 ;
        RECT 94.670 178.880 94.950 179.160 ;
        RECT 65.705 176.160 65.985 176.440 ;
        RECT 66.105 176.160 66.385 176.440 ;
        RECT 66.505 176.160 66.785 176.440 ;
        RECT 66.905 176.160 67.185 176.440 ;
        RECT 84.215 176.160 84.495 176.440 ;
        RECT 84.615 176.160 84.895 176.440 ;
        RECT 85.015 176.160 85.295 176.440 ;
        RECT 85.415 176.160 85.695 176.440 ;
        RECT 102.725 176.160 103.005 176.440 ;
        RECT 103.125 176.160 103.405 176.440 ;
        RECT 103.525 176.160 103.805 176.440 ;
        RECT 103.925 176.160 104.205 176.440 ;
        RECT 74.960 173.440 75.240 173.720 ;
        RECT 75.360 173.440 75.640 173.720 ;
        RECT 75.760 173.440 76.040 173.720 ;
        RECT 76.160 173.440 76.440 173.720 ;
        RECT 93.470 173.440 93.750 173.720 ;
        RECT 93.870 173.440 94.150 173.720 ;
        RECT 94.270 173.440 94.550 173.720 ;
        RECT 94.670 173.440 94.950 173.720 ;
        RECT 65.705 170.720 65.985 171.000 ;
        RECT 66.105 170.720 66.385 171.000 ;
        RECT 66.505 170.720 66.785 171.000 ;
        RECT 66.905 170.720 67.185 171.000 ;
        RECT 84.215 170.720 84.495 171.000 ;
        RECT 84.615 170.720 84.895 171.000 ;
        RECT 85.015 170.720 85.295 171.000 ;
        RECT 85.415 170.720 85.695 171.000 ;
        RECT 102.725 170.720 103.005 171.000 ;
        RECT 103.125 170.720 103.405 171.000 ;
        RECT 103.525 170.720 103.805 171.000 ;
        RECT 103.925 170.720 104.205 171.000 ;
        RECT 74.960 168.000 75.240 168.280 ;
        RECT 75.360 168.000 75.640 168.280 ;
        RECT 75.760 168.000 76.040 168.280 ;
        RECT 76.160 168.000 76.440 168.280 ;
        RECT 93.470 168.000 93.750 168.280 ;
        RECT 93.870 168.000 94.150 168.280 ;
        RECT 94.270 168.000 94.550 168.280 ;
        RECT 94.670 168.000 94.950 168.280 ;
        RECT 65.705 165.280 65.985 165.560 ;
        RECT 66.105 165.280 66.385 165.560 ;
        RECT 66.505 165.280 66.785 165.560 ;
        RECT 66.905 165.280 67.185 165.560 ;
        RECT 84.215 165.280 84.495 165.560 ;
        RECT 84.615 165.280 84.895 165.560 ;
        RECT 85.015 165.280 85.295 165.560 ;
        RECT 85.415 165.280 85.695 165.560 ;
        RECT 102.725 165.280 103.005 165.560 ;
        RECT 103.125 165.280 103.405 165.560 ;
        RECT 103.525 165.280 103.805 165.560 ;
        RECT 103.925 165.280 104.205 165.560 ;
        RECT 74.960 162.560 75.240 162.840 ;
        RECT 75.360 162.560 75.640 162.840 ;
        RECT 75.760 162.560 76.040 162.840 ;
        RECT 76.160 162.560 76.440 162.840 ;
        RECT 93.470 162.560 93.750 162.840 ;
        RECT 93.870 162.560 94.150 162.840 ;
        RECT 94.270 162.560 94.550 162.840 ;
        RECT 94.670 162.560 94.950 162.840 ;
        RECT 121.235 197.920 121.515 198.200 ;
        RECT 121.635 197.920 121.915 198.200 ;
        RECT 122.035 197.920 122.315 198.200 ;
        RECT 122.435 197.920 122.715 198.200 ;
        RECT 111.980 195.200 112.260 195.480 ;
        RECT 112.380 195.200 112.660 195.480 ;
        RECT 112.780 195.200 113.060 195.480 ;
        RECT 113.180 195.200 113.460 195.480 ;
        RECT 121.235 192.480 121.515 192.760 ;
        RECT 121.635 192.480 121.915 192.760 ;
        RECT 122.035 192.480 122.315 192.760 ;
        RECT 122.435 192.480 122.715 192.760 ;
        RECT 111.980 189.760 112.260 190.040 ;
        RECT 112.380 189.760 112.660 190.040 ;
        RECT 112.780 189.760 113.060 190.040 ;
        RECT 113.180 189.760 113.460 190.040 ;
        RECT 130.490 200.640 130.770 200.920 ;
        RECT 130.890 200.640 131.170 200.920 ;
        RECT 131.290 200.640 131.570 200.920 ;
        RECT 131.690 200.640 131.970 200.920 ;
        RECT 130.490 195.200 130.770 195.480 ;
        RECT 130.890 195.200 131.170 195.480 ;
        RECT 131.290 195.200 131.570 195.480 ;
        RECT 131.690 195.200 131.970 195.480 ;
        RECT 130.490 189.760 130.770 190.040 ;
        RECT 130.890 189.760 131.170 190.040 ;
        RECT 131.290 189.760 131.570 190.040 ;
        RECT 131.690 189.760 131.970 190.040 ;
        RECT 121.235 187.040 121.515 187.320 ;
        RECT 121.635 187.040 121.915 187.320 ;
        RECT 122.035 187.040 122.315 187.320 ;
        RECT 122.435 187.040 122.715 187.320 ;
        RECT 128.120 186.020 128.400 186.300 ;
        RECT 111.980 184.320 112.260 184.600 ;
        RECT 112.380 184.320 112.660 184.600 ;
        RECT 112.780 184.320 113.060 184.600 ;
        RECT 113.180 184.320 113.460 184.600 ;
        RECT 130.490 184.320 130.770 184.600 ;
        RECT 130.890 184.320 131.170 184.600 ;
        RECT 131.290 184.320 131.570 184.600 ;
        RECT 131.690 184.320 131.970 184.600 ;
        RECT 121.235 181.600 121.515 181.880 ;
        RECT 121.635 181.600 121.915 181.880 ;
        RECT 122.035 181.600 122.315 181.880 ;
        RECT 122.435 181.600 122.715 181.880 ;
        RECT 111.980 178.880 112.260 179.160 ;
        RECT 112.380 178.880 112.660 179.160 ;
        RECT 112.780 178.880 113.060 179.160 ;
        RECT 113.180 178.880 113.460 179.160 ;
        RECT 130.490 178.880 130.770 179.160 ;
        RECT 130.890 178.880 131.170 179.160 ;
        RECT 131.290 178.880 131.570 179.160 ;
        RECT 131.690 178.880 131.970 179.160 ;
        RECT 121.235 176.160 121.515 176.440 ;
        RECT 121.635 176.160 121.915 176.440 ;
        RECT 122.035 176.160 122.315 176.440 ;
        RECT 122.435 176.160 122.715 176.440 ;
        RECT 111.980 173.440 112.260 173.720 ;
        RECT 112.380 173.440 112.660 173.720 ;
        RECT 112.780 173.440 113.060 173.720 ;
        RECT 113.180 173.440 113.460 173.720 ;
        RECT 130.490 173.440 130.770 173.720 ;
        RECT 130.890 173.440 131.170 173.720 ;
        RECT 131.290 173.440 131.570 173.720 ;
        RECT 131.690 173.440 131.970 173.720 ;
        RECT 121.235 170.720 121.515 171.000 ;
        RECT 121.635 170.720 121.915 171.000 ;
        RECT 122.035 170.720 122.315 171.000 ;
        RECT 122.435 170.720 122.715 171.000 ;
        RECT 111.980 168.000 112.260 168.280 ;
        RECT 112.380 168.000 112.660 168.280 ;
        RECT 112.780 168.000 113.060 168.280 ;
        RECT 113.180 168.000 113.460 168.280 ;
        RECT 130.490 168.000 130.770 168.280 ;
        RECT 130.890 168.000 131.170 168.280 ;
        RECT 131.290 168.000 131.570 168.280 ;
        RECT 131.690 168.000 131.970 168.280 ;
        RECT 121.235 165.280 121.515 165.560 ;
        RECT 121.635 165.280 121.915 165.560 ;
        RECT 122.035 165.280 122.315 165.560 ;
        RECT 122.435 165.280 122.715 165.560 ;
        RECT 111.980 162.560 112.260 162.840 ;
        RECT 112.380 162.560 112.660 162.840 ;
        RECT 112.780 162.560 113.060 162.840 ;
        RECT 113.180 162.560 113.460 162.840 ;
        RECT 130.490 162.560 130.770 162.840 ;
        RECT 130.890 162.560 131.170 162.840 ;
        RECT 131.290 162.560 131.570 162.840 ;
        RECT 131.690 162.560 131.970 162.840 ;
        RECT 65.705 159.840 65.985 160.120 ;
        RECT 66.105 159.840 66.385 160.120 ;
        RECT 66.505 159.840 66.785 160.120 ;
        RECT 66.905 159.840 67.185 160.120 ;
        RECT 84.215 159.840 84.495 160.120 ;
        RECT 84.615 159.840 84.895 160.120 ;
        RECT 85.015 159.840 85.295 160.120 ;
        RECT 85.415 159.840 85.695 160.120 ;
        RECT 102.725 159.840 103.005 160.120 ;
        RECT 103.125 159.840 103.405 160.120 ;
        RECT 103.525 159.840 103.805 160.120 ;
        RECT 103.925 159.840 104.205 160.120 ;
        RECT 74.960 157.120 75.240 157.400 ;
        RECT 75.360 157.120 75.640 157.400 ;
        RECT 75.760 157.120 76.040 157.400 ;
        RECT 76.160 157.120 76.440 157.400 ;
        RECT 93.470 157.120 93.750 157.400 ;
        RECT 93.870 157.120 94.150 157.400 ;
        RECT 94.270 157.120 94.550 157.400 ;
        RECT 94.670 157.120 94.950 157.400 ;
        RECT 65.705 154.400 65.985 154.680 ;
        RECT 66.105 154.400 66.385 154.680 ;
        RECT 66.505 154.400 66.785 154.680 ;
        RECT 66.905 154.400 67.185 154.680 ;
        RECT 84.215 154.400 84.495 154.680 ;
        RECT 84.615 154.400 84.895 154.680 ;
        RECT 85.015 154.400 85.295 154.680 ;
        RECT 85.415 154.400 85.695 154.680 ;
        RECT 102.725 154.400 103.005 154.680 ;
        RECT 103.125 154.400 103.405 154.680 ;
        RECT 103.525 154.400 103.805 154.680 ;
        RECT 103.925 154.400 104.205 154.680 ;
        RECT 74.960 151.680 75.240 151.960 ;
        RECT 75.360 151.680 75.640 151.960 ;
        RECT 75.760 151.680 76.040 151.960 ;
        RECT 76.160 151.680 76.440 151.960 ;
        RECT 93.470 151.680 93.750 151.960 ;
        RECT 93.870 151.680 94.150 151.960 ;
        RECT 94.270 151.680 94.550 151.960 ;
        RECT 94.670 151.680 94.950 151.960 ;
        RECT 121.235 159.840 121.515 160.120 ;
        RECT 121.635 159.840 121.915 160.120 ;
        RECT 122.035 159.840 122.315 160.120 ;
        RECT 122.435 159.840 122.715 160.120 ;
        RECT 111.980 157.120 112.260 157.400 ;
        RECT 112.380 157.120 112.660 157.400 ;
        RECT 112.780 157.120 113.060 157.400 ;
        RECT 113.180 157.120 113.460 157.400 ;
        RECT 130.490 157.120 130.770 157.400 ;
        RECT 130.890 157.120 131.170 157.400 ;
        RECT 131.290 157.120 131.570 157.400 ;
        RECT 131.690 157.120 131.970 157.400 ;
        RECT 121.235 154.400 121.515 154.680 ;
        RECT 121.635 154.400 121.915 154.680 ;
        RECT 122.035 154.400 122.315 154.680 ;
        RECT 122.435 154.400 122.715 154.680 ;
        RECT 111.980 151.680 112.260 151.960 ;
        RECT 112.380 151.680 112.660 151.960 ;
        RECT 112.780 151.680 113.060 151.960 ;
        RECT 113.180 151.680 113.460 151.960 ;
        RECT 130.490 151.680 130.770 151.960 ;
        RECT 130.890 151.680 131.170 151.960 ;
        RECT 131.290 151.680 131.570 151.960 ;
        RECT 131.690 151.680 131.970 151.960 ;
        RECT 65.705 148.960 65.985 149.240 ;
        RECT 66.105 148.960 66.385 149.240 ;
        RECT 66.505 148.960 66.785 149.240 ;
        RECT 66.905 148.960 67.185 149.240 ;
        RECT 84.215 148.960 84.495 149.240 ;
        RECT 84.615 148.960 84.895 149.240 ;
        RECT 85.015 148.960 85.295 149.240 ;
        RECT 85.415 148.960 85.695 149.240 ;
        RECT 102.725 148.960 103.005 149.240 ;
        RECT 103.125 148.960 103.405 149.240 ;
        RECT 103.525 148.960 103.805 149.240 ;
        RECT 103.925 148.960 104.205 149.240 ;
        RECT 121.235 148.960 121.515 149.240 ;
        RECT 121.635 148.960 121.915 149.240 ;
        RECT 122.035 148.960 122.315 149.240 ;
        RECT 122.435 148.960 122.715 149.240 ;
        RECT 110.640 147.940 110.920 148.220 ;
        RECT 74.960 146.240 75.240 146.520 ;
        RECT 75.360 146.240 75.640 146.520 ;
        RECT 75.760 146.240 76.040 146.520 ;
        RECT 76.160 146.240 76.440 146.520 ;
        RECT 93.470 146.240 93.750 146.520 ;
        RECT 93.870 146.240 94.150 146.520 ;
        RECT 94.270 146.240 94.550 146.520 ;
        RECT 94.670 146.240 94.950 146.520 ;
        RECT 111.980 146.240 112.260 146.520 ;
        RECT 112.380 146.240 112.660 146.520 ;
        RECT 112.780 146.240 113.060 146.520 ;
        RECT 113.180 146.240 113.460 146.520 ;
        RECT 130.490 146.240 130.770 146.520 ;
        RECT 130.890 146.240 131.170 146.520 ;
        RECT 131.290 146.240 131.570 146.520 ;
        RECT 131.690 146.240 131.970 146.520 ;
        RECT 65.705 143.520 65.985 143.800 ;
        RECT 66.105 143.520 66.385 143.800 ;
        RECT 66.505 143.520 66.785 143.800 ;
        RECT 66.905 143.520 67.185 143.800 ;
        RECT 84.215 143.520 84.495 143.800 ;
        RECT 84.615 143.520 84.895 143.800 ;
        RECT 85.015 143.520 85.295 143.800 ;
        RECT 85.415 143.520 85.695 143.800 ;
        RECT 102.725 143.520 103.005 143.800 ;
        RECT 103.125 143.520 103.405 143.800 ;
        RECT 103.525 143.520 103.805 143.800 ;
        RECT 103.925 143.520 104.205 143.800 ;
        RECT 121.235 143.520 121.515 143.800 ;
        RECT 121.635 143.520 121.915 143.800 ;
        RECT 122.035 143.520 122.315 143.800 ;
        RECT 122.435 143.520 122.715 143.800 ;
        RECT 74.960 140.800 75.240 141.080 ;
        RECT 75.360 140.800 75.640 141.080 ;
        RECT 75.760 140.800 76.040 141.080 ;
        RECT 76.160 140.800 76.440 141.080 ;
        RECT 93.470 140.800 93.750 141.080 ;
        RECT 93.870 140.800 94.150 141.080 ;
        RECT 94.270 140.800 94.550 141.080 ;
        RECT 94.670 140.800 94.950 141.080 ;
        RECT 111.980 140.800 112.260 141.080 ;
        RECT 112.380 140.800 112.660 141.080 ;
        RECT 112.780 140.800 113.060 141.080 ;
        RECT 113.180 140.800 113.460 141.080 ;
        RECT 130.490 140.800 130.770 141.080 ;
        RECT 130.890 140.800 131.170 141.080 ;
        RECT 131.290 140.800 131.570 141.080 ;
        RECT 131.690 140.800 131.970 141.080 ;
        RECT 65.705 138.080 65.985 138.360 ;
        RECT 66.105 138.080 66.385 138.360 ;
        RECT 66.505 138.080 66.785 138.360 ;
        RECT 66.905 138.080 67.185 138.360 ;
        RECT 84.215 138.080 84.495 138.360 ;
        RECT 84.615 138.080 84.895 138.360 ;
        RECT 85.015 138.080 85.295 138.360 ;
        RECT 85.415 138.080 85.695 138.360 ;
        RECT 102.725 138.080 103.005 138.360 ;
        RECT 103.125 138.080 103.405 138.360 ;
        RECT 103.525 138.080 103.805 138.360 ;
        RECT 103.925 138.080 104.205 138.360 ;
        RECT 121.235 138.080 121.515 138.360 ;
        RECT 121.635 138.080 121.915 138.360 ;
        RECT 122.035 138.080 122.315 138.360 ;
        RECT 122.435 138.080 122.715 138.360 ;
        RECT 74.960 135.360 75.240 135.640 ;
        RECT 75.360 135.360 75.640 135.640 ;
        RECT 75.760 135.360 76.040 135.640 ;
        RECT 76.160 135.360 76.440 135.640 ;
        RECT 93.470 135.360 93.750 135.640 ;
        RECT 93.870 135.360 94.150 135.640 ;
        RECT 94.270 135.360 94.550 135.640 ;
        RECT 94.670 135.360 94.950 135.640 ;
        RECT 111.980 135.360 112.260 135.640 ;
        RECT 112.380 135.360 112.660 135.640 ;
        RECT 112.780 135.360 113.060 135.640 ;
        RECT 113.180 135.360 113.460 135.640 ;
        RECT 130.490 135.360 130.770 135.640 ;
        RECT 130.890 135.360 131.170 135.640 ;
        RECT 131.290 135.360 131.570 135.640 ;
        RECT 131.690 135.360 131.970 135.640 ;
        RECT 65.705 132.640 65.985 132.920 ;
        RECT 66.105 132.640 66.385 132.920 ;
        RECT 66.505 132.640 66.785 132.920 ;
        RECT 66.905 132.640 67.185 132.920 ;
        RECT 84.215 132.640 84.495 132.920 ;
        RECT 84.615 132.640 84.895 132.920 ;
        RECT 85.015 132.640 85.295 132.920 ;
        RECT 85.415 132.640 85.695 132.920 ;
        RECT 102.725 132.640 103.005 132.920 ;
        RECT 103.125 132.640 103.405 132.920 ;
        RECT 103.525 132.640 103.805 132.920 ;
        RECT 103.925 132.640 104.205 132.920 ;
        RECT 121.235 132.640 121.515 132.920 ;
        RECT 121.635 132.640 121.915 132.920 ;
        RECT 122.035 132.640 122.315 132.920 ;
        RECT 122.435 132.640 122.715 132.920 ;
        RECT 74.960 129.920 75.240 130.200 ;
        RECT 75.360 129.920 75.640 130.200 ;
        RECT 75.760 129.920 76.040 130.200 ;
        RECT 76.160 129.920 76.440 130.200 ;
        RECT 93.470 129.920 93.750 130.200 ;
        RECT 93.870 129.920 94.150 130.200 ;
        RECT 94.270 129.920 94.550 130.200 ;
        RECT 94.670 129.920 94.950 130.200 ;
        RECT 111.980 129.920 112.260 130.200 ;
        RECT 112.380 129.920 112.660 130.200 ;
        RECT 112.780 129.920 113.060 130.200 ;
        RECT 113.180 129.920 113.460 130.200 ;
        RECT 130.490 129.920 130.770 130.200 ;
        RECT 130.890 129.920 131.170 130.200 ;
        RECT 131.290 129.920 131.570 130.200 ;
        RECT 131.690 129.920 131.970 130.200 ;
        RECT 138.570 86.620 140.120 87.020 ;
        RECT 150.920 86.670 152.520 86.970 ;
        RECT 144.920 84.170 145.220 84.470 ;
        RECT 134.000 79.000 136.000 80.000 ;
        RECT 147.920 80.220 148.470 80.570 ;
        RECT 145.770 77.020 146.470 77.620 ;
        RECT 156.000 79.000 158.000 80.000 ;
        RECT 145.770 72.670 146.470 73.420 ;
      LAYER met3 ;
        RECT 128.950 224.500 129.550 225.000 ;
        RECT 132.950 224.500 133.550 225.000 ;
        RECT 136.450 224.500 137.050 225.000 ;
        RECT 139.950 224.500 140.550 225.000 ;
        RECT 143.950 224.500 144.550 225.000 ;
        RECT 147.450 224.500 148.050 225.000 ;
        RECT 150.950 224.500 151.550 225.000 ;
        RECT 154.750 224.540 155.310 224.690 ;
        RECT 129.000 215.525 129.500 224.500 ;
        RECT 128.950 214.975 129.550 215.525 ;
        RECT 133.000 214.525 133.500 224.500 ;
        RECT 132.950 213.975 133.550 214.525 ;
        RECT 136.500 213.525 137.000 224.500 ;
        RECT 136.450 212.975 137.050 213.525 ;
        RECT 140.000 212.525 140.500 224.500 ;
        RECT 139.950 211.975 140.550 212.525 ;
        RECT 144.000 211.525 144.500 224.500 ;
        RECT 143.950 210.975 144.550 211.525 ;
        RECT 147.500 210.525 148.000 224.500 ;
        RECT 147.450 209.975 148.050 210.525 ;
        RECT 151.000 209.525 151.500 224.500 ;
        RECT 154.720 224.160 155.310 224.540 ;
        RECT 150.950 208.975 151.550 209.525 ;
        RECT 154.720 207.750 155.305 224.160 ;
        RECT 65.655 203.335 67.235 203.665 ;
        RECT 84.165 203.335 85.745 203.665 ;
        RECT 102.675 203.335 104.255 203.665 ;
        RECT 121.185 203.335 122.765 203.665 ;
        RECT 74.910 200.615 76.490 200.945 ;
        RECT 93.420 200.615 95.000 200.945 ;
        RECT 111.930 200.615 113.510 200.945 ;
        RECT 130.440 200.615 132.020 200.945 ;
        RECT 65.655 197.895 67.235 198.225 ;
        RECT 84.165 197.895 85.745 198.225 ;
        RECT 102.675 197.895 104.255 198.225 ;
        RECT 121.185 197.895 122.765 198.225 ;
        RECT 74.910 195.175 76.490 195.505 ;
        RECT 93.420 195.175 95.000 195.505 ;
        RECT 111.930 195.175 113.510 195.505 ;
        RECT 130.440 195.175 132.020 195.505 ;
        RECT 65.655 192.455 67.235 192.785 ;
        RECT 84.165 192.455 85.745 192.785 ;
        RECT 102.675 192.455 104.255 192.785 ;
        RECT 121.185 192.455 122.765 192.785 ;
        RECT 74.910 189.735 76.490 190.065 ;
        RECT 93.420 189.735 95.000 190.065 ;
        RECT 111.930 189.735 113.510 190.065 ;
        RECT 130.440 189.735 132.020 190.065 ;
        RECT 65.655 187.015 67.235 187.345 ;
        RECT 84.165 187.015 85.745 187.345 ;
        RECT 102.675 187.015 104.255 187.345 ;
        RECT 121.185 187.015 122.765 187.345 ;
        RECT 137.950 187.000 139.050 187.025 ;
        RECT 134.000 186.460 139.050 187.000 ;
        RECT 128.095 186.310 128.425 186.325 ;
        RECT 132.430 186.310 139.050 186.460 ;
        RECT 128.095 186.010 139.050 186.310 ;
        RECT 128.095 185.995 128.425 186.010 ;
        RECT 132.430 185.860 139.050 186.010 ;
        RECT 134.000 185.000 139.050 185.860 ;
        RECT 137.950 184.975 139.050 185.000 ;
        RECT 74.910 184.295 76.490 184.625 ;
        RECT 93.420 184.295 95.000 184.625 ;
        RECT 111.930 184.295 113.510 184.625 ;
        RECT 130.440 184.295 132.020 184.625 ;
        RECT 65.655 181.575 67.235 181.905 ;
        RECT 84.165 181.575 85.745 181.905 ;
        RECT 102.675 181.575 104.255 181.905 ;
        RECT 121.185 181.575 122.765 181.905 ;
        RECT 74.910 178.855 76.490 179.185 ;
        RECT 93.420 178.855 95.000 179.185 ;
        RECT 111.930 178.855 113.510 179.185 ;
        RECT 130.440 178.855 132.020 179.185 ;
        RECT 65.655 176.135 67.235 176.465 ;
        RECT 84.165 176.135 85.745 176.465 ;
        RECT 102.675 176.135 104.255 176.465 ;
        RECT 121.185 176.135 122.765 176.465 ;
        RECT 74.910 173.415 76.490 173.745 ;
        RECT 93.420 173.415 95.000 173.745 ;
        RECT 111.930 173.415 113.510 173.745 ;
        RECT 130.440 173.415 132.020 173.745 ;
        RECT 65.655 170.695 67.235 171.025 ;
        RECT 84.165 170.695 85.745 171.025 ;
        RECT 102.675 170.695 104.255 171.025 ;
        RECT 121.185 170.695 122.765 171.025 ;
        RECT 74.910 167.975 76.490 168.305 ;
        RECT 93.420 167.975 95.000 168.305 ;
        RECT 111.930 167.975 113.510 168.305 ;
        RECT 130.440 167.975 132.020 168.305 ;
        RECT 65.655 165.255 67.235 165.585 ;
        RECT 84.165 165.255 85.745 165.585 ;
        RECT 102.675 165.255 104.255 165.585 ;
        RECT 121.185 165.255 122.765 165.585 ;
        RECT 74.910 162.535 76.490 162.865 ;
        RECT 93.420 162.535 95.000 162.865 ;
        RECT 111.930 162.535 113.510 162.865 ;
        RECT 130.440 162.535 132.020 162.865 ;
        RECT 65.655 159.815 67.235 160.145 ;
        RECT 84.165 159.815 85.745 160.145 ;
        RECT 102.675 159.815 104.255 160.145 ;
        RECT 121.185 159.815 122.765 160.145 ;
        RECT 74.910 157.095 76.490 157.425 ;
        RECT 93.420 157.095 95.000 157.425 ;
        RECT 111.930 157.095 113.510 157.425 ;
        RECT 130.440 157.095 132.020 157.425 ;
        RECT 65.655 154.375 67.235 154.705 ;
        RECT 84.165 154.375 85.745 154.705 ;
        RECT 102.675 154.375 104.255 154.705 ;
        RECT 121.185 154.375 122.765 154.705 ;
        RECT 74.910 151.655 76.490 151.985 ;
        RECT 93.420 151.655 95.000 151.985 ;
        RECT 111.930 151.655 113.510 151.985 ;
        RECT 130.440 151.655 132.020 151.985 ;
        RECT 65.655 148.935 67.235 149.265 ;
        RECT 84.165 148.935 85.745 149.265 ;
        RECT 102.675 148.935 104.255 149.265 ;
        RECT 121.185 148.935 122.765 149.265 ;
        RECT 110.615 148.230 110.945 148.245 ;
        RECT 110.615 148.190 132.320 148.230 ;
        RECT 110.615 147.930 134.160 148.190 ;
        RECT 110.615 147.915 110.945 147.930 ;
        RECT 132.020 147.890 134.160 147.930 ;
        RECT 133.860 147.020 134.160 147.890 ;
        RECT 132.430 147.000 134.430 147.020 ;
        RECT 136.950 147.000 138.050 147.025 ;
        RECT 74.910 146.215 76.490 146.545 ;
        RECT 93.420 146.215 95.000 146.545 ;
        RECT 111.930 146.215 113.510 146.545 ;
        RECT 130.440 146.215 132.020 146.545 ;
        RECT 132.430 146.420 138.050 147.000 ;
        RECT 133.000 145.000 138.050 146.420 ;
        RECT 136.950 144.975 138.050 145.000 ;
        RECT 65.655 143.495 67.235 143.825 ;
        RECT 84.165 143.495 85.745 143.825 ;
        RECT 102.675 143.495 104.255 143.825 ;
        RECT 121.185 143.495 122.765 143.825 ;
        RECT 74.910 140.775 76.490 141.105 ;
        RECT 93.420 140.775 95.000 141.105 ;
        RECT 111.930 140.775 113.510 141.105 ;
        RECT 130.440 140.775 132.020 141.105 ;
        RECT 65.655 138.055 67.235 138.385 ;
        RECT 84.165 138.055 85.745 138.385 ;
        RECT 102.675 138.055 104.255 138.385 ;
        RECT 121.185 138.055 122.765 138.385 ;
        RECT 74.910 135.335 76.490 135.665 ;
        RECT 93.420 135.335 95.000 135.665 ;
        RECT 111.930 135.335 113.510 135.665 ;
        RECT 130.440 135.335 132.020 135.665 ;
        RECT 65.655 132.615 67.235 132.945 ;
        RECT 84.165 132.615 85.745 132.945 ;
        RECT 102.675 132.615 104.255 132.945 ;
        RECT 121.185 132.615 122.765 132.945 ;
        RECT 74.910 129.895 76.490 130.225 ;
        RECT 93.420 129.895 95.000 130.225 ;
        RECT 111.930 129.895 113.510 130.225 ;
        RECT 130.440 129.895 132.020 130.225 ;
        RECT 1.005 121.640 2.495 121.665 ;
        RECT 65.630 121.640 67.130 124.760 ;
        RECT 84.050 121.640 85.550 124.730 ;
        RECT 102.760 121.640 104.260 124.760 ;
        RECT 121.180 121.640 122.680 124.760 ;
        RECT 1.000 120.140 122.680 121.640 ;
        RECT 1.005 120.115 2.495 120.140 ;
        RECT 137.950 101.000 139.050 101.025 ;
        RECT 134.950 99.000 139.050 101.000 ;
        RECT 137.950 98.975 139.050 99.000 ;
        RECT 137.950 97.000 139.050 97.025 ;
        RECT 134.950 95.000 139.050 97.000 ;
        RECT 137.950 94.975 139.050 95.000 ;
        RECT 9.950 92.025 121.000 93.000 ;
        RECT 9.950 87.975 121.050 92.025 ;
        RECT 9.950 87.000 121.000 87.975 ;
        RECT 138.470 86.570 140.220 87.070 ;
        RECT 150.820 86.570 152.620 87.070 ;
        RECT 138.470 86.070 152.620 86.570 ;
        RECT 145.620 84.570 146.670 86.070 ;
        RECT 144.820 84.070 146.670 84.570 ;
        RECT 145.620 80.620 146.670 84.070 ;
        RECT 145.620 80.170 148.620 80.620 ;
        RECT 133.950 78.975 136.050 80.025 ;
        RECT 134.000 78.000 136.000 78.975 ;
        RECT 133.950 77.000 136.050 78.000 ;
        RECT 59.950 74.025 121.000 75.000 ;
        RECT 59.950 69.975 121.050 74.025 ;
        RECT 145.620 72.570 146.670 80.170 ;
        RECT 155.950 78.975 158.050 80.025 ;
        RECT 156.000 78.000 158.000 78.975 ;
        RECT 155.950 77.000 158.050 78.000 ;
        RECT 59.950 69.000 121.000 69.975 ;
      LAYER via3 ;
        RECT 129.000 224.500 129.500 225.000 ;
        RECT 133.000 224.500 133.500 225.000 ;
        RECT 136.500 224.500 137.000 225.000 ;
        RECT 140.000 224.500 140.500 225.000 ;
        RECT 144.000 224.500 144.500 225.000 ;
        RECT 147.500 224.500 148.000 225.000 ;
        RECT 151.000 224.500 151.500 225.000 ;
        RECT 154.800 224.330 155.250 224.660 ;
        RECT 65.685 203.340 66.005 203.660 ;
        RECT 66.085 203.340 66.405 203.660 ;
        RECT 66.485 203.340 66.805 203.660 ;
        RECT 66.885 203.340 67.205 203.660 ;
        RECT 84.195 203.340 84.515 203.660 ;
        RECT 84.595 203.340 84.915 203.660 ;
        RECT 84.995 203.340 85.315 203.660 ;
        RECT 85.395 203.340 85.715 203.660 ;
        RECT 102.705 203.340 103.025 203.660 ;
        RECT 103.105 203.340 103.425 203.660 ;
        RECT 103.505 203.340 103.825 203.660 ;
        RECT 103.905 203.340 104.225 203.660 ;
        RECT 121.215 203.340 121.535 203.660 ;
        RECT 121.615 203.340 121.935 203.660 ;
        RECT 122.015 203.340 122.335 203.660 ;
        RECT 122.415 203.340 122.735 203.660 ;
        RECT 74.940 200.620 75.260 200.940 ;
        RECT 75.340 200.620 75.660 200.940 ;
        RECT 75.740 200.620 76.060 200.940 ;
        RECT 76.140 200.620 76.460 200.940 ;
        RECT 93.450 200.620 93.770 200.940 ;
        RECT 93.850 200.620 94.170 200.940 ;
        RECT 94.250 200.620 94.570 200.940 ;
        RECT 94.650 200.620 94.970 200.940 ;
        RECT 111.960 200.620 112.280 200.940 ;
        RECT 112.360 200.620 112.680 200.940 ;
        RECT 112.760 200.620 113.080 200.940 ;
        RECT 113.160 200.620 113.480 200.940 ;
        RECT 130.470 200.620 130.790 200.940 ;
        RECT 130.870 200.620 131.190 200.940 ;
        RECT 131.270 200.620 131.590 200.940 ;
        RECT 131.670 200.620 131.990 200.940 ;
        RECT 65.685 197.900 66.005 198.220 ;
        RECT 66.085 197.900 66.405 198.220 ;
        RECT 66.485 197.900 66.805 198.220 ;
        RECT 66.885 197.900 67.205 198.220 ;
        RECT 84.195 197.900 84.515 198.220 ;
        RECT 84.595 197.900 84.915 198.220 ;
        RECT 84.995 197.900 85.315 198.220 ;
        RECT 85.395 197.900 85.715 198.220 ;
        RECT 102.705 197.900 103.025 198.220 ;
        RECT 103.105 197.900 103.425 198.220 ;
        RECT 103.505 197.900 103.825 198.220 ;
        RECT 103.905 197.900 104.225 198.220 ;
        RECT 121.215 197.900 121.535 198.220 ;
        RECT 121.615 197.900 121.935 198.220 ;
        RECT 122.015 197.900 122.335 198.220 ;
        RECT 122.415 197.900 122.735 198.220 ;
        RECT 74.940 195.180 75.260 195.500 ;
        RECT 75.340 195.180 75.660 195.500 ;
        RECT 75.740 195.180 76.060 195.500 ;
        RECT 76.140 195.180 76.460 195.500 ;
        RECT 93.450 195.180 93.770 195.500 ;
        RECT 93.850 195.180 94.170 195.500 ;
        RECT 94.250 195.180 94.570 195.500 ;
        RECT 94.650 195.180 94.970 195.500 ;
        RECT 111.960 195.180 112.280 195.500 ;
        RECT 112.360 195.180 112.680 195.500 ;
        RECT 112.760 195.180 113.080 195.500 ;
        RECT 113.160 195.180 113.480 195.500 ;
        RECT 130.470 195.180 130.790 195.500 ;
        RECT 130.870 195.180 131.190 195.500 ;
        RECT 131.270 195.180 131.590 195.500 ;
        RECT 131.670 195.180 131.990 195.500 ;
        RECT 65.685 192.460 66.005 192.780 ;
        RECT 66.085 192.460 66.405 192.780 ;
        RECT 66.485 192.460 66.805 192.780 ;
        RECT 66.885 192.460 67.205 192.780 ;
        RECT 84.195 192.460 84.515 192.780 ;
        RECT 84.595 192.460 84.915 192.780 ;
        RECT 84.995 192.460 85.315 192.780 ;
        RECT 85.395 192.460 85.715 192.780 ;
        RECT 102.705 192.460 103.025 192.780 ;
        RECT 103.105 192.460 103.425 192.780 ;
        RECT 103.505 192.460 103.825 192.780 ;
        RECT 103.905 192.460 104.225 192.780 ;
        RECT 121.215 192.460 121.535 192.780 ;
        RECT 121.615 192.460 121.935 192.780 ;
        RECT 122.015 192.460 122.335 192.780 ;
        RECT 122.415 192.460 122.735 192.780 ;
        RECT 74.940 189.740 75.260 190.060 ;
        RECT 75.340 189.740 75.660 190.060 ;
        RECT 75.740 189.740 76.060 190.060 ;
        RECT 76.140 189.740 76.460 190.060 ;
        RECT 93.450 189.740 93.770 190.060 ;
        RECT 93.850 189.740 94.170 190.060 ;
        RECT 94.250 189.740 94.570 190.060 ;
        RECT 94.650 189.740 94.970 190.060 ;
        RECT 111.960 189.740 112.280 190.060 ;
        RECT 112.360 189.740 112.680 190.060 ;
        RECT 112.760 189.740 113.080 190.060 ;
        RECT 113.160 189.740 113.480 190.060 ;
        RECT 130.470 189.740 130.790 190.060 ;
        RECT 130.870 189.740 131.190 190.060 ;
        RECT 131.270 189.740 131.590 190.060 ;
        RECT 131.670 189.740 131.990 190.060 ;
        RECT 65.685 187.020 66.005 187.340 ;
        RECT 66.085 187.020 66.405 187.340 ;
        RECT 66.485 187.020 66.805 187.340 ;
        RECT 66.885 187.020 67.205 187.340 ;
        RECT 84.195 187.020 84.515 187.340 ;
        RECT 84.595 187.020 84.915 187.340 ;
        RECT 84.995 187.020 85.315 187.340 ;
        RECT 85.395 187.020 85.715 187.340 ;
        RECT 102.705 187.020 103.025 187.340 ;
        RECT 103.105 187.020 103.425 187.340 ;
        RECT 103.505 187.020 103.825 187.340 ;
        RECT 103.905 187.020 104.225 187.340 ;
        RECT 121.215 187.020 121.535 187.340 ;
        RECT 121.615 187.020 121.935 187.340 ;
        RECT 122.015 187.020 122.335 187.340 ;
        RECT 122.415 187.020 122.735 187.340 ;
        RECT 74.940 184.300 75.260 184.620 ;
        RECT 75.340 184.300 75.660 184.620 ;
        RECT 75.740 184.300 76.060 184.620 ;
        RECT 76.140 184.300 76.460 184.620 ;
        RECT 93.450 184.300 93.770 184.620 ;
        RECT 93.850 184.300 94.170 184.620 ;
        RECT 94.250 184.300 94.570 184.620 ;
        RECT 94.650 184.300 94.970 184.620 ;
        RECT 111.960 184.300 112.280 184.620 ;
        RECT 112.360 184.300 112.680 184.620 ;
        RECT 112.760 184.300 113.080 184.620 ;
        RECT 113.160 184.300 113.480 184.620 ;
        RECT 130.470 184.300 130.790 184.620 ;
        RECT 130.870 184.300 131.190 184.620 ;
        RECT 131.270 184.300 131.590 184.620 ;
        RECT 131.670 184.300 131.990 184.620 ;
        RECT 65.685 181.580 66.005 181.900 ;
        RECT 66.085 181.580 66.405 181.900 ;
        RECT 66.485 181.580 66.805 181.900 ;
        RECT 66.885 181.580 67.205 181.900 ;
        RECT 84.195 181.580 84.515 181.900 ;
        RECT 84.595 181.580 84.915 181.900 ;
        RECT 84.995 181.580 85.315 181.900 ;
        RECT 85.395 181.580 85.715 181.900 ;
        RECT 102.705 181.580 103.025 181.900 ;
        RECT 103.105 181.580 103.425 181.900 ;
        RECT 103.505 181.580 103.825 181.900 ;
        RECT 103.905 181.580 104.225 181.900 ;
        RECT 121.215 181.580 121.535 181.900 ;
        RECT 121.615 181.580 121.935 181.900 ;
        RECT 122.015 181.580 122.335 181.900 ;
        RECT 122.415 181.580 122.735 181.900 ;
        RECT 74.940 178.860 75.260 179.180 ;
        RECT 75.340 178.860 75.660 179.180 ;
        RECT 75.740 178.860 76.060 179.180 ;
        RECT 76.140 178.860 76.460 179.180 ;
        RECT 93.450 178.860 93.770 179.180 ;
        RECT 93.850 178.860 94.170 179.180 ;
        RECT 94.250 178.860 94.570 179.180 ;
        RECT 94.650 178.860 94.970 179.180 ;
        RECT 111.960 178.860 112.280 179.180 ;
        RECT 112.360 178.860 112.680 179.180 ;
        RECT 112.760 178.860 113.080 179.180 ;
        RECT 113.160 178.860 113.480 179.180 ;
        RECT 130.470 178.860 130.790 179.180 ;
        RECT 130.870 178.860 131.190 179.180 ;
        RECT 131.270 178.860 131.590 179.180 ;
        RECT 131.670 178.860 131.990 179.180 ;
        RECT 65.685 176.140 66.005 176.460 ;
        RECT 66.085 176.140 66.405 176.460 ;
        RECT 66.485 176.140 66.805 176.460 ;
        RECT 66.885 176.140 67.205 176.460 ;
        RECT 84.195 176.140 84.515 176.460 ;
        RECT 84.595 176.140 84.915 176.460 ;
        RECT 84.995 176.140 85.315 176.460 ;
        RECT 85.395 176.140 85.715 176.460 ;
        RECT 102.705 176.140 103.025 176.460 ;
        RECT 103.105 176.140 103.425 176.460 ;
        RECT 103.505 176.140 103.825 176.460 ;
        RECT 103.905 176.140 104.225 176.460 ;
        RECT 121.215 176.140 121.535 176.460 ;
        RECT 121.615 176.140 121.935 176.460 ;
        RECT 122.015 176.140 122.335 176.460 ;
        RECT 122.415 176.140 122.735 176.460 ;
        RECT 74.940 173.420 75.260 173.740 ;
        RECT 75.340 173.420 75.660 173.740 ;
        RECT 75.740 173.420 76.060 173.740 ;
        RECT 76.140 173.420 76.460 173.740 ;
        RECT 93.450 173.420 93.770 173.740 ;
        RECT 93.850 173.420 94.170 173.740 ;
        RECT 94.250 173.420 94.570 173.740 ;
        RECT 94.650 173.420 94.970 173.740 ;
        RECT 111.960 173.420 112.280 173.740 ;
        RECT 112.360 173.420 112.680 173.740 ;
        RECT 112.760 173.420 113.080 173.740 ;
        RECT 113.160 173.420 113.480 173.740 ;
        RECT 130.470 173.420 130.790 173.740 ;
        RECT 130.870 173.420 131.190 173.740 ;
        RECT 131.270 173.420 131.590 173.740 ;
        RECT 131.670 173.420 131.990 173.740 ;
        RECT 65.685 170.700 66.005 171.020 ;
        RECT 66.085 170.700 66.405 171.020 ;
        RECT 66.485 170.700 66.805 171.020 ;
        RECT 66.885 170.700 67.205 171.020 ;
        RECT 84.195 170.700 84.515 171.020 ;
        RECT 84.595 170.700 84.915 171.020 ;
        RECT 84.995 170.700 85.315 171.020 ;
        RECT 85.395 170.700 85.715 171.020 ;
        RECT 102.705 170.700 103.025 171.020 ;
        RECT 103.105 170.700 103.425 171.020 ;
        RECT 103.505 170.700 103.825 171.020 ;
        RECT 103.905 170.700 104.225 171.020 ;
        RECT 121.215 170.700 121.535 171.020 ;
        RECT 121.615 170.700 121.935 171.020 ;
        RECT 122.015 170.700 122.335 171.020 ;
        RECT 122.415 170.700 122.735 171.020 ;
        RECT 74.940 167.980 75.260 168.300 ;
        RECT 75.340 167.980 75.660 168.300 ;
        RECT 75.740 167.980 76.060 168.300 ;
        RECT 76.140 167.980 76.460 168.300 ;
        RECT 93.450 167.980 93.770 168.300 ;
        RECT 93.850 167.980 94.170 168.300 ;
        RECT 94.250 167.980 94.570 168.300 ;
        RECT 94.650 167.980 94.970 168.300 ;
        RECT 111.960 167.980 112.280 168.300 ;
        RECT 112.360 167.980 112.680 168.300 ;
        RECT 112.760 167.980 113.080 168.300 ;
        RECT 113.160 167.980 113.480 168.300 ;
        RECT 130.470 167.980 130.790 168.300 ;
        RECT 130.870 167.980 131.190 168.300 ;
        RECT 131.270 167.980 131.590 168.300 ;
        RECT 131.670 167.980 131.990 168.300 ;
        RECT 65.685 165.260 66.005 165.580 ;
        RECT 66.085 165.260 66.405 165.580 ;
        RECT 66.485 165.260 66.805 165.580 ;
        RECT 66.885 165.260 67.205 165.580 ;
        RECT 84.195 165.260 84.515 165.580 ;
        RECT 84.595 165.260 84.915 165.580 ;
        RECT 84.995 165.260 85.315 165.580 ;
        RECT 85.395 165.260 85.715 165.580 ;
        RECT 102.705 165.260 103.025 165.580 ;
        RECT 103.105 165.260 103.425 165.580 ;
        RECT 103.505 165.260 103.825 165.580 ;
        RECT 103.905 165.260 104.225 165.580 ;
        RECT 121.215 165.260 121.535 165.580 ;
        RECT 121.615 165.260 121.935 165.580 ;
        RECT 122.015 165.260 122.335 165.580 ;
        RECT 122.415 165.260 122.735 165.580 ;
        RECT 74.940 162.540 75.260 162.860 ;
        RECT 75.340 162.540 75.660 162.860 ;
        RECT 75.740 162.540 76.060 162.860 ;
        RECT 76.140 162.540 76.460 162.860 ;
        RECT 93.450 162.540 93.770 162.860 ;
        RECT 93.850 162.540 94.170 162.860 ;
        RECT 94.250 162.540 94.570 162.860 ;
        RECT 94.650 162.540 94.970 162.860 ;
        RECT 111.960 162.540 112.280 162.860 ;
        RECT 112.360 162.540 112.680 162.860 ;
        RECT 112.760 162.540 113.080 162.860 ;
        RECT 113.160 162.540 113.480 162.860 ;
        RECT 130.470 162.540 130.790 162.860 ;
        RECT 130.870 162.540 131.190 162.860 ;
        RECT 131.270 162.540 131.590 162.860 ;
        RECT 131.670 162.540 131.990 162.860 ;
        RECT 65.685 159.820 66.005 160.140 ;
        RECT 66.085 159.820 66.405 160.140 ;
        RECT 66.485 159.820 66.805 160.140 ;
        RECT 66.885 159.820 67.205 160.140 ;
        RECT 84.195 159.820 84.515 160.140 ;
        RECT 84.595 159.820 84.915 160.140 ;
        RECT 84.995 159.820 85.315 160.140 ;
        RECT 85.395 159.820 85.715 160.140 ;
        RECT 102.705 159.820 103.025 160.140 ;
        RECT 103.105 159.820 103.425 160.140 ;
        RECT 103.505 159.820 103.825 160.140 ;
        RECT 103.905 159.820 104.225 160.140 ;
        RECT 121.215 159.820 121.535 160.140 ;
        RECT 121.615 159.820 121.935 160.140 ;
        RECT 122.015 159.820 122.335 160.140 ;
        RECT 122.415 159.820 122.735 160.140 ;
        RECT 74.940 157.100 75.260 157.420 ;
        RECT 75.340 157.100 75.660 157.420 ;
        RECT 75.740 157.100 76.060 157.420 ;
        RECT 76.140 157.100 76.460 157.420 ;
        RECT 93.450 157.100 93.770 157.420 ;
        RECT 93.850 157.100 94.170 157.420 ;
        RECT 94.250 157.100 94.570 157.420 ;
        RECT 94.650 157.100 94.970 157.420 ;
        RECT 111.960 157.100 112.280 157.420 ;
        RECT 112.360 157.100 112.680 157.420 ;
        RECT 112.760 157.100 113.080 157.420 ;
        RECT 113.160 157.100 113.480 157.420 ;
        RECT 130.470 157.100 130.790 157.420 ;
        RECT 130.870 157.100 131.190 157.420 ;
        RECT 131.270 157.100 131.590 157.420 ;
        RECT 131.670 157.100 131.990 157.420 ;
        RECT 65.685 154.380 66.005 154.700 ;
        RECT 66.085 154.380 66.405 154.700 ;
        RECT 66.485 154.380 66.805 154.700 ;
        RECT 66.885 154.380 67.205 154.700 ;
        RECT 84.195 154.380 84.515 154.700 ;
        RECT 84.595 154.380 84.915 154.700 ;
        RECT 84.995 154.380 85.315 154.700 ;
        RECT 85.395 154.380 85.715 154.700 ;
        RECT 102.705 154.380 103.025 154.700 ;
        RECT 103.105 154.380 103.425 154.700 ;
        RECT 103.505 154.380 103.825 154.700 ;
        RECT 103.905 154.380 104.225 154.700 ;
        RECT 121.215 154.380 121.535 154.700 ;
        RECT 121.615 154.380 121.935 154.700 ;
        RECT 122.015 154.380 122.335 154.700 ;
        RECT 122.415 154.380 122.735 154.700 ;
        RECT 74.940 151.660 75.260 151.980 ;
        RECT 75.340 151.660 75.660 151.980 ;
        RECT 75.740 151.660 76.060 151.980 ;
        RECT 76.140 151.660 76.460 151.980 ;
        RECT 93.450 151.660 93.770 151.980 ;
        RECT 93.850 151.660 94.170 151.980 ;
        RECT 94.250 151.660 94.570 151.980 ;
        RECT 94.650 151.660 94.970 151.980 ;
        RECT 111.960 151.660 112.280 151.980 ;
        RECT 112.360 151.660 112.680 151.980 ;
        RECT 112.760 151.660 113.080 151.980 ;
        RECT 113.160 151.660 113.480 151.980 ;
        RECT 130.470 151.660 130.790 151.980 ;
        RECT 130.870 151.660 131.190 151.980 ;
        RECT 131.270 151.660 131.590 151.980 ;
        RECT 131.670 151.660 131.990 151.980 ;
        RECT 65.685 148.940 66.005 149.260 ;
        RECT 66.085 148.940 66.405 149.260 ;
        RECT 66.485 148.940 66.805 149.260 ;
        RECT 66.885 148.940 67.205 149.260 ;
        RECT 84.195 148.940 84.515 149.260 ;
        RECT 84.595 148.940 84.915 149.260 ;
        RECT 84.995 148.940 85.315 149.260 ;
        RECT 85.395 148.940 85.715 149.260 ;
        RECT 102.705 148.940 103.025 149.260 ;
        RECT 103.105 148.940 103.425 149.260 ;
        RECT 103.505 148.940 103.825 149.260 ;
        RECT 103.905 148.940 104.225 149.260 ;
        RECT 121.215 148.940 121.535 149.260 ;
        RECT 121.615 148.940 121.935 149.260 ;
        RECT 122.015 148.940 122.335 149.260 ;
        RECT 122.415 148.940 122.735 149.260 ;
        RECT 74.940 146.220 75.260 146.540 ;
        RECT 75.340 146.220 75.660 146.540 ;
        RECT 75.740 146.220 76.060 146.540 ;
        RECT 76.140 146.220 76.460 146.540 ;
        RECT 93.450 146.220 93.770 146.540 ;
        RECT 93.850 146.220 94.170 146.540 ;
        RECT 94.250 146.220 94.570 146.540 ;
        RECT 94.650 146.220 94.970 146.540 ;
        RECT 111.960 146.220 112.280 146.540 ;
        RECT 112.360 146.220 112.680 146.540 ;
        RECT 112.760 146.220 113.080 146.540 ;
        RECT 113.160 146.220 113.480 146.540 ;
        RECT 130.470 146.220 130.790 146.540 ;
        RECT 130.870 146.220 131.190 146.540 ;
        RECT 131.270 146.220 131.590 146.540 ;
        RECT 131.670 146.220 131.990 146.540 ;
        RECT 65.685 143.500 66.005 143.820 ;
        RECT 66.085 143.500 66.405 143.820 ;
        RECT 66.485 143.500 66.805 143.820 ;
        RECT 66.885 143.500 67.205 143.820 ;
        RECT 84.195 143.500 84.515 143.820 ;
        RECT 84.595 143.500 84.915 143.820 ;
        RECT 84.995 143.500 85.315 143.820 ;
        RECT 85.395 143.500 85.715 143.820 ;
        RECT 102.705 143.500 103.025 143.820 ;
        RECT 103.105 143.500 103.425 143.820 ;
        RECT 103.505 143.500 103.825 143.820 ;
        RECT 103.905 143.500 104.225 143.820 ;
        RECT 121.215 143.500 121.535 143.820 ;
        RECT 121.615 143.500 121.935 143.820 ;
        RECT 122.015 143.500 122.335 143.820 ;
        RECT 122.415 143.500 122.735 143.820 ;
        RECT 74.940 140.780 75.260 141.100 ;
        RECT 75.340 140.780 75.660 141.100 ;
        RECT 75.740 140.780 76.060 141.100 ;
        RECT 76.140 140.780 76.460 141.100 ;
        RECT 93.450 140.780 93.770 141.100 ;
        RECT 93.850 140.780 94.170 141.100 ;
        RECT 94.250 140.780 94.570 141.100 ;
        RECT 94.650 140.780 94.970 141.100 ;
        RECT 111.960 140.780 112.280 141.100 ;
        RECT 112.360 140.780 112.680 141.100 ;
        RECT 112.760 140.780 113.080 141.100 ;
        RECT 113.160 140.780 113.480 141.100 ;
        RECT 130.470 140.780 130.790 141.100 ;
        RECT 130.870 140.780 131.190 141.100 ;
        RECT 131.270 140.780 131.590 141.100 ;
        RECT 131.670 140.780 131.990 141.100 ;
        RECT 65.685 138.060 66.005 138.380 ;
        RECT 66.085 138.060 66.405 138.380 ;
        RECT 66.485 138.060 66.805 138.380 ;
        RECT 66.885 138.060 67.205 138.380 ;
        RECT 84.195 138.060 84.515 138.380 ;
        RECT 84.595 138.060 84.915 138.380 ;
        RECT 84.995 138.060 85.315 138.380 ;
        RECT 85.395 138.060 85.715 138.380 ;
        RECT 102.705 138.060 103.025 138.380 ;
        RECT 103.105 138.060 103.425 138.380 ;
        RECT 103.505 138.060 103.825 138.380 ;
        RECT 103.905 138.060 104.225 138.380 ;
        RECT 121.215 138.060 121.535 138.380 ;
        RECT 121.615 138.060 121.935 138.380 ;
        RECT 122.015 138.060 122.335 138.380 ;
        RECT 122.415 138.060 122.735 138.380 ;
        RECT 74.940 135.340 75.260 135.660 ;
        RECT 75.340 135.340 75.660 135.660 ;
        RECT 75.740 135.340 76.060 135.660 ;
        RECT 76.140 135.340 76.460 135.660 ;
        RECT 93.450 135.340 93.770 135.660 ;
        RECT 93.850 135.340 94.170 135.660 ;
        RECT 94.250 135.340 94.570 135.660 ;
        RECT 94.650 135.340 94.970 135.660 ;
        RECT 111.960 135.340 112.280 135.660 ;
        RECT 112.360 135.340 112.680 135.660 ;
        RECT 112.760 135.340 113.080 135.660 ;
        RECT 113.160 135.340 113.480 135.660 ;
        RECT 130.470 135.340 130.790 135.660 ;
        RECT 130.870 135.340 131.190 135.660 ;
        RECT 131.270 135.340 131.590 135.660 ;
        RECT 131.670 135.340 131.990 135.660 ;
        RECT 65.685 132.620 66.005 132.940 ;
        RECT 66.085 132.620 66.405 132.940 ;
        RECT 66.485 132.620 66.805 132.940 ;
        RECT 66.885 132.620 67.205 132.940 ;
        RECT 84.195 132.620 84.515 132.940 ;
        RECT 84.595 132.620 84.915 132.940 ;
        RECT 84.995 132.620 85.315 132.940 ;
        RECT 85.395 132.620 85.715 132.940 ;
        RECT 102.705 132.620 103.025 132.940 ;
        RECT 103.105 132.620 103.425 132.940 ;
        RECT 103.505 132.620 103.825 132.940 ;
        RECT 103.905 132.620 104.225 132.940 ;
        RECT 121.215 132.620 121.535 132.940 ;
        RECT 121.615 132.620 121.935 132.940 ;
        RECT 122.015 132.620 122.335 132.940 ;
        RECT 122.415 132.620 122.735 132.940 ;
        RECT 74.940 129.900 75.260 130.220 ;
        RECT 75.340 129.900 75.660 130.220 ;
        RECT 75.740 129.900 76.060 130.220 ;
        RECT 76.140 129.900 76.460 130.220 ;
        RECT 93.450 129.900 93.770 130.220 ;
        RECT 93.850 129.900 94.170 130.220 ;
        RECT 94.250 129.900 94.570 130.220 ;
        RECT 94.650 129.900 94.970 130.220 ;
        RECT 111.960 129.900 112.280 130.220 ;
        RECT 112.360 129.900 112.680 130.220 ;
        RECT 112.760 129.900 113.080 130.220 ;
        RECT 113.160 129.900 113.480 130.220 ;
        RECT 130.470 129.900 130.790 130.220 ;
        RECT 130.870 129.900 131.190 130.220 ;
        RECT 131.270 129.900 131.590 130.220 ;
        RECT 131.670 129.900 131.990 130.220 ;
        RECT 65.630 123.230 67.130 124.730 ;
        RECT 84.050 123.170 85.550 124.670 ;
        RECT 102.760 123.230 104.260 124.730 ;
        RECT 121.180 123.230 122.680 124.730 ;
        RECT 1.005 120.145 2.495 121.635 ;
        RECT 135.000 99.000 136.000 101.000 ;
        RECT 135.000 95.000 136.000 97.000 ;
        RECT 10.000 87.000 11.000 93.000 ;
        RECT 134.000 77.000 136.000 78.000 ;
        RECT 60.000 69.000 61.000 75.000 ;
        RECT 156.000 77.000 158.000 78.000 ;
      LAYER met4 ;
        RECT 3.000 224.760 3.990 225.000 ;
        RECT 4.290 224.760 7.670 225.000 ;
        RECT 7.970 224.760 11.350 225.000 ;
        RECT 11.650 224.760 15.030 225.000 ;
        RECT 15.330 224.760 18.710 225.000 ;
        RECT 19.010 224.760 22.390 225.000 ;
        RECT 22.690 224.760 26.070 225.000 ;
        RECT 26.370 224.760 29.750 225.000 ;
        RECT 30.050 224.760 33.430 225.000 ;
        RECT 33.730 224.760 37.110 225.000 ;
        RECT 37.410 224.760 40.790 225.000 ;
        RECT 41.090 224.760 44.470 225.000 ;
        RECT 44.770 224.760 48.150 225.000 ;
        RECT 48.450 224.760 51.830 225.000 ;
        RECT 52.130 224.760 55.510 225.000 ;
        RECT 55.810 224.760 59.190 225.000 ;
        RECT 59.490 224.760 62.870 225.000 ;
        RECT 63.170 224.760 66.550 225.000 ;
        RECT 66.850 224.760 70.230 225.000 ;
        RECT 70.530 224.760 73.910 225.000 ;
        RECT 74.210 224.760 77.590 225.000 ;
        RECT 77.890 224.760 81.270 225.000 ;
        RECT 81.570 224.760 84.950 225.000 ;
        RECT 85.250 224.760 88.630 225.000 ;
        RECT 88.930 224.760 89.000 225.000 ;
        RECT 128.995 224.760 129.110 225.005 ;
        RECT 129.410 224.760 129.505 225.005 ;
        RECT 3.000 224.000 89.000 224.760 ;
        RECT 121.750 224.750 122.050 224.760 ;
        RECT 128.995 224.495 129.505 224.760 ;
        RECT 132.500 224.760 132.790 225.000 ;
        RECT 133.090 224.760 133.505 225.005 ;
        RECT 132.500 224.500 133.505 224.760 ;
        RECT 136.000 224.760 136.470 225.000 ;
        RECT 136.770 224.760 137.005 225.005 ;
        RECT 136.000 224.500 137.005 224.760 ;
        RECT 132.995 224.495 133.505 224.500 ;
        RECT 136.495 224.495 137.005 224.500 ;
        RECT 139.995 224.760 140.150 225.005 ;
        RECT 140.450 224.760 140.505 225.005 ;
        RECT 139.995 224.495 140.505 224.760 ;
        RECT 143.500 224.760 143.830 225.000 ;
        RECT 144.130 224.760 144.505 225.005 ;
        RECT 143.500 224.500 144.505 224.760 ;
        RECT 143.995 224.495 144.505 224.500 ;
        RECT 147.495 224.760 147.510 225.005 ;
        RECT 147.810 224.760 148.005 225.005 ;
        RECT 147.495 224.495 148.005 224.760 ;
        RECT 150.980 224.760 151.190 225.010 ;
        RECT 151.490 225.005 151.500 225.010 ;
        RECT 151.490 224.760 151.505 225.005 ;
        RECT 150.980 224.495 151.505 224.760 ;
        RECT 154.870 224.695 155.170 224.760 ;
        RECT 150.980 224.480 151.500 224.495 ;
        RECT 154.765 224.285 155.315 224.695 ;
        RECT 49.000 222.760 51.000 224.000 ;
        RECT 48.950 222.300 51.000 222.760 ;
        RECT 48.950 220.760 50.970 222.300 ;
        RECT 48.950 219.970 49.000 220.760 ;
        RECT 50.500 219.970 50.970 220.760 ;
        RECT 65.645 131.030 67.245 203.740 ;
        RECT 65.630 129.820 67.245 131.030 ;
        RECT 74.900 129.820 76.500 203.740 ;
        RECT 84.155 130.810 85.755 203.740 ;
        RECT 84.050 129.820 85.755 130.810 ;
        RECT 93.410 129.820 95.010 203.740 ;
        RECT 102.665 129.820 104.265 203.740 ;
        RECT 111.920 129.820 113.520 203.740 ;
        RECT 121.175 129.820 122.775 203.740 ;
        RECT 130.430 130.970 132.030 203.740 ;
        RECT 130.410 129.820 132.030 130.970 ;
        RECT 65.630 124.735 67.130 129.820 ;
        RECT 65.625 123.225 67.135 124.735 ;
        RECT 50.500 118.750 51.950 118.830 ;
        RECT 74.950 118.750 76.450 129.820 ;
        RECT 84.050 124.675 85.550 129.820 ;
        RECT 84.045 123.165 85.555 124.675 ;
        RECT 93.450 118.750 94.950 129.820 ;
        RECT 102.760 124.735 104.260 129.820 ;
        RECT 102.755 123.225 104.265 124.735 ;
        RECT 111.930 118.750 113.430 129.820 ;
        RECT 121.180 124.735 122.680 129.820 ;
        RECT 130.410 128.510 131.910 129.820 ;
        RECT 130.320 127.640 131.910 128.510 ;
        RECT 121.175 123.225 122.685 124.735 ;
        RECT 130.320 118.750 131.820 127.640 ;
        RECT 50.500 117.250 131.820 118.750 ;
        RECT 50.500 117.240 51.950 117.250 ;
        RECT 111.930 117.240 113.430 117.250 ;
        RECT 134.995 101.000 136.005 101.005 ;
        RECT 99.000 99.000 136.005 101.000 ;
        RECT 9.995 93.000 11.005 93.005 ;
        RECT 2.500 87.000 11.005 93.000 ;
        RECT 9.995 86.995 11.005 87.000 ;
        RECT 50.500 75.000 52.330 75.430 ;
        RECT 59.995 75.000 61.005 75.005 ;
        RECT 50.500 69.000 61.005 75.000 ;
        RECT 50.500 68.220 52.330 69.000 ;
        RECT 59.995 68.995 61.005 69.000 ;
        RECT 99.000 16.000 101.000 99.000 ;
        RECT 134.995 98.995 136.005 99.000 ;
        RECT 134.995 97.000 136.005 97.005 ;
        RECT 90.000 14.000 101.000 16.000 ;
        RECT 103.000 95.000 136.005 97.000 ;
        RECT 103.000 16.000 105.000 95.000 ;
        RECT 134.995 94.995 136.005 95.000 ;
        RECT 133.995 76.995 136.005 78.005 ;
        RECT 155.995 76.995 158.005 78.005 ;
        RECT 134.000 67.000 136.000 76.995 ;
        RECT 156.000 67.000 158.000 76.995 ;
        RECT 134.000 65.000 145.000 67.000 ;
        RECT 143.000 16.000 145.000 65.000 ;
        RECT 103.000 14.000 114.000 16.000 ;
        RECT 90.000 2.150 92.000 14.000 ;
        RECT 112.000 2.150 114.000 14.000 ;
        RECT 134.000 14.000 145.000 16.000 ;
        RECT 147.000 65.000 158.000 67.000 ;
        RECT 147.000 16.000 149.000 65.000 ;
        RECT 147.000 14.000 158.000 16.000 ;
        RECT 134.000 2.170 136.000 14.000 ;
        RECT 156.000 2.170 158.000 14.000 ;
        RECT 134.320 2.160 136.000 2.170 ;
        RECT 156.400 2.160 158.000 2.170 ;
        RECT 90.160 1.380 91.070 2.150 ;
        RECT 90.170 1.000 91.070 1.380 ;
        RECT 112.250 1.000 113.150 2.150 ;
        RECT 134.330 1.000 135.230 2.160 ;
        RECT 156.410 2.150 158.000 2.160 ;
        RECT 156.410 1.000 157.310 2.150 ;
  END
END tt_um_KolosKoblasz_mixer
END LIBRARY

