module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \top_I.branch[0].block[0].um_I.ana[2] ;
 wire \top_I.branch[0].block[0].um_I.ana[3] ;
 wire \top_I.branch[0].block[0].um_I.ana[4] ;
 wire \top_I.branch[0].block[0].um_I.ana[5] ;
 wire \top_I.branch[0].block[0].um_I.ana[6] ;
 wire \top_I.branch[0].block[0].um_I.ana[7] ;
 wire \top_I.branch[0].block[0].um_I.clk ;
 wire \top_I.branch[0].block[0].um_I.ena ;
 wire \top_I.branch[0].block[0].um_I.iw[10] ;
 wire \top_I.branch[0].block[0].um_I.iw[11] ;
 wire \top_I.branch[0].block[0].um_I.iw[12] ;
 wire \top_I.branch[0].block[0].um_I.iw[13] ;
 wire \top_I.branch[0].block[0].um_I.iw[14] ;
 wire \top_I.branch[0].block[0].um_I.iw[15] ;
 wire \top_I.branch[0].block[0].um_I.iw[16] ;
 wire \top_I.branch[0].block[0].um_I.iw[17] ;
 wire \top_I.branch[0].block[0].um_I.iw[1] ;
 wire \top_I.branch[0].block[0].um_I.iw[2] ;
 wire \top_I.branch[0].block[0].um_I.iw[3] ;
 wire \top_I.branch[0].block[0].um_I.iw[4] ;
 wire \top_I.branch[0].block[0].um_I.iw[5] ;
 wire \top_I.branch[0].block[0].um_I.iw[6] ;
 wire \top_I.branch[0].block[0].um_I.iw[7] ;
 wire \top_I.branch[0].block[0].um_I.iw[8] ;
 wire \top_I.branch[0].block[0].um_I.iw[9] ;
 wire \top_I.branch[0].block[0].um_I.k_zero ;
 wire \top_I.branch[0].block[0].um_I.ow[0] ;
 wire \top_I.branch[0].block[0].um_I.ow[10] ;
 wire \top_I.branch[0].block[0].um_I.ow[11] ;
 wire \top_I.branch[0].block[0].um_I.ow[12] ;
 wire \top_I.branch[0].block[0].um_I.ow[13] ;
 wire \top_I.branch[0].block[0].um_I.ow[14] ;
 wire \top_I.branch[0].block[0].um_I.ow[15] ;
 wire \top_I.branch[0].block[0].um_I.ow[16] ;
 wire \top_I.branch[0].block[0].um_I.ow[17] ;
 wire \top_I.branch[0].block[0].um_I.ow[18] ;
 wire \top_I.branch[0].block[0].um_I.ow[19] ;
 wire \top_I.branch[0].block[0].um_I.ow[1] ;
 wire \top_I.branch[0].block[0].um_I.ow[20] ;
 wire \top_I.branch[0].block[0].um_I.ow[21] ;
 wire \top_I.branch[0].block[0].um_I.ow[22] ;
 wire \top_I.branch[0].block[0].um_I.ow[23] ;
 wire \top_I.branch[0].block[0].um_I.ow[2] ;
 wire \top_I.branch[0].block[0].um_I.ow[3] ;
 wire \top_I.branch[0].block[0].um_I.ow[4] ;
 wire \top_I.branch[0].block[0].um_I.ow[5] ;
 wire \top_I.branch[0].block[0].um_I.ow[6] ;
 wire \top_I.branch[0].block[0].um_I.ow[7] ;
 wire \top_I.branch[0].block[0].um_I.ow[8] ;
 wire \top_I.branch[0].block[0].um_I.ow[9] ;
 wire \top_I.branch[0].block[0].um_I.pg_vdd ;
 wire \top_I.branch[0].block[10].um_I.ana[2] ;
 wire \top_I.branch[0].block[10].um_I.ana[3] ;
 wire \top_I.branch[0].block[10].um_I.ana[4] ;
 wire \top_I.branch[0].block[10].um_I.ana[5] ;
 wire \top_I.branch[0].block[10].um_I.ana[6] ;
 wire \top_I.branch[0].block[10].um_I.ana[7] ;
 wire \top_I.branch[0].block[10].um_I.clk ;
 wire \top_I.branch[0].block[10].um_I.ena ;
 wire \top_I.branch[0].block[10].um_I.iw[10] ;
 wire \top_I.branch[0].block[10].um_I.iw[11] ;
 wire \top_I.branch[0].block[10].um_I.iw[12] ;
 wire \top_I.branch[0].block[10].um_I.iw[13] ;
 wire \top_I.branch[0].block[10].um_I.iw[14] ;
 wire \top_I.branch[0].block[10].um_I.iw[15] ;
 wire \top_I.branch[0].block[10].um_I.iw[16] ;
 wire \top_I.branch[0].block[10].um_I.iw[17] ;
 wire \top_I.branch[0].block[10].um_I.iw[1] ;
 wire \top_I.branch[0].block[10].um_I.iw[2] ;
 wire \top_I.branch[0].block[10].um_I.iw[3] ;
 wire \top_I.branch[0].block[10].um_I.iw[4] ;
 wire \top_I.branch[0].block[10].um_I.iw[5] ;
 wire \top_I.branch[0].block[10].um_I.iw[6] ;
 wire \top_I.branch[0].block[10].um_I.iw[7] ;
 wire \top_I.branch[0].block[10].um_I.iw[8] ;
 wire \top_I.branch[0].block[10].um_I.iw[9] ;
 wire \top_I.branch[0].block[10].um_I.k_zero ;
 wire \top_I.branch[0].block[10].um_I.pg_vdd ;
 wire \top_I.branch[0].block[11].um_I.ana[2] ;
 wire \top_I.branch[0].block[11].um_I.ana[3] ;
 wire \top_I.branch[0].block[11].um_I.ana[4] ;
 wire \top_I.branch[0].block[11].um_I.ana[5] ;
 wire \top_I.branch[0].block[11].um_I.ana[6] ;
 wire \top_I.branch[0].block[11].um_I.ana[7] ;
 wire \top_I.branch[0].block[11].um_I.clk ;
 wire \top_I.branch[0].block[11].um_I.ena ;
 wire \top_I.branch[0].block[11].um_I.iw[10] ;
 wire \top_I.branch[0].block[11].um_I.iw[11] ;
 wire \top_I.branch[0].block[11].um_I.iw[12] ;
 wire \top_I.branch[0].block[11].um_I.iw[13] ;
 wire \top_I.branch[0].block[11].um_I.iw[14] ;
 wire \top_I.branch[0].block[11].um_I.iw[15] ;
 wire \top_I.branch[0].block[11].um_I.iw[16] ;
 wire \top_I.branch[0].block[11].um_I.iw[17] ;
 wire \top_I.branch[0].block[11].um_I.iw[1] ;
 wire \top_I.branch[0].block[11].um_I.iw[2] ;
 wire \top_I.branch[0].block[11].um_I.iw[3] ;
 wire \top_I.branch[0].block[11].um_I.iw[4] ;
 wire \top_I.branch[0].block[11].um_I.iw[5] ;
 wire \top_I.branch[0].block[11].um_I.iw[6] ;
 wire \top_I.branch[0].block[11].um_I.iw[7] ;
 wire \top_I.branch[0].block[11].um_I.iw[8] ;
 wire \top_I.branch[0].block[11].um_I.iw[9] ;
 wire \top_I.branch[0].block[11].um_I.k_zero ;
 wire \top_I.branch[0].block[11].um_I.pg_vdd ;
 wire \top_I.branch[0].block[12].um_I.ana[2] ;
 wire \top_I.branch[0].block[12].um_I.ana[3] ;
 wire \top_I.branch[0].block[12].um_I.ana[4] ;
 wire \top_I.branch[0].block[12].um_I.ana[5] ;
 wire \top_I.branch[0].block[12].um_I.ana[6] ;
 wire \top_I.branch[0].block[12].um_I.ana[7] ;
 wire \top_I.branch[0].block[12].um_I.clk ;
 wire \top_I.branch[0].block[12].um_I.ena ;
 wire \top_I.branch[0].block[12].um_I.iw[10] ;
 wire \top_I.branch[0].block[12].um_I.iw[11] ;
 wire \top_I.branch[0].block[12].um_I.iw[12] ;
 wire \top_I.branch[0].block[12].um_I.iw[13] ;
 wire \top_I.branch[0].block[12].um_I.iw[14] ;
 wire \top_I.branch[0].block[12].um_I.iw[15] ;
 wire \top_I.branch[0].block[12].um_I.iw[16] ;
 wire \top_I.branch[0].block[12].um_I.iw[17] ;
 wire \top_I.branch[0].block[12].um_I.iw[1] ;
 wire \top_I.branch[0].block[12].um_I.iw[2] ;
 wire \top_I.branch[0].block[12].um_I.iw[3] ;
 wire \top_I.branch[0].block[12].um_I.iw[4] ;
 wire \top_I.branch[0].block[12].um_I.iw[5] ;
 wire \top_I.branch[0].block[12].um_I.iw[6] ;
 wire \top_I.branch[0].block[12].um_I.iw[7] ;
 wire \top_I.branch[0].block[12].um_I.iw[8] ;
 wire \top_I.branch[0].block[12].um_I.iw[9] ;
 wire \top_I.branch[0].block[12].um_I.k_zero ;
 wire \top_I.branch[0].block[12].um_I.pg_vdd ;
 wire \top_I.branch[0].block[13].um_I.ana[2] ;
 wire \top_I.branch[0].block[13].um_I.ana[3] ;
 wire \top_I.branch[0].block[13].um_I.ana[4] ;
 wire \top_I.branch[0].block[13].um_I.ana[5] ;
 wire \top_I.branch[0].block[13].um_I.ana[6] ;
 wire \top_I.branch[0].block[13].um_I.ana[7] ;
 wire \top_I.branch[0].block[13].um_I.clk ;
 wire \top_I.branch[0].block[13].um_I.ena ;
 wire \top_I.branch[0].block[13].um_I.iw[10] ;
 wire \top_I.branch[0].block[13].um_I.iw[11] ;
 wire \top_I.branch[0].block[13].um_I.iw[12] ;
 wire \top_I.branch[0].block[13].um_I.iw[13] ;
 wire \top_I.branch[0].block[13].um_I.iw[14] ;
 wire \top_I.branch[0].block[13].um_I.iw[15] ;
 wire \top_I.branch[0].block[13].um_I.iw[16] ;
 wire \top_I.branch[0].block[13].um_I.iw[17] ;
 wire \top_I.branch[0].block[13].um_I.iw[1] ;
 wire \top_I.branch[0].block[13].um_I.iw[2] ;
 wire \top_I.branch[0].block[13].um_I.iw[3] ;
 wire \top_I.branch[0].block[13].um_I.iw[4] ;
 wire \top_I.branch[0].block[13].um_I.iw[5] ;
 wire \top_I.branch[0].block[13].um_I.iw[6] ;
 wire \top_I.branch[0].block[13].um_I.iw[7] ;
 wire \top_I.branch[0].block[13].um_I.iw[8] ;
 wire \top_I.branch[0].block[13].um_I.iw[9] ;
 wire \top_I.branch[0].block[13].um_I.k_zero ;
 wire \top_I.branch[0].block[13].um_I.pg_vdd ;
 wire \top_I.branch[0].block[14].um_I.ana[2] ;
 wire \top_I.branch[0].block[14].um_I.ana[3] ;
 wire \top_I.branch[0].block[14].um_I.ana[4] ;
 wire \top_I.branch[0].block[14].um_I.ana[5] ;
 wire \top_I.branch[0].block[14].um_I.ana[6] ;
 wire \top_I.branch[0].block[14].um_I.ana[7] ;
 wire \top_I.branch[0].block[14].um_I.clk ;
 wire \top_I.branch[0].block[14].um_I.ena ;
 wire \top_I.branch[0].block[14].um_I.iw[10] ;
 wire \top_I.branch[0].block[14].um_I.iw[11] ;
 wire \top_I.branch[0].block[14].um_I.iw[12] ;
 wire \top_I.branch[0].block[14].um_I.iw[13] ;
 wire \top_I.branch[0].block[14].um_I.iw[14] ;
 wire \top_I.branch[0].block[14].um_I.iw[15] ;
 wire \top_I.branch[0].block[14].um_I.iw[16] ;
 wire \top_I.branch[0].block[14].um_I.iw[17] ;
 wire \top_I.branch[0].block[14].um_I.iw[1] ;
 wire \top_I.branch[0].block[14].um_I.iw[2] ;
 wire \top_I.branch[0].block[14].um_I.iw[3] ;
 wire \top_I.branch[0].block[14].um_I.iw[4] ;
 wire \top_I.branch[0].block[14].um_I.iw[5] ;
 wire \top_I.branch[0].block[14].um_I.iw[6] ;
 wire \top_I.branch[0].block[14].um_I.iw[7] ;
 wire \top_I.branch[0].block[14].um_I.iw[8] ;
 wire \top_I.branch[0].block[14].um_I.iw[9] ;
 wire \top_I.branch[0].block[14].um_I.k_zero ;
 wire \top_I.branch[0].block[14].um_I.pg_vdd ;
 wire \top_I.branch[0].block[15].um_I.ana[2] ;
 wire \top_I.branch[0].block[15].um_I.ana[3] ;
 wire \top_I.branch[0].block[15].um_I.ana[4] ;
 wire \top_I.branch[0].block[15].um_I.ana[5] ;
 wire \top_I.branch[0].block[15].um_I.ana[6] ;
 wire \top_I.branch[0].block[15].um_I.ana[7] ;
 wire \top_I.branch[0].block[15].um_I.clk ;
 wire \top_I.branch[0].block[15].um_I.ena ;
 wire \top_I.branch[0].block[15].um_I.iw[10] ;
 wire \top_I.branch[0].block[15].um_I.iw[11] ;
 wire \top_I.branch[0].block[15].um_I.iw[12] ;
 wire \top_I.branch[0].block[15].um_I.iw[13] ;
 wire \top_I.branch[0].block[15].um_I.iw[14] ;
 wire \top_I.branch[0].block[15].um_I.iw[15] ;
 wire \top_I.branch[0].block[15].um_I.iw[16] ;
 wire \top_I.branch[0].block[15].um_I.iw[17] ;
 wire \top_I.branch[0].block[15].um_I.iw[1] ;
 wire \top_I.branch[0].block[15].um_I.iw[2] ;
 wire \top_I.branch[0].block[15].um_I.iw[3] ;
 wire \top_I.branch[0].block[15].um_I.iw[4] ;
 wire \top_I.branch[0].block[15].um_I.iw[5] ;
 wire \top_I.branch[0].block[15].um_I.iw[6] ;
 wire \top_I.branch[0].block[15].um_I.iw[7] ;
 wire \top_I.branch[0].block[15].um_I.iw[8] ;
 wire \top_I.branch[0].block[15].um_I.iw[9] ;
 wire \top_I.branch[0].block[15].um_I.k_zero ;
 wire \top_I.branch[0].block[15].um_I.pg_vdd ;
 wire \top_I.branch[0].block[1].um_I.ana[2] ;
 wire \top_I.branch[0].block[1].um_I.ana[3] ;
 wire \top_I.branch[0].block[1].um_I.ana[4] ;
 wire \top_I.branch[0].block[1].um_I.ana[5] ;
 wire \top_I.branch[0].block[1].um_I.ana[6] ;
 wire \top_I.branch[0].block[1].um_I.ana[7] ;
 wire \top_I.branch[0].block[1].um_I.clk ;
 wire \top_I.branch[0].block[1].um_I.ena ;
 wire \top_I.branch[0].block[1].um_I.iw[10] ;
 wire \top_I.branch[0].block[1].um_I.iw[11] ;
 wire \top_I.branch[0].block[1].um_I.iw[12] ;
 wire \top_I.branch[0].block[1].um_I.iw[13] ;
 wire \top_I.branch[0].block[1].um_I.iw[14] ;
 wire \top_I.branch[0].block[1].um_I.iw[15] ;
 wire \top_I.branch[0].block[1].um_I.iw[16] ;
 wire \top_I.branch[0].block[1].um_I.iw[17] ;
 wire \top_I.branch[0].block[1].um_I.iw[1] ;
 wire \top_I.branch[0].block[1].um_I.iw[2] ;
 wire \top_I.branch[0].block[1].um_I.iw[3] ;
 wire \top_I.branch[0].block[1].um_I.iw[4] ;
 wire \top_I.branch[0].block[1].um_I.iw[5] ;
 wire \top_I.branch[0].block[1].um_I.iw[6] ;
 wire \top_I.branch[0].block[1].um_I.iw[7] ;
 wire \top_I.branch[0].block[1].um_I.iw[8] ;
 wire \top_I.branch[0].block[1].um_I.iw[9] ;
 wire \top_I.branch[0].block[1].um_I.k_zero ;
 wire \top_I.branch[0].block[1].um_I.ow[0] ;
 wire \top_I.branch[0].block[1].um_I.ow[10] ;
 wire \top_I.branch[0].block[1].um_I.ow[11] ;
 wire \top_I.branch[0].block[1].um_I.ow[12] ;
 wire \top_I.branch[0].block[1].um_I.ow[13] ;
 wire \top_I.branch[0].block[1].um_I.ow[14] ;
 wire \top_I.branch[0].block[1].um_I.ow[15] ;
 wire \top_I.branch[0].block[1].um_I.ow[16] ;
 wire \top_I.branch[0].block[1].um_I.ow[17] ;
 wire \top_I.branch[0].block[1].um_I.ow[18] ;
 wire \top_I.branch[0].block[1].um_I.ow[19] ;
 wire \top_I.branch[0].block[1].um_I.ow[1] ;
 wire \top_I.branch[0].block[1].um_I.ow[20] ;
 wire \top_I.branch[0].block[1].um_I.ow[21] ;
 wire \top_I.branch[0].block[1].um_I.ow[22] ;
 wire \top_I.branch[0].block[1].um_I.ow[23] ;
 wire \top_I.branch[0].block[1].um_I.ow[2] ;
 wire \top_I.branch[0].block[1].um_I.ow[3] ;
 wire \top_I.branch[0].block[1].um_I.ow[4] ;
 wire \top_I.branch[0].block[1].um_I.ow[5] ;
 wire \top_I.branch[0].block[1].um_I.ow[6] ;
 wire \top_I.branch[0].block[1].um_I.ow[7] ;
 wire \top_I.branch[0].block[1].um_I.ow[8] ;
 wire \top_I.branch[0].block[1].um_I.ow[9] ;
 wire \top_I.branch[0].block[1].um_I.pg_vdd ;
 wire \top_I.branch[0].block[2].um_I.ana[2] ;
 wire \top_I.branch[0].block[2].um_I.ana[3] ;
 wire \top_I.branch[0].block[2].um_I.ana[4] ;
 wire \top_I.branch[0].block[2].um_I.ana[5] ;
 wire \top_I.branch[0].block[2].um_I.ana[6] ;
 wire \top_I.branch[0].block[2].um_I.ana[7] ;
 wire \top_I.branch[0].block[2].um_I.clk ;
 wire \top_I.branch[0].block[2].um_I.ena ;
 wire \top_I.branch[0].block[2].um_I.iw[10] ;
 wire \top_I.branch[0].block[2].um_I.iw[11] ;
 wire \top_I.branch[0].block[2].um_I.iw[12] ;
 wire \top_I.branch[0].block[2].um_I.iw[13] ;
 wire \top_I.branch[0].block[2].um_I.iw[14] ;
 wire \top_I.branch[0].block[2].um_I.iw[15] ;
 wire \top_I.branch[0].block[2].um_I.iw[16] ;
 wire \top_I.branch[0].block[2].um_I.iw[17] ;
 wire \top_I.branch[0].block[2].um_I.iw[1] ;
 wire \top_I.branch[0].block[2].um_I.iw[2] ;
 wire \top_I.branch[0].block[2].um_I.iw[3] ;
 wire \top_I.branch[0].block[2].um_I.iw[4] ;
 wire \top_I.branch[0].block[2].um_I.iw[5] ;
 wire \top_I.branch[0].block[2].um_I.iw[6] ;
 wire \top_I.branch[0].block[2].um_I.iw[7] ;
 wire \top_I.branch[0].block[2].um_I.iw[8] ;
 wire \top_I.branch[0].block[2].um_I.iw[9] ;
 wire \top_I.branch[0].block[2].um_I.k_zero ;
 wire \top_I.branch[0].block[2].um_I.pg_vdd ;
 wire \top_I.branch[0].block[3].um_I.ana[2] ;
 wire \top_I.branch[0].block[3].um_I.ana[3] ;
 wire \top_I.branch[0].block[3].um_I.ana[4] ;
 wire \top_I.branch[0].block[3].um_I.ana[5] ;
 wire \top_I.branch[0].block[3].um_I.ana[6] ;
 wire \top_I.branch[0].block[3].um_I.ana[7] ;
 wire \top_I.branch[0].block[3].um_I.clk ;
 wire \top_I.branch[0].block[3].um_I.ena ;
 wire \top_I.branch[0].block[3].um_I.iw[10] ;
 wire \top_I.branch[0].block[3].um_I.iw[11] ;
 wire \top_I.branch[0].block[3].um_I.iw[12] ;
 wire \top_I.branch[0].block[3].um_I.iw[13] ;
 wire \top_I.branch[0].block[3].um_I.iw[14] ;
 wire \top_I.branch[0].block[3].um_I.iw[15] ;
 wire \top_I.branch[0].block[3].um_I.iw[16] ;
 wire \top_I.branch[0].block[3].um_I.iw[17] ;
 wire \top_I.branch[0].block[3].um_I.iw[1] ;
 wire \top_I.branch[0].block[3].um_I.iw[2] ;
 wire \top_I.branch[0].block[3].um_I.iw[3] ;
 wire \top_I.branch[0].block[3].um_I.iw[4] ;
 wire \top_I.branch[0].block[3].um_I.iw[5] ;
 wire \top_I.branch[0].block[3].um_I.iw[6] ;
 wire \top_I.branch[0].block[3].um_I.iw[7] ;
 wire \top_I.branch[0].block[3].um_I.iw[8] ;
 wire \top_I.branch[0].block[3].um_I.iw[9] ;
 wire \top_I.branch[0].block[3].um_I.k_zero ;
 wire \top_I.branch[0].block[3].um_I.pg_vdd ;
 wire \top_I.branch[0].block[4].um_I.ana[2] ;
 wire \top_I.branch[0].block[4].um_I.ana[3] ;
 wire \top_I.branch[0].block[4].um_I.ana[4] ;
 wire \top_I.branch[0].block[4].um_I.ana[5] ;
 wire \top_I.branch[0].block[4].um_I.ana[6] ;
 wire \top_I.branch[0].block[4].um_I.ana[7] ;
 wire \top_I.branch[0].block[4].um_I.clk ;
 wire \top_I.branch[0].block[4].um_I.ena ;
 wire \top_I.branch[0].block[4].um_I.iw[10] ;
 wire \top_I.branch[0].block[4].um_I.iw[11] ;
 wire \top_I.branch[0].block[4].um_I.iw[12] ;
 wire \top_I.branch[0].block[4].um_I.iw[13] ;
 wire \top_I.branch[0].block[4].um_I.iw[14] ;
 wire \top_I.branch[0].block[4].um_I.iw[15] ;
 wire \top_I.branch[0].block[4].um_I.iw[16] ;
 wire \top_I.branch[0].block[4].um_I.iw[17] ;
 wire \top_I.branch[0].block[4].um_I.iw[1] ;
 wire \top_I.branch[0].block[4].um_I.iw[2] ;
 wire \top_I.branch[0].block[4].um_I.iw[3] ;
 wire \top_I.branch[0].block[4].um_I.iw[4] ;
 wire \top_I.branch[0].block[4].um_I.iw[5] ;
 wire \top_I.branch[0].block[4].um_I.iw[6] ;
 wire \top_I.branch[0].block[4].um_I.iw[7] ;
 wire \top_I.branch[0].block[4].um_I.iw[8] ;
 wire \top_I.branch[0].block[4].um_I.iw[9] ;
 wire \top_I.branch[0].block[4].um_I.k_zero ;
 wire \top_I.branch[0].block[4].um_I.pg_vdd ;
 wire \top_I.branch[0].block[5].um_I.ana[2] ;
 wire \top_I.branch[0].block[5].um_I.ana[3] ;
 wire \top_I.branch[0].block[5].um_I.ana[4] ;
 wire \top_I.branch[0].block[5].um_I.ana[5] ;
 wire \top_I.branch[0].block[5].um_I.ana[6] ;
 wire \top_I.branch[0].block[5].um_I.ana[7] ;
 wire \top_I.branch[0].block[5].um_I.clk ;
 wire \top_I.branch[0].block[5].um_I.ena ;
 wire \top_I.branch[0].block[5].um_I.iw[10] ;
 wire \top_I.branch[0].block[5].um_I.iw[11] ;
 wire \top_I.branch[0].block[5].um_I.iw[12] ;
 wire \top_I.branch[0].block[5].um_I.iw[13] ;
 wire \top_I.branch[0].block[5].um_I.iw[14] ;
 wire \top_I.branch[0].block[5].um_I.iw[15] ;
 wire \top_I.branch[0].block[5].um_I.iw[16] ;
 wire \top_I.branch[0].block[5].um_I.iw[17] ;
 wire \top_I.branch[0].block[5].um_I.iw[1] ;
 wire \top_I.branch[0].block[5].um_I.iw[2] ;
 wire \top_I.branch[0].block[5].um_I.iw[3] ;
 wire \top_I.branch[0].block[5].um_I.iw[4] ;
 wire \top_I.branch[0].block[5].um_I.iw[5] ;
 wire \top_I.branch[0].block[5].um_I.iw[6] ;
 wire \top_I.branch[0].block[5].um_I.iw[7] ;
 wire \top_I.branch[0].block[5].um_I.iw[8] ;
 wire \top_I.branch[0].block[5].um_I.iw[9] ;
 wire \top_I.branch[0].block[5].um_I.k_zero ;
 wire \top_I.branch[0].block[5].um_I.pg_vdd ;
 wire \top_I.branch[0].block[6].um_I.ana[2] ;
 wire \top_I.branch[0].block[6].um_I.ana[3] ;
 wire \top_I.branch[0].block[6].um_I.ana[4] ;
 wire \top_I.branch[0].block[6].um_I.ana[5] ;
 wire \top_I.branch[0].block[6].um_I.ana[6] ;
 wire \top_I.branch[0].block[6].um_I.ana[7] ;
 wire \top_I.branch[0].block[6].um_I.clk ;
 wire \top_I.branch[0].block[6].um_I.ena ;
 wire \top_I.branch[0].block[6].um_I.iw[10] ;
 wire \top_I.branch[0].block[6].um_I.iw[11] ;
 wire \top_I.branch[0].block[6].um_I.iw[12] ;
 wire \top_I.branch[0].block[6].um_I.iw[13] ;
 wire \top_I.branch[0].block[6].um_I.iw[14] ;
 wire \top_I.branch[0].block[6].um_I.iw[15] ;
 wire \top_I.branch[0].block[6].um_I.iw[16] ;
 wire \top_I.branch[0].block[6].um_I.iw[17] ;
 wire \top_I.branch[0].block[6].um_I.iw[1] ;
 wire \top_I.branch[0].block[6].um_I.iw[2] ;
 wire \top_I.branch[0].block[6].um_I.iw[3] ;
 wire \top_I.branch[0].block[6].um_I.iw[4] ;
 wire \top_I.branch[0].block[6].um_I.iw[5] ;
 wire \top_I.branch[0].block[6].um_I.iw[6] ;
 wire \top_I.branch[0].block[6].um_I.iw[7] ;
 wire \top_I.branch[0].block[6].um_I.iw[8] ;
 wire \top_I.branch[0].block[6].um_I.iw[9] ;
 wire \top_I.branch[0].block[6].um_I.k_zero ;
 wire \top_I.branch[0].block[6].um_I.pg_vdd ;
 wire \top_I.branch[0].block[7].um_I.ana[2] ;
 wire \top_I.branch[0].block[7].um_I.ana[3] ;
 wire \top_I.branch[0].block[7].um_I.ana[4] ;
 wire \top_I.branch[0].block[7].um_I.ana[5] ;
 wire \top_I.branch[0].block[7].um_I.ana[6] ;
 wire \top_I.branch[0].block[7].um_I.ana[7] ;
 wire \top_I.branch[0].block[7].um_I.clk ;
 wire \top_I.branch[0].block[7].um_I.ena ;
 wire \top_I.branch[0].block[7].um_I.iw[10] ;
 wire \top_I.branch[0].block[7].um_I.iw[11] ;
 wire \top_I.branch[0].block[7].um_I.iw[12] ;
 wire \top_I.branch[0].block[7].um_I.iw[13] ;
 wire \top_I.branch[0].block[7].um_I.iw[14] ;
 wire \top_I.branch[0].block[7].um_I.iw[15] ;
 wire \top_I.branch[0].block[7].um_I.iw[16] ;
 wire \top_I.branch[0].block[7].um_I.iw[17] ;
 wire \top_I.branch[0].block[7].um_I.iw[1] ;
 wire \top_I.branch[0].block[7].um_I.iw[2] ;
 wire \top_I.branch[0].block[7].um_I.iw[3] ;
 wire \top_I.branch[0].block[7].um_I.iw[4] ;
 wire \top_I.branch[0].block[7].um_I.iw[5] ;
 wire \top_I.branch[0].block[7].um_I.iw[6] ;
 wire \top_I.branch[0].block[7].um_I.iw[7] ;
 wire \top_I.branch[0].block[7].um_I.iw[8] ;
 wire \top_I.branch[0].block[7].um_I.iw[9] ;
 wire \top_I.branch[0].block[7].um_I.k_zero ;
 wire \top_I.branch[0].block[7].um_I.pg_vdd ;
 wire \top_I.branch[0].block[8].um_I.ana[2] ;
 wire \top_I.branch[0].block[8].um_I.ana[3] ;
 wire \top_I.branch[0].block[8].um_I.ana[4] ;
 wire \top_I.branch[0].block[8].um_I.ana[5] ;
 wire \top_I.branch[0].block[8].um_I.ana[6] ;
 wire \top_I.branch[0].block[8].um_I.ana[7] ;
 wire \top_I.branch[0].block[8].um_I.clk ;
 wire \top_I.branch[0].block[8].um_I.ena ;
 wire \top_I.branch[0].block[8].um_I.iw[10] ;
 wire \top_I.branch[0].block[8].um_I.iw[11] ;
 wire \top_I.branch[0].block[8].um_I.iw[12] ;
 wire \top_I.branch[0].block[8].um_I.iw[13] ;
 wire \top_I.branch[0].block[8].um_I.iw[14] ;
 wire \top_I.branch[0].block[8].um_I.iw[15] ;
 wire \top_I.branch[0].block[8].um_I.iw[16] ;
 wire \top_I.branch[0].block[8].um_I.iw[17] ;
 wire \top_I.branch[0].block[8].um_I.iw[1] ;
 wire \top_I.branch[0].block[8].um_I.iw[2] ;
 wire \top_I.branch[0].block[8].um_I.iw[3] ;
 wire \top_I.branch[0].block[8].um_I.iw[4] ;
 wire \top_I.branch[0].block[8].um_I.iw[5] ;
 wire \top_I.branch[0].block[8].um_I.iw[6] ;
 wire \top_I.branch[0].block[8].um_I.iw[7] ;
 wire \top_I.branch[0].block[8].um_I.iw[8] ;
 wire \top_I.branch[0].block[8].um_I.iw[9] ;
 wire \top_I.branch[0].block[8].um_I.k_zero ;
 wire \top_I.branch[0].block[8].um_I.pg_vdd ;
 wire \top_I.branch[0].block[9].um_I.ana[2] ;
 wire \top_I.branch[0].block[9].um_I.ana[3] ;
 wire \top_I.branch[0].block[9].um_I.ana[4] ;
 wire \top_I.branch[0].block[9].um_I.ana[5] ;
 wire \top_I.branch[0].block[9].um_I.ana[6] ;
 wire \top_I.branch[0].block[9].um_I.ana[7] ;
 wire \top_I.branch[0].block[9].um_I.clk ;
 wire \top_I.branch[0].block[9].um_I.ena ;
 wire \top_I.branch[0].block[9].um_I.iw[10] ;
 wire \top_I.branch[0].block[9].um_I.iw[11] ;
 wire \top_I.branch[0].block[9].um_I.iw[12] ;
 wire \top_I.branch[0].block[9].um_I.iw[13] ;
 wire \top_I.branch[0].block[9].um_I.iw[14] ;
 wire \top_I.branch[0].block[9].um_I.iw[15] ;
 wire \top_I.branch[0].block[9].um_I.iw[16] ;
 wire \top_I.branch[0].block[9].um_I.iw[17] ;
 wire \top_I.branch[0].block[9].um_I.iw[1] ;
 wire \top_I.branch[0].block[9].um_I.iw[2] ;
 wire \top_I.branch[0].block[9].um_I.iw[3] ;
 wire \top_I.branch[0].block[9].um_I.iw[4] ;
 wire \top_I.branch[0].block[9].um_I.iw[5] ;
 wire \top_I.branch[0].block[9].um_I.iw[6] ;
 wire \top_I.branch[0].block[9].um_I.iw[7] ;
 wire \top_I.branch[0].block[9].um_I.iw[8] ;
 wire \top_I.branch[0].block[9].um_I.iw[9] ;
 wire \top_I.branch[0].block[9].um_I.k_zero ;
 wire \top_I.branch[0].block[9].um_I.pg_vdd ;
 wire \top_I.branch[0].l_addr[0] ;
 wire \top_I.branch[0].l_k_one ;
 wire \top_I.branch[0].l_spine_iw[0] ;
 wire \top_I.branch[0].l_spine_iw[10] ;
 wire \top_I.branch[0].l_spine_iw[11] ;
 wire \top_I.branch[0].l_spine_iw[12] ;
 wire \top_I.branch[0].l_spine_iw[13] ;
 wire \top_I.branch[0].l_spine_iw[14] ;
 wire \top_I.branch[0].l_spine_iw[15] ;
 wire \top_I.branch[0].l_spine_iw[16] ;
 wire \top_I.branch[0].l_spine_iw[17] ;
 wire \top_I.branch[0].l_spine_iw[18] ;
 wire \top_I.branch[0].l_spine_iw[19] ;
 wire \top_I.branch[0].l_spine_iw[1] ;
 wire \top_I.branch[0].l_spine_iw[20] ;
 wire \top_I.branch[0].l_spine_iw[21] ;
 wire \top_I.branch[0].l_spine_iw[22] ;
 wire \top_I.branch[0].l_spine_iw[23] ;
 wire \top_I.branch[0].l_spine_iw[24] ;
 wire \top_I.branch[0].l_spine_iw[25] ;
 wire \top_I.branch[0].l_spine_iw[26] ;
 wire \top_I.branch[0].l_spine_iw[27] ;
 wire \top_I.branch[0].l_spine_iw[28] ;
 wire \top_I.branch[0].l_spine_iw[29] ;
 wire \top_I.branch[0].l_spine_iw[2] ;
 wire \top_I.branch[0].l_spine_iw[3] ;
 wire \top_I.branch[0].l_spine_iw[4] ;
 wire \top_I.branch[0].l_spine_iw[5] ;
 wire \top_I.branch[0].l_spine_iw[6] ;
 wire \top_I.branch[0].l_spine_iw[7] ;
 wire \top_I.branch[0].l_spine_iw[8] ;
 wire \top_I.branch[0].l_spine_iw[9] ;
 wire \top_I.branch[0].l_spine_ow[0] ;
 wire \top_I.branch[0].l_spine_ow[10] ;
 wire \top_I.branch[0].l_spine_ow[11] ;
 wire \top_I.branch[0].l_spine_ow[12] ;
 wire \top_I.branch[0].l_spine_ow[13] ;
 wire \top_I.branch[0].l_spine_ow[14] ;
 wire \top_I.branch[0].l_spine_ow[15] ;
 wire \top_I.branch[0].l_spine_ow[16] ;
 wire \top_I.branch[0].l_spine_ow[17] ;
 wire \top_I.branch[0].l_spine_ow[18] ;
 wire \top_I.branch[0].l_spine_ow[19] ;
 wire \top_I.branch[0].l_spine_ow[1] ;
 wire \top_I.branch[0].l_spine_ow[20] ;
 wire \top_I.branch[0].l_spine_ow[21] ;
 wire \top_I.branch[0].l_spine_ow[22] ;
 wire \top_I.branch[0].l_spine_ow[23] ;
 wire \top_I.branch[0].l_spine_ow[24] ;
 wire \top_I.branch[0].l_spine_ow[25] ;
 wire \top_I.branch[0].l_spine_ow[2] ;
 wire \top_I.branch[0].l_spine_ow[3] ;
 wire \top_I.branch[0].l_spine_ow[4] ;
 wire \top_I.branch[0].l_spine_ow[5] ;
 wire \top_I.branch[0].l_spine_ow[6] ;
 wire \top_I.branch[0].l_spine_ow[7] ;
 wire \top_I.branch[0].l_spine_ow[8] ;
 wire \top_I.branch[0].l_spine_ow[9] ;
 wire \top_I.branch[10].block[0].um_I.ana[2] ;
 wire \top_I.branch[10].block[0].um_I.ana[3] ;
 wire \top_I.branch[10].block[0].um_I.ana[4] ;
 wire \top_I.branch[10].block[0].um_I.ana[5] ;
 wire \top_I.branch[10].block[0].um_I.ana[6] ;
 wire \top_I.branch[10].block[0].um_I.ana[7] ;
 wire \top_I.branch[10].block[0].um_I.clk ;
 wire \top_I.branch[10].block[0].um_I.ena ;
 wire \top_I.branch[10].block[0].um_I.iw[10] ;
 wire \top_I.branch[10].block[0].um_I.iw[11] ;
 wire \top_I.branch[10].block[0].um_I.iw[12] ;
 wire \top_I.branch[10].block[0].um_I.iw[13] ;
 wire \top_I.branch[10].block[0].um_I.iw[14] ;
 wire \top_I.branch[10].block[0].um_I.iw[15] ;
 wire \top_I.branch[10].block[0].um_I.iw[16] ;
 wire \top_I.branch[10].block[0].um_I.iw[17] ;
 wire \top_I.branch[10].block[0].um_I.iw[1] ;
 wire \top_I.branch[10].block[0].um_I.iw[2] ;
 wire \top_I.branch[10].block[0].um_I.iw[3] ;
 wire \top_I.branch[10].block[0].um_I.iw[4] ;
 wire \top_I.branch[10].block[0].um_I.iw[5] ;
 wire \top_I.branch[10].block[0].um_I.iw[6] ;
 wire \top_I.branch[10].block[0].um_I.iw[7] ;
 wire \top_I.branch[10].block[0].um_I.iw[8] ;
 wire \top_I.branch[10].block[0].um_I.iw[9] ;
 wire \top_I.branch[10].block[0].um_I.k_zero ;
 wire \top_I.branch[10].block[0].um_I.pg_vdd ;
 wire \top_I.branch[10].block[10].um_I.ana[2] ;
 wire \top_I.branch[10].block[10].um_I.ana[3] ;
 wire \top_I.branch[10].block[10].um_I.ana[4] ;
 wire \top_I.branch[10].block[10].um_I.ana[5] ;
 wire \top_I.branch[10].block[10].um_I.ana[6] ;
 wire \top_I.branch[10].block[10].um_I.ana[7] ;
 wire \top_I.branch[10].block[10].um_I.clk ;
 wire \top_I.branch[10].block[10].um_I.ena ;
 wire \top_I.branch[10].block[10].um_I.iw[10] ;
 wire \top_I.branch[10].block[10].um_I.iw[11] ;
 wire \top_I.branch[10].block[10].um_I.iw[12] ;
 wire \top_I.branch[10].block[10].um_I.iw[13] ;
 wire \top_I.branch[10].block[10].um_I.iw[14] ;
 wire \top_I.branch[10].block[10].um_I.iw[15] ;
 wire \top_I.branch[10].block[10].um_I.iw[16] ;
 wire \top_I.branch[10].block[10].um_I.iw[17] ;
 wire \top_I.branch[10].block[10].um_I.iw[1] ;
 wire \top_I.branch[10].block[10].um_I.iw[2] ;
 wire \top_I.branch[10].block[10].um_I.iw[3] ;
 wire \top_I.branch[10].block[10].um_I.iw[4] ;
 wire \top_I.branch[10].block[10].um_I.iw[5] ;
 wire \top_I.branch[10].block[10].um_I.iw[6] ;
 wire \top_I.branch[10].block[10].um_I.iw[7] ;
 wire \top_I.branch[10].block[10].um_I.iw[8] ;
 wire \top_I.branch[10].block[10].um_I.iw[9] ;
 wire \top_I.branch[10].block[10].um_I.k_zero ;
 wire \top_I.branch[10].block[10].um_I.pg_vdd ;
 wire \top_I.branch[10].block[11].um_I.ana[2] ;
 wire \top_I.branch[10].block[11].um_I.ana[3] ;
 wire \top_I.branch[10].block[11].um_I.ana[4] ;
 wire \top_I.branch[10].block[11].um_I.ana[5] ;
 wire \top_I.branch[10].block[11].um_I.ana[6] ;
 wire \top_I.branch[10].block[11].um_I.ana[7] ;
 wire \top_I.branch[10].block[11].um_I.clk ;
 wire \top_I.branch[10].block[11].um_I.ena ;
 wire \top_I.branch[10].block[11].um_I.iw[10] ;
 wire \top_I.branch[10].block[11].um_I.iw[11] ;
 wire \top_I.branch[10].block[11].um_I.iw[12] ;
 wire \top_I.branch[10].block[11].um_I.iw[13] ;
 wire \top_I.branch[10].block[11].um_I.iw[14] ;
 wire \top_I.branch[10].block[11].um_I.iw[15] ;
 wire \top_I.branch[10].block[11].um_I.iw[16] ;
 wire \top_I.branch[10].block[11].um_I.iw[17] ;
 wire \top_I.branch[10].block[11].um_I.iw[1] ;
 wire \top_I.branch[10].block[11].um_I.iw[2] ;
 wire \top_I.branch[10].block[11].um_I.iw[3] ;
 wire \top_I.branch[10].block[11].um_I.iw[4] ;
 wire \top_I.branch[10].block[11].um_I.iw[5] ;
 wire \top_I.branch[10].block[11].um_I.iw[6] ;
 wire \top_I.branch[10].block[11].um_I.iw[7] ;
 wire \top_I.branch[10].block[11].um_I.iw[8] ;
 wire \top_I.branch[10].block[11].um_I.iw[9] ;
 wire \top_I.branch[10].block[11].um_I.k_zero ;
 wire \top_I.branch[10].block[11].um_I.pg_vdd ;
 wire \top_I.branch[10].block[12].um_I.ana[2] ;
 wire \top_I.branch[10].block[12].um_I.ana[3] ;
 wire \top_I.branch[10].block[12].um_I.ana[4] ;
 wire \top_I.branch[10].block[12].um_I.ana[5] ;
 wire \top_I.branch[10].block[12].um_I.ana[6] ;
 wire \top_I.branch[10].block[12].um_I.ana[7] ;
 wire \top_I.branch[10].block[12].um_I.clk ;
 wire \top_I.branch[10].block[12].um_I.ena ;
 wire \top_I.branch[10].block[12].um_I.iw[10] ;
 wire \top_I.branch[10].block[12].um_I.iw[11] ;
 wire \top_I.branch[10].block[12].um_I.iw[12] ;
 wire \top_I.branch[10].block[12].um_I.iw[13] ;
 wire \top_I.branch[10].block[12].um_I.iw[14] ;
 wire \top_I.branch[10].block[12].um_I.iw[15] ;
 wire \top_I.branch[10].block[12].um_I.iw[16] ;
 wire \top_I.branch[10].block[12].um_I.iw[17] ;
 wire \top_I.branch[10].block[12].um_I.iw[1] ;
 wire \top_I.branch[10].block[12].um_I.iw[2] ;
 wire \top_I.branch[10].block[12].um_I.iw[3] ;
 wire \top_I.branch[10].block[12].um_I.iw[4] ;
 wire \top_I.branch[10].block[12].um_I.iw[5] ;
 wire \top_I.branch[10].block[12].um_I.iw[6] ;
 wire \top_I.branch[10].block[12].um_I.iw[7] ;
 wire \top_I.branch[10].block[12].um_I.iw[8] ;
 wire \top_I.branch[10].block[12].um_I.iw[9] ;
 wire \top_I.branch[10].block[12].um_I.k_zero ;
 wire \top_I.branch[10].block[12].um_I.pg_vdd ;
 wire \top_I.branch[10].block[13].um_I.ana[2] ;
 wire \top_I.branch[10].block[13].um_I.ana[3] ;
 wire \top_I.branch[10].block[13].um_I.ana[4] ;
 wire \top_I.branch[10].block[13].um_I.ana[5] ;
 wire \top_I.branch[10].block[13].um_I.ana[6] ;
 wire \top_I.branch[10].block[13].um_I.ana[7] ;
 wire \top_I.branch[10].block[13].um_I.clk ;
 wire \top_I.branch[10].block[13].um_I.ena ;
 wire \top_I.branch[10].block[13].um_I.iw[10] ;
 wire \top_I.branch[10].block[13].um_I.iw[11] ;
 wire \top_I.branch[10].block[13].um_I.iw[12] ;
 wire \top_I.branch[10].block[13].um_I.iw[13] ;
 wire \top_I.branch[10].block[13].um_I.iw[14] ;
 wire \top_I.branch[10].block[13].um_I.iw[15] ;
 wire \top_I.branch[10].block[13].um_I.iw[16] ;
 wire \top_I.branch[10].block[13].um_I.iw[17] ;
 wire \top_I.branch[10].block[13].um_I.iw[1] ;
 wire \top_I.branch[10].block[13].um_I.iw[2] ;
 wire \top_I.branch[10].block[13].um_I.iw[3] ;
 wire \top_I.branch[10].block[13].um_I.iw[4] ;
 wire \top_I.branch[10].block[13].um_I.iw[5] ;
 wire \top_I.branch[10].block[13].um_I.iw[6] ;
 wire \top_I.branch[10].block[13].um_I.iw[7] ;
 wire \top_I.branch[10].block[13].um_I.iw[8] ;
 wire \top_I.branch[10].block[13].um_I.iw[9] ;
 wire \top_I.branch[10].block[13].um_I.k_zero ;
 wire \top_I.branch[10].block[13].um_I.pg_vdd ;
 wire \top_I.branch[10].block[14].um_I.ana[2] ;
 wire \top_I.branch[10].block[14].um_I.ana[3] ;
 wire \top_I.branch[10].block[14].um_I.ana[4] ;
 wire \top_I.branch[10].block[14].um_I.ana[5] ;
 wire \top_I.branch[10].block[14].um_I.ana[6] ;
 wire \top_I.branch[10].block[14].um_I.ana[7] ;
 wire \top_I.branch[10].block[14].um_I.clk ;
 wire \top_I.branch[10].block[14].um_I.ena ;
 wire \top_I.branch[10].block[14].um_I.iw[10] ;
 wire \top_I.branch[10].block[14].um_I.iw[11] ;
 wire \top_I.branch[10].block[14].um_I.iw[12] ;
 wire \top_I.branch[10].block[14].um_I.iw[13] ;
 wire \top_I.branch[10].block[14].um_I.iw[14] ;
 wire \top_I.branch[10].block[14].um_I.iw[15] ;
 wire \top_I.branch[10].block[14].um_I.iw[16] ;
 wire \top_I.branch[10].block[14].um_I.iw[17] ;
 wire \top_I.branch[10].block[14].um_I.iw[1] ;
 wire \top_I.branch[10].block[14].um_I.iw[2] ;
 wire \top_I.branch[10].block[14].um_I.iw[3] ;
 wire \top_I.branch[10].block[14].um_I.iw[4] ;
 wire \top_I.branch[10].block[14].um_I.iw[5] ;
 wire \top_I.branch[10].block[14].um_I.iw[6] ;
 wire \top_I.branch[10].block[14].um_I.iw[7] ;
 wire \top_I.branch[10].block[14].um_I.iw[8] ;
 wire \top_I.branch[10].block[14].um_I.iw[9] ;
 wire \top_I.branch[10].block[14].um_I.k_zero ;
 wire \top_I.branch[10].block[14].um_I.pg_vdd ;
 wire \top_I.branch[10].block[15].um_I.ana[2] ;
 wire \top_I.branch[10].block[15].um_I.ana[3] ;
 wire \top_I.branch[10].block[15].um_I.ana[4] ;
 wire \top_I.branch[10].block[15].um_I.ana[5] ;
 wire \top_I.branch[10].block[15].um_I.ana[6] ;
 wire \top_I.branch[10].block[15].um_I.ana[7] ;
 wire \top_I.branch[10].block[15].um_I.clk ;
 wire \top_I.branch[10].block[15].um_I.ena ;
 wire \top_I.branch[10].block[15].um_I.iw[10] ;
 wire \top_I.branch[10].block[15].um_I.iw[11] ;
 wire \top_I.branch[10].block[15].um_I.iw[12] ;
 wire \top_I.branch[10].block[15].um_I.iw[13] ;
 wire \top_I.branch[10].block[15].um_I.iw[14] ;
 wire \top_I.branch[10].block[15].um_I.iw[15] ;
 wire \top_I.branch[10].block[15].um_I.iw[16] ;
 wire \top_I.branch[10].block[15].um_I.iw[17] ;
 wire \top_I.branch[10].block[15].um_I.iw[1] ;
 wire \top_I.branch[10].block[15].um_I.iw[2] ;
 wire \top_I.branch[10].block[15].um_I.iw[3] ;
 wire \top_I.branch[10].block[15].um_I.iw[4] ;
 wire \top_I.branch[10].block[15].um_I.iw[5] ;
 wire \top_I.branch[10].block[15].um_I.iw[6] ;
 wire \top_I.branch[10].block[15].um_I.iw[7] ;
 wire \top_I.branch[10].block[15].um_I.iw[8] ;
 wire \top_I.branch[10].block[15].um_I.iw[9] ;
 wire \top_I.branch[10].block[15].um_I.k_zero ;
 wire \top_I.branch[10].block[15].um_I.pg_vdd ;
 wire \top_I.branch[10].block[1].um_I.ana[2] ;
 wire \top_I.branch[10].block[1].um_I.ana[3] ;
 wire \top_I.branch[10].block[1].um_I.ana[4] ;
 wire \top_I.branch[10].block[1].um_I.ana[5] ;
 wire \top_I.branch[10].block[1].um_I.ana[6] ;
 wire \top_I.branch[10].block[1].um_I.ana[7] ;
 wire \top_I.branch[10].block[1].um_I.clk ;
 wire \top_I.branch[10].block[1].um_I.ena ;
 wire \top_I.branch[10].block[1].um_I.iw[10] ;
 wire \top_I.branch[10].block[1].um_I.iw[11] ;
 wire \top_I.branch[10].block[1].um_I.iw[12] ;
 wire \top_I.branch[10].block[1].um_I.iw[13] ;
 wire \top_I.branch[10].block[1].um_I.iw[14] ;
 wire \top_I.branch[10].block[1].um_I.iw[15] ;
 wire \top_I.branch[10].block[1].um_I.iw[16] ;
 wire \top_I.branch[10].block[1].um_I.iw[17] ;
 wire \top_I.branch[10].block[1].um_I.iw[1] ;
 wire \top_I.branch[10].block[1].um_I.iw[2] ;
 wire \top_I.branch[10].block[1].um_I.iw[3] ;
 wire \top_I.branch[10].block[1].um_I.iw[4] ;
 wire \top_I.branch[10].block[1].um_I.iw[5] ;
 wire \top_I.branch[10].block[1].um_I.iw[6] ;
 wire \top_I.branch[10].block[1].um_I.iw[7] ;
 wire \top_I.branch[10].block[1].um_I.iw[8] ;
 wire \top_I.branch[10].block[1].um_I.iw[9] ;
 wire \top_I.branch[10].block[1].um_I.k_zero ;
 wire \top_I.branch[10].block[1].um_I.pg_vdd ;
 wire \top_I.branch[10].block[2].um_I.ana[2] ;
 wire \top_I.branch[10].block[2].um_I.ana[3] ;
 wire \top_I.branch[10].block[2].um_I.ana[4] ;
 wire \top_I.branch[10].block[2].um_I.ana[5] ;
 wire \top_I.branch[10].block[2].um_I.ana[6] ;
 wire \top_I.branch[10].block[2].um_I.ana[7] ;
 wire \top_I.branch[10].block[2].um_I.clk ;
 wire \top_I.branch[10].block[2].um_I.ena ;
 wire \top_I.branch[10].block[2].um_I.iw[10] ;
 wire \top_I.branch[10].block[2].um_I.iw[11] ;
 wire \top_I.branch[10].block[2].um_I.iw[12] ;
 wire \top_I.branch[10].block[2].um_I.iw[13] ;
 wire \top_I.branch[10].block[2].um_I.iw[14] ;
 wire \top_I.branch[10].block[2].um_I.iw[15] ;
 wire \top_I.branch[10].block[2].um_I.iw[16] ;
 wire \top_I.branch[10].block[2].um_I.iw[17] ;
 wire \top_I.branch[10].block[2].um_I.iw[1] ;
 wire \top_I.branch[10].block[2].um_I.iw[2] ;
 wire \top_I.branch[10].block[2].um_I.iw[3] ;
 wire \top_I.branch[10].block[2].um_I.iw[4] ;
 wire \top_I.branch[10].block[2].um_I.iw[5] ;
 wire \top_I.branch[10].block[2].um_I.iw[6] ;
 wire \top_I.branch[10].block[2].um_I.iw[7] ;
 wire \top_I.branch[10].block[2].um_I.iw[8] ;
 wire \top_I.branch[10].block[2].um_I.iw[9] ;
 wire \top_I.branch[10].block[2].um_I.k_zero ;
 wire \top_I.branch[10].block[2].um_I.pg_vdd ;
 wire \top_I.branch[10].block[3].um_I.ana[2] ;
 wire \top_I.branch[10].block[3].um_I.ana[3] ;
 wire \top_I.branch[10].block[3].um_I.ana[4] ;
 wire \top_I.branch[10].block[3].um_I.ana[5] ;
 wire \top_I.branch[10].block[3].um_I.ana[6] ;
 wire \top_I.branch[10].block[3].um_I.ana[7] ;
 wire \top_I.branch[10].block[3].um_I.clk ;
 wire \top_I.branch[10].block[3].um_I.ena ;
 wire \top_I.branch[10].block[3].um_I.iw[10] ;
 wire \top_I.branch[10].block[3].um_I.iw[11] ;
 wire \top_I.branch[10].block[3].um_I.iw[12] ;
 wire \top_I.branch[10].block[3].um_I.iw[13] ;
 wire \top_I.branch[10].block[3].um_I.iw[14] ;
 wire \top_I.branch[10].block[3].um_I.iw[15] ;
 wire \top_I.branch[10].block[3].um_I.iw[16] ;
 wire \top_I.branch[10].block[3].um_I.iw[17] ;
 wire \top_I.branch[10].block[3].um_I.iw[1] ;
 wire \top_I.branch[10].block[3].um_I.iw[2] ;
 wire \top_I.branch[10].block[3].um_I.iw[3] ;
 wire \top_I.branch[10].block[3].um_I.iw[4] ;
 wire \top_I.branch[10].block[3].um_I.iw[5] ;
 wire \top_I.branch[10].block[3].um_I.iw[6] ;
 wire \top_I.branch[10].block[3].um_I.iw[7] ;
 wire \top_I.branch[10].block[3].um_I.iw[8] ;
 wire \top_I.branch[10].block[3].um_I.iw[9] ;
 wire \top_I.branch[10].block[3].um_I.k_zero ;
 wire \top_I.branch[10].block[3].um_I.pg_vdd ;
 wire \top_I.branch[10].block[4].um_I.ana[2] ;
 wire \top_I.branch[10].block[4].um_I.ana[3] ;
 wire \top_I.branch[10].block[4].um_I.ana[4] ;
 wire \top_I.branch[10].block[4].um_I.ana[5] ;
 wire \top_I.branch[10].block[4].um_I.ana[6] ;
 wire \top_I.branch[10].block[4].um_I.ana[7] ;
 wire \top_I.branch[10].block[4].um_I.clk ;
 wire \top_I.branch[10].block[4].um_I.ena ;
 wire \top_I.branch[10].block[4].um_I.iw[10] ;
 wire \top_I.branch[10].block[4].um_I.iw[11] ;
 wire \top_I.branch[10].block[4].um_I.iw[12] ;
 wire \top_I.branch[10].block[4].um_I.iw[13] ;
 wire \top_I.branch[10].block[4].um_I.iw[14] ;
 wire \top_I.branch[10].block[4].um_I.iw[15] ;
 wire \top_I.branch[10].block[4].um_I.iw[16] ;
 wire \top_I.branch[10].block[4].um_I.iw[17] ;
 wire \top_I.branch[10].block[4].um_I.iw[1] ;
 wire \top_I.branch[10].block[4].um_I.iw[2] ;
 wire \top_I.branch[10].block[4].um_I.iw[3] ;
 wire \top_I.branch[10].block[4].um_I.iw[4] ;
 wire \top_I.branch[10].block[4].um_I.iw[5] ;
 wire \top_I.branch[10].block[4].um_I.iw[6] ;
 wire \top_I.branch[10].block[4].um_I.iw[7] ;
 wire \top_I.branch[10].block[4].um_I.iw[8] ;
 wire \top_I.branch[10].block[4].um_I.iw[9] ;
 wire \top_I.branch[10].block[4].um_I.k_zero ;
 wire \top_I.branch[10].block[4].um_I.pg_vdd ;
 wire \top_I.branch[10].block[5].um_I.ana[2] ;
 wire \top_I.branch[10].block[5].um_I.ana[3] ;
 wire \top_I.branch[10].block[5].um_I.ana[4] ;
 wire \top_I.branch[10].block[5].um_I.ana[5] ;
 wire \top_I.branch[10].block[5].um_I.ana[6] ;
 wire \top_I.branch[10].block[5].um_I.ana[7] ;
 wire \top_I.branch[10].block[5].um_I.clk ;
 wire \top_I.branch[10].block[5].um_I.ena ;
 wire \top_I.branch[10].block[5].um_I.iw[10] ;
 wire \top_I.branch[10].block[5].um_I.iw[11] ;
 wire \top_I.branch[10].block[5].um_I.iw[12] ;
 wire \top_I.branch[10].block[5].um_I.iw[13] ;
 wire \top_I.branch[10].block[5].um_I.iw[14] ;
 wire \top_I.branch[10].block[5].um_I.iw[15] ;
 wire \top_I.branch[10].block[5].um_I.iw[16] ;
 wire \top_I.branch[10].block[5].um_I.iw[17] ;
 wire \top_I.branch[10].block[5].um_I.iw[1] ;
 wire \top_I.branch[10].block[5].um_I.iw[2] ;
 wire \top_I.branch[10].block[5].um_I.iw[3] ;
 wire \top_I.branch[10].block[5].um_I.iw[4] ;
 wire \top_I.branch[10].block[5].um_I.iw[5] ;
 wire \top_I.branch[10].block[5].um_I.iw[6] ;
 wire \top_I.branch[10].block[5].um_I.iw[7] ;
 wire \top_I.branch[10].block[5].um_I.iw[8] ;
 wire \top_I.branch[10].block[5].um_I.iw[9] ;
 wire \top_I.branch[10].block[5].um_I.k_zero ;
 wire \top_I.branch[10].block[5].um_I.pg_vdd ;
 wire \top_I.branch[10].block[6].um_I.ana[2] ;
 wire \top_I.branch[10].block[6].um_I.ana[3] ;
 wire \top_I.branch[10].block[6].um_I.ana[4] ;
 wire \top_I.branch[10].block[6].um_I.ana[5] ;
 wire \top_I.branch[10].block[6].um_I.ana[6] ;
 wire \top_I.branch[10].block[6].um_I.ana[7] ;
 wire \top_I.branch[10].block[6].um_I.clk ;
 wire \top_I.branch[10].block[6].um_I.ena ;
 wire \top_I.branch[10].block[6].um_I.iw[10] ;
 wire \top_I.branch[10].block[6].um_I.iw[11] ;
 wire \top_I.branch[10].block[6].um_I.iw[12] ;
 wire \top_I.branch[10].block[6].um_I.iw[13] ;
 wire \top_I.branch[10].block[6].um_I.iw[14] ;
 wire \top_I.branch[10].block[6].um_I.iw[15] ;
 wire \top_I.branch[10].block[6].um_I.iw[16] ;
 wire \top_I.branch[10].block[6].um_I.iw[17] ;
 wire \top_I.branch[10].block[6].um_I.iw[1] ;
 wire \top_I.branch[10].block[6].um_I.iw[2] ;
 wire \top_I.branch[10].block[6].um_I.iw[3] ;
 wire \top_I.branch[10].block[6].um_I.iw[4] ;
 wire \top_I.branch[10].block[6].um_I.iw[5] ;
 wire \top_I.branch[10].block[6].um_I.iw[6] ;
 wire \top_I.branch[10].block[6].um_I.iw[7] ;
 wire \top_I.branch[10].block[6].um_I.iw[8] ;
 wire \top_I.branch[10].block[6].um_I.iw[9] ;
 wire \top_I.branch[10].block[6].um_I.k_zero ;
 wire \top_I.branch[10].block[6].um_I.pg_vdd ;
 wire \top_I.branch[10].block[7].um_I.ana[2] ;
 wire \top_I.branch[10].block[7].um_I.ana[3] ;
 wire \top_I.branch[10].block[7].um_I.ana[4] ;
 wire \top_I.branch[10].block[7].um_I.ana[5] ;
 wire \top_I.branch[10].block[7].um_I.ana[6] ;
 wire \top_I.branch[10].block[7].um_I.ana[7] ;
 wire \top_I.branch[10].block[7].um_I.clk ;
 wire \top_I.branch[10].block[7].um_I.ena ;
 wire \top_I.branch[10].block[7].um_I.iw[10] ;
 wire \top_I.branch[10].block[7].um_I.iw[11] ;
 wire \top_I.branch[10].block[7].um_I.iw[12] ;
 wire \top_I.branch[10].block[7].um_I.iw[13] ;
 wire \top_I.branch[10].block[7].um_I.iw[14] ;
 wire \top_I.branch[10].block[7].um_I.iw[15] ;
 wire \top_I.branch[10].block[7].um_I.iw[16] ;
 wire \top_I.branch[10].block[7].um_I.iw[17] ;
 wire \top_I.branch[10].block[7].um_I.iw[1] ;
 wire \top_I.branch[10].block[7].um_I.iw[2] ;
 wire \top_I.branch[10].block[7].um_I.iw[3] ;
 wire \top_I.branch[10].block[7].um_I.iw[4] ;
 wire \top_I.branch[10].block[7].um_I.iw[5] ;
 wire \top_I.branch[10].block[7].um_I.iw[6] ;
 wire \top_I.branch[10].block[7].um_I.iw[7] ;
 wire \top_I.branch[10].block[7].um_I.iw[8] ;
 wire \top_I.branch[10].block[7].um_I.iw[9] ;
 wire \top_I.branch[10].block[7].um_I.k_zero ;
 wire \top_I.branch[10].block[7].um_I.pg_vdd ;
 wire \top_I.branch[10].block[8].um_I.ana[2] ;
 wire \top_I.branch[10].block[8].um_I.ana[3] ;
 wire \top_I.branch[10].block[8].um_I.ana[4] ;
 wire \top_I.branch[10].block[8].um_I.ana[5] ;
 wire \top_I.branch[10].block[8].um_I.ana[6] ;
 wire \top_I.branch[10].block[8].um_I.ana[7] ;
 wire \top_I.branch[10].block[8].um_I.clk ;
 wire \top_I.branch[10].block[8].um_I.ena ;
 wire \top_I.branch[10].block[8].um_I.iw[10] ;
 wire \top_I.branch[10].block[8].um_I.iw[11] ;
 wire \top_I.branch[10].block[8].um_I.iw[12] ;
 wire \top_I.branch[10].block[8].um_I.iw[13] ;
 wire \top_I.branch[10].block[8].um_I.iw[14] ;
 wire \top_I.branch[10].block[8].um_I.iw[15] ;
 wire \top_I.branch[10].block[8].um_I.iw[16] ;
 wire \top_I.branch[10].block[8].um_I.iw[17] ;
 wire \top_I.branch[10].block[8].um_I.iw[1] ;
 wire \top_I.branch[10].block[8].um_I.iw[2] ;
 wire \top_I.branch[10].block[8].um_I.iw[3] ;
 wire \top_I.branch[10].block[8].um_I.iw[4] ;
 wire \top_I.branch[10].block[8].um_I.iw[5] ;
 wire \top_I.branch[10].block[8].um_I.iw[6] ;
 wire \top_I.branch[10].block[8].um_I.iw[7] ;
 wire \top_I.branch[10].block[8].um_I.iw[8] ;
 wire \top_I.branch[10].block[8].um_I.iw[9] ;
 wire \top_I.branch[10].block[8].um_I.k_zero ;
 wire \top_I.branch[10].block[8].um_I.pg_vdd ;
 wire \top_I.branch[10].block[9].um_I.ana[2] ;
 wire \top_I.branch[10].block[9].um_I.ana[3] ;
 wire \top_I.branch[10].block[9].um_I.ana[4] ;
 wire \top_I.branch[10].block[9].um_I.ana[5] ;
 wire \top_I.branch[10].block[9].um_I.ana[6] ;
 wire \top_I.branch[10].block[9].um_I.ana[7] ;
 wire \top_I.branch[10].block[9].um_I.clk ;
 wire \top_I.branch[10].block[9].um_I.ena ;
 wire \top_I.branch[10].block[9].um_I.iw[10] ;
 wire \top_I.branch[10].block[9].um_I.iw[11] ;
 wire \top_I.branch[10].block[9].um_I.iw[12] ;
 wire \top_I.branch[10].block[9].um_I.iw[13] ;
 wire \top_I.branch[10].block[9].um_I.iw[14] ;
 wire \top_I.branch[10].block[9].um_I.iw[15] ;
 wire \top_I.branch[10].block[9].um_I.iw[16] ;
 wire \top_I.branch[10].block[9].um_I.iw[17] ;
 wire \top_I.branch[10].block[9].um_I.iw[1] ;
 wire \top_I.branch[10].block[9].um_I.iw[2] ;
 wire \top_I.branch[10].block[9].um_I.iw[3] ;
 wire \top_I.branch[10].block[9].um_I.iw[4] ;
 wire \top_I.branch[10].block[9].um_I.iw[5] ;
 wire \top_I.branch[10].block[9].um_I.iw[6] ;
 wire \top_I.branch[10].block[9].um_I.iw[7] ;
 wire \top_I.branch[10].block[9].um_I.iw[8] ;
 wire \top_I.branch[10].block[9].um_I.iw[9] ;
 wire \top_I.branch[10].block[9].um_I.k_zero ;
 wire \top_I.branch[10].block[9].um_I.pg_vdd ;
 wire \top_I.branch[10].l_addr[0] ;
 wire \top_I.branch[10].l_addr[1] ;
 wire \top_I.branch[11].block[0].um_I.ana[2] ;
 wire \top_I.branch[11].block[0].um_I.ana[3] ;
 wire \top_I.branch[11].block[0].um_I.ana[4] ;
 wire \top_I.branch[11].block[0].um_I.ana[5] ;
 wire \top_I.branch[11].block[0].um_I.ana[6] ;
 wire \top_I.branch[11].block[0].um_I.ana[7] ;
 wire \top_I.branch[11].block[0].um_I.clk ;
 wire \top_I.branch[11].block[0].um_I.ena ;
 wire \top_I.branch[11].block[0].um_I.iw[10] ;
 wire \top_I.branch[11].block[0].um_I.iw[11] ;
 wire \top_I.branch[11].block[0].um_I.iw[12] ;
 wire \top_I.branch[11].block[0].um_I.iw[13] ;
 wire \top_I.branch[11].block[0].um_I.iw[14] ;
 wire \top_I.branch[11].block[0].um_I.iw[15] ;
 wire \top_I.branch[11].block[0].um_I.iw[16] ;
 wire \top_I.branch[11].block[0].um_I.iw[17] ;
 wire \top_I.branch[11].block[0].um_I.iw[1] ;
 wire \top_I.branch[11].block[0].um_I.iw[2] ;
 wire \top_I.branch[11].block[0].um_I.iw[3] ;
 wire \top_I.branch[11].block[0].um_I.iw[4] ;
 wire \top_I.branch[11].block[0].um_I.iw[5] ;
 wire \top_I.branch[11].block[0].um_I.iw[6] ;
 wire \top_I.branch[11].block[0].um_I.iw[7] ;
 wire \top_I.branch[11].block[0].um_I.iw[8] ;
 wire \top_I.branch[11].block[0].um_I.iw[9] ;
 wire \top_I.branch[11].block[0].um_I.k_zero ;
 wire \top_I.branch[11].block[0].um_I.pg_vdd ;
 wire \top_I.branch[11].block[10].um_I.ana[2] ;
 wire \top_I.branch[11].block[10].um_I.ana[3] ;
 wire \top_I.branch[11].block[10].um_I.ana[4] ;
 wire \top_I.branch[11].block[10].um_I.ana[5] ;
 wire \top_I.branch[11].block[10].um_I.ana[6] ;
 wire \top_I.branch[11].block[10].um_I.ana[7] ;
 wire \top_I.branch[11].block[10].um_I.clk ;
 wire \top_I.branch[11].block[10].um_I.ena ;
 wire \top_I.branch[11].block[10].um_I.iw[10] ;
 wire \top_I.branch[11].block[10].um_I.iw[11] ;
 wire \top_I.branch[11].block[10].um_I.iw[12] ;
 wire \top_I.branch[11].block[10].um_I.iw[13] ;
 wire \top_I.branch[11].block[10].um_I.iw[14] ;
 wire \top_I.branch[11].block[10].um_I.iw[15] ;
 wire \top_I.branch[11].block[10].um_I.iw[16] ;
 wire \top_I.branch[11].block[10].um_I.iw[17] ;
 wire \top_I.branch[11].block[10].um_I.iw[1] ;
 wire \top_I.branch[11].block[10].um_I.iw[2] ;
 wire \top_I.branch[11].block[10].um_I.iw[3] ;
 wire \top_I.branch[11].block[10].um_I.iw[4] ;
 wire \top_I.branch[11].block[10].um_I.iw[5] ;
 wire \top_I.branch[11].block[10].um_I.iw[6] ;
 wire \top_I.branch[11].block[10].um_I.iw[7] ;
 wire \top_I.branch[11].block[10].um_I.iw[8] ;
 wire \top_I.branch[11].block[10].um_I.iw[9] ;
 wire \top_I.branch[11].block[10].um_I.k_zero ;
 wire \top_I.branch[11].block[10].um_I.pg_vdd ;
 wire \top_I.branch[11].block[11].um_I.ana[2] ;
 wire \top_I.branch[11].block[11].um_I.ana[3] ;
 wire \top_I.branch[11].block[11].um_I.ana[4] ;
 wire \top_I.branch[11].block[11].um_I.ana[5] ;
 wire \top_I.branch[11].block[11].um_I.ana[6] ;
 wire \top_I.branch[11].block[11].um_I.ana[7] ;
 wire \top_I.branch[11].block[11].um_I.clk ;
 wire \top_I.branch[11].block[11].um_I.ena ;
 wire \top_I.branch[11].block[11].um_I.iw[10] ;
 wire \top_I.branch[11].block[11].um_I.iw[11] ;
 wire \top_I.branch[11].block[11].um_I.iw[12] ;
 wire \top_I.branch[11].block[11].um_I.iw[13] ;
 wire \top_I.branch[11].block[11].um_I.iw[14] ;
 wire \top_I.branch[11].block[11].um_I.iw[15] ;
 wire \top_I.branch[11].block[11].um_I.iw[16] ;
 wire \top_I.branch[11].block[11].um_I.iw[17] ;
 wire \top_I.branch[11].block[11].um_I.iw[1] ;
 wire \top_I.branch[11].block[11].um_I.iw[2] ;
 wire \top_I.branch[11].block[11].um_I.iw[3] ;
 wire \top_I.branch[11].block[11].um_I.iw[4] ;
 wire \top_I.branch[11].block[11].um_I.iw[5] ;
 wire \top_I.branch[11].block[11].um_I.iw[6] ;
 wire \top_I.branch[11].block[11].um_I.iw[7] ;
 wire \top_I.branch[11].block[11].um_I.iw[8] ;
 wire \top_I.branch[11].block[11].um_I.iw[9] ;
 wire \top_I.branch[11].block[11].um_I.k_zero ;
 wire \top_I.branch[11].block[11].um_I.pg_vdd ;
 wire \top_I.branch[11].block[12].um_I.ana[2] ;
 wire \top_I.branch[11].block[12].um_I.ana[3] ;
 wire \top_I.branch[11].block[12].um_I.ana[4] ;
 wire \top_I.branch[11].block[12].um_I.ana[5] ;
 wire \top_I.branch[11].block[12].um_I.ana[6] ;
 wire \top_I.branch[11].block[12].um_I.ana[7] ;
 wire \top_I.branch[11].block[12].um_I.clk ;
 wire \top_I.branch[11].block[12].um_I.ena ;
 wire \top_I.branch[11].block[12].um_I.iw[10] ;
 wire \top_I.branch[11].block[12].um_I.iw[11] ;
 wire \top_I.branch[11].block[12].um_I.iw[12] ;
 wire \top_I.branch[11].block[12].um_I.iw[13] ;
 wire \top_I.branch[11].block[12].um_I.iw[14] ;
 wire \top_I.branch[11].block[12].um_I.iw[15] ;
 wire \top_I.branch[11].block[12].um_I.iw[16] ;
 wire \top_I.branch[11].block[12].um_I.iw[17] ;
 wire \top_I.branch[11].block[12].um_I.iw[1] ;
 wire \top_I.branch[11].block[12].um_I.iw[2] ;
 wire \top_I.branch[11].block[12].um_I.iw[3] ;
 wire \top_I.branch[11].block[12].um_I.iw[4] ;
 wire \top_I.branch[11].block[12].um_I.iw[5] ;
 wire \top_I.branch[11].block[12].um_I.iw[6] ;
 wire \top_I.branch[11].block[12].um_I.iw[7] ;
 wire \top_I.branch[11].block[12].um_I.iw[8] ;
 wire \top_I.branch[11].block[12].um_I.iw[9] ;
 wire \top_I.branch[11].block[12].um_I.k_zero ;
 wire \top_I.branch[11].block[12].um_I.pg_vdd ;
 wire \top_I.branch[11].block[13].um_I.ana[2] ;
 wire \top_I.branch[11].block[13].um_I.ana[3] ;
 wire \top_I.branch[11].block[13].um_I.ana[4] ;
 wire \top_I.branch[11].block[13].um_I.ana[5] ;
 wire \top_I.branch[11].block[13].um_I.ana[6] ;
 wire \top_I.branch[11].block[13].um_I.ana[7] ;
 wire \top_I.branch[11].block[13].um_I.clk ;
 wire \top_I.branch[11].block[13].um_I.ena ;
 wire \top_I.branch[11].block[13].um_I.iw[10] ;
 wire \top_I.branch[11].block[13].um_I.iw[11] ;
 wire \top_I.branch[11].block[13].um_I.iw[12] ;
 wire \top_I.branch[11].block[13].um_I.iw[13] ;
 wire \top_I.branch[11].block[13].um_I.iw[14] ;
 wire \top_I.branch[11].block[13].um_I.iw[15] ;
 wire \top_I.branch[11].block[13].um_I.iw[16] ;
 wire \top_I.branch[11].block[13].um_I.iw[17] ;
 wire \top_I.branch[11].block[13].um_I.iw[1] ;
 wire \top_I.branch[11].block[13].um_I.iw[2] ;
 wire \top_I.branch[11].block[13].um_I.iw[3] ;
 wire \top_I.branch[11].block[13].um_I.iw[4] ;
 wire \top_I.branch[11].block[13].um_I.iw[5] ;
 wire \top_I.branch[11].block[13].um_I.iw[6] ;
 wire \top_I.branch[11].block[13].um_I.iw[7] ;
 wire \top_I.branch[11].block[13].um_I.iw[8] ;
 wire \top_I.branch[11].block[13].um_I.iw[9] ;
 wire \top_I.branch[11].block[13].um_I.k_zero ;
 wire \top_I.branch[11].block[13].um_I.pg_vdd ;
 wire \top_I.branch[11].block[14].um_I.ana[2] ;
 wire \top_I.branch[11].block[14].um_I.ana[3] ;
 wire \top_I.branch[11].block[14].um_I.ana[4] ;
 wire \top_I.branch[11].block[14].um_I.ana[5] ;
 wire \top_I.branch[11].block[14].um_I.ana[6] ;
 wire \top_I.branch[11].block[14].um_I.ana[7] ;
 wire \top_I.branch[11].block[14].um_I.clk ;
 wire \top_I.branch[11].block[14].um_I.ena ;
 wire \top_I.branch[11].block[14].um_I.iw[10] ;
 wire \top_I.branch[11].block[14].um_I.iw[11] ;
 wire \top_I.branch[11].block[14].um_I.iw[12] ;
 wire \top_I.branch[11].block[14].um_I.iw[13] ;
 wire \top_I.branch[11].block[14].um_I.iw[14] ;
 wire \top_I.branch[11].block[14].um_I.iw[15] ;
 wire \top_I.branch[11].block[14].um_I.iw[16] ;
 wire \top_I.branch[11].block[14].um_I.iw[17] ;
 wire \top_I.branch[11].block[14].um_I.iw[1] ;
 wire \top_I.branch[11].block[14].um_I.iw[2] ;
 wire \top_I.branch[11].block[14].um_I.iw[3] ;
 wire \top_I.branch[11].block[14].um_I.iw[4] ;
 wire \top_I.branch[11].block[14].um_I.iw[5] ;
 wire \top_I.branch[11].block[14].um_I.iw[6] ;
 wire \top_I.branch[11].block[14].um_I.iw[7] ;
 wire \top_I.branch[11].block[14].um_I.iw[8] ;
 wire \top_I.branch[11].block[14].um_I.iw[9] ;
 wire \top_I.branch[11].block[14].um_I.k_zero ;
 wire \top_I.branch[11].block[14].um_I.pg_vdd ;
 wire \top_I.branch[11].block[15].um_I.ana[2] ;
 wire \top_I.branch[11].block[15].um_I.ana[3] ;
 wire \top_I.branch[11].block[15].um_I.ana[4] ;
 wire \top_I.branch[11].block[15].um_I.ana[5] ;
 wire \top_I.branch[11].block[15].um_I.ana[6] ;
 wire \top_I.branch[11].block[15].um_I.ana[7] ;
 wire \top_I.branch[11].block[15].um_I.clk ;
 wire \top_I.branch[11].block[15].um_I.ena ;
 wire \top_I.branch[11].block[15].um_I.iw[10] ;
 wire \top_I.branch[11].block[15].um_I.iw[11] ;
 wire \top_I.branch[11].block[15].um_I.iw[12] ;
 wire \top_I.branch[11].block[15].um_I.iw[13] ;
 wire \top_I.branch[11].block[15].um_I.iw[14] ;
 wire \top_I.branch[11].block[15].um_I.iw[15] ;
 wire \top_I.branch[11].block[15].um_I.iw[16] ;
 wire \top_I.branch[11].block[15].um_I.iw[17] ;
 wire \top_I.branch[11].block[15].um_I.iw[1] ;
 wire \top_I.branch[11].block[15].um_I.iw[2] ;
 wire \top_I.branch[11].block[15].um_I.iw[3] ;
 wire \top_I.branch[11].block[15].um_I.iw[4] ;
 wire \top_I.branch[11].block[15].um_I.iw[5] ;
 wire \top_I.branch[11].block[15].um_I.iw[6] ;
 wire \top_I.branch[11].block[15].um_I.iw[7] ;
 wire \top_I.branch[11].block[15].um_I.iw[8] ;
 wire \top_I.branch[11].block[15].um_I.iw[9] ;
 wire \top_I.branch[11].block[15].um_I.k_zero ;
 wire \top_I.branch[11].block[15].um_I.pg_vdd ;
 wire \top_I.branch[11].block[1].um_I.ana[2] ;
 wire \top_I.branch[11].block[1].um_I.ana[3] ;
 wire \top_I.branch[11].block[1].um_I.ana[4] ;
 wire \top_I.branch[11].block[1].um_I.ana[5] ;
 wire \top_I.branch[11].block[1].um_I.ana[6] ;
 wire \top_I.branch[11].block[1].um_I.ana[7] ;
 wire \top_I.branch[11].block[1].um_I.clk ;
 wire \top_I.branch[11].block[1].um_I.ena ;
 wire \top_I.branch[11].block[1].um_I.iw[10] ;
 wire \top_I.branch[11].block[1].um_I.iw[11] ;
 wire \top_I.branch[11].block[1].um_I.iw[12] ;
 wire \top_I.branch[11].block[1].um_I.iw[13] ;
 wire \top_I.branch[11].block[1].um_I.iw[14] ;
 wire \top_I.branch[11].block[1].um_I.iw[15] ;
 wire \top_I.branch[11].block[1].um_I.iw[16] ;
 wire \top_I.branch[11].block[1].um_I.iw[17] ;
 wire \top_I.branch[11].block[1].um_I.iw[1] ;
 wire \top_I.branch[11].block[1].um_I.iw[2] ;
 wire \top_I.branch[11].block[1].um_I.iw[3] ;
 wire \top_I.branch[11].block[1].um_I.iw[4] ;
 wire \top_I.branch[11].block[1].um_I.iw[5] ;
 wire \top_I.branch[11].block[1].um_I.iw[6] ;
 wire \top_I.branch[11].block[1].um_I.iw[7] ;
 wire \top_I.branch[11].block[1].um_I.iw[8] ;
 wire \top_I.branch[11].block[1].um_I.iw[9] ;
 wire \top_I.branch[11].block[1].um_I.k_zero ;
 wire \top_I.branch[11].block[1].um_I.pg_vdd ;
 wire \top_I.branch[11].block[2].um_I.ana[2] ;
 wire \top_I.branch[11].block[2].um_I.ana[3] ;
 wire \top_I.branch[11].block[2].um_I.ana[4] ;
 wire \top_I.branch[11].block[2].um_I.ana[5] ;
 wire \top_I.branch[11].block[2].um_I.ana[6] ;
 wire \top_I.branch[11].block[2].um_I.ana[7] ;
 wire \top_I.branch[11].block[2].um_I.clk ;
 wire \top_I.branch[11].block[2].um_I.ena ;
 wire \top_I.branch[11].block[2].um_I.iw[10] ;
 wire \top_I.branch[11].block[2].um_I.iw[11] ;
 wire \top_I.branch[11].block[2].um_I.iw[12] ;
 wire \top_I.branch[11].block[2].um_I.iw[13] ;
 wire \top_I.branch[11].block[2].um_I.iw[14] ;
 wire \top_I.branch[11].block[2].um_I.iw[15] ;
 wire \top_I.branch[11].block[2].um_I.iw[16] ;
 wire \top_I.branch[11].block[2].um_I.iw[17] ;
 wire \top_I.branch[11].block[2].um_I.iw[1] ;
 wire \top_I.branch[11].block[2].um_I.iw[2] ;
 wire \top_I.branch[11].block[2].um_I.iw[3] ;
 wire \top_I.branch[11].block[2].um_I.iw[4] ;
 wire \top_I.branch[11].block[2].um_I.iw[5] ;
 wire \top_I.branch[11].block[2].um_I.iw[6] ;
 wire \top_I.branch[11].block[2].um_I.iw[7] ;
 wire \top_I.branch[11].block[2].um_I.iw[8] ;
 wire \top_I.branch[11].block[2].um_I.iw[9] ;
 wire \top_I.branch[11].block[2].um_I.k_zero ;
 wire \top_I.branch[11].block[2].um_I.pg_vdd ;
 wire \top_I.branch[11].block[3].um_I.ana[2] ;
 wire \top_I.branch[11].block[3].um_I.ana[3] ;
 wire \top_I.branch[11].block[3].um_I.ana[4] ;
 wire \top_I.branch[11].block[3].um_I.ana[5] ;
 wire \top_I.branch[11].block[3].um_I.ana[6] ;
 wire \top_I.branch[11].block[3].um_I.ana[7] ;
 wire \top_I.branch[11].block[3].um_I.clk ;
 wire \top_I.branch[11].block[3].um_I.ena ;
 wire \top_I.branch[11].block[3].um_I.iw[10] ;
 wire \top_I.branch[11].block[3].um_I.iw[11] ;
 wire \top_I.branch[11].block[3].um_I.iw[12] ;
 wire \top_I.branch[11].block[3].um_I.iw[13] ;
 wire \top_I.branch[11].block[3].um_I.iw[14] ;
 wire \top_I.branch[11].block[3].um_I.iw[15] ;
 wire \top_I.branch[11].block[3].um_I.iw[16] ;
 wire \top_I.branch[11].block[3].um_I.iw[17] ;
 wire \top_I.branch[11].block[3].um_I.iw[1] ;
 wire \top_I.branch[11].block[3].um_I.iw[2] ;
 wire \top_I.branch[11].block[3].um_I.iw[3] ;
 wire \top_I.branch[11].block[3].um_I.iw[4] ;
 wire \top_I.branch[11].block[3].um_I.iw[5] ;
 wire \top_I.branch[11].block[3].um_I.iw[6] ;
 wire \top_I.branch[11].block[3].um_I.iw[7] ;
 wire \top_I.branch[11].block[3].um_I.iw[8] ;
 wire \top_I.branch[11].block[3].um_I.iw[9] ;
 wire \top_I.branch[11].block[3].um_I.k_zero ;
 wire \top_I.branch[11].block[3].um_I.pg_vdd ;
 wire \top_I.branch[11].block[4].um_I.ana[2] ;
 wire \top_I.branch[11].block[4].um_I.ana[3] ;
 wire \top_I.branch[11].block[4].um_I.ana[4] ;
 wire \top_I.branch[11].block[4].um_I.ana[5] ;
 wire \top_I.branch[11].block[4].um_I.ana[6] ;
 wire \top_I.branch[11].block[4].um_I.ana[7] ;
 wire \top_I.branch[11].block[4].um_I.clk ;
 wire \top_I.branch[11].block[4].um_I.ena ;
 wire \top_I.branch[11].block[4].um_I.iw[10] ;
 wire \top_I.branch[11].block[4].um_I.iw[11] ;
 wire \top_I.branch[11].block[4].um_I.iw[12] ;
 wire \top_I.branch[11].block[4].um_I.iw[13] ;
 wire \top_I.branch[11].block[4].um_I.iw[14] ;
 wire \top_I.branch[11].block[4].um_I.iw[15] ;
 wire \top_I.branch[11].block[4].um_I.iw[16] ;
 wire \top_I.branch[11].block[4].um_I.iw[17] ;
 wire \top_I.branch[11].block[4].um_I.iw[1] ;
 wire \top_I.branch[11].block[4].um_I.iw[2] ;
 wire \top_I.branch[11].block[4].um_I.iw[3] ;
 wire \top_I.branch[11].block[4].um_I.iw[4] ;
 wire \top_I.branch[11].block[4].um_I.iw[5] ;
 wire \top_I.branch[11].block[4].um_I.iw[6] ;
 wire \top_I.branch[11].block[4].um_I.iw[7] ;
 wire \top_I.branch[11].block[4].um_I.iw[8] ;
 wire \top_I.branch[11].block[4].um_I.iw[9] ;
 wire \top_I.branch[11].block[4].um_I.k_zero ;
 wire \top_I.branch[11].block[4].um_I.pg_vdd ;
 wire \top_I.branch[11].block[5].um_I.ana[2] ;
 wire \top_I.branch[11].block[5].um_I.ana[3] ;
 wire \top_I.branch[11].block[5].um_I.ana[4] ;
 wire \top_I.branch[11].block[5].um_I.ana[5] ;
 wire \top_I.branch[11].block[5].um_I.ana[6] ;
 wire \top_I.branch[11].block[5].um_I.ana[7] ;
 wire \top_I.branch[11].block[5].um_I.clk ;
 wire \top_I.branch[11].block[5].um_I.ena ;
 wire \top_I.branch[11].block[5].um_I.iw[10] ;
 wire \top_I.branch[11].block[5].um_I.iw[11] ;
 wire \top_I.branch[11].block[5].um_I.iw[12] ;
 wire \top_I.branch[11].block[5].um_I.iw[13] ;
 wire \top_I.branch[11].block[5].um_I.iw[14] ;
 wire \top_I.branch[11].block[5].um_I.iw[15] ;
 wire \top_I.branch[11].block[5].um_I.iw[16] ;
 wire \top_I.branch[11].block[5].um_I.iw[17] ;
 wire \top_I.branch[11].block[5].um_I.iw[1] ;
 wire \top_I.branch[11].block[5].um_I.iw[2] ;
 wire \top_I.branch[11].block[5].um_I.iw[3] ;
 wire \top_I.branch[11].block[5].um_I.iw[4] ;
 wire \top_I.branch[11].block[5].um_I.iw[5] ;
 wire \top_I.branch[11].block[5].um_I.iw[6] ;
 wire \top_I.branch[11].block[5].um_I.iw[7] ;
 wire \top_I.branch[11].block[5].um_I.iw[8] ;
 wire \top_I.branch[11].block[5].um_I.iw[9] ;
 wire \top_I.branch[11].block[5].um_I.k_zero ;
 wire \top_I.branch[11].block[5].um_I.pg_vdd ;
 wire \top_I.branch[11].block[6].um_I.ana[2] ;
 wire \top_I.branch[11].block[6].um_I.ana[3] ;
 wire \top_I.branch[11].block[6].um_I.ana[4] ;
 wire \top_I.branch[11].block[6].um_I.ana[5] ;
 wire \top_I.branch[11].block[6].um_I.ana[6] ;
 wire \top_I.branch[11].block[6].um_I.ana[7] ;
 wire \top_I.branch[11].block[6].um_I.clk ;
 wire \top_I.branch[11].block[6].um_I.ena ;
 wire \top_I.branch[11].block[6].um_I.iw[10] ;
 wire \top_I.branch[11].block[6].um_I.iw[11] ;
 wire \top_I.branch[11].block[6].um_I.iw[12] ;
 wire \top_I.branch[11].block[6].um_I.iw[13] ;
 wire \top_I.branch[11].block[6].um_I.iw[14] ;
 wire \top_I.branch[11].block[6].um_I.iw[15] ;
 wire \top_I.branch[11].block[6].um_I.iw[16] ;
 wire \top_I.branch[11].block[6].um_I.iw[17] ;
 wire \top_I.branch[11].block[6].um_I.iw[1] ;
 wire \top_I.branch[11].block[6].um_I.iw[2] ;
 wire \top_I.branch[11].block[6].um_I.iw[3] ;
 wire \top_I.branch[11].block[6].um_I.iw[4] ;
 wire \top_I.branch[11].block[6].um_I.iw[5] ;
 wire \top_I.branch[11].block[6].um_I.iw[6] ;
 wire \top_I.branch[11].block[6].um_I.iw[7] ;
 wire \top_I.branch[11].block[6].um_I.iw[8] ;
 wire \top_I.branch[11].block[6].um_I.iw[9] ;
 wire \top_I.branch[11].block[6].um_I.k_zero ;
 wire \top_I.branch[11].block[6].um_I.pg_vdd ;
 wire \top_I.branch[11].block[7].um_I.ana[2] ;
 wire \top_I.branch[11].block[7].um_I.ana[3] ;
 wire \top_I.branch[11].block[7].um_I.ana[4] ;
 wire \top_I.branch[11].block[7].um_I.ana[5] ;
 wire \top_I.branch[11].block[7].um_I.ana[6] ;
 wire \top_I.branch[11].block[7].um_I.ana[7] ;
 wire \top_I.branch[11].block[7].um_I.clk ;
 wire \top_I.branch[11].block[7].um_I.ena ;
 wire \top_I.branch[11].block[7].um_I.iw[10] ;
 wire \top_I.branch[11].block[7].um_I.iw[11] ;
 wire \top_I.branch[11].block[7].um_I.iw[12] ;
 wire \top_I.branch[11].block[7].um_I.iw[13] ;
 wire \top_I.branch[11].block[7].um_I.iw[14] ;
 wire \top_I.branch[11].block[7].um_I.iw[15] ;
 wire \top_I.branch[11].block[7].um_I.iw[16] ;
 wire \top_I.branch[11].block[7].um_I.iw[17] ;
 wire \top_I.branch[11].block[7].um_I.iw[1] ;
 wire \top_I.branch[11].block[7].um_I.iw[2] ;
 wire \top_I.branch[11].block[7].um_I.iw[3] ;
 wire \top_I.branch[11].block[7].um_I.iw[4] ;
 wire \top_I.branch[11].block[7].um_I.iw[5] ;
 wire \top_I.branch[11].block[7].um_I.iw[6] ;
 wire \top_I.branch[11].block[7].um_I.iw[7] ;
 wire \top_I.branch[11].block[7].um_I.iw[8] ;
 wire \top_I.branch[11].block[7].um_I.iw[9] ;
 wire \top_I.branch[11].block[7].um_I.k_zero ;
 wire \top_I.branch[11].block[7].um_I.pg_vdd ;
 wire \top_I.branch[11].block[8].um_I.ana[2] ;
 wire \top_I.branch[11].block[8].um_I.ana[3] ;
 wire \top_I.branch[11].block[8].um_I.ana[4] ;
 wire \top_I.branch[11].block[8].um_I.ana[5] ;
 wire \top_I.branch[11].block[8].um_I.ana[6] ;
 wire \top_I.branch[11].block[8].um_I.ana[7] ;
 wire \top_I.branch[11].block[8].um_I.clk ;
 wire \top_I.branch[11].block[8].um_I.ena ;
 wire \top_I.branch[11].block[8].um_I.iw[10] ;
 wire \top_I.branch[11].block[8].um_I.iw[11] ;
 wire \top_I.branch[11].block[8].um_I.iw[12] ;
 wire \top_I.branch[11].block[8].um_I.iw[13] ;
 wire \top_I.branch[11].block[8].um_I.iw[14] ;
 wire \top_I.branch[11].block[8].um_I.iw[15] ;
 wire \top_I.branch[11].block[8].um_I.iw[16] ;
 wire \top_I.branch[11].block[8].um_I.iw[17] ;
 wire \top_I.branch[11].block[8].um_I.iw[1] ;
 wire \top_I.branch[11].block[8].um_I.iw[2] ;
 wire \top_I.branch[11].block[8].um_I.iw[3] ;
 wire \top_I.branch[11].block[8].um_I.iw[4] ;
 wire \top_I.branch[11].block[8].um_I.iw[5] ;
 wire \top_I.branch[11].block[8].um_I.iw[6] ;
 wire \top_I.branch[11].block[8].um_I.iw[7] ;
 wire \top_I.branch[11].block[8].um_I.iw[8] ;
 wire \top_I.branch[11].block[8].um_I.iw[9] ;
 wire \top_I.branch[11].block[8].um_I.k_zero ;
 wire \top_I.branch[11].block[8].um_I.pg_vdd ;
 wire \top_I.branch[11].block[9].um_I.ana[2] ;
 wire \top_I.branch[11].block[9].um_I.ana[3] ;
 wire \top_I.branch[11].block[9].um_I.ana[4] ;
 wire \top_I.branch[11].block[9].um_I.ana[5] ;
 wire \top_I.branch[11].block[9].um_I.ana[6] ;
 wire \top_I.branch[11].block[9].um_I.ana[7] ;
 wire \top_I.branch[11].block[9].um_I.clk ;
 wire \top_I.branch[11].block[9].um_I.ena ;
 wire \top_I.branch[11].block[9].um_I.iw[10] ;
 wire \top_I.branch[11].block[9].um_I.iw[11] ;
 wire \top_I.branch[11].block[9].um_I.iw[12] ;
 wire \top_I.branch[11].block[9].um_I.iw[13] ;
 wire \top_I.branch[11].block[9].um_I.iw[14] ;
 wire \top_I.branch[11].block[9].um_I.iw[15] ;
 wire \top_I.branch[11].block[9].um_I.iw[16] ;
 wire \top_I.branch[11].block[9].um_I.iw[17] ;
 wire \top_I.branch[11].block[9].um_I.iw[1] ;
 wire \top_I.branch[11].block[9].um_I.iw[2] ;
 wire \top_I.branch[11].block[9].um_I.iw[3] ;
 wire \top_I.branch[11].block[9].um_I.iw[4] ;
 wire \top_I.branch[11].block[9].um_I.iw[5] ;
 wire \top_I.branch[11].block[9].um_I.iw[6] ;
 wire \top_I.branch[11].block[9].um_I.iw[7] ;
 wire \top_I.branch[11].block[9].um_I.iw[8] ;
 wire \top_I.branch[11].block[9].um_I.iw[9] ;
 wire \top_I.branch[11].block[9].um_I.k_zero ;
 wire \top_I.branch[11].block[9].um_I.pg_vdd ;
 wire \top_I.branch[11].l_addr[0] ;
 wire \top_I.branch[11].l_addr[1] ;
 wire \top_I.branch[11].l_spine_iw[0] ;
 wire \top_I.branch[11].l_spine_iw[10] ;
 wire \top_I.branch[11].l_spine_iw[11] ;
 wire \top_I.branch[11].l_spine_iw[12] ;
 wire \top_I.branch[11].l_spine_iw[13] ;
 wire \top_I.branch[11].l_spine_iw[14] ;
 wire \top_I.branch[11].l_spine_iw[15] ;
 wire \top_I.branch[11].l_spine_iw[16] ;
 wire \top_I.branch[11].l_spine_iw[17] ;
 wire \top_I.branch[11].l_spine_iw[18] ;
 wire \top_I.branch[11].l_spine_iw[19] ;
 wire \top_I.branch[11].l_spine_iw[1] ;
 wire \top_I.branch[11].l_spine_iw[20] ;
 wire \top_I.branch[11].l_spine_iw[21] ;
 wire \top_I.branch[11].l_spine_iw[22] ;
 wire \top_I.branch[11].l_spine_iw[23] ;
 wire \top_I.branch[11].l_spine_iw[24] ;
 wire \top_I.branch[11].l_spine_iw[25] ;
 wire \top_I.branch[11].l_spine_iw[26] ;
 wire \top_I.branch[11].l_spine_iw[27] ;
 wire \top_I.branch[11].l_spine_iw[28] ;
 wire \top_I.branch[11].l_spine_iw[29] ;
 wire \top_I.branch[11].l_spine_iw[2] ;
 wire \top_I.branch[11].l_spine_iw[3] ;
 wire \top_I.branch[11].l_spine_iw[4] ;
 wire \top_I.branch[11].l_spine_iw[5] ;
 wire \top_I.branch[11].l_spine_iw[6] ;
 wire \top_I.branch[11].l_spine_iw[7] ;
 wire \top_I.branch[11].l_spine_iw[8] ;
 wire \top_I.branch[11].l_spine_iw[9] ;
 wire \top_I.branch[11].l_spine_ow[0] ;
 wire \top_I.branch[11].l_spine_ow[10] ;
 wire \top_I.branch[11].l_spine_ow[11] ;
 wire \top_I.branch[11].l_spine_ow[12] ;
 wire \top_I.branch[11].l_spine_ow[13] ;
 wire \top_I.branch[11].l_spine_ow[14] ;
 wire \top_I.branch[11].l_spine_ow[15] ;
 wire \top_I.branch[11].l_spine_ow[16] ;
 wire \top_I.branch[11].l_spine_ow[17] ;
 wire \top_I.branch[11].l_spine_ow[18] ;
 wire \top_I.branch[11].l_spine_ow[19] ;
 wire \top_I.branch[11].l_spine_ow[1] ;
 wire \top_I.branch[11].l_spine_ow[20] ;
 wire \top_I.branch[11].l_spine_ow[21] ;
 wire \top_I.branch[11].l_spine_ow[22] ;
 wire \top_I.branch[11].l_spine_ow[23] ;
 wire \top_I.branch[11].l_spine_ow[24] ;
 wire \top_I.branch[11].l_spine_ow[25] ;
 wire \top_I.branch[11].l_spine_ow[2] ;
 wire \top_I.branch[11].l_spine_ow[3] ;
 wire \top_I.branch[11].l_spine_ow[4] ;
 wire \top_I.branch[11].l_spine_ow[5] ;
 wire \top_I.branch[11].l_spine_ow[6] ;
 wire \top_I.branch[11].l_spine_ow[7] ;
 wire \top_I.branch[11].l_spine_ow[8] ;
 wire \top_I.branch[11].l_spine_ow[9] ;
 wire \top_I.branch[12].block[0].um_I.ana[2] ;
 wire \top_I.branch[12].block[0].um_I.ana[3] ;
 wire \top_I.branch[12].block[0].um_I.ana[4] ;
 wire \top_I.branch[12].block[0].um_I.ana[5] ;
 wire \top_I.branch[12].block[0].um_I.ana[6] ;
 wire \top_I.branch[12].block[0].um_I.ana[7] ;
 wire \top_I.branch[12].block[0].um_I.clk ;
 wire \top_I.branch[12].block[0].um_I.ena ;
 wire \top_I.branch[12].block[0].um_I.iw[10] ;
 wire \top_I.branch[12].block[0].um_I.iw[11] ;
 wire \top_I.branch[12].block[0].um_I.iw[12] ;
 wire \top_I.branch[12].block[0].um_I.iw[13] ;
 wire \top_I.branch[12].block[0].um_I.iw[14] ;
 wire \top_I.branch[12].block[0].um_I.iw[15] ;
 wire \top_I.branch[12].block[0].um_I.iw[16] ;
 wire \top_I.branch[12].block[0].um_I.iw[17] ;
 wire \top_I.branch[12].block[0].um_I.iw[1] ;
 wire \top_I.branch[12].block[0].um_I.iw[2] ;
 wire \top_I.branch[12].block[0].um_I.iw[3] ;
 wire \top_I.branch[12].block[0].um_I.iw[4] ;
 wire \top_I.branch[12].block[0].um_I.iw[5] ;
 wire \top_I.branch[12].block[0].um_I.iw[6] ;
 wire \top_I.branch[12].block[0].um_I.iw[7] ;
 wire \top_I.branch[12].block[0].um_I.iw[8] ;
 wire \top_I.branch[12].block[0].um_I.iw[9] ;
 wire \top_I.branch[12].block[0].um_I.k_zero ;
 wire \top_I.branch[12].block[0].um_I.pg_vdd ;
 wire \top_I.branch[12].block[10].um_I.ana[2] ;
 wire \top_I.branch[12].block[10].um_I.ana[3] ;
 wire \top_I.branch[12].block[10].um_I.ana[4] ;
 wire \top_I.branch[12].block[10].um_I.ana[5] ;
 wire \top_I.branch[12].block[10].um_I.ana[6] ;
 wire \top_I.branch[12].block[10].um_I.ana[7] ;
 wire \top_I.branch[12].block[10].um_I.clk ;
 wire \top_I.branch[12].block[10].um_I.ena ;
 wire \top_I.branch[12].block[10].um_I.iw[10] ;
 wire \top_I.branch[12].block[10].um_I.iw[11] ;
 wire \top_I.branch[12].block[10].um_I.iw[12] ;
 wire \top_I.branch[12].block[10].um_I.iw[13] ;
 wire \top_I.branch[12].block[10].um_I.iw[14] ;
 wire \top_I.branch[12].block[10].um_I.iw[15] ;
 wire \top_I.branch[12].block[10].um_I.iw[16] ;
 wire \top_I.branch[12].block[10].um_I.iw[17] ;
 wire \top_I.branch[12].block[10].um_I.iw[1] ;
 wire \top_I.branch[12].block[10].um_I.iw[2] ;
 wire \top_I.branch[12].block[10].um_I.iw[3] ;
 wire \top_I.branch[12].block[10].um_I.iw[4] ;
 wire \top_I.branch[12].block[10].um_I.iw[5] ;
 wire \top_I.branch[12].block[10].um_I.iw[6] ;
 wire \top_I.branch[12].block[10].um_I.iw[7] ;
 wire \top_I.branch[12].block[10].um_I.iw[8] ;
 wire \top_I.branch[12].block[10].um_I.iw[9] ;
 wire \top_I.branch[12].block[10].um_I.k_zero ;
 wire \top_I.branch[12].block[10].um_I.pg_vdd ;
 wire \top_I.branch[12].block[11].um_I.ana[2] ;
 wire \top_I.branch[12].block[11].um_I.ana[3] ;
 wire \top_I.branch[12].block[11].um_I.ana[4] ;
 wire \top_I.branch[12].block[11].um_I.ana[5] ;
 wire \top_I.branch[12].block[11].um_I.ana[6] ;
 wire \top_I.branch[12].block[11].um_I.ana[7] ;
 wire \top_I.branch[12].block[11].um_I.clk ;
 wire \top_I.branch[12].block[11].um_I.ena ;
 wire \top_I.branch[12].block[11].um_I.iw[10] ;
 wire \top_I.branch[12].block[11].um_I.iw[11] ;
 wire \top_I.branch[12].block[11].um_I.iw[12] ;
 wire \top_I.branch[12].block[11].um_I.iw[13] ;
 wire \top_I.branch[12].block[11].um_I.iw[14] ;
 wire \top_I.branch[12].block[11].um_I.iw[15] ;
 wire \top_I.branch[12].block[11].um_I.iw[16] ;
 wire \top_I.branch[12].block[11].um_I.iw[17] ;
 wire \top_I.branch[12].block[11].um_I.iw[1] ;
 wire \top_I.branch[12].block[11].um_I.iw[2] ;
 wire \top_I.branch[12].block[11].um_I.iw[3] ;
 wire \top_I.branch[12].block[11].um_I.iw[4] ;
 wire \top_I.branch[12].block[11].um_I.iw[5] ;
 wire \top_I.branch[12].block[11].um_I.iw[6] ;
 wire \top_I.branch[12].block[11].um_I.iw[7] ;
 wire \top_I.branch[12].block[11].um_I.iw[8] ;
 wire \top_I.branch[12].block[11].um_I.iw[9] ;
 wire \top_I.branch[12].block[11].um_I.k_zero ;
 wire \top_I.branch[12].block[11].um_I.pg_vdd ;
 wire \top_I.branch[12].block[12].um_I.ana[2] ;
 wire \top_I.branch[12].block[12].um_I.ana[3] ;
 wire \top_I.branch[12].block[12].um_I.ana[4] ;
 wire \top_I.branch[12].block[12].um_I.ana[5] ;
 wire \top_I.branch[12].block[12].um_I.ana[6] ;
 wire \top_I.branch[12].block[12].um_I.ana[7] ;
 wire \top_I.branch[12].block[12].um_I.clk ;
 wire \top_I.branch[12].block[12].um_I.ena ;
 wire \top_I.branch[12].block[12].um_I.iw[10] ;
 wire \top_I.branch[12].block[12].um_I.iw[11] ;
 wire \top_I.branch[12].block[12].um_I.iw[12] ;
 wire \top_I.branch[12].block[12].um_I.iw[13] ;
 wire \top_I.branch[12].block[12].um_I.iw[14] ;
 wire \top_I.branch[12].block[12].um_I.iw[15] ;
 wire \top_I.branch[12].block[12].um_I.iw[16] ;
 wire \top_I.branch[12].block[12].um_I.iw[17] ;
 wire \top_I.branch[12].block[12].um_I.iw[1] ;
 wire \top_I.branch[12].block[12].um_I.iw[2] ;
 wire \top_I.branch[12].block[12].um_I.iw[3] ;
 wire \top_I.branch[12].block[12].um_I.iw[4] ;
 wire \top_I.branch[12].block[12].um_I.iw[5] ;
 wire \top_I.branch[12].block[12].um_I.iw[6] ;
 wire \top_I.branch[12].block[12].um_I.iw[7] ;
 wire \top_I.branch[12].block[12].um_I.iw[8] ;
 wire \top_I.branch[12].block[12].um_I.iw[9] ;
 wire \top_I.branch[12].block[12].um_I.k_zero ;
 wire \top_I.branch[12].block[12].um_I.pg_vdd ;
 wire \top_I.branch[12].block[13].um_I.ana[2] ;
 wire \top_I.branch[12].block[13].um_I.ana[3] ;
 wire \top_I.branch[12].block[13].um_I.ana[4] ;
 wire \top_I.branch[12].block[13].um_I.ana[5] ;
 wire \top_I.branch[12].block[13].um_I.ana[6] ;
 wire \top_I.branch[12].block[13].um_I.ana[7] ;
 wire \top_I.branch[12].block[13].um_I.clk ;
 wire \top_I.branch[12].block[13].um_I.ena ;
 wire \top_I.branch[12].block[13].um_I.iw[10] ;
 wire \top_I.branch[12].block[13].um_I.iw[11] ;
 wire \top_I.branch[12].block[13].um_I.iw[12] ;
 wire \top_I.branch[12].block[13].um_I.iw[13] ;
 wire \top_I.branch[12].block[13].um_I.iw[14] ;
 wire \top_I.branch[12].block[13].um_I.iw[15] ;
 wire \top_I.branch[12].block[13].um_I.iw[16] ;
 wire \top_I.branch[12].block[13].um_I.iw[17] ;
 wire \top_I.branch[12].block[13].um_I.iw[1] ;
 wire \top_I.branch[12].block[13].um_I.iw[2] ;
 wire \top_I.branch[12].block[13].um_I.iw[3] ;
 wire \top_I.branch[12].block[13].um_I.iw[4] ;
 wire \top_I.branch[12].block[13].um_I.iw[5] ;
 wire \top_I.branch[12].block[13].um_I.iw[6] ;
 wire \top_I.branch[12].block[13].um_I.iw[7] ;
 wire \top_I.branch[12].block[13].um_I.iw[8] ;
 wire \top_I.branch[12].block[13].um_I.iw[9] ;
 wire \top_I.branch[12].block[13].um_I.k_zero ;
 wire \top_I.branch[12].block[13].um_I.pg_vdd ;
 wire \top_I.branch[12].block[14].um_I.ana[2] ;
 wire \top_I.branch[12].block[14].um_I.ana[3] ;
 wire \top_I.branch[12].block[14].um_I.ana[4] ;
 wire \top_I.branch[12].block[14].um_I.ana[5] ;
 wire \top_I.branch[12].block[14].um_I.ana[6] ;
 wire \top_I.branch[12].block[14].um_I.ana[7] ;
 wire \top_I.branch[12].block[14].um_I.clk ;
 wire \top_I.branch[12].block[14].um_I.ena ;
 wire \top_I.branch[12].block[14].um_I.iw[10] ;
 wire \top_I.branch[12].block[14].um_I.iw[11] ;
 wire \top_I.branch[12].block[14].um_I.iw[12] ;
 wire \top_I.branch[12].block[14].um_I.iw[13] ;
 wire \top_I.branch[12].block[14].um_I.iw[14] ;
 wire \top_I.branch[12].block[14].um_I.iw[15] ;
 wire \top_I.branch[12].block[14].um_I.iw[16] ;
 wire \top_I.branch[12].block[14].um_I.iw[17] ;
 wire \top_I.branch[12].block[14].um_I.iw[1] ;
 wire \top_I.branch[12].block[14].um_I.iw[2] ;
 wire \top_I.branch[12].block[14].um_I.iw[3] ;
 wire \top_I.branch[12].block[14].um_I.iw[4] ;
 wire \top_I.branch[12].block[14].um_I.iw[5] ;
 wire \top_I.branch[12].block[14].um_I.iw[6] ;
 wire \top_I.branch[12].block[14].um_I.iw[7] ;
 wire \top_I.branch[12].block[14].um_I.iw[8] ;
 wire \top_I.branch[12].block[14].um_I.iw[9] ;
 wire \top_I.branch[12].block[14].um_I.k_zero ;
 wire \top_I.branch[12].block[14].um_I.pg_vdd ;
 wire \top_I.branch[12].block[15].um_I.ana[2] ;
 wire \top_I.branch[12].block[15].um_I.ana[3] ;
 wire \top_I.branch[12].block[15].um_I.ana[4] ;
 wire \top_I.branch[12].block[15].um_I.ana[5] ;
 wire \top_I.branch[12].block[15].um_I.ana[6] ;
 wire \top_I.branch[12].block[15].um_I.ana[7] ;
 wire \top_I.branch[12].block[15].um_I.clk ;
 wire \top_I.branch[12].block[15].um_I.ena ;
 wire \top_I.branch[12].block[15].um_I.iw[10] ;
 wire \top_I.branch[12].block[15].um_I.iw[11] ;
 wire \top_I.branch[12].block[15].um_I.iw[12] ;
 wire \top_I.branch[12].block[15].um_I.iw[13] ;
 wire \top_I.branch[12].block[15].um_I.iw[14] ;
 wire \top_I.branch[12].block[15].um_I.iw[15] ;
 wire \top_I.branch[12].block[15].um_I.iw[16] ;
 wire \top_I.branch[12].block[15].um_I.iw[17] ;
 wire \top_I.branch[12].block[15].um_I.iw[1] ;
 wire \top_I.branch[12].block[15].um_I.iw[2] ;
 wire \top_I.branch[12].block[15].um_I.iw[3] ;
 wire \top_I.branch[12].block[15].um_I.iw[4] ;
 wire \top_I.branch[12].block[15].um_I.iw[5] ;
 wire \top_I.branch[12].block[15].um_I.iw[6] ;
 wire \top_I.branch[12].block[15].um_I.iw[7] ;
 wire \top_I.branch[12].block[15].um_I.iw[8] ;
 wire \top_I.branch[12].block[15].um_I.iw[9] ;
 wire \top_I.branch[12].block[15].um_I.k_zero ;
 wire \top_I.branch[12].block[15].um_I.pg_vdd ;
 wire \top_I.branch[12].block[1].um_I.ana[2] ;
 wire \top_I.branch[12].block[1].um_I.ana[3] ;
 wire \top_I.branch[12].block[1].um_I.ana[4] ;
 wire \top_I.branch[12].block[1].um_I.ana[5] ;
 wire \top_I.branch[12].block[1].um_I.ana[6] ;
 wire \top_I.branch[12].block[1].um_I.ana[7] ;
 wire \top_I.branch[12].block[1].um_I.clk ;
 wire \top_I.branch[12].block[1].um_I.ena ;
 wire \top_I.branch[12].block[1].um_I.iw[10] ;
 wire \top_I.branch[12].block[1].um_I.iw[11] ;
 wire \top_I.branch[12].block[1].um_I.iw[12] ;
 wire \top_I.branch[12].block[1].um_I.iw[13] ;
 wire \top_I.branch[12].block[1].um_I.iw[14] ;
 wire \top_I.branch[12].block[1].um_I.iw[15] ;
 wire \top_I.branch[12].block[1].um_I.iw[16] ;
 wire \top_I.branch[12].block[1].um_I.iw[17] ;
 wire \top_I.branch[12].block[1].um_I.iw[1] ;
 wire \top_I.branch[12].block[1].um_I.iw[2] ;
 wire \top_I.branch[12].block[1].um_I.iw[3] ;
 wire \top_I.branch[12].block[1].um_I.iw[4] ;
 wire \top_I.branch[12].block[1].um_I.iw[5] ;
 wire \top_I.branch[12].block[1].um_I.iw[6] ;
 wire \top_I.branch[12].block[1].um_I.iw[7] ;
 wire \top_I.branch[12].block[1].um_I.iw[8] ;
 wire \top_I.branch[12].block[1].um_I.iw[9] ;
 wire \top_I.branch[12].block[1].um_I.k_zero ;
 wire \top_I.branch[12].block[1].um_I.pg_vdd ;
 wire \top_I.branch[12].block[2].um_I.ana[2] ;
 wire \top_I.branch[12].block[2].um_I.ana[3] ;
 wire \top_I.branch[12].block[2].um_I.ana[4] ;
 wire \top_I.branch[12].block[2].um_I.ana[5] ;
 wire \top_I.branch[12].block[2].um_I.ana[6] ;
 wire \top_I.branch[12].block[2].um_I.ana[7] ;
 wire \top_I.branch[12].block[2].um_I.clk ;
 wire \top_I.branch[12].block[2].um_I.ena ;
 wire \top_I.branch[12].block[2].um_I.iw[10] ;
 wire \top_I.branch[12].block[2].um_I.iw[11] ;
 wire \top_I.branch[12].block[2].um_I.iw[12] ;
 wire \top_I.branch[12].block[2].um_I.iw[13] ;
 wire \top_I.branch[12].block[2].um_I.iw[14] ;
 wire \top_I.branch[12].block[2].um_I.iw[15] ;
 wire \top_I.branch[12].block[2].um_I.iw[16] ;
 wire \top_I.branch[12].block[2].um_I.iw[17] ;
 wire \top_I.branch[12].block[2].um_I.iw[1] ;
 wire \top_I.branch[12].block[2].um_I.iw[2] ;
 wire \top_I.branch[12].block[2].um_I.iw[3] ;
 wire \top_I.branch[12].block[2].um_I.iw[4] ;
 wire \top_I.branch[12].block[2].um_I.iw[5] ;
 wire \top_I.branch[12].block[2].um_I.iw[6] ;
 wire \top_I.branch[12].block[2].um_I.iw[7] ;
 wire \top_I.branch[12].block[2].um_I.iw[8] ;
 wire \top_I.branch[12].block[2].um_I.iw[9] ;
 wire \top_I.branch[12].block[2].um_I.k_zero ;
 wire \top_I.branch[12].block[2].um_I.pg_vdd ;
 wire \top_I.branch[12].block[3].um_I.ana[2] ;
 wire \top_I.branch[12].block[3].um_I.ana[3] ;
 wire \top_I.branch[12].block[3].um_I.ana[4] ;
 wire \top_I.branch[12].block[3].um_I.ana[5] ;
 wire \top_I.branch[12].block[3].um_I.ana[6] ;
 wire \top_I.branch[12].block[3].um_I.ana[7] ;
 wire \top_I.branch[12].block[3].um_I.clk ;
 wire \top_I.branch[12].block[3].um_I.ena ;
 wire \top_I.branch[12].block[3].um_I.iw[10] ;
 wire \top_I.branch[12].block[3].um_I.iw[11] ;
 wire \top_I.branch[12].block[3].um_I.iw[12] ;
 wire \top_I.branch[12].block[3].um_I.iw[13] ;
 wire \top_I.branch[12].block[3].um_I.iw[14] ;
 wire \top_I.branch[12].block[3].um_I.iw[15] ;
 wire \top_I.branch[12].block[3].um_I.iw[16] ;
 wire \top_I.branch[12].block[3].um_I.iw[17] ;
 wire \top_I.branch[12].block[3].um_I.iw[1] ;
 wire \top_I.branch[12].block[3].um_I.iw[2] ;
 wire \top_I.branch[12].block[3].um_I.iw[3] ;
 wire \top_I.branch[12].block[3].um_I.iw[4] ;
 wire \top_I.branch[12].block[3].um_I.iw[5] ;
 wire \top_I.branch[12].block[3].um_I.iw[6] ;
 wire \top_I.branch[12].block[3].um_I.iw[7] ;
 wire \top_I.branch[12].block[3].um_I.iw[8] ;
 wire \top_I.branch[12].block[3].um_I.iw[9] ;
 wire \top_I.branch[12].block[3].um_I.k_zero ;
 wire \top_I.branch[12].block[3].um_I.pg_vdd ;
 wire \top_I.branch[12].block[4].um_I.ana[2] ;
 wire \top_I.branch[12].block[4].um_I.ana[3] ;
 wire \top_I.branch[12].block[4].um_I.ana[4] ;
 wire \top_I.branch[12].block[4].um_I.ana[5] ;
 wire \top_I.branch[12].block[4].um_I.ana[6] ;
 wire \top_I.branch[12].block[4].um_I.ana[7] ;
 wire \top_I.branch[12].block[4].um_I.clk ;
 wire \top_I.branch[12].block[4].um_I.ena ;
 wire \top_I.branch[12].block[4].um_I.iw[10] ;
 wire \top_I.branch[12].block[4].um_I.iw[11] ;
 wire \top_I.branch[12].block[4].um_I.iw[12] ;
 wire \top_I.branch[12].block[4].um_I.iw[13] ;
 wire \top_I.branch[12].block[4].um_I.iw[14] ;
 wire \top_I.branch[12].block[4].um_I.iw[15] ;
 wire \top_I.branch[12].block[4].um_I.iw[16] ;
 wire \top_I.branch[12].block[4].um_I.iw[17] ;
 wire \top_I.branch[12].block[4].um_I.iw[1] ;
 wire \top_I.branch[12].block[4].um_I.iw[2] ;
 wire \top_I.branch[12].block[4].um_I.iw[3] ;
 wire \top_I.branch[12].block[4].um_I.iw[4] ;
 wire \top_I.branch[12].block[4].um_I.iw[5] ;
 wire \top_I.branch[12].block[4].um_I.iw[6] ;
 wire \top_I.branch[12].block[4].um_I.iw[7] ;
 wire \top_I.branch[12].block[4].um_I.iw[8] ;
 wire \top_I.branch[12].block[4].um_I.iw[9] ;
 wire \top_I.branch[12].block[4].um_I.k_zero ;
 wire \top_I.branch[12].block[4].um_I.pg_vdd ;
 wire \top_I.branch[12].block[5].um_I.ana[2] ;
 wire \top_I.branch[12].block[5].um_I.ana[3] ;
 wire \top_I.branch[12].block[5].um_I.ana[4] ;
 wire \top_I.branch[12].block[5].um_I.ana[5] ;
 wire \top_I.branch[12].block[5].um_I.ana[6] ;
 wire \top_I.branch[12].block[5].um_I.ana[7] ;
 wire \top_I.branch[12].block[5].um_I.clk ;
 wire \top_I.branch[12].block[5].um_I.ena ;
 wire \top_I.branch[12].block[5].um_I.iw[10] ;
 wire \top_I.branch[12].block[5].um_I.iw[11] ;
 wire \top_I.branch[12].block[5].um_I.iw[12] ;
 wire \top_I.branch[12].block[5].um_I.iw[13] ;
 wire \top_I.branch[12].block[5].um_I.iw[14] ;
 wire \top_I.branch[12].block[5].um_I.iw[15] ;
 wire \top_I.branch[12].block[5].um_I.iw[16] ;
 wire \top_I.branch[12].block[5].um_I.iw[17] ;
 wire \top_I.branch[12].block[5].um_I.iw[1] ;
 wire \top_I.branch[12].block[5].um_I.iw[2] ;
 wire \top_I.branch[12].block[5].um_I.iw[3] ;
 wire \top_I.branch[12].block[5].um_I.iw[4] ;
 wire \top_I.branch[12].block[5].um_I.iw[5] ;
 wire \top_I.branch[12].block[5].um_I.iw[6] ;
 wire \top_I.branch[12].block[5].um_I.iw[7] ;
 wire \top_I.branch[12].block[5].um_I.iw[8] ;
 wire \top_I.branch[12].block[5].um_I.iw[9] ;
 wire \top_I.branch[12].block[5].um_I.k_zero ;
 wire \top_I.branch[12].block[5].um_I.pg_vdd ;
 wire \top_I.branch[12].block[6].um_I.ana[2] ;
 wire \top_I.branch[12].block[6].um_I.ana[3] ;
 wire \top_I.branch[12].block[6].um_I.ana[4] ;
 wire \top_I.branch[12].block[6].um_I.ana[5] ;
 wire \top_I.branch[12].block[6].um_I.ana[6] ;
 wire \top_I.branch[12].block[6].um_I.ana[7] ;
 wire \top_I.branch[12].block[6].um_I.clk ;
 wire \top_I.branch[12].block[6].um_I.ena ;
 wire \top_I.branch[12].block[6].um_I.iw[10] ;
 wire \top_I.branch[12].block[6].um_I.iw[11] ;
 wire \top_I.branch[12].block[6].um_I.iw[12] ;
 wire \top_I.branch[12].block[6].um_I.iw[13] ;
 wire \top_I.branch[12].block[6].um_I.iw[14] ;
 wire \top_I.branch[12].block[6].um_I.iw[15] ;
 wire \top_I.branch[12].block[6].um_I.iw[16] ;
 wire \top_I.branch[12].block[6].um_I.iw[17] ;
 wire \top_I.branch[12].block[6].um_I.iw[1] ;
 wire \top_I.branch[12].block[6].um_I.iw[2] ;
 wire \top_I.branch[12].block[6].um_I.iw[3] ;
 wire \top_I.branch[12].block[6].um_I.iw[4] ;
 wire \top_I.branch[12].block[6].um_I.iw[5] ;
 wire \top_I.branch[12].block[6].um_I.iw[6] ;
 wire \top_I.branch[12].block[6].um_I.iw[7] ;
 wire \top_I.branch[12].block[6].um_I.iw[8] ;
 wire \top_I.branch[12].block[6].um_I.iw[9] ;
 wire \top_I.branch[12].block[6].um_I.k_zero ;
 wire \top_I.branch[12].block[6].um_I.pg_vdd ;
 wire \top_I.branch[12].block[7].um_I.ana[2] ;
 wire \top_I.branch[12].block[7].um_I.ana[3] ;
 wire \top_I.branch[12].block[7].um_I.ana[4] ;
 wire \top_I.branch[12].block[7].um_I.ana[5] ;
 wire \top_I.branch[12].block[7].um_I.ana[6] ;
 wire \top_I.branch[12].block[7].um_I.ana[7] ;
 wire \top_I.branch[12].block[7].um_I.clk ;
 wire \top_I.branch[12].block[7].um_I.ena ;
 wire \top_I.branch[12].block[7].um_I.iw[10] ;
 wire \top_I.branch[12].block[7].um_I.iw[11] ;
 wire \top_I.branch[12].block[7].um_I.iw[12] ;
 wire \top_I.branch[12].block[7].um_I.iw[13] ;
 wire \top_I.branch[12].block[7].um_I.iw[14] ;
 wire \top_I.branch[12].block[7].um_I.iw[15] ;
 wire \top_I.branch[12].block[7].um_I.iw[16] ;
 wire \top_I.branch[12].block[7].um_I.iw[17] ;
 wire \top_I.branch[12].block[7].um_I.iw[1] ;
 wire \top_I.branch[12].block[7].um_I.iw[2] ;
 wire \top_I.branch[12].block[7].um_I.iw[3] ;
 wire \top_I.branch[12].block[7].um_I.iw[4] ;
 wire \top_I.branch[12].block[7].um_I.iw[5] ;
 wire \top_I.branch[12].block[7].um_I.iw[6] ;
 wire \top_I.branch[12].block[7].um_I.iw[7] ;
 wire \top_I.branch[12].block[7].um_I.iw[8] ;
 wire \top_I.branch[12].block[7].um_I.iw[9] ;
 wire \top_I.branch[12].block[7].um_I.k_zero ;
 wire \top_I.branch[12].block[7].um_I.pg_vdd ;
 wire \top_I.branch[12].block[8].um_I.ana[2] ;
 wire \top_I.branch[12].block[8].um_I.ana[3] ;
 wire \top_I.branch[12].block[8].um_I.ana[4] ;
 wire \top_I.branch[12].block[8].um_I.ana[5] ;
 wire \top_I.branch[12].block[8].um_I.ana[6] ;
 wire \top_I.branch[12].block[8].um_I.ana[7] ;
 wire \top_I.branch[12].block[8].um_I.clk ;
 wire \top_I.branch[12].block[8].um_I.ena ;
 wire \top_I.branch[12].block[8].um_I.iw[10] ;
 wire \top_I.branch[12].block[8].um_I.iw[11] ;
 wire \top_I.branch[12].block[8].um_I.iw[12] ;
 wire \top_I.branch[12].block[8].um_I.iw[13] ;
 wire \top_I.branch[12].block[8].um_I.iw[14] ;
 wire \top_I.branch[12].block[8].um_I.iw[15] ;
 wire \top_I.branch[12].block[8].um_I.iw[16] ;
 wire \top_I.branch[12].block[8].um_I.iw[17] ;
 wire \top_I.branch[12].block[8].um_I.iw[1] ;
 wire \top_I.branch[12].block[8].um_I.iw[2] ;
 wire \top_I.branch[12].block[8].um_I.iw[3] ;
 wire \top_I.branch[12].block[8].um_I.iw[4] ;
 wire \top_I.branch[12].block[8].um_I.iw[5] ;
 wire \top_I.branch[12].block[8].um_I.iw[6] ;
 wire \top_I.branch[12].block[8].um_I.iw[7] ;
 wire \top_I.branch[12].block[8].um_I.iw[8] ;
 wire \top_I.branch[12].block[8].um_I.iw[9] ;
 wire \top_I.branch[12].block[8].um_I.k_zero ;
 wire \top_I.branch[12].block[8].um_I.pg_vdd ;
 wire \top_I.branch[12].block[9].um_I.ana[2] ;
 wire \top_I.branch[12].block[9].um_I.ana[3] ;
 wire \top_I.branch[12].block[9].um_I.ana[4] ;
 wire \top_I.branch[12].block[9].um_I.ana[5] ;
 wire \top_I.branch[12].block[9].um_I.ana[6] ;
 wire \top_I.branch[12].block[9].um_I.ana[7] ;
 wire \top_I.branch[12].block[9].um_I.clk ;
 wire \top_I.branch[12].block[9].um_I.ena ;
 wire \top_I.branch[12].block[9].um_I.iw[10] ;
 wire \top_I.branch[12].block[9].um_I.iw[11] ;
 wire \top_I.branch[12].block[9].um_I.iw[12] ;
 wire \top_I.branch[12].block[9].um_I.iw[13] ;
 wire \top_I.branch[12].block[9].um_I.iw[14] ;
 wire \top_I.branch[12].block[9].um_I.iw[15] ;
 wire \top_I.branch[12].block[9].um_I.iw[16] ;
 wire \top_I.branch[12].block[9].um_I.iw[17] ;
 wire \top_I.branch[12].block[9].um_I.iw[1] ;
 wire \top_I.branch[12].block[9].um_I.iw[2] ;
 wire \top_I.branch[12].block[9].um_I.iw[3] ;
 wire \top_I.branch[12].block[9].um_I.iw[4] ;
 wire \top_I.branch[12].block[9].um_I.iw[5] ;
 wire \top_I.branch[12].block[9].um_I.iw[6] ;
 wire \top_I.branch[12].block[9].um_I.iw[7] ;
 wire \top_I.branch[12].block[9].um_I.iw[8] ;
 wire \top_I.branch[12].block[9].um_I.iw[9] ;
 wire \top_I.branch[12].block[9].um_I.k_zero ;
 wire \top_I.branch[12].block[9].um_I.pg_vdd ;
 wire \top_I.branch[12].l_addr[0] ;
 wire \top_I.branch[12].l_addr[1] ;
 wire \top_I.branch[13].block[0].um_I.ana[2] ;
 wire \top_I.branch[13].block[0].um_I.ana[3] ;
 wire \top_I.branch[13].block[0].um_I.ana[4] ;
 wire \top_I.branch[13].block[0].um_I.ana[5] ;
 wire \top_I.branch[13].block[0].um_I.ana[6] ;
 wire \top_I.branch[13].block[0].um_I.ana[7] ;
 wire \top_I.branch[13].block[0].um_I.clk ;
 wire \top_I.branch[13].block[0].um_I.ena ;
 wire \top_I.branch[13].block[0].um_I.iw[10] ;
 wire \top_I.branch[13].block[0].um_I.iw[11] ;
 wire \top_I.branch[13].block[0].um_I.iw[12] ;
 wire \top_I.branch[13].block[0].um_I.iw[13] ;
 wire \top_I.branch[13].block[0].um_I.iw[14] ;
 wire \top_I.branch[13].block[0].um_I.iw[15] ;
 wire \top_I.branch[13].block[0].um_I.iw[16] ;
 wire \top_I.branch[13].block[0].um_I.iw[17] ;
 wire \top_I.branch[13].block[0].um_I.iw[1] ;
 wire \top_I.branch[13].block[0].um_I.iw[2] ;
 wire \top_I.branch[13].block[0].um_I.iw[3] ;
 wire \top_I.branch[13].block[0].um_I.iw[4] ;
 wire \top_I.branch[13].block[0].um_I.iw[5] ;
 wire \top_I.branch[13].block[0].um_I.iw[6] ;
 wire \top_I.branch[13].block[0].um_I.iw[7] ;
 wire \top_I.branch[13].block[0].um_I.iw[8] ;
 wire \top_I.branch[13].block[0].um_I.iw[9] ;
 wire \top_I.branch[13].block[0].um_I.k_zero ;
 wire \top_I.branch[13].block[0].um_I.pg_vdd ;
 wire \top_I.branch[13].block[10].um_I.ana[2] ;
 wire \top_I.branch[13].block[10].um_I.ana[3] ;
 wire \top_I.branch[13].block[10].um_I.ana[4] ;
 wire \top_I.branch[13].block[10].um_I.ana[5] ;
 wire \top_I.branch[13].block[10].um_I.ana[6] ;
 wire \top_I.branch[13].block[10].um_I.ana[7] ;
 wire \top_I.branch[13].block[10].um_I.clk ;
 wire \top_I.branch[13].block[10].um_I.ena ;
 wire \top_I.branch[13].block[10].um_I.iw[10] ;
 wire \top_I.branch[13].block[10].um_I.iw[11] ;
 wire \top_I.branch[13].block[10].um_I.iw[12] ;
 wire \top_I.branch[13].block[10].um_I.iw[13] ;
 wire \top_I.branch[13].block[10].um_I.iw[14] ;
 wire \top_I.branch[13].block[10].um_I.iw[15] ;
 wire \top_I.branch[13].block[10].um_I.iw[16] ;
 wire \top_I.branch[13].block[10].um_I.iw[17] ;
 wire \top_I.branch[13].block[10].um_I.iw[1] ;
 wire \top_I.branch[13].block[10].um_I.iw[2] ;
 wire \top_I.branch[13].block[10].um_I.iw[3] ;
 wire \top_I.branch[13].block[10].um_I.iw[4] ;
 wire \top_I.branch[13].block[10].um_I.iw[5] ;
 wire \top_I.branch[13].block[10].um_I.iw[6] ;
 wire \top_I.branch[13].block[10].um_I.iw[7] ;
 wire \top_I.branch[13].block[10].um_I.iw[8] ;
 wire \top_I.branch[13].block[10].um_I.iw[9] ;
 wire \top_I.branch[13].block[10].um_I.k_zero ;
 wire \top_I.branch[13].block[10].um_I.pg_vdd ;
 wire \top_I.branch[13].block[11].um_I.ana[2] ;
 wire \top_I.branch[13].block[11].um_I.ana[3] ;
 wire \top_I.branch[13].block[11].um_I.ana[4] ;
 wire \top_I.branch[13].block[11].um_I.ana[5] ;
 wire \top_I.branch[13].block[11].um_I.ana[6] ;
 wire \top_I.branch[13].block[11].um_I.ana[7] ;
 wire \top_I.branch[13].block[11].um_I.clk ;
 wire \top_I.branch[13].block[11].um_I.ena ;
 wire \top_I.branch[13].block[11].um_I.iw[10] ;
 wire \top_I.branch[13].block[11].um_I.iw[11] ;
 wire \top_I.branch[13].block[11].um_I.iw[12] ;
 wire \top_I.branch[13].block[11].um_I.iw[13] ;
 wire \top_I.branch[13].block[11].um_I.iw[14] ;
 wire \top_I.branch[13].block[11].um_I.iw[15] ;
 wire \top_I.branch[13].block[11].um_I.iw[16] ;
 wire \top_I.branch[13].block[11].um_I.iw[17] ;
 wire \top_I.branch[13].block[11].um_I.iw[1] ;
 wire \top_I.branch[13].block[11].um_I.iw[2] ;
 wire \top_I.branch[13].block[11].um_I.iw[3] ;
 wire \top_I.branch[13].block[11].um_I.iw[4] ;
 wire \top_I.branch[13].block[11].um_I.iw[5] ;
 wire \top_I.branch[13].block[11].um_I.iw[6] ;
 wire \top_I.branch[13].block[11].um_I.iw[7] ;
 wire \top_I.branch[13].block[11].um_I.iw[8] ;
 wire \top_I.branch[13].block[11].um_I.iw[9] ;
 wire \top_I.branch[13].block[11].um_I.k_zero ;
 wire \top_I.branch[13].block[11].um_I.pg_vdd ;
 wire \top_I.branch[13].block[12].um_I.ana[2] ;
 wire \top_I.branch[13].block[12].um_I.ana[3] ;
 wire \top_I.branch[13].block[12].um_I.ana[4] ;
 wire \top_I.branch[13].block[12].um_I.ana[5] ;
 wire \top_I.branch[13].block[12].um_I.ana[6] ;
 wire \top_I.branch[13].block[12].um_I.ana[7] ;
 wire \top_I.branch[13].block[12].um_I.clk ;
 wire \top_I.branch[13].block[12].um_I.ena ;
 wire \top_I.branch[13].block[12].um_I.iw[10] ;
 wire \top_I.branch[13].block[12].um_I.iw[11] ;
 wire \top_I.branch[13].block[12].um_I.iw[12] ;
 wire \top_I.branch[13].block[12].um_I.iw[13] ;
 wire \top_I.branch[13].block[12].um_I.iw[14] ;
 wire \top_I.branch[13].block[12].um_I.iw[15] ;
 wire \top_I.branch[13].block[12].um_I.iw[16] ;
 wire \top_I.branch[13].block[12].um_I.iw[17] ;
 wire \top_I.branch[13].block[12].um_I.iw[1] ;
 wire \top_I.branch[13].block[12].um_I.iw[2] ;
 wire \top_I.branch[13].block[12].um_I.iw[3] ;
 wire \top_I.branch[13].block[12].um_I.iw[4] ;
 wire \top_I.branch[13].block[12].um_I.iw[5] ;
 wire \top_I.branch[13].block[12].um_I.iw[6] ;
 wire \top_I.branch[13].block[12].um_I.iw[7] ;
 wire \top_I.branch[13].block[12].um_I.iw[8] ;
 wire \top_I.branch[13].block[12].um_I.iw[9] ;
 wire \top_I.branch[13].block[12].um_I.k_zero ;
 wire \top_I.branch[13].block[12].um_I.pg_vdd ;
 wire \top_I.branch[13].block[13].um_I.ana[2] ;
 wire \top_I.branch[13].block[13].um_I.ana[3] ;
 wire \top_I.branch[13].block[13].um_I.ana[4] ;
 wire \top_I.branch[13].block[13].um_I.ana[5] ;
 wire \top_I.branch[13].block[13].um_I.ana[6] ;
 wire \top_I.branch[13].block[13].um_I.ana[7] ;
 wire \top_I.branch[13].block[13].um_I.clk ;
 wire \top_I.branch[13].block[13].um_I.ena ;
 wire \top_I.branch[13].block[13].um_I.iw[10] ;
 wire \top_I.branch[13].block[13].um_I.iw[11] ;
 wire \top_I.branch[13].block[13].um_I.iw[12] ;
 wire \top_I.branch[13].block[13].um_I.iw[13] ;
 wire \top_I.branch[13].block[13].um_I.iw[14] ;
 wire \top_I.branch[13].block[13].um_I.iw[15] ;
 wire \top_I.branch[13].block[13].um_I.iw[16] ;
 wire \top_I.branch[13].block[13].um_I.iw[17] ;
 wire \top_I.branch[13].block[13].um_I.iw[1] ;
 wire \top_I.branch[13].block[13].um_I.iw[2] ;
 wire \top_I.branch[13].block[13].um_I.iw[3] ;
 wire \top_I.branch[13].block[13].um_I.iw[4] ;
 wire \top_I.branch[13].block[13].um_I.iw[5] ;
 wire \top_I.branch[13].block[13].um_I.iw[6] ;
 wire \top_I.branch[13].block[13].um_I.iw[7] ;
 wire \top_I.branch[13].block[13].um_I.iw[8] ;
 wire \top_I.branch[13].block[13].um_I.iw[9] ;
 wire \top_I.branch[13].block[13].um_I.k_zero ;
 wire \top_I.branch[13].block[13].um_I.pg_vdd ;
 wire \top_I.branch[13].block[14].um_I.ana[2] ;
 wire \top_I.branch[13].block[14].um_I.ana[3] ;
 wire \top_I.branch[13].block[14].um_I.ana[4] ;
 wire \top_I.branch[13].block[14].um_I.ana[5] ;
 wire \top_I.branch[13].block[14].um_I.ana[6] ;
 wire \top_I.branch[13].block[14].um_I.ana[7] ;
 wire \top_I.branch[13].block[14].um_I.clk ;
 wire \top_I.branch[13].block[14].um_I.ena ;
 wire \top_I.branch[13].block[14].um_I.iw[10] ;
 wire \top_I.branch[13].block[14].um_I.iw[11] ;
 wire \top_I.branch[13].block[14].um_I.iw[12] ;
 wire \top_I.branch[13].block[14].um_I.iw[13] ;
 wire \top_I.branch[13].block[14].um_I.iw[14] ;
 wire \top_I.branch[13].block[14].um_I.iw[15] ;
 wire \top_I.branch[13].block[14].um_I.iw[16] ;
 wire \top_I.branch[13].block[14].um_I.iw[17] ;
 wire \top_I.branch[13].block[14].um_I.iw[1] ;
 wire \top_I.branch[13].block[14].um_I.iw[2] ;
 wire \top_I.branch[13].block[14].um_I.iw[3] ;
 wire \top_I.branch[13].block[14].um_I.iw[4] ;
 wire \top_I.branch[13].block[14].um_I.iw[5] ;
 wire \top_I.branch[13].block[14].um_I.iw[6] ;
 wire \top_I.branch[13].block[14].um_I.iw[7] ;
 wire \top_I.branch[13].block[14].um_I.iw[8] ;
 wire \top_I.branch[13].block[14].um_I.iw[9] ;
 wire \top_I.branch[13].block[14].um_I.k_zero ;
 wire \top_I.branch[13].block[14].um_I.pg_vdd ;
 wire \top_I.branch[13].block[15].um_I.ana[2] ;
 wire \top_I.branch[13].block[15].um_I.ana[3] ;
 wire \top_I.branch[13].block[15].um_I.ana[4] ;
 wire \top_I.branch[13].block[15].um_I.ana[5] ;
 wire \top_I.branch[13].block[15].um_I.ana[6] ;
 wire \top_I.branch[13].block[15].um_I.ana[7] ;
 wire \top_I.branch[13].block[15].um_I.clk ;
 wire \top_I.branch[13].block[15].um_I.ena ;
 wire \top_I.branch[13].block[15].um_I.iw[10] ;
 wire \top_I.branch[13].block[15].um_I.iw[11] ;
 wire \top_I.branch[13].block[15].um_I.iw[12] ;
 wire \top_I.branch[13].block[15].um_I.iw[13] ;
 wire \top_I.branch[13].block[15].um_I.iw[14] ;
 wire \top_I.branch[13].block[15].um_I.iw[15] ;
 wire \top_I.branch[13].block[15].um_I.iw[16] ;
 wire \top_I.branch[13].block[15].um_I.iw[17] ;
 wire \top_I.branch[13].block[15].um_I.iw[1] ;
 wire \top_I.branch[13].block[15].um_I.iw[2] ;
 wire \top_I.branch[13].block[15].um_I.iw[3] ;
 wire \top_I.branch[13].block[15].um_I.iw[4] ;
 wire \top_I.branch[13].block[15].um_I.iw[5] ;
 wire \top_I.branch[13].block[15].um_I.iw[6] ;
 wire \top_I.branch[13].block[15].um_I.iw[7] ;
 wire \top_I.branch[13].block[15].um_I.iw[8] ;
 wire \top_I.branch[13].block[15].um_I.iw[9] ;
 wire \top_I.branch[13].block[15].um_I.k_zero ;
 wire \top_I.branch[13].block[15].um_I.pg_vdd ;
 wire \top_I.branch[13].block[1].um_I.ana[2] ;
 wire \top_I.branch[13].block[1].um_I.ana[3] ;
 wire \top_I.branch[13].block[1].um_I.ana[4] ;
 wire \top_I.branch[13].block[1].um_I.ana[5] ;
 wire \top_I.branch[13].block[1].um_I.ana[6] ;
 wire \top_I.branch[13].block[1].um_I.ana[7] ;
 wire \top_I.branch[13].block[1].um_I.clk ;
 wire \top_I.branch[13].block[1].um_I.ena ;
 wire \top_I.branch[13].block[1].um_I.iw[10] ;
 wire \top_I.branch[13].block[1].um_I.iw[11] ;
 wire \top_I.branch[13].block[1].um_I.iw[12] ;
 wire \top_I.branch[13].block[1].um_I.iw[13] ;
 wire \top_I.branch[13].block[1].um_I.iw[14] ;
 wire \top_I.branch[13].block[1].um_I.iw[15] ;
 wire \top_I.branch[13].block[1].um_I.iw[16] ;
 wire \top_I.branch[13].block[1].um_I.iw[17] ;
 wire \top_I.branch[13].block[1].um_I.iw[1] ;
 wire \top_I.branch[13].block[1].um_I.iw[2] ;
 wire \top_I.branch[13].block[1].um_I.iw[3] ;
 wire \top_I.branch[13].block[1].um_I.iw[4] ;
 wire \top_I.branch[13].block[1].um_I.iw[5] ;
 wire \top_I.branch[13].block[1].um_I.iw[6] ;
 wire \top_I.branch[13].block[1].um_I.iw[7] ;
 wire \top_I.branch[13].block[1].um_I.iw[8] ;
 wire \top_I.branch[13].block[1].um_I.iw[9] ;
 wire \top_I.branch[13].block[1].um_I.k_zero ;
 wire \top_I.branch[13].block[1].um_I.pg_vdd ;
 wire \top_I.branch[13].block[2].um_I.ana[2] ;
 wire \top_I.branch[13].block[2].um_I.ana[3] ;
 wire \top_I.branch[13].block[2].um_I.ana[4] ;
 wire \top_I.branch[13].block[2].um_I.ana[5] ;
 wire \top_I.branch[13].block[2].um_I.ana[6] ;
 wire \top_I.branch[13].block[2].um_I.ana[7] ;
 wire \top_I.branch[13].block[2].um_I.clk ;
 wire \top_I.branch[13].block[2].um_I.ena ;
 wire \top_I.branch[13].block[2].um_I.iw[10] ;
 wire \top_I.branch[13].block[2].um_I.iw[11] ;
 wire \top_I.branch[13].block[2].um_I.iw[12] ;
 wire \top_I.branch[13].block[2].um_I.iw[13] ;
 wire \top_I.branch[13].block[2].um_I.iw[14] ;
 wire \top_I.branch[13].block[2].um_I.iw[15] ;
 wire \top_I.branch[13].block[2].um_I.iw[16] ;
 wire \top_I.branch[13].block[2].um_I.iw[17] ;
 wire \top_I.branch[13].block[2].um_I.iw[1] ;
 wire \top_I.branch[13].block[2].um_I.iw[2] ;
 wire \top_I.branch[13].block[2].um_I.iw[3] ;
 wire \top_I.branch[13].block[2].um_I.iw[4] ;
 wire \top_I.branch[13].block[2].um_I.iw[5] ;
 wire \top_I.branch[13].block[2].um_I.iw[6] ;
 wire \top_I.branch[13].block[2].um_I.iw[7] ;
 wire \top_I.branch[13].block[2].um_I.iw[8] ;
 wire \top_I.branch[13].block[2].um_I.iw[9] ;
 wire \top_I.branch[13].block[2].um_I.k_zero ;
 wire \top_I.branch[13].block[2].um_I.pg_vdd ;
 wire \top_I.branch[13].block[3].um_I.ana[2] ;
 wire \top_I.branch[13].block[3].um_I.ana[3] ;
 wire \top_I.branch[13].block[3].um_I.ana[4] ;
 wire \top_I.branch[13].block[3].um_I.ana[5] ;
 wire \top_I.branch[13].block[3].um_I.ana[6] ;
 wire \top_I.branch[13].block[3].um_I.ana[7] ;
 wire \top_I.branch[13].block[3].um_I.clk ;
 wire \top_I.branch[13].block[3].um_I.ena ;
 wire \top_I.branch[13].block[3].um_I.iw[10] ;
 wire \top_I.branch[13].block[3].um_I.iw[11] ;
 wire \top_I.branch[13].block[3].um_I.iw[12] ;
 wire \top_I.branch[13].block[3].um_I.iw[13] ;
 wire \top_I.branch[13].block[3].um_I.iw[14] ;
 wire \top_I.branch[13].block[3].um_I.iw[15] ;
 wire \top_I.branch[13].block[3].um_I.iw[16] ;
 wire \top_I.branch[13].block[3].um_I.iw[17] ;
 wire \top_I.branch[13].block[3].um_I.iw[1] ;
 wire \top_I.branch[13].block[3].um_I.iw[2] ;
 wire \top_I.branch[13].block[3].um_I.iw[3] ;
 wire \top_I.branch[13].block[3].um_I.iw[4] ;
 wire \top_I.branch[13].block[3].um_I.iw[5] ;
 wire \top_I.branch[13].block[3].um_I.iw[6] ;
 wire \top_I.branch[13].block[3].um_I.iw[7] ;
 wire \top_I.branch[13].block[3].um_I.iw[8] ;
 wire \top_I.branch[13].block[3].um_I.iw[9] ;
 wire \top_I.branch[13].block[3].um_I.k_zero ;
 wire \top_I.branch[13].block[3].um_I.pg_vdd ;
 wire \top_I.branch[13].block[4].um_I.ana[2] ;
 wire \top_I.branch[13].block[4].um_I.ana[3] ;
 wire \top_I.branch[13].block[4].um_I.ana[4] ;
 wire \top_I.branch[13].block[4].um_I.ana[5] ;
 wire \top_I.branch[13].block[4].um_I.ana[6] ;
 wire \top_I.branch[13].block[4].um_I.ana[7] ;
 wire \top_I.branch[13].block[4].um_I.clk ;
 wire \top_I.branch[13].block[4].um_I.ena ;
 wire \top_I.branch[13].block[4].um_I.iw[10] ;
 wire \top_I.branch[13].block[4].um_I.iw[11] ;
 wire \top_I.branch[13].block[4].um_I.iw[12] ;
 wire \top_I.branch[13].block[4].um_I.iw[13] ;
 wire \top_I.branch[13].block[4].um_I.iw[14] ;
 wire \top_I.branch[13].block[4].um_I.iw[15] ;
 wire \top_I.branch[13].block[4].um_I.iw[16] ;
 wire \top_I.branch[13].block[4].um_I.iw[17] ;
 wire \top_I.branch[13].block[4].um_I.iw[1] ;
 wire \top_I.branch[13].block[4].um_I.iw[2] ;
 wire \top_I.branch[13].block[4].um_I.iw[3] ;
 wire \top_I.branch[13].block[4].um_I.iw[4] ;
 wire \top_I.branch[13].block[4].um_I.iw[5] ;
 wire \top_I.branch[13].block[4].um_I.iw[6] ;
 wire \top_I.branch[13].block[4].um_I.iw[7] ;
 wire \top_I.branch[13].block[4].um_I.iw[8] ;
 wire \top_I.branch[13].block[4].um_I.iw[9] ;
 wire \top_I.branch[13].block[4].um_I.k_zero ;
 wire \top_I.branch[13].block[4].um_I.pg_vdd ;
 wire \top_I.branch[13].block[5].um_I.ana[2] ;
 wire \top_I.branch[13].block[5].um_I.ana[3] ;
 wire \top_I.branch[13].block[5].um_I.ana[4] ;
 wire \top_I.branch[13].block[5].um_I.ana[5] ;
 wire \top_I.branch[13].block[5].um_I.ana[6] ;
 wire \top_I.branch[13].block[5].um_I.ana[7] ;
 wire \top_I.branch[13].block[5].um_I.clk ;
 wire \top_I.branch[13].block[5].um_I.ena ;
 wire \top_I.branch[13].block[5].um_I.iw[10] ;
 wire \top_I.branch[13].block[5].um_I.iw[11] ;
 wire \top_I.branch[13].block[5].um_I.iw[12] ;
 wire \top_I.branch[13].block[5].um_I.iw[13] ;
 wire \top_I.branch[13].block[5].um_I.iw[14] ;
 wire \top_I.branch[13].block[5].um_I.iw[15] ;
 wire \top_I.branch[13].block[5].um_I.iw[16] ;
 wire \top_I.branch[13].block[5].um_I.iw[17] ;
 wire \top_I.branch[13].block[5].um_I.iw[1] ;
 wire \top_I.branch[13].block[5].um_I.iw[2] ;
 wire \top_I.branch[13].block[5].um_I.iw[3] ;
 wire \top_I.branch[13].block[5].um_I.iw[4] ;
 wire \top_I.branch[13].block[5].um_I.iw[5] ;
 wire \top_I.branch[13].block[5].um_I.iw[6] ;
 wire \top_I.branch[13].block[5].um_I.iw[7] ;
 wire \top_I.branch[13].block[5].um_I.iw[8] ;
 wire \top_I.branch[13].block[5].um_I.iw[9] ;
 wire \top_I.branch[13].block[5].um_I.k_zero ;
 wire \top_I.branch[13].block[5].um_I.pg_vdd ;
 wire \top_I.branch[13].block[6].um_I.ana[2] ;
 wire \top_I.branch[13].block[6].um_I.ana[3] ;
 wire \top_I.branch[13].block[6].um_I.ana[4] ;
 wire \top_I.branch[13].block[6].um_I.ana[5] ;
 wire \top_I.branch[13].block[6].um_I.ana[6] ;
 wire \top_I.branch[13].block[6].um_I.ana[7] ;
 wire \top_I.branch[13].block[6].um_I.clk ;
 wire \top_I.branch[13].block[6].um_I.ena ;
 wire \top_I.branch[13].block[6].um_I.iw[10] ;
 wire \top_I.branch[13].block[6].um_I.iw[11] ;
 wire \top_I.branch[13].block[6].um_I.iw[12] ;
 wire \top_I.branch[13].block[6].um_I.iw[13] ;
 wire \top_I.branch[13].block[6].um_I.iw[14] ;
 wire \top_I.branch[13].block[6].um_I.iw[15] ;
 wire \top_I.branch[13].block[6].um_I.iw[16] ;
 wire \top_I.branch[13].block[6].um_I.iw[17] ;
 wire \top_I.branch[13].block[6].um_I.iw[1] ;
 wire \top_I.branch[13].block[6].um_I.iw[2] ;
 wire \top_I.branch[13].block[6].um_I.iw[3] ;
 wire \top_I.branch[13].block[6].um_I.iw[4] ;
 wire \top_I.branch[13].block[6].um_I.iw[5] ;
 wire \top_I.branch[13].block[6].um_I.iw[6] ;
 wire \top_I.branch[13].block[6].um_I.iw[7] ;
 wire \top_I.branch[13].block[6].um_I.iw[8] ;
 wire \top_I.branch[13].block[6].um_I.iw[9] ;
 wire \top_I.branch[13].block[6].um_I.k_zero ;
 wire \top_I.branch[13].block[6].um_I.pg_vdd ;
 wire \top_I.branch[13].block[7].um_I.ana[2] ;
 wire \top_I.branch[13].block[7].um_I.ana[3] ;
 wire \top_I.branch[13].block[7].um_I.ana[4] ;
 wire \top_I.branch[13].block[7].um_I.ana[5] ;
 wire \top_I.branch[13].block[7].um_I.ana[6] ;
 wire \top_I.branch[13].block[7].um_I.ana[7] ;
 wire \top_I.branch[13].block[7].um_I.clk ;
 wire \top_I.branch[13].block[7].um_I.ena ;
 wire \top_I.branch[13].block[7].um_I.iw[10] ;
 wire \top_I.branch[13].block[7].um_I.iw[11] ;
 wire \top_I.branch[13].block[7].um_I.iw[12] ;
 wire \top_I.branch[13].block[7].um_I.iw[13] ;
 wire \top_I.branch[13].block[7].um_I.iw[14] ;
 wire \top_I.branch[13].block[7].um_I.iw[15] ;
 wire \top_I.branch[13].block[7].um_I.iw[16] ;
 wire \top_I.branch[13].block[7].um_I.iw[17] ;
 wire \top_I.branch[13].block[7].um_I.iw[1] ;
 wire \top_I.branch[13].block[7].um_I.iw[2] ;
 wire \top_I.branch[13].block[7].um_I.iw[3] ;
 wire \top_I.branch[13].block[7].um_I.iw[4] ;
 wire \top_I.branch[13].block[7].um_I.iw[5] ;
 wire \top_I.branch[13].block[7].um_I.iw[6] ;
 wire \top_I.branch[13].block[7].um_I.iw[7] ;
 wire \top_I.branch[13].block[7].um_I.iw[8] ;
 wire \top_I.branch[13].block[7].um_I.iw[9] ;
 wire \top_I.branch[13].block[7].um_I.k_zero ;
 wire \top_I.branch[13].block[7].um_I.pg_vdd ;
 wire \top_I.branch[13].block[8].um_I.ana[2] ;
 wire \top_I.branch[13].block[8].um_I.ana[3] ;
 wire \top_I.branch[13].block[8].um_I.ana[4] ;
 wire \top_I.branch[13].block[8].um_I.ana[5] ;
 wire \top_I.branch[13].block[8].um_I.ana[6] ;
 wire \top_I.branch[13].block[8].um_I.ana[7] ;
 wire \top_I.branch[13].block[8].um_I.clk ;
 wire \top_I.branch[13].block[8].um_I.ena ;
 wire \top_I.branch[13].block[8].um_I.iw[10] ;
 wire \top_I.branch[13].block[8].um_I.iw[11] ;
 wire \top_I.branch[13].block[8].um_I.iw[12] ;
 wire \top_I.branch[13].block[8].um_I.iw[13] ;
 wire \top_I.branch[13].block[8].um_I.iw[14] ;
 wire \top_I.branch[13].block[8].um_I.iw[15] ;
 wire \top_I.branch[13].block[8].um_I.iw[16] ;
 wire \top_I.branch[13].block[8].um_I.iw[17] ;
 wire \top_I.branch[13].block[8].um_I.iw[1] ;
 wire \top_I.branch[13].block[8].um_I.iw[2] ;
 wire \top_I.branch[13].block[8].um_I.iw[3] ;
 wire \top_I.branch[13].block[8].um_I.iw[4] ;
 wire \top_I.branch[13].block[8].um_I.iw[5] ;
 wire \top_I.branch[13].block[8].um_I.iw[6] ;
 wire \top_I.branch[13].block[8].um_I.iw[7] ;
 wire \top_I.branch[13].block[8].um_I.iw[8] ;
 wire \top_I.branch[13].block[8].um_I.iw[9] ;
 wire \top_I.branch[13].block[8].um_I.k_zero ;
 wire \top_I.branch[13].block[8].um_I.pg_vdd ;
 wire \top_I.branch[13].block[9].um_I.ana[2] ;
 wire \top_I.branch[13].block[9].um_I.ana[3] ;
 wire \top_I.branch[13].block[9].um_I.ana[4] ;
 wire \top_I.branch[13].block[9].um_I.ana[5] ;
 wire \top_I.branch[13].block[9].um_I.ana[6] ;
 wire \top_I.branch[13].block[9].um_I.ana[7] ;
 wire \top_I.branch[13].block[9].um_I.clk ;
 wire \top_I.branch[13].block[9].um_I.ena ;
 wire \top_I.branch[13].block[9].um_I.iw[10] ;
 wire \top_I.branch[13].block[9].um_I.iw[11] ;
 wire \top_I.branch[13].block[9].um_I.iw[12] ;
 wire \top_I.branch[13].block[9].um_I.iw[13] ;
 wire \top_I.branch[13].block[9].um_I.iw[14] ;
 wire \top_I.branch[13].block[9].um_I.iw[15] ;
 wire \top_I.branch[13].block[9].um_I.iw[16] ;
 wire \top_I.branch[13].block[9].um_I.iw[17] ;
 wire \top_I.branch[13].block[9].um_I.iw[1] ;
 wire \top_I.branch[13].block[9].um_I.iw[2] ;
 wire \top_I.branch[13].block[9].um_I.iw[3] ;
 wire \top_I.branch[13].block[9].um_I.iw[4] ;
 wire \top_I.branch[13].block[9].um_I.iw[5] ;
 wire \top_I.branch[13].block[9].um_I.iw[6] ;
 wire \top_I.branch[13].block[9].um_I.iw[7] ;
 wire \top_I.branch[13].block[9].um_I.iw[8] ;
 wire \top_I.branch[13].block[9].um_I.iw[9] ;
 wire \top_I.branch[13].block[9].um_I.k_zero ;
 wire \top_I.branch[13].block[9].um_I.pg_vdd ;
 wire \top_I.branch[13].l_addr[0] ;
 wire \top_I.branch[13].l_addr[1] ;
 wire \top_I.branch[14].block[0].um_I.ana[2] ;
 wire \top_I.branch[14].block[0].um_I.ana[3] ;
 wire \top_I.branch[14].block[0].um_I.ana[4] ;
 wire \top_I.branch[14].block[0].um_I.ana[5] ;
 wire \top_I.branch[14].block[0].um_I.ana[6] ;
 wire \top_I.branch[14].block[0].um_I.ana[7] ;
 wire \top_I.branch[14].block[0].um_I.clk ;
 wire \top_I.branch[14].block[0].um_I.ena ;
 wire \top_I.branch[14].block[0].um_I.iw[10] ;
 wire \top_I.branch[14].block[0].um_I.iw[11] ;
 wire \top_I.branch[14].block[0].um_I.iw[12] ;
 wire \top_I.branch[14].block[0].um_I.iw[13] ;
 wire \top_I.branch[14].block[0].um_I.iw[14] ;
 wire \top_I.branch[14].block[0].um_I.iw[15] ;
 wire \top_I.branch[14].block[0].um_I.iw[16] ;
 wire \top_I.branch[14].block[0].um_I.iw[17] ;
 wire \top_I.branch[14].block[0].um_I.iw[1] ;
 wire \top_I.branch[14].block[0].um_I.iw[2] ;
 wire \top_I.branch[14].block[0].um_I.iw[3] ;
 wire \top_I.branch[14].block[0].um_I.iw[4] ;
 wire \top_I.branch[14].block[0].um_I.iw[5] ;
 wire \top_I.branch[14].block[0].um_I.iw[6] ;
 wire \top_I.branch[14].block[0].um_I.iw[7] ;
 wire \top_I.branch[14].block[0].um_I.iw[8] ;
 wire \top_I.branch[14].block[0].um_I.iw[9] ;
 wire \top_I.branch[14].block[0].um_I.k_zero ;
 wire \top_I.branch[14].block[0].um_I.pg_vdd ;
 wire \top_I.branch[14].block[10].um_I.ana[2] ;
 wire \top_I.branch[14].block[10].um_I.ana[3] ;
 wire \top_I.branch[14].block[10].um_I.ana[4] ;
 wire \top_I.branch[14].block[10].um_I.ana[5] ;
 wire \top_I.branch[14].block[10].um_I.ana[6] ;
 wire \top_I.branch[14].block[10].um_I.ana[7] ;
 wire \top_I.branch[14].block[10].um_I.clk ;
 wire \top_I.branch[14].block[10].um_I.ena ;
 wire \top_I.branch[14].block[10].um_I.iw[10] ;
 wire \top_I.branch[14].block[10].um_I.iw[11] ;
 wire \top_I.branch[14].block[10].um_I.iw[12] ;
 wire \top_I.branch[14].block[10].um_I.iw[13] ;
 wire \top_I.branch[14].block[10].um_I.iw[14] ;
 wire \top_I.branch[14].block[10].um_I.iw[15] ;
 wire \top_I.branch[14].block[10].um_I.iw[16] ;
 wire \top_I.branch[14].block[10].um_I.iw[17] ;
 wire \top_I.branch[14].block[10].um_I.iw[1] ;
 wire \top_I.branch[14].block[10].um_I.iw[2] ;
 wire \top_I.branch[14].block[10].um_I.iw[3] ;
 wire \top_I.branch[14].block[10].um_I.iw[4] ;
 wire \top_I.branch[14].block[10].um_I.iw[5] ;
 wire \top_I.branch[14].block[10].um_I.iw[6] ;
 wire \top_I.branch[14].block[10].um_I.iw[7] ;
 wire \top_I.branch[14].block[10].um_I.iw[8] ;
 wire \top_I.branch[14].block[10].um_I.iw[9] ;
 wire \top_I.branch[14].block[10].um_I.k_zero ;
 wire \top_I.branch[14].block[10].um_I.pg_vdd ;
 wire \top_I.branch[14].block[11].um_I.ana[2] ;
 wire \top_I.branch[14].block[11].um_I.ana[3] ;
 wire \top_I.branch[14].block[11].um_I.ana[4] ;
 wire \top_I.branch[14].block[11].um_I.ana[5] ;
 wire \top_I.branch[14].block[11].um_I.ana[6] ;
 wire \top_I.branch[14].block[11].um_I.ana[7] ;
 wire \top_I.branch[14].block[11].um_I.clk ;
 wire \top_I.branch[14].block[11].um_I.ena ;
 wire \top_I.branch[14].block[11].um_I.iw[10] ;
 wire \top_I.branch[14].block[11].um_I.iw[11] ;
 wire \top_I.branch[14].block[11].um_I.iw[12] ;
 wire \top_I.branch[14].block[11].um_I.iw[13] ;
 wire \top_I.branch[14].block[11].um_I.iw[14] ;
 wire \top_I.branch[14].block[11].um_I.iw[15] ;
 wire \top_I.branch[14].block[11].um_I.iw[16] ;
 wire \top_I.branch[14].block[11].um_I.iw[17] ;
 wire \top_I.branch[14].block[11].um_I.iw[1] ;
 wire \top_I.branch[14].block[11].um_I.iw[2] ;
 wire \top_I.branch[14].block[11].um_I.iw[3] ;
 wire \top_I.branch[14].block[11].um_I.iw[4] ;
 wire \top_I.branch[14].block[11].um_I.iw[5] ;
 wire \top_I.branch[14].block[11].um_I.iw[6] ;
 wire \top_I.branch[14].block[11].um_I.iw[7] ;
 wire \top_I.branch[14].block[11].um_I.iw[8] ;
 wire \top_I.branch[14].block[11].um_I.iw[9] ;
 wire \top_I.branch[14].block[11].um_I.k_zero ;
 wire \top_I.branch[14].block[11].um_I.pg_vdd ;
 wire \top_I.branch[14].block[12].um_I.ana[2] ;
 wire \top_I.branch[14].block[12].um_I.ana[3] ;
 wire \top_I.branch[14].block[12].um_I.ana[4] ;
 wire \top_I.branch[14].block[12].um_I.ana[5] ;
 wire \top_I.branch[14].block[12].um_I.ana[6] ;
 wire \top_I.branch[14].block[12].um_I.ana[7] ;
 wire \top_I.branch[14].block[12].um_I.clk ;
 wire \top_I.branch[14].block[12].um_I.ena ;
 wire \top_I.branch[14].block[12].um_I.iw[10] ;
 wire \top_I.branch[14].block[12].um_I.iw[11] ;
 wire \top_I.branch[14].block[12].um_I.iw[12] ;
 wire \top_I.branch[14].block[12].um_I.iw[13] ;
 wire \top_I.branch[14].block[12].um_I.iw[14] ;
 wire \top_I.branch[14].block[12].um_I.iw[15] ;
 wire \top_I.branch[14].block[12].um_I.iw[16] ;
 wire \top_I.branch[14].block[12].um_I.iw[17] ;
 wire \top_I.branch[14].block[12].um_I.iw[1] ;
 wire \top_I.branch[14].block[12].um_I.iw[2] ;
 wire \top_I.branch[14].block[12].um_I.iw[3] ;
 wire \top_I.branch[14].block[12].um_I.iw[4] ;
 wire \top_I.branch[14].block[12].um_I.iw[5] ;
 wire \top_I.branch[14].block[12].um_I.iw[6] ;
 wire \top_I.branch[14].block[12].um_I.iw[7] ;
 wire \top_I.branch[14].block[12].um_I.iw[8] ;
 wire \top_I.branch[14].block[12].um_I.iw[9] ;
 wire \top_I.branch[14].block[12].um_I.k_zero ;
 wire \top_I.branch[14].block[12].um_I.pg_vdd ;
 wire \top_I.branch[14].block[13].um_I.ana[2] ;
 wire \top_I.branch[14].block[13].um_I.ana[3] ;
 wire \top_I.branch[14].block[13].um_I.ana[4] ;
 wire \top_I.branch[14].block[13].um_I.ana[5] ;
 wire \top_I.branch[14].block[13].um_I.ana[6] ;
 wire \top_I.branch[14].block[13].um_I.ana[7] ;
 wire \top_I.branch[14].block[13].um_I.clk ;
 wire \top_I.branch[14].block[13].um_I.ena ;
 wire \top_I.branch[14].block[13].um_I.iw[10] ;
 wire \top_I.branch[14].block[13].um_I.iw[11] ;
 wire \top_I.branch[14].block[13].um_I.iw[12] ;
 wire \top_I.branch[14].block[13].um_I.iw[13] ;
 wire \top_I.branch[14].block[13].um_I.iw[14] ;
 wire \top_I.branch[14].block[13].um_I.iw[15] ;
 wire \top_I.branch[14].block[13].um_I.iw[16] ;
 wire \top_I.branch[14].block[13].um_I.iw[17] ;
 wire \top_I.branch[14].block[13].um_I.iw[1] ;
 wire \top_I.branch[14].block[13].um_I.iw[2] ;
 wire \top_I.branch[14].block[13].um_I.iw[3] ;
 wire \top_I.branch[14].block[13].um_I.iw[4] ;
 wire \top_I.branch[14].block[13].um_I.iw[5] ;
 wire \top_I.branch[14].block[13].um_I.iw[6] ;
 wire \top_I.branch[14].block[13].um_I.iw[7] ;
 wire \top_I.branch[14].block[13].um_I.iw[8] ;
 wire \top_I.branch[14].block[13].um_I.iw[9] ;
 wire \top_I.branch[14].block[13].um_I.k_zero ;
 wire \top_I.branch[14].block[13].um_I.pg_vdd ;
 wire \top_I.branch[14].block[14].um_I.ana[2] ;
 wire \top_I.branch[14].block[14].um_I.ana[3] ;
 wire \top_I.branch[14].block[14].um_I.ana[4] ;
 wire \top_I.branch[14].block[14].um_I.ana[5] ;
 wire \top_I.branch[14].block[14].um_I.ana[6] ;
 wire \top_I.branch[14].block[14].um_I.ana[7] ;
 wire \top_I.branch[14].block[14].um_I.clk ;
 wire \top_I.branch[14].block[14].um_I.ena ;
 wire \top_I.branch[14].block[14].um_I.iw[10] ;
 wire \top_I.branch[14].block[14].um_I.iw[11] ;
 wire \top_I.branch[14].block[14].um_I.iw[12] ;
 wire \top_I.branch[14].block[14].um_I.iw[13] ;
 wire \top_I.branch[14].block[14].um_I.iw[14] ;
 wire \top_I.branch[14].block[14].um_I.iw[15] ;
 wire \top_I.branch[14].block[14].um_I.iw[16] ;
 wire \top_I.branch[14].block[14].um_I.iw[17] ;
 wire \top_I.branch[14].block[14].um_I.iw[1] ;
 wire \top_I.branch[14].block[14].um_I.iw[2] ;
 wire \top_I.branch[14].block[14].um_I.iw[3] ;
 wire \top_I.branch[14].block[14].um_I.iw[4] ;
 wire \top_I.branch[14].block[14].um_I.iw[5] ;
 wire \top_I.branch[14].block[14].um_I.iw[6] ;
 wire \top_I.branch[14].block[14].um_I.iw[7] ;
 wire \top_I.branch[14].block[14].um_I.iw[8] ;
 wire \top_I.branch[14].block[14].um_I.iw[9] ;
 wire \top_I.branch[14].block[14].um_I.k_zero ;
 wire \top_I.branch[14].block[14].um_I.pg_vdd ;
 wire \top_I.branch[14].block[15].um_I.ana[2] ;
 wire \top_I.branch[14].block[15].um_I.ana[3] ;
 wire \top_I.branch[14].block[15].um_I.ana[4] ;
 wire \top_I.branch[14].block[15].um_I.ana[5] ;
 wire \top_I.branch[14].block[15].um_I.ana[6] ;
 wire \top_I.branch[14].block[15].um_I.ana[7] ;
 wire \top_I.branch[14].block[15].um_I.clk ;
 wire \top_I.branch[14].block[15].um_I.ena ;
 wire \top_I.branch[14].block[15].um_I.iw[10] ;
 wire \top_I.branch[14].block[15].um_I.iw[11] ;
 wire \top_I.branch[14].block[15].um_I.iw[12] ;
 wire \top_I.branch[14].block[15].um_I.iw[13] ;
 wire \top_I.branch[14].block[15].um_I.iw[14] ;
 wire \top_I.branch[14].block[15].um_I.iw[15] ;
 wire \top_I.branch[14].block[15].um_I.iw[16] ;
 wire \top_I.branch[14].block[15].um_I.iw[17] ;
 wire \top_I.branch[14].block[15].um_I.iw[1] ;
 wire \top_I.branch[14].block[15].um_I.iw[2] ;
 wire \top_I.branch[14].block[15].um_I.iw[3] ;
 wire \top_I.branch[14].block[15].um_I.iw[4] ;
 wire \top_I.branch[14].block[15].um_I.iw[5] ;
 wire \top_I.branch[14].block[15].um_I.iw[6] ;
 wire \top_I.branch[14].block[15].um_I.iw[7] ;
 wire \top_I.branch[14].block[15].um_I.iw[8] ;
 wire \top_I.branch[14].block[15].um_I.iw[9] ;
 wire \top_I.branch[14].block[15].um_I.k_zero ;
 wire \top_I.branch[14].block[15].um_I.pg_vdd ;
 wire \top_I.branch[14].block[1].um_I.ana[2] ;
 wire \top_I.branch[14].block[1].um_I.ana[3] ;
 wire \top_I.branch[14].block[1].um_I.ana[4] ;
 wire \top_I.branch[14].block[1].um_I.ana[5] ;
 wire \top_I.branch[14].block[1].um_I.ana[6] ;
 wire \top_I.branch[14].block[1].um_I.ana[7] ;
 wire \top_I.branch[14].block[1].um_I.clk ;
 wire \top_I.branch[14].block[1].um_I.ena ;
 wire \top_I.branch[14].block[1].um_I.iw[10] ;
 wire \top_I.branch[14].block[1].um_I.iw[11] ;
 wire \top_I.branch[14].block[1].um_I.iw[12] ;
 wire \top_I.branch[14].block[1].um_I.iw[13] ;
 wire \top_I.branch[14].block[1].um_I.iw[14] ;
 wire \top_I.branch[14].block[1].um_I.iw[15] ;
 wire \top_I.branch[14].block[1].um_I.iw[16] ;
 wire \top_I.branch[14].block[1].um_I.iw[17] ;
 wire \top_I.branch[14].block[1].um_I.iw[1] ;
 wire \top_I.branch[14].block[1].um_I.iw[2] ;
 wire \top_I.branch[14].block[1].um_I.iw[3] ;
 wire \top_I.branch[14].block[1].um_I.iw[4] ;
 wire \top_I.branch[14].block[1].um_I.iw[5] ;
 wire \top_I.branch[14].block[1].um_I.iw[6] ;
 wire \top_I.branch[14].block[1].um_I.iw[7] ;
 wire \top_I.branch[14].block[1].um_I.iw[8] ;
 wire \top_I.branch[14].block[1].um_I.iw[9] ;
 wire \top_I.branch[14].block[1].um_I.k_zero ;
 wire \top_I.branch[14].block[1].um_I.pg_vdd ;
 wire \top_I.branch[14].block[2].um_I.ana[2] ;
 wire \top_I.branch[14].block[2].um_I.ana[3] ;
 wire \top_I.branch[14].block[2].um_I.ana[4] ;
 wire \top_I.branch[14].block[2].um_I.ana[5] ;
 wire \top_I.branch[14].block[2].um_I.ana[6] ;
 wire \top_I.branch[14].block[2].um_I.ana[7] ;
 wire \top_I.branch[14].block[2].um_I.clk ;
 wire \top_I.branch[14].block[2].um_I.ena ;
 wire \top_I.branch[14].block[2].um_I.iw[10] ;
 wire \top_I.branch[14].block[2].um_I.iw[11] ;
 wire \top_I.branch[14].block[2].um_I.iw[12] ;
 wire \top_I.branch[14].block[2].um_I.iw[13] ;
 wire \top_I.branch[14].block[2].um_I.iw[14] ;
 wire \top_I.branch[14].block[2].um_I.iw[15] ;
 wire \top_I.branch[14].block[2].um_I.iw[16] ;
 wire \top_I.branch[14].block[2].um_I.iw[17] ;
 wire \top_I.branch[14].block[2].um_I.iw[1] ;
 wire \top_I.branch[14].block[2].um_I.iw[2] ;
 wire \top_I.branch[14].block[2].um_I.iw[3] ;
 wire \top_I.branch[14].block[2].um_I.iw[4] ;
 wire \top_I.branch[14].block[2].um_I.iw[5] ;
 wire \top_I.branch[14].block[2].um_I.iw[6] ;
 wire \top_I.branch[14].block[2].um_I.iw[7] ;
 wire \top_I.branch[14].block[2].um_I.iw[8] ;
 wire \top_I.branch[14].block[2].um_I.iw[9] ;
 wire \top_I.branch[14].block[2].um_I.k_zero ;
 wire \top_I.branch[14].block[2].um_I.pg_vdd ;
 wire \top_I.branch[14].block[3].um_I.ana[2] ;
 wire \top_I.branch[14].block[3].um_I.ana[3] ;
 wire \top_I.branch[14].block[3].um_I.ana[4] ;
 wire \top_I.branch[14].block[3].um_I.ana[5] ;
 wire \top_I.branch[14].block[3].um_I.ana[6] ;
 wire \top_I.branch[14].block[3].um_I.ana[7] ;
 wire \top_I.branch[14].block[3].um_I.clk ;
 wire \top_I.branch[14].block[3].um_I.ena ;
 wire \top_I.branch[14].block[3].um_I.iw[10] ;
 wire \top_I.branch[14].block[3].um_I.iw[11] ;
 wire \top_I.branch[14].block[3].um_I.iw[12] ;
 wire \top_I.branch[14].block[3].um_I.iw[13] ;
 wire \top_I.branch[14].block[3].um_I.iw[14] ;
 wire \top_I.branch[14].block[3].um_I.iw[15] ;
 wire \top_I.branch[14].block[3].um_I.iw[16] ;
 wire \top_I.branch[14].block[3].um_I.iw[17] ;
 wire \top_I.branch[14].block[3].um_I.iw[1] ;
 wire \top_I.branch[14].block[3].um_I.iw[2] ;
 wire \top_I.branch[14].block[3].um_I.iw[3] ;
 wire \top_I.branch[14].block[3].um_I.iw[4] ;
 wire \top_I.branch[14].block[3].um_I.iw[5] ;
 wire \top_I.branch[14].block[3].um_I.iw[6] ;
 wire \top_I.branch[14].block[3].um_I.iw[7] ;
 wire \top_I.branch[14].block[3].um_I.iw[8] ;
 wire \top_I.branch[14].block[3].um_I.iw[9] ;
 wire \top_I.branch[14].block[3].um_I.k_zero ;
 wire \top_I.branch[14].block[3].um_I.pg_vdd ;
 wire \top_I.branch[14].block[4].um_I.ana[2] ;
 wire \top_I.branch[14].block[4].um_I.ana[3] ;
 wire \top_I.branch[14].block[4].um_I.ana[4] ;
 wire \top_I.branch[14].block[4].um_I.ana[5] ;
 wire \top_I.branch[14].block[4].um_I.ana[6] ;
 wire \top_I.branch[14].block[4].um_I.ana[7] ;
 wire \top_I.branch[14].block[4].um_I.clk ;
 wire \top_I.branch[14].block[4].um_I.ena ;
 wire \top_I.branch[14].block[4].um_I.iw[10] ;
 wire \top_I.branch[14].block[4].um_I.iw[11] ;
 wire \top_I.branch[14].block[4].um_I.iw[12] ;
 wire \top_I.branch[14].block[4].um_I.iw[13] ;
 wire \top_I.branch[14].block[4].um_I.iw[14] ;
 wire \top_I.branch[14].block[4].um_I.iw[15] ;
 wire \top_I.branch[14].block[4].um_I.iw[16] ;
 wire \top_I.branch[14].block[4].um_I.iw[17] ;
 wire \top_I.branch[14].block[4].um_I.iw[1] ;
 wire \top_I.branch[14].block[4].um_I.iw[2] ;
 wire \top_I.branch[14].block[4].um_I.iw[3] ;
 wire \top_I.branch[14].block[4].um_I.iw[4] ;
 wire \top_I.branch[14].block[4].um_I.iw[5] ;
 wire \top_I.branch[14].block[4].um_I.iw[6] ;
 wire \top_I.branch[14].block[4].um_I.iw[7] ;
 wire \top_I.branch[14].block[4].um_I.iw[8] ;
 wire \top_I.branch[14].block[4].um_I.iw[9] ;
 wire \top_I.branch[14].block[4].um_I.k_zero ;
 wire \top_I.branch[14].block[4].um_I.pg_vdd ;
 wire \top_I.branch[14].block[5].um_I.ana[2] ;
 wire \top_I.branch[14].block[5].um_I.ana[3] ;
 wire \top_I.branch[14].block[5].um_I.ana[4] ;
 wire \top_I.branch[14].block[5].um_I.ana[5] ;
 wire \top_I.branch[14].block[5].um_I.ana[6] ;
 wire \top_I.branch[14].block[5].um_I.ana[7] ;
 wire \top_I.branch[14].block[5].um_I.clk ;
 wire \top_I.branch[14].block[5].um_I.ena ;
 wire \top_I.branch[14].block[5].um_I.iw[10] ;
 wire \top_I.branch[14].block[5].um_I.iw[11] ;
 wire \top_I.branch[14].block[5].um_I.iw[12] ;
 wire \top_I.branch[14].block[5].um_I.iw[13] ;
 wire \top_I.branch[14].block[5].um_I.iw[14] ;
 wire \top_I.branch[14].block[5].um_I.iw[15] ;
 wire \top_I.branch[14].block[5].um_I.iw[16] ;
 wire \top_I.branch[14].block[5].um_I.iw[17] ;
 wire \top_I.branch[14].block[5].um_I.iw[1] ;
 wire \top_I.branch[14].block[5].um_I.iw[2] ;
 wire \top_I.branch[14].block[5].um_I.iw[3] ;
 wire \top_I.branch[14].block[5].um_I.iw[4] ;
 wire \top_I.branch[14].block[5].um_I.iw[5] ;
 wire \top_I.branch[14].block[5].um_I.iw[6] ;
 wire \top_I.branch[14].block[5].um_I.iw[7] ;
 wire \top_I.branch[14].block[5].um_I.iw[8] ;
 wire \top_I.branch[14].block[5].um_I.iw[9] ;
 wire \top_I.branch[14].block[5].um_I.k_zero ;
 wire \top_I.branch[14].block[5].um_I.pg_vdd ;
 wire \top_I.branch[14].block[6].um_I.ana[2] ;
 wire \top_I.branch[14].block[6].um_I.ana[3] ;
 wire \top_I.branch[14].block[6].um_I.ana[4] ;
 wire \top_I.branch[14].block[6].um_I.ana[5] ;
 wire \top_I.branch[14].block[6].um_I.ana[6] ;
 wire \top_I.branch[14].block[6].um_I.ana[7] ;
 wire \top_I.branch[14].block[6].um_I.clk ;
 wire \top_I.branch[14].block[6].um_I.ena ;
 wire \top_I.branch[14].block[6].um_I.iw[10] ;
 wire \top_I.branch[14].block[6].um_I.iw[11] ;
 wire \top_I.branch[14].block[6].um_I.iw[12] ;
 wire \top_I.branch[14].block[6].um_I.iw[13] ;
 wire \top_I.branch[14].block[6].um_I.iw[14] ;
 wire \top_I.branch[14].block[6].um_I.iw[15] ;
 wire \top_I.branch[14].block[6].um_I.iw[16] ;
 wire \top_I.branch[14].block[6].um_I.iw[17] ;
 wire \top_I.branch[14].block[6].um_I.iw[1] ;
 wire \top_I.branch[14].block[6].um_I.iw[2] ;
 wire \top_I.branch[14].block[6].um_I.iw[3] ;
 wire \top_I.branch[14].block[6].um_I.iw[4] ;
 wire \top_I.branch[14].block[6].um_I.iw[5] ;
 wire \top_I.branch[14].block[6].um_I.iw[6] ;
 wire \top_I.branch[14].block[6].um_I.iw[7] ;
 wire \top_I.branch[14].block[6].um_I.iw[8] ;
 wire \top_I.branch[14].block[6].um_I.iw[9] ;
 wire \top_I.branch[14].block[6].um_I.k_zero ;
 wire \top_I.branch[14].block[6].um_I.pg_vdd ;
 wire \top_I.branch[14].block[7].um_I.ana[2] ;
 wire \top_I.branch[14].block[7].um_I.ana[3] ;
 wire \top_I.branch[14].block[7].um_I.ana[4] ;
 wire \top_I.branch[14].block[7].um_I.ana[5] ;
 wire \top_I.branch[14].block[7].um_I.ana[6] ;
 wire \top_I.branch[14].block[7].um_I.ana[7] ;
 wire \top_I.branch[14].block[7].um_I.clk ;
 wire \top_I.branch[14].block[7].um_I.ena ;
 wire \top_I.branch[14].block[7].um_I.iw[10] ;
 wire \top_I.branch[14].block[7].um_I.iw[11] ;
 wire \top_I.branch[14].block[7].um_I.iw[12] ;
 wire \top_I.branch[14].block[7].um_I.iw[13] ;
 wire \top_I.branch[14].block[7].um_I.iw[14] ;
 wire \top_I.branch[14].block[7].um_I.iw[15] ;
 wire \top_I.branch[14].block[7].um_I.iw[16] ;
 wire \top_I.branch[14].block[7].um_I.iw[17] ;
 wire \top_I.branch[14].block[7].um_I.iw[1] ;
 wire \top_I.branch[14].block[7].um_I.iw[2] ;
 wire \top_I.branch[14].block[7].um_I.iw[3] ;
 wire \top_I.branch[14].block[7].um_I.iw[4] ;
 wire \top_I.branch[14].block[7].um_I.iw[5] ;
 wire \top_I.branch[14].block[7].um_I.iw[6] ;
 wire \top_I.branch[14].block[7].um_I.iw[7] ;
 wire \top_I.branch[14].block[7].um_I.iw[8] ;
 wire \top_I.branch[14].block[7].um_I.iw[9] ;
 wire \top_I.branch[14].block[7].um_I.k_zero ;
 wire \top_I.branch[14].block[7].um_I.pg_vdd ;
 wire \top_I.branch[14].block[8].um_I.ana[2] ;
 wire \top_I.branch[14].block[8].um_I.ana[3] ;
 wire \top_I.branch[14].block[8].um_I.ana[4] ;
 wire \top_I.branch[14].block[8].um_I.ana[5] ;
 wire \top_I.branch[14].block[8].um_I.ana[6] ;
 wire \top_I.branch[14].block[8].um_I.ana[7] ;
 wire \top_I.branch[14].block[8].um_I.clk ;
 wire \top_I.branch[14].block[8].um_I.ena ;
 wire \top_I.branch[14].block[8].um_I.iw[10] ;
 wire \top_I.branch[14].block[8].um_I.iw[11] ;
 wire \top_I.branch[14].block[8].um_I.iw[12] ;
 wire \top_I.branch[14].block[8].um_I.iw[13] ;
 wire \top_I.branch[14].block[8].um_I.iw[14] ;
 wire \top_I.branch[14].block[8].um_I.iw[15] ;
 wire \top_I.branch[14].block[8].um_I.iw[16] ;
 wire \top_I.branch[14].block[8].um_I.iw[17] ;
 wire \top_I.branch[14].block[8].um_I.iw[1] ;
 wire \top_I.branch[14].block[8].um_I.iw[2] ;
 wire \top_I.branch[14].block[8].um_I.iw[3] ;
 wire \top_I.branch[14].block[8].um_I.iw[4] ;
 wire \top_I.branch[14].block[8].um_I.iw[5] ;
 wire \top_I.branch[14].block[8].um_I.iw[6] ;
 wire \top_I.branch[14].block[8].um_I.iw[7] ;
 wire \top_I.branch[14].block[8].um_I.iw[8] ;
 wire \top_I.branch[14].block[8].um_I.iw[9] ;
 wire \top_I.branch[14].block[8].um_I.k_zero ;
 wire \top_I.branch[14].block[8].um_I.pg_vdd ;
 wire \top_I.branch[14].block[9].um_I.ana[2] ;
 wire \top_I.branch[14].block[9].um_I.ana[3] ;
 wire \top_I.branch[14].block[9].um_I.ana[4] ;
 wire \top_I.branch[14].block[9].um_I.ana[5] ;
 wire \top_I.branch[14].block[9].um_I.ana[6] ;
 wire \top_I.branch[14].block[9].um_I.ana[7] ;
 wire \top_I.branch[14].block[9].um_I.clk ;
 wire \top_I.branch[14].block[9].um_I.ena ;
 wire \top_I.branch[14].block[9].um_I.iw[10] ;
 wire \top_I.branch[14].block[9].um_I.iw[11] ;
 wire \top_I.branch[14].block[9].um_I.iw[12] ;
 wire \top_I.branch[14].block[9].um_I.iw[13] ;
 wire \top_I.branch[14].block[9].um_I.iw[14] ;
 wire \top_I.branch[14].block[9].um_I.iw[15] ;
 wire \top_I.branch[14].block[9].um_I.iw[16] ;
 wire \top_I.branch[14].block[9].um_I.iw[17] ;
 wire \top_I.branch[14].block[9].um_I.iw[1] ;
 wire \top_I.branch[14].block[9].um_I.iw[2] ;
 wire \top_I.branch[14].block[9].um_I.iw[3] ;
 wire \top_I.branch[14].block[9].um_I.iw[4] ;
 wire \top_I.branch[14].block[9].um_I.iw[5] ;
 wire \top_I.branch[14].block[9].um_I.iw[6] ;
 wire \top_I.branch[14].block[9].um_I.iw[7] ;
 wire \top_I.branch[14].block[9].um_I.iw[8] ;
 wire \top_I.branch[14].block[9].um_I.iw[9] ;
 wire \top_I.branch[14].block[9].um_I.k_zero ;
 wire \top_I.branch[14].block[9].um_I.pg_vdd ;
 wire \top_I.branch[14].l_addr[0] ;
 wire \top_I.branch[14].l_addr[3] ;
 wire \top_I.branch[15].block[0].um_I.ana[2] ;
 wire \top_I.branch[15].block[0].um_I.ana[3] ;
 wire \top_I.branch[15].block[0].um_I.ana[4] ;
 wire \top_I.branch[15].block[0].um_I.ana[5] ;
 wire \top_I.branch[15].block[0].um_I.ana[6] ;
 wire \top_I.branch[15].block[0].um_I.ana[7] ;
 wire \top_I.branch[15].block[0].um_I.clk ;
 wire \top_I.branch[15].block[0].um_I.ena ;
 wire \top_I.branch[15].block[0].um_I.iw[10] ;
 wire \top_I.branch[15].block[0].um_I.iw[11] ;
 wire \top_I.branch[15].block[0].um_I.iw[12] ;
 wire \top_I.branch[15].block[0].um_I.iw[13] ;
 wire \top_I.branch[15].block[0].um_I.iw[14] ;
 wire \top_I.branch[15].block[0].um_I.iw[15] ;
 wire \top_I.branch[15].block[0].um_I.iw[16] ;
 wire \top_I.branch[15].block[0].um_I.iw[17] ;
 wire \top_I.branch[15].block[0].um_I.iw[1] ;
 wire \top_I.branch[15].block[0].um_I.iw[2] ;
 wire \top_I.branch[15].block[0].um_I.iw[3] ;
 wire \top_I.branch[15].block[0].um_I.iw[4] ;
 wire \top_I.branch[15].block[0].um_I.iw[5] ;
 wire \top_I.branch[15].block[0].um_I.iw[6] ;
 wire \top_I.branch[15].block[0].um_I.iw[7] ;
 wire \top_I.branch[15].block[0].um_I.iw[8] ;
 wire \top_I.branch[15].block[0].um_I.iw[9] ;
 wire \top_I.branch[15].block[0].um_I.k_zero ;
 wire \top_I.branch[15].block[0].um_I.pg_vdd ;
 wire \top_I.branch[15].block[10].um_I.ana[2] ;
 wire \top_I.branch[15].block[10].um_I.ana[3] ;
 wire \top_I.branch[15].block[10].um_I.ana[4] ;
 wire \top_I.branch[15].block[10].um_I.ana[5] ;
 wire \top_I.branch[15].block[10].um_I.ana[6] ;
 wire \top_I.branch[15].block[10].um_I.ana[7] ;
 wire \top_I.branch[15].block[10].um_I.clk ;
 wire \top_I.branch[15].block[10].um_I.ena ;
 wire \top_I.branch[15].block[10].um_I.iw[10] ;
 wire \top_I.branch[15].block[10].um_I.iw[11] ;
 wire \top_I.branch[15].block[10].um_I.iw[12] ;
 wire \top_I.branch[15].block[10].um_I.iw[13] ;
 wire \top_I.branch[15].block[10].um_I.iw[14] ;
 wire \top_I.branch[15].block[10].um_I.iw[15] ;
 wire \top_I.branch[15].block[10].um_I.iw[16] ;
 wire \top_I.branch[15].block[10].um_I.iw[17] ;
 wire \top_I.branch[15].block[10].um_I.iw[1] ;
 wire \top_I.branch[15].block[10].um_I.iw[2] ;
 wire \top_I.branch[15].block[10].um_I.iw[3] ;
 wire \top_I.branch[15].block[10].um_I.iw[4] ;
 wire \top_I.branch[15].block[10].um_I.iw[5] ;
 wire \top_I.branch[15].block[10].um_I.iw[6] ;
 wire \top_I.branch[15].block[10].um_I.iw[7] ;
 wire \top_I.branch[15].block[10].um_I.iw[8] ;
 wire \top_I.branch[15].block[10].um_I.iw[9] ;
 wire \top_I.branch[15].block[10].um_I.k_zero ;
 wire \top_I.branch[15].block[10].um_I.pg_vdd ;
 wire \top_I.branch[15].block[11].um_I.ana[2] ;
 wire \top_I.branch[15].block[11].um_I.ana[3] ;
 wire \top_I.branch[15].block[11].um_I.ana[4] ;
 wire \top_I.branch[15].block[11].um_I.ana[5] ;
 wire \top_I.branch[15].block[11].um_I.ana[6] ;
 wire \top_I.branch[15].block[11].um_I.ana[7] ;
 wire \top_I.branch[15].block[11].um_I.clk ;
 wire \top_I.branch[15].block[11].um_I.ena ;
 wire \top_I.branch[15].block[11].um_I.iw[10] ;
 wire \top_I.branch[15].block[11].um_I.iw[11] ;
 wire \top_I.branch[15].block[11].um_I.iw[12] ;
 wire \top_I.branch[15].block[11].um_I.iw[13] ;
 wire \top_I.branch[15].block[11].um_I.iw[14] ;
 wire \top_I.branch[15].block[11].um_I.iw[15] ;
 wire \top_I.branch[15].block[11].um_I.iw[16] ;
 wire \top_I.branch[15].block[11].um_I.iw[17] ;
 wire \top_I.branch[15].block[11].um_I.iw[1] ;
 wire \top_I.branch[15].block[11].um_I.iw[2] ;
 wire \top_I.branch[15].block[11].um_I.iw[3] ;
 wire \top_I.branch[15].block[11].um_I.iw[4] ;
 wire \top_I.branch[15].block[11].um_I.iw[5] ;
 wire \top_I.branch[15].block[11].um_I.iw[6] ;
 wire \top_I.branch[15].block[11].um_I.iw[7] ;
 wire \top_I.branch[15].block[11].um_I.iw[8] ;
 wire \top_I.branch[15].block[11].um_I.iw[9] ;
 wire \top_I.branch[15].block[11].um_I.k_zero ;
 wire \top_I.branch[15].block[11].um_I.pg_vdd ;
 wire \top_I.branch[15].block[12].um_I.ana[2] ;
 wire \top_I.branch[15].block[12].um_I.ana[3] ;
 wire \top_I.branch[15].block[12].um_I.ana[4] ;
 wire \top_I.branch[15].block[12].um_I.ana[5] ;
 wire \top_I.branch[15].block[12].um_I.ana[6] ;
 wire \top_I.branch[15].block[12].um_I.ana[7] ;
 wire \top_I.branch[15].block[12].um_I.clk ;
 wire \top_I.branch[15].block[12].um_I.ena ;
 wire \top_I.branch[15].block[12].um_I.iw[10] ;
 wire \top_I.branch[15].block[12].um_I.iw[11] ;
 wire \top_I.branch[15].block[12].um_I.iw[12] ;
 wire \top_I.branch[15].block[12].um_I.iw[13] ;
 wire \top_I.branch[15].block[12].um_I.iw[14] ;
 wire \top_I.branch[15].block[12].um_I.iw[15] ;
 wire \top_I.branch[15].block[12].um_I.iw[16] ;
 wire \top_I.branch[15].block[12].um_I.iw[17] ;
 wire \top_I.branch[15].block[12].um_I.iw[1] ;
 wire \top_I.branch[15].block[12].um_I.iw[2] ;
 wire \top_I.branch[15].block[12].um_I.iw[3] ;
 wire \top_I.branch[15].block[12].um_I.iw[4] ;
 wire \top_I.branch[15].block[12].um_I.iw[5] ;
 wire \top_I.branch[15].block[12].um_I.iw[6] ;
 wire \top_I.branch[15].block[12].um_I.iw[7] ;
 wire \top_I.branch[15].block[12].um_I.iw[8] ;
 wire \top_I.branch[15].block[12].um_I.iw[9] ;
 wire \top_I.branch[15].block[12].um_I.k_zero ;
 wire \top_I.branch[15].block[12].um_I.pg_vdd ;
 wire \top_I.branch[15].block[13].um_I.ana[2] ;
 wire \top_I.branch[15].block[13].um_I.ana[3] ;
 wire \top_I.branch[15].block[13].um_I.ana[4] ;
 wire \top_I.branch[15].block[13].um_I.ana[5] ;
 wire \top_I.branch[15].block[13].um_I.ana[6] ;
 wire \top_I.branch[15].block[13].um_I.ana[7] ;
 wire \top_I.branch[15].block[13].um_I.clk ;
 wire \top_I.branch[15].block[13].um_I.ena ;
 wire \top_I.branch[15].block[13].um_I.iw[10] ;
 wire \top_I.branch[15].block[13].um_I.iw[11] ;
 wire \top_I.branch[15].block[13].um_I.iw[12] ;
 wire \top_I.branch[15].block[13].um_I.iw[13] ;
 wire \top_I.branch[15].block[13].um_I.iw[14] ;
 wire \top_I.branch[15].block[13].um_I.iw[15] ;
 wire \top_I.branch[15].block[13].um_I.iw[16] ;
 wire \top_I.branch[15].block[13].um_I.iw[17] ;
 wire \top_I.branch[15].block[13].um_I.iw[1] ;
 wire \top_I.branch[15].block[13].um_I.iw[2] ;
 wire \top_I.branch[15].block[13].um_I.iw[3] ;
 wire \top_I.branch[15].block[13].um_I.iw[4] ;
 wire \top_I.branch[15].block[13].um_I.iw[5] ;
 wire \top_I.branch[15].block[13].um_I.iw[6] ;
 wire \top_I.branch[15].block[13].um_I.iw[7] ;
 wire \top_I.branch[15].block[13].um_I.iw[8] ;
 wire \top_I.branch[15].block[13].um_I.iw[9] ;
 wire \top_I.branch[15].block[13].um_I.k_zero ;
 wire \top_I.branch[15].block[13].um_I.pg_vdd ;
 wire \top_I.branch[15].block[14].um_I.ana[2] ;
 wire \top_I.branch[15].block[14].um_I.ana[3] ;
 wire \top_I.branch[15].block[14].um_I.ana[4] ;
 wire \top_I.branch[15].block[14].um_I.ana[5] ;
 wire \top_I.branch[15].block[14].um_I.ana[6] ;
 wire \top_I.branch[15].block[14].um_I.ana[7] ;
 wire \top_I.branch[15].block[14].um_I.clk ;
 wire \top_I.branch[15].block[14].um_I.ena ;
 wire \top_I.branch[15].block[14].um_I.iw[10] ;
 wire \top_I.branch[15].block[14].um_I.iw[11] ;
 wire \top_I.branch[15].block[14].um_I.iw[12] ;
 wire \top_I.branch[15].block[14].um_I.iw[13] ;
 wire \top_I.branch[15].block[14].um_I.iw[14] ;
 wire \top_I.branch[15].block[14].um_I.iw[15] ;
 wire \top_I.branch[15].block[14].um_I.iw[16] ;
 wire \top_I.branch[15].block[14].um_I.iw[17] ;
 wire \top_I.branch[15].block[14].um_I.iw[1] ;
 wire \top_I.branch[15].block[14].um_I.iw[2] ;
 wire \top_I.branch[15].block[14].um_I.iw[3] ;
 wire \top_I.branch[15].block[14].um_I.iw[4] ;
 wire \top_I.branch[15].block[14].um_I.iw[5] ;
 wire \top_I.branch[15].block[14].um_I.iw[6] ;
 wire \top_I.branch[15].block[14].um_I.iw[7] ;
 wire \top_I.branch[15].block[14].um_I.iw[8] ;
 wire \top_I.branch[15].block[14].um_I.iw[9] ;
 wire \top_I.branch[15].block[14].um_I.k_zero ;
 wire \top_I.branch[15].block[14].um_I.pg_vdd ;
 wire \top_I.branch[15].block[15].um_I.ana[2] ;
 wire \top_I.branch[15].block[15].um_I.ana[3] ;
 wire \top_I.branch[15].block[15].um_I.ana[4] ;
 wire \top_I.branch[15].block[15].um_I.ana[5] ;
 wire \top_I.branch[15].block[15].um_I.ana[6] ;
 wire \top_I.branch[15].block[15].um_I.ana[7] ;
 wire \top_I.branch[15].block[15].um_I.clk ;
 wire \top_I.branch[15].block[15].um_I.ena ;
 wire \top_I.branch[15].block[15].um_I.iw[10] ;
 wire \top_I.branch[15].block[15].um_I.iw[11] ;
 wire \top_I.branch[15].block[15].um_I.iw[12] ;
 wire \top_I.branch[15].block[15].um_I.iw[13] ;
 wire \top_I.branch[15].block[15].um_I.iw[14] ;
 wire \top_I.branch[15].block[15].um_I.iw[15] ;
 wire \top_I.branch[15].block[15].um_I.iw[16] ;
 wire \top_I.branch[15].block[15].um_I.iw[17] ;
 wire \top_I.branch[15].block[15].um_I.iw[1] ;
 wire \top_I.branch[15].block[15].um_I.iw[2] ;
 wire \top_I.branch[15].block[15].um_I.iw[3] ;
 wire \top_I.branch[15].block[15].um_I.iw[4] ;
 wire \top_I.branch[15].block[15].um_I.iw[5] ;
 wire \top_I.branch[15].block[15].um_I.iw[6] ;
 wire \top_I.branch[15].block[15].um_I.iw[7] ;
 wire \top_I.branch[15].block[15].um_I.iw[8] ;
 wire \top_I.branch[15].block[15].um_I.iw[9] ;
 wire \top_I.branch[15].block[15].um_I.k_zero ;
 wire \top_I.branch[15].block[15].um_I.pg_vdd ;
 wire \top_I.branch[15].block[1].um_I.ana[2] ;
 wire \top_I.branch[15].block[1].um_I.ana[3] ;
 wire \top_I.branch[15].block[1].um_I.ana[4] ;
 wire \top_I.branch[15].block[1].um_I.ana[5] ;
 wire \top_I.branch[15].block[1].um_I.ana[6] ;
 wire \top_I.branch[15].block[1].um_I.ana[7] ;
 wire \top_I.branch[15].block[1].um_I.clk ;
 wire \top_I.branch[15].block[1].um_I.ena ;
 wire \top_I.branch[15].block[1].um_I.iw[10] ;
 wire \top_I.branch[15].block[1].um_I.iw[11] ;
 wire \top_I.branch[15].block[1].um_I.iw[12] ;
 wire \top_I.branch[15].block[1].um_I.iw[13] ;
 wire \top_I.branch[15].block[1].um_I.iw[14] ;
 wire \top_I.branch[15].block[1].um_I.iw[15] ;
 wire \top_I.branch[15].block[1].um_I.iw[16] ;
 wire \top_I.branch[15].block[1].um_I.iw[17] ;
 wire \top_I.branch[15].block[1].um_I.iw[1] ;
 wire \top_I.branch[15].block[1].um_I.iw[2] ;
 wire \top_I.branch[15].block[1].um_I.iw[3] ;
 wire \top_I.branch[15].block[1].um_I.iw[4] ;
 wire \top_I.branch[15].block[1].um_I.iw[5] ;
 wire \top_I.branch[15].block[1].um_I.iw[6] ;
 wire \top_I.branch[15].block[1].um_I.iw[7] ;
 wire \top_I.branch[15].block[1].um_I.iw[8] ;
 wire \top_I.branch[15].block[1].um_I.iw[9] ;
 wire \top_I.branch[15].block[1].um_I.k_zero ;
 wire \top_I.branch[15].block[1].um_I.pg_vdd ;
 wire \top_I.branch[15].block[2].um_I.ana[2] ;
 wire \top_I.branch[15].block[2].um_I.ana[3] ;
 wire \top_I.branch[15].block[2].um_I.ana[4] ;
 wire \top_I.branch[15].block[2].um_I.ana[5] ;
 wire \top_I.branch[15].block[2].um_I.ana[6] ;
 wire \top_I.branch[15].block[2].um_I.ana[7] ;
 wire \top_I.branch[15].block[2].um_I.clk ;
 wire \top_I.branch[15].block[2].um_I.ena ;
 wire \top_I.branch[15].block[2].um_I.iw[10] ;
 wire \top_I.branch[15].block[2].um_I.iw[11] ;
 wire \top_I.branch[15].block[2].um_I.iw[12] ;
 wire \top_I.branch[15].block[2].um_I.iw[13] ;
 wire \top_I.branch[15].block[2].um_I.iw[14] ;
 wire \top_I.branch[15].block[2].um_I.iw[15] ;
 wire \top_I.branch[15].block[2].um_I.iw[16] ;
 wire \top_I.branch[15].block[2].um_I.iw[17] ;
 wire \top_I.branch[15].block[2].um_I.iw[1] ;
 wire \top_I.branch[15].block[2].um_I.iw[2] ;
 wire \top_I.branch[15].block[2].um_I.iw[3] ;
 wire \top_I.branch[15].block[2].um_I.iw[4] ;
 wire \top_I.branch[15].block[2].um_I.iw[5] ;
 wire \top_I.branch[15].block[2].um_I.iw[6] ;
 wire \top_I.branch[15].block[2].um_I.iw[7] ;
 wire \top_I.branch[15].block[2].um_I.iw[8] ;
 wire \top_I.branch[15].block[2].um_I.iw[9] ;
 wire \top_I.branch[15].block[2].um_I.k_zero ;
 wire \top_I.branch[15].block[2].um_I.pg_vdd ;
 wire \top_I.branch[15].block[3].um_I.ana[2] ;
 wire \top_I.branch[15].block[3].um_I.ana[3] ;
 wire \top_I.branch[15].block[3].um_I.ana[4] ;
 wire \top_I.branch[15].block[3].um_I.ana[5] ;
 wire \top_I.branch[15].block[3].um_I.ana[6] ;
 wire \top_I.branch[15].block[3].um_I.ana[7] ;
 wire \top_I.branch[15].block[3].um_I.clk ;
 wire \top_I.branch[15].block[3].um_I.ena ;
 wire \top_I.branch[15].block[3].um_I.iw[10] ;
 wire \top_I.branch[15].block[3].um_I.iw[11] ;
 wire \top_I.branch[15].block[3].um_I.iw[12] ;
 wire \top_I.branch[15].block[3].um_I.iw[13] ;
 wire \top_I.branch[15].block[3].um_I.iw[14] ;
 wire \top_I.branch[15].block[3].um_I.iw[15] ;
 wire \top_I.branch[15].block[3].um_I.iw[16] ;
 wire \top_I.branch[15].block[3].um_I.iw[17] ;
 wire \top_I.branch[15].block[3].um_I.iw[1] ;
 wire \top_I.branch[15].block[3].um_I.iw[2] ;
 wire \top_I.branch[15].block[3].um_I.iw[3] ;
 wire \top_I.branch[15].block[3].um_I.iw[4] ;
 wire \top_I.branch[15].block[3].um_I.iw[5] ;
 wire \top_I.branch[15].block[3].um_I.iw[6] ;
 wire \top_I.branch[15].block[3].um_I.iw[7] ;
 wire \top_I.branch[15].block[3].um_I.iw[8] ;
 wire \top_I.branch[15].block[3].um_I.iw[9] ;
 wire \top_I.branch[15].block[3].um_I.k_zero ;
 wire \top_I.branch[15].block[3].um_I.pg_vdd ;
 wire \top_I.branch[15].block[4].um_I.ana[2] ;
 wire \top_I.branch[15].block[4].um_I.ana[3] ;
 wire \top_I.branch[15].block[4].um_I.ana[4] ;
 wire \top_I.branch[15].block[4].um_I.ana[5] ;
 wire \top_I.branch[15].block[4].um_I.ana[6] ;
 wire \top_I.branch[15].block[4].um_I.ana[7] ;
 wire \top_I.branch[15].block[4].um_I.clk ;
 wire \top_I.branch[15].block[4].um_I.ena ;
 wire \top_I.branch[15].block[4].um_I.iw[10] ;
 wire \top_I.branch[15].block[4].um_I.iw[11] ;
 wire \top_I.branch[15].block[4].um_I.iw[12] ;
 wire \top_I.branch[15].block[4].um_I.iw[13] ;
 wire \top_I.branch[15].block[4].um_I.iw[14] ;
 wire \top_I.branch[15].block[4].um_I.iw[15] ;
 wire \top_I.branch[15].block[4].um_I.iw[16] ;
 wire \top_I.branch[15].block[4].um_I.iw[17] ;
 wire \top_I.branch[15].block[4].um_I.iw[1] ;
 wire \top_I.branch[15].block[4].um_I.iw[2] ;
 wire \top_I.branch[15].block[4].um_I.iw[3] ;
 wire \top_I.branch[15].block[4].um_I.iw[4] ;
 wire \top_I.branch[15].block[4].um_I.iw[5] ;
 wire \top_I.branch[15].block[4].um_I.iw[6] ;
 wire \top_I.branch[15].block[4].um_I.iw[7] ;
 wire \top_I.branch[15].block[4].um_I.iw[8] ;
 wire \top_I.branch[15].block[4].um_I.iw[9] ;
 wire \top_I.branch[15].block[4].um_I.k_zero ;
 wire \top_I.branch[15].block[4].um_I.pg_vdd ;
 wire \top_I.branch[15].block[5].um_I.ana[2] ;
 wire \top_I.branch[15].block[5].um_I.ana[3] ;
 wire \top_I.branch[15].block[5].um_I.ana[4] ;
 wire \top_I.branch[15].block[5].um_I.ana[5] ;
 wire \top_I.branch[15].block[5].um_I.ana[6] ;
 wire \top_I.branch[15].block[5].um_I.ana[7] ;
 wire \top_I.branch[15].block[5].um_I.clk ;
 wire \top_I.branch[15].block[5].um_I.ena ;
 wire \top_I.branch[15].block[5].um_I.iw[10] ;
 wire \top_I.branch[15].block[5].um_I.iw[11] ;
 wire \top_I.branch[15].block[5].um_I.iw[12] ;
 wire \top_I.branch[15].block[5].um_I.iw[13] ;
 wire \top_I.branch[15].block[5].um_I.iw[14] ;
 wire \top_I.branch[15].block[5].um_I.iw[15] ;
 wire \top_I.branch[15].block[5].um_I.iw[16] ;
 wire \top_I.branch[15].block[5].um_I.iw[17] ;
 wire \top_I.branch[15].block[5].um_I.iw[1] ;
 wire \top_I.branch[15].block[5].um_I.iw[2] ;
 wire \top_I.branch[15].block[5].um_I.iw[3] ;
 wire \top_I.branch[15].block[5].um_I.iw[4] ;
 wire \top_I.branch[15].block[5].um_I.iw[5] ;
 wire \top_I.branch[15].block[5].um_I.iw[6] ;
 wire \top_I.branch[15].block[5].um_I.iw[7] ;
 wire \top_I.branch[15].block[5].um_I.iw[8] ;
 wire \top_I.branch[15].block[5].um_I.iw[9] ;
 wire \top_I.branch[15].block[5].um_I.k_zero ;
 wire \top_I.branch[15].block[5].um_I.pg_vdd ;
 wire \top_I.branch[15].block[6].um_I.ana[2] ;
 wire \top_I.branch[15].block[6].um_I.ana[3] ;
 wire \top_I.branch[15].block[6].um_I.ana[4] ;
 wire \top_I.branch[15].block[6].um_I.ana[5] ;
 wire \top_I.branch[15].block[6].um_I.ana[6] ;
 wire \top_I.branch[15].block[6].um_I.ana[7] ;
 wire \top_I.branch[15].block[6].um_I.clk ;
 wire \top_I.branch[15].block[6].um_I.ena ;
 wire \top_I.branch[15].block[6].um_I.iw[10] ;
 wire \top_I.branch[15].block[6].um_I.iw[11] ;
 wire \top_I.branch[15].block[6].um_I.iw[12] ;
 wire \top_I.branch[15].block[6].um_I.iw[13] ;
 wire \top_I.branch[15].block[6].um_I.iw[14] ;
 wire \top_I.branch[15].block[6].um_I.iw[15] ;
 wire \top_I.branch[15].block[6].um_I.iw[16] ;
 wire \top_I.branch[15].block[6].um_I.iw[17] ;
 wire \top_I.branch[15].block[6].um_I.iw[1] ;
 wire \top_I.branch[15].block[6].um_I.iw[2] ;
 wire \top_I.branch[15].block[6].um_I.iw[3] ;
 wire \top_I.branch[15].block[6].um_I.iw[4] ;
 wire \top_I.branch[15].block[6].um_I.iw[5] ;
 wire \top_I.branch[15].block[6].um_I.iw[6] ;
 wire \top_I.branch[15].block[6].um_I.iw[7] ;
 wire \top_I.branch[15].block[6].um_I.iw[8] ;
 wire \top_I.branch[15].block[6].um_I.iw[9] ;
 wire \top_I.branch[15].block[6].um_I.k_zero ;
 wire \top_I.branch[15].block[6].um_I.pg_vdd ;
 wire \top_I.branch[15].block[7].um_I.ana[2] ;
 wire \top_I.branch[15].block[7].um_I.ana[3] ;
 wire \top_I.branch[15].block[7].um_I.ana[4] ;
 wire \top_I.branch[15].block[7].um_I.ana[5] ;
 wire \top_I.branch[15].block[7].um_I.ana[6] ;
 wire \top_I.branch[15].block[7].um_I.ana[7] ;
 wire \top_I.branch[15].block[7].um_I.clk ;
 wire \top_I.branch[15].block[7].um_I.ena ;
 wire \top_I.branch[15].block[7].um_I.iw[10] ;
 wire \top_I.branch[15].block[7].um_I.iw[11] ;
 wire \top_I.branch[15].block[7].um_I.iw[12] ;
 wire \top_I.branch[15].block[7].um_I.iw[13] ;
 wire \top_I.branch[15].block[7].um_I.iw[14] ;
 wire \top_I.branch[15].block[7].um_I.iw[15] ;
 wire \top_I.branch[15].block[7].um_I.iw[16] ;
 wire \top_I.branch[15].block[7].um_I.iw[17] ;
 wire \top_I.branch[15].block[7].um_I.iw[1] ;
 wire \top_I.branch[15].block[7].um_I.iw[2] ;
 wire \top_I.branch[15].block[7].um_I.iw[3] ;
 wire \top_I.branch[15].block[7].um_I.iw[4] ;
 wire \top_I.branch[15].block[7].um_I.iw[5] ;
 wire \top_I.branch[15].block[7].um_I.iw[6] ;
 wire \top_I.branch[15].block[7].um_I.iw[7] ;
 wire \top_I.branch[15].block[7].um_I.iw[8] ;
 wire \top_I.branch[15].block[7].um_I.iw[9] ;
 wire \top_I.branch[15].block[7].um_I.k_zero ;
 wire \top_I.branch[15].block[7].um_I.pg_vdd ;
 wire \top_I.branch[15].block[8].um_I.ana[2] ;
 wire \top_I.branch[15].block[8].um_I.ana[3] ;
 wire \top_I.branch[15].block[8].um_I.ana[4] ;
 wire \top_I.branch[15].block[8].um_I.ana[5] ;
 wire \top_I.branch[15].block[8].um_I.ana[6] ;
 wire \top_I.branch[15].block[8].um_I.ana[7] ;
 wire \top_I.branch[15].block[8].um_I.clk ;
 wire \top_I.branch[15].block[8].um_I.ena ;
 wire \top_I.branch[15].block[8].um_I.iw[10] ;
 wire \top_I.branch[15].block[8].um_I.iw[11] ;
 wire \top_I.branch[15].block[8].um_I.iw[12] ;
 wire \top_I.branch[15].block[8].um_I.iw[13] ;
 wire \top_I.branch[15].block[8].um_I.iw[14] ;
 wire \top_I.branch[15].block[8].um_I.iw[15] ;
 wire \top_I.branch[15].block[8].um_I.iw[16] ;
 wire \top_I.branch[15].block[8].um_I.iw[17] ;
 wire \top_I.branch[15].block[8].um_I.iw[1] ;
 wire \top_I.branch[15].block[8].um_I.iw[2] ;
 wire \top_I.branch[15].block[8].um_I.iw[3] ;
 wire \top_I.branch[15].block[8].um_I.iw[4] ;
 wire \top_I.branch[15].block[8].um_I.iw[5] ;
 wire \top_I.branch[15].block[8].um_I.iw[6] ;
 wire \top_I.branch[15].block[8].um_I.iw[7] ;
 wire \top_I.branch[15].block[8].um_I.iw[8] ;
 wire \top_I.branch[15].block[8].um_I.iw[9] ;
 wire \top_I.branch[15].block[8].um_I.k_zero ;
 wire \top_I.branch[15].block[8].um_I.pg_vdd ;
 wire \top_I.branch[15].block[9].um_I.ana[2] ;
 wire \top_I.branch[15].block[9].um_I.ana[3] ;
 wire \top_I.branch[15].block[9].um_I.ana[4] ;
 wire \top_I.branch[15].block[9].um_I.ana[5] ;
 wire \top_I.branch[15].block[9].um_I.ana[6] ;
 wire \top_I.branch[15].block[9].um_I.ana[7] ;
 wire \top_I.branch[15].block[9].um_I.clk ;
 wire \top_I.branch[15].block[9].um_I.ena ;
 wire \top_I.branch[15].block[9].um_I.iw[10] ;
 wire \top_I.branch[15].block[9].um_I.iw[11] ;
 wire \top_I.branch[15].block[9].um_I.iw[12] ;
 wire \top_I.branch[15].block[9].um_I.iw[13] ;
 wire \top_I.branch[15].block[9].um_I.iw[14] ;
 wire \top_I.branch[15].block[9].um_I.iw[15] ;
 wire \top_I.branch[15].block[9].um_I.iw[16] ;
 wire \top_I.branch[15].block[9].um_I.iw[17] ;
 wire \top_I.branch[15].block[9].um_I.iw[1] ;
 wire \top_I.branch[15].block[9].um_I.iw[2] ;
 wire \top_I.branch[15].block[9].um_I.iw[3] ;
 wire \top_I.branch[15].block[9].um_I.iw[4] ;
 wire \top_I.branch[15].block[9].um_I.iw[5] ;
 wire \top_I.branch[15].block[9].um_I.iw[6] ;
 wire \top_I.branch[15].block[9].um_I.iw[7] ;
 wire \top_I.branch[15].block[9].um_I.iw[8] ;
 wire \top_I.branch[15].block[9].um_I.iw[9] ;
 wire \top_I.branch[15].block[9].um_I.k_zero ;
 wire \top_I.branch[15].block[9].um_I.pg_vdd ;
 wire \top_I.branch[15].l_addr[0] ;
 wire \top_I.branch[15].l_addr[3] ;
 wire \top_I.branch[16].block[0].um_I.ana[2] ;
 wire \top_I.branch[16].block[0].um_I.ana[3] ;
 wire \top_I.branch[16].block[0].um_I.ana[4] ;
 wire \top_I.branch[16].block[0].um_I.ana[5] ;
 wire \top_I.branch[16].block[0].um_I.ana[6] ;
 wire \top_I.branch[16].block[0].um_I.ana[7] ;
 wire \top_I.branch[16].block[0].um_I.clk ;
 wire \top_I.branch[16].block[0].um_I.ena ;
 wire \top_I.branch[16].block[0].um_I.iw[10] ;
 wire \top_I.branch[16].block[0].um_I.iw[11] ;
 wire \top_I.branch[16].block[0].um_I.iw[12] ;
 wire \top_I.branch[16].block[0].um_I.iw[13] ;
 wire \top_I.branch[16].block[0].um_I.iw[14] ;
 wire \top_I.branch[16].block[0].um_I.iw[15] ;
 wire \top_I.branch[16].block[0].um_I.iw[16] ;
 wire \top_I.branch[16].block[0].um_I.iw[17] ;
 wire \top_I.branch[16].block[0].um_I.iw[1] ;
 wire \top_I.branch[16].block[0].um_I.iw[2] ;
 wire \top_I.branch[16].block[0].um_I.iw[3] ;
 wire \top_I.branch[16].block[0].um_I.iw[4] ;
 wire \top_I.branch[16].block[0].um_I.iw[5] ;
 wire \top_I.branch[16].block[0].um_I.iw[6] ;
 wire \top_I.branch[16].block[0].um_I.iw[7] ;
 wire \top_I.branch[16].block[0].um_I.iw[8] ;
 wire \top_I.branch[16].block[0].um_I.iw[9] ;
 wire \top_I.branch[16].block[0].um_I.k_zero ;
 wire \top_I.branch[16].block[0].um_I.pg_vdd ;
 wire \top_I.branch[16].block[10].um_I.ana[2] ;
 wire \top_I.branch[16].block[10].um_I.ana[3] ;
 wire \top_I.branch[16].block[10].um_I.ana[4] ;
 wire \top_I.branch[16].block[10].um_I.ana[5] ;
 wire \top_I.branch[16].block[10].um_I.ana[6] ;
 wire \top_I.branch[16].block[10].um_I.ana[7] ;
 wire \top_I.branch[16].block[10].um_I.clk ;
 wire \top_I.branch[16].block[10].um_I.ena ;
 wire \top_I.branch[16].block[10].um_I.iw[10] ;
 wire \top_I.branch[16].block[10].um_I.iw[11] ;
 wire \top_I.branch[16].block[10].um_I.iw[12] ;
 wire \top_I.branch[16].block[10].um_I.iw[13] ;
 wire \top_I.branch[16].block[10].um_I.iw[14] ;
 wire \top_I.branch[16].block[10].um_I.iw[15] ;
 wire \top_I.branch[16].block[10].um_I.iw[16] ;
 wire \top_I.branch[16].block[10].um_I.iw[17] ;
 wire \top_I.branch[16].block[10].um_I.iw[1] ;
 wire \top_I.branch[16].block[10].um_I.iw[2] ;
 wire \top_I.branch[16].block[10].um_I.iw[3] ;
 wire \top_I.branch[16].block[10].um_I.iw[4] ;
 wire \top_I.branch[16].block[10].um_I.iw[5] ;
 wire \top_I.branch[16].block[10].um_I.iw[6] ;
 wire \top_I.branch[16].block[10].um_I.iw[7] ;
 wire \top_I.branch[16].block[10].um_I.iw[8] ;
 wire \top_I.branch[16].block[10].um_I.iw[9] ;
 wire \top_I.branch[16].block[10].um_I.k_zero ;
 wire \top_I.branch[16].block[10].um_I.pg_vdd ;
 wire \top_I.branch[16].block[11].um_I.ana[2] ;
 wire \top_I.branch[16].block[11].um_I.ana[3] ;
 wire \top_I.branch[16].block[11].um_I.ana[4] ;
 wire \top_I.branch[16].block[11].um_I.ana[5] ;
 wire \top_I.branch[16].block[11].um_I.ana[6] ;
 wire \top_I.branch[16].block[11].um_I.ana[7] ;
 wire \top_I.branch[16].block[11].um_I.clk ;
 wire \top_I.branch[16].block[11].um_I.ena ;
 wire \top_I.branch[16].block[11].um_I.iw[10] ;
 wire \top_I.branch[16].block[11].um_I.iw[11] ;
 wire \top_I.branch[16].block[11].um_I.iw[12] ;
 wire \top_I.branch[16].block[11].um_I.iw[13] ;
 wire \top_I.branch[16].block[11].um_I.iw[14] ;
 wire \top_I.branch[16].block[11].um_I.iw[15] ;
 wire \top_I.branch[16].block[11].um_I.iw[16] ;
 wire \top_I.branch[16].block[11].um_I.iw[17] ;
 wire \top_I.branch[16].block[11].um_I.iw[1] ;
 wire \top_I.branch[16].block[11].um_I.iw[2] ;
 wire \top_I.branch[16].block[11].um_I.iw[3] ;
 wire \top_I.branch[16].block[11].um_I.iw[4] ;
 wire \top_I.branch[16].block[11].um_I.iw[5] ;
 wire \top_I.branch[16].block[11].um_I.iw[6] ;
 wire \top_I.branch[16].block[11].um_I.iw[7] ;
 wire \top_I.branch[16].block[11].um_I.iw[8] ;
 wire \top_I.branch[16].block[11].um_I.iw[9] ;
 wire \top_I.branch[16].block[11].um_I.k_zero ;
 wire \top_I.branch[16].block[11].um_I.pg_vdd ;
 wire \top_I.branch[16].block[12].um_I.ana[2] ;
 wire \top_I.branch[16].block[12].um_I.ana[3] ;
 wire \top_I.branch[16].block[12].um_I.ana[4] ;
 wire \top_I.branch[16].block[12].um_I.ana[5] ;
 wire \top_I.branch[16].block[12].um_I.ana[6] ;
 wire \top_I.branch[16].block[12].um_I.ana[7] ;
 wire \top_I.branch[16].block[12].um_I.clk ;
 wire \top_I.branch[16].block[12].um_I.ena ;
 wire \top_I.branch[16].block[12].um_I.iw[10] ;
 wire \top_I.branch[16].block[12].um_I.iw[11] ;
 wire \top_I.branch[16].block[12].um_I.iw[12] ;
 wire \top_I.branch[16].block[12].um_I.iw[13] ;
 wire \top_I.branch[16].block[12].um_I.iw[14] ;
 wire \top_I.branch[16].block[12].um_I.iw[15] ;
 wire \top_I.branch[16].block[12].um_I.iw[16] ;
 wire \top_I.branch[16].block[12].um_I.iw[17] ;
 wire \top_I.branch[16].block[12].um_I.iw[1] ;
 wire \top_I.branch[16].block[12].um_I.iw[2] ;
 wire \top_I.branch[16].block[12].um_I.iw[3] ;
 wire \top_I.branch[16].block[12].um_I.iw[4] ;
 wire \top_I.branch[16].block[12].um_I.iw[5] ;
 wire \top_I.branch[16].block[12].um_I.iw[6] ;
 wire \top_I.branch[16].block[12].um_I.iw[7] ;
 wire \top_I.branch[16].block[12].um_I.iw[8] ;
 wire \top_I.branch[16].block[12].um_I.iw[9] ;
 wire \top_I.branch[16].block[12].um_I.k_zero ;
 wire \top_I.branch[16].block[12].um_I.pg_vdd ;
 wire \top_I.branch[16].block[13].um_I.ana[2] ;
 wire \top_I.branch[16].block[13].um_I.ana[3] ;
 wire \top_I.branch[16].block[13].um_I.ana[4] ;
 wire \top_I.branch[16].block[13].um_I.ana[5] ;
 wire \top_I.branch[16].block[13].um_I.ana[6] ;
 wire \top_I.branch[16].block[13].um_I.ana[7] ;
 wire \top_I.branch[16].block[13].um_I.clk ;
 wire \top_I.branch[16].block[13].um_I.ena ;
 wire \top_I.branch[16].block[13].um_I.iw[10] ;
 wire \top_I.branch[16].block[13].um_I.iw[11] ;
 wire \top_I.branch[16].block[13].um_I.iw[12] ;
 wire \top_I.branch[16].block[13].um_I.iw[13] ;
 wire \top_I.branch[16].block[13].um_I.iw[14] ;
 wire \top_I.branch[16].block[13].um_I.iw[15] ;
 wire \top_I.branch[16].block[13].um_I.iw[16] ;
 wire \top_I.branch[16].block[13].um_I.iw[17] ;
 wire \top_I.branch[16].block[13].um_I.iw[1] ;
 wire \top_I.branch[16].block[13].um_I.iw[2] ;
 wire \top_I.branch[16].block[13].um_I.iw[3] ;
 wire \top_I.branch[16].block[13].um_I.iw[4] ;
 wire \top_I.branch[16].block[13].um_I.iw[5] ;
 wire \top_I.branch[16].block[13].um_I.iw[6] ;
 wire \top_I.branch[16].block[13].um_I.iw[7] ;
 wire \top_I.branch[16].block[13].um_I.iw[8] ;
 wire \top_I.branch[16].block[13].um_I.iw[9] ;
 wire \top_I.branch[16].block[13].um_I.k_zero ;
 wire \top_I.branch[16].block[13].um_I.pg_vdd ;
 wire \top_I.branch[16].block[14].um_I.ana[2] ;
 wire \top_I.branch[16].block[14].um_I.ana[3] ;
 wire \top_I.branch[16].block[14].um_I.ana[4] ;
 wire \top_I.branch[16].block[14].um_I.ana[5] ;
 wire \top_I.branch[16].block[14].um_I.ana[6] ;
 wire \top_I.branch[16].block[14].um_I.ana[7] ;
 wire \top_I.branch[16].block[14].um_I.clk ;
 wire \top_I.branch[16].block[14].um_I.ena ;
 wire \top_I.branch[16].block[14].um_I.iw[10] ;
 wire \top_I.branch[16].block[14].um_I.iw[11] ;
 wire \top_I.branch[16].block[14].um_I.iw[12] ;
 wire \top_I.branch[16].block[14].um_I.iw[13] ;
 wire \top_I.branch[16].block[14].um_I.iw[14] ;
 wire \top_I.branch[16].block[14].um_I.iw[15] ;
 wire \top_I.branch[16].block[14].um_I.iw[16] ;
 wire \top_I.branch[16].block[14].um_I.iw[17] ;
 wire \top_I.branch[16].block[14].um_I.iw[1] ;
 wire \top_I.branch[16].block[14].um_I.iw[2] ;
 wire \top_I.branch[16].block[14].um_I.iw[3] ;
 wire \top_I.branch[16].block[14].um_I.iw[4] ;
 wire \top_I.branch[16].block[14].um_I.iw[5] ;
 wire \top_I.branch[16].block[14].um_I.iw[6] ;
 wire \top_I.branch[16].block[14].um_I.iw[7] ;
 wire \top_I.branch[16].block[14].um_I.iw[8] ;
 wire \top_I.branch[16].block[14].um_I.iw[9] ;
 wire \top_I.branch[16].block[14].um_I.k_zero ;
 wire \top_I.branch[16].block[14].um_I.pg_vdd ;
 wire \top_I.branch[16].block[15].um_I.ana[2] ;
 wire \top_I.branch[16].block[15].um_I.ana[3] ;
 wire \top_I.branch[16].block[15].um_I.ana[4] ;
 wire \top_I.branch[16].block[15].um_I.ana[5] ;
 wire \top_I.branch[16].block[15].um_I.ana[6] ;
 wire \top_I.branch[16].block[15].um_I.ana[7] ;
 wire \top_I.branch[16].block[15].um_I.clk ;
 wire \top_I.branch[16].block[15].um_I.ena ;
 wire \top_I.branch[16].block[15].um_I.iw[10] ;
 wire \top_I.branch[16].block[15].um_I.iw[11] ;
 wire \top_I.branch[16].block[15].um_I.iw[12] ;
 wire \top_I.branch[16].block[15].um_I.iw[13] ;
 wire \top_I.branch[16].block[15].um_I.iw[14] ;
 wire \top_I.branch[16].block[15].um_I.iw[15] ;
 wire \top_I.branch[16].block[15].um_I.iw[16] ;
 wire \top_I.branch[16].block[15].um_I.iw[17] ;
 wire \top_I.branch[16].block[15].um_I.iw[1] ;
 wire \top_I.branch[16].block[15].um_I.iw[2] ;
 wire \top_I.branch[16].block[15].um_I.iw[3] ;
 wire \top_I.branch[16].block[15].um_I.iw[4] ;
 wire \top_I.branch[16].block[15].um_I.iw[5] ;
 wire \top_I.branch[16].block[15].um_I.iw[6] ;
 wire \top_I.branch[16].block[15].um_I.iw[7] ;
 wire \top_I.branch[16].block[15].um_I.iw[8] ;
 wire \top_I.branch[16].block[15].um_I.iw[9] ;
 wire \top_I.branch[16].block[15].um_I.k_zero ;
 wire \top_I.branch[16].block[15].um_I.pg_vdd ;
 wire \top_I.branch[16].block[1].um_I.ana[2] ;
 wire \top_I.branch[16].block[1].um_I.ana[3] ;
 wire \top_I.branch[16].block[1].um_I.ana[4] ;
 wire \top_I.branch[16].block[1].um_I.ana[5] ;
 wire \top_I.branch[16].block[1].um_I.ana[6] ;
 wire \top_I.branch[16].block[1].um_I.ana[7] ;
 wire \top_I.branch[16].block[1].um_I.clk ;
 wire \top_I.branch[16].block[1].um_I.ena ;
 wire \top_I.branch[16].block[1].um_I.iw[10] ;
 wire \top_I.branch[16].block[1].um_I.iw[11] ;
 wire \top_I.branch[16].block[1].um_I.iw[12] ;
 wire \top_I.branch[16].block[1].um_I.iw[13] ;
 wire \top_I.branch[16].block[1].um_I.iw[14] ;
 wire \top_I.branch[16].block[1].um_I.iw[15] ;
 wire \top_I.branch[16].block[1].um_I.iw[16] ;
 wire \top_I.branch[16].block[1].um_I.iw[17] ;
 wire \top_I.branch[16].block[1].um_I.iw[1] ;
 wire \top_I.branch[16].block[1].um_I.iw[2] ;
 wire \top_I.branch[16].block[1].um_I.iw[3] ;
 wire \top_I.branch[16].block[1].um_I.iw[4] ;
 wire \top_I.branch[16].block[1].um_I.iw[5] ;
 wire \top_I.branch[16].block[1].um_I.iw[6] ;
 wire \top_I.branch[16].block[1].um_I.iw[7] ;
 wire \top_I.branch[16].block[1].um_I.iw[8] ;
 wire \top_I.branch[16].block[1].um_I.iw[9] ;
 wire \top_I.branch[16].block[1].um_I.k_zero ;
 wire \top_I.branch[16].block[1].um_I.pg_vdd ;
 wire \top_I.branch[16].block[2].um_I.ana[2] ;
 wire \top_I.branch[16].block[2].um_I.ana[3] ;
 wire \top_I.branch[16].block[2].um_I.ana[4] ;
 wire \top_I.branch[16].block[2].um_I.ana[5] ;
 wire \top_I.branch[16].block[2].um_I.ana[6] ;
 wire \top_I.branch[16].block[2].um_I.ana[7] ;
 wire \top_I.branch[16].block[2].um_I.clk ;
 wire \top_I.branch[16].block[2].um_I.ena ;
 wire \top_I.branch[16].block[2].um_I.iw[10] ;
 wire \top_I.branch[16].block[2].um_I.iw[11] ;
 wire \top_I.branch[16].block[2].um_I.iw[12] ;
 wire \top_I.branch[16].block[2].um_I.iw[13] ;
 wire \top_I.branch[16].block[2].um_I.iw[14] ;
 wire \top_I.branch[16].block[2].um_I.iw[15] ;
 wire \top_I.branch[16].block[2].um_I.iw[16] ;
 wire \top_I.branch[16].block[2].um_I.iw[17] ;
 wire \top_I.branch[16].block[2].um_I.iw[1] ;
 wire \top_I.branch[16].block[2].um_I.iw[2] ;
 wire \top_I.branch[16].block[2].um_I.iw[3] ;
 wire \top_I.branch[16].block[2].um_I.iw[4] ;
 wire \top_I.branch[16].block[2].um_I.iw[5] ;
 wire \top_I.branch[16].block[2].um_I.iw[6] ;
 wire \top_I.branch[16].block[2].um_I.iw[7] ;
 wire \top_I.branch[16].block[2].um_I.iw[8] ;
 wire \top_I.branch[16].block[2].um_I.iw[9] ;
 wire \top_I.branch[16].block[2].um_I.k_zero ;
 wire \top_I.branch[16].block[2].um_I.pg_vdd ;
 wire \top_I.branch[16].block[3].um_I.ana[2] ;
 wire \top_I.branch[16].block[3].um_I.ana[3] ;
 wire \top_I.branch[16].block[3].um_I.ana[4] ;
 wire \top_I.branch[16].block[3].um_I.ana[5] ;
 wire \top_I.branch[16].block[3].um_I.ana[6] ;
 wire \top_I.branch[16].block[3].um_I.ana[7] ;
 wire \top_I.branch[16].block[3].um_I.clk ;
 wire \top_I.branch[16].block[3].um_I.ena ;
 wire \top_I.branch[16].block[3].um_I.iw[10] ;
 wire \top_I.branch[16].block[3].um_I.iw[11] ;
 wire \top_I.branch[16].block[3].um_I.iw[12] ;
 wire \top_I.branch[16].block[3].um_I.iw[13] ;
 wire \top_I.branch[16].block[3].um_I.iw[14] ;
 wire \top_I.branch[16].block[3].um_I.iw[15] ;
 wire \top_I.branch[16].block[3].um_I.iw[16] ;
 wire \top_I.branch[16].block[3].um_I.iw[17] ;
 wire \top_I.branch[16].block[3].um_I.iw[1] ;
 wire \top_I.branch[16].block[3].um_I.iw[2] ;
 wire \top_I.branch[16].block[3].um_I.iw[3] ;
 wire \top_I.branch[16].block[3].um_I.iw[4] ;
 wire \top_I.branch[16].block[3].um_I.iw[5] ;
 wire \top_I.branch[16].block[3].um_I.iw[6] ;
 wire \top_I.branch[16].block[3].um_I.iw[7] ;
 wire \top_I.branch[16].block[3].um_I.iw[8] ;
 wire \top_I.branch[16].block[3].um_I.iw[9] ;
 wire \top_I.branch[16].block[3].um_I.k_zero ;
 wire \top_I.branch[16].block[3].um_I.pg_vdd ;
 wire \top_I.branch[16].block[4].um_I.ana[2] ;
 wire \top_I.branch[16].block[4].um_I.ana[3] ;
 wire \top_I.branch[16].block[4].um_I.ana[4] ;
 wire \top_I.branch[16].block[4].um_I.ana[5] ;
 wire \top_I.branch[16].block[4].um_I.ana[6] ;
 wire \top_I.branch[16].block[4].um_I.ana[7] ;
 wire \top_I.branch[16].block[4].um_I.clk ;
 wire \top_I.branch[16].block[4].um_I.ena ;
 wire \top_I.branch[16].block[4].um_I.iw[10] ;
 wire \top_I.branch[16].block[4].um_I.iw[11] ;
 wire \top_I.branch[16].block[4].um_I.iw[12] ;
 wire \top_I.branch[16].block[4].um_I.iw[13] ;
 wire \top_I.branch[16].block[4].um_I.iw[14] ;
 wire \top_I.branch[16].block[4].um_I.iw[15] ;
 wire \top_I.branch[16].block[4].um_I.iw[16] ;
 wire \top_I.branch[16].block[4].um_I.iw[17] ;
 wire \top_I.branch[16].block[4].um_I.iw[1] ;
 wire \top_I.branch[16].block[4].um_I.iw[2] ;
 wire \top_I.branch[16].block[4].um_I.iw[3] ;
 wire \top_I.branch[16].block[4].um_I.iw[4] ;
 wire \top_I.branch[16].block[4].um_I.iw[5] ;
 wire \top_I.branch[16].block[4].um_I.iw[6] ;
 wire \top_I.branch[16].block[4].um_I.iw[7] ;
 wire \top_I.branch[16].block[4].um_I.iw[8] ;
 wire \top_I.branch[16].block[4].um_I.iw[9] ;
 wire \top_I.branch[16].block[4].um_I.k_zero ;
 wire \top_I.branch[16].block[4].um_I.ow[0] ;
 wire \top_I.branch[16].block[4].um_I.ow[10] ;
 wire \top_I.branch[16].block[4].um_I.ow[11] ;
 wire \top_I.branch[16].block[4].um_I.ow[12] ;
 wire \top_I.branch[16].block[4].um_I.ow[13] ;
 wire \top_I.branch[16].block[4].um_I.ow[14] ;
 wire \top_I.branch[16].block[4].um_I.ow[15] ;
 wire \top_I.branch[16].block[4].um_I.ow[16] ;
 wire \top_I.branch[16].block[4].um_I.ow[17] ;
 wire \top_I.branch[16].block[4].um_I.ow[18] ;
 wire \top_I.branch[16].block[4].um_I.ow[19] ;
 wire \top_I.branch[16].block[4].um_I.ow[1] ;
 wire \top_I.branch[16].block[4].um_I.ow[20] ;
 wire \top_I.branch[16].block[4].um_I.ow[21] ;
 wire \top_I.branch[16].block[4].um_I.ow[22] ;
 wire \top_I.branch[16].block[4].um_I.ow[23] ;
 wire \top_I.branch[16].block[4].um_I.ow[2] ;
 wire \top_I.branch[16].block[4].um_I.ow[3] ;
 wire \top_I.branch[16].block[4].um_I.ow[4] ;
 wire \top_I.branch[16].block[4].um_I.ow[5] ;
 wire \top_I.branch[16].block[4].um_I.ow[6] ;
 wire \top_I.branch[16].block[4].um_I.ow[7] ;
 wire \top_I.branch[16].block[4].um_I.ow[8] ;
 wire \top_I.branch[16].block[4].um_I.ow[9] ;
 wire \top_I.branch[16].block[4].um_I.pg_vdd ;
 wire \top_I.branch[16].block[5].um_I.ana[2] ;
 wire \top_I.branch[16].block[5].um_I.ana[3] ;
 wire \top_I.branch[16].block[5].um_I.ana[4] ;
 wire \top_I.branch[16].block[5].um_I.ana[5] ;
 wire \top_I.branch[16].block[5].um_I.ana[6] ;
 wire \top_I.branch[16].block[5].um_I.ana[7] ;
 wire \top_I.branch[16].block[5].um_I.clk ;
 wire \top_I.branch[16].block[5].um_I.ena ;
 wire \top_I.branch[16].block[5].um_I.iw[10] ;
 wire \top_I.branch[16].block[5].um_I.iw[11] ;
 wire \top_I.branch[16].block[5].um_I.iw[12] ;
 wire \top_I.branch[16].block[5].um_I.iw[13] ;
 wire \top_I.branch[16].block[5].um_I.iw[14] ;
 wire \top_I.branch[16].block[5].um_I.iw[15] ;
 wire \top_I.branch[16].block[5].um_I.iw[16] ;
 wire \top_I.branch[16].block[5].um_I.iw[17] ;
 wire \top_I.branch[16].block[5].um_I.iw[1] ;
 wire \top_I.branch[16].block[5].um_I.iw[2] ;
 wire \top_I.branch[16].block[5].um_I.iw[3] ;
 wire \top_I.branch[16].block[5].um_I.iw[4] ;
 wire \top_I.branch[16].block[5].um_I.iw[5] ;
 wire \top_I.branch[16].block[5].um_I.iw[6] ;
 wire \top_I.branch[16].block[5].um_I.iw[7] ;
 wire \top_I.branch[16].block[5].um_I.iw[8] ;
 wire \top_I.branch[16].block[5].um_I.iw[9] ;
 wire \top_I.branch[16].block[5].um_I.k_zero ;
 wire \top_I.branch[16].block[5].um_I.pg_vdd ;
 wire \top_I.branch[16].block[6].um_I.ana[2] ;
 wire \top_I.branch[16].block[6].um_I.ana[3] ;
 wire \top_I.branch[16].block[6].um_I.ana[4] ;
 wire \top_I.branch[16].block[6].um_I.ana[5] ;
 wire \top_I.branch[16].block[6].um_I.ana[6] ;
 wire \top_I.branch[16].block[6].um_I.ana[7] ;
 wire \top_I.branch[16].block[6].um_I.clk ;
 wire \top_I.branch[16].block[6].um_I.ena ;
 wire \top_I.branch[16].block[6].um_I.iw[10] ;
 wire \top_I.branch[16].block[6].um_I.iw[11] ;
 wire \top_I.branch[16].block[6].um_I.iw[12] ;
 wire \top_I.branch[16].block[6].um_I.iw[13] ;
 wire \top_I.branch[16].block[6].um_I.iw[14] ;
 wire \top_I.branch[16].block[6].um_I.iw[15] ;
 wire \top_I.branch[16].block[6].um_I.iw[16] ;
 wire \top_I.branch[16].block[6].um_I.iw[17] ;
 wire \top_I.branch[16].block[6].um_I.iw[1] ;
 wire \top_I.branch[16].block[6].um_I.iw[2] ;
 wire \top_I.branch[16].block[6].um_I.iw[3] ;
 wire \top_I.branch[16].block[6].um_I.iw[4] ;
 wire \top_I.branch[16].block[6].um_I.iw[5] ;
 wire \top_I.branch[16].block[6].um_I.iw[6] ;
 wire \top_I.branch[16].block[6].um_I.iw[7] ;
 wire \top_I.branch[16].block[6].um_I.iw[8] ;
 wire \top_I.branch[16].block[6].um_I.iw[9] ;
 wire \top_I.branch[16].block[6].um_I.k_zero ;
 wire \top_I.branch[16].block[6].um_I.pg_vdd ;
 wire \top_I.branch[16].block[7].um_I.ana[2] ;
 wire \top_I.branch[16].block[7].um_I.ana[3] ;
 wire \top_I.branch[16].block[7].um_I.ana[4] ;
 wire \top_I.branch[16].block[7].um_I.ana[5] ;
 wire \top_I.branch[16].block[7].um_I.ana[6] ;
 wire \top_I.branch[16].block[7].um_I.ana[7] ;
 wire \top_I.branch[16].block[7].um_I.clk ;
 wire \top_I.branch[16].block[7].um_I.ena ;
 wire \top_I.branch[16].block[7].um_I.iw[10] ;
 wire \top_I.branch[16].block[7].um_I.iw[11] ;
 wire \top_I.branch[16].block[7].um_I.iw[12] ;
 wire \top_I.branch[16].block[7].um_I.iw[13] ;
 wire \top_I.branch[16].block[7].um_I.iw[14] ;
 wire \top_I.branch[16].block[7].um_I.iw[15] ;
 wire \top_I.branch[16].block[7].um_I.iw[16] ;
 wire \top_I.branch[16].block[7].um_I.iw[17] ;
 wire \top_I.branch[16].block[7].um_I.iw[1] ;
 wire \top_I.branch[16].block[7].um_I.iw[2] ;
 wire \top_I.branch[16].block[7].um_I.iw[3] ;
 wire \top_I.branch[16].block[7].um_I.iw[4] ;
 wire \top_I.branch[16].block[7].um_I.iw[5] ;
 wire \top_I.branch[16].block[7].um_I.iw[6] ;
 wire \top_I.branch[16].block[7].um_I.iw[7] ;
 wire \top_I.branch[16].block[7].um_I.iw[8] ;
 wire \top_I.branch[16].block[7].um_I.iw[9] ;
 wire \top_I.branch[16].block[7].um_I.k_zero ;
 wire \top_I.branch[16].block[7].um_I.pg_vdd ;
 wire \top_I.branch[16].block[8].um_I.ana[2] ;
 wire \top_I.branch[16].block[8].um_I.ana[3] ;
 wire \top_I.branch[16].block[8].um_I.ana[4] ;
 wire \top_I.branch[16].block[8].um_I.ana[5] ;
 wire \top_I.branch[16].block[8].um_I.ana[6] ;
 wire \top_I.branch[16].block[8].um_I.ana[7] ;
 wire \top_I.branch[16].block[8].um_I.clk ;
 wire \top_I.branch[16].block[8].um_I.ena ;
 wire \top_I.branch[16].block[8].um_I.iw[10] ;
 wire \top_I.branch[16].block[8].um_I.iw[11] ;
 wire \top_I.branch[16].block[8].um_I.iw[12] ;
 wire \top_I.branch[16].block[8].um_I.iw[13] ;
 wire \top_I.branch[16].block[8].um_I.iw[14] ;
 wire \top_I.branch[16].block[8].um_I.iw[15] ;
 wire \top_I.branch[16].block[8].um_I.iw[16] ;
 wire \top_I.branch[16].block[8].um_I.iw[17] ;
 wire \top_I.branch[16].block[8].um_I.iw[1] ;
 wire \top_I.branch[16].block[8].um_I.iw[2] ;
 wire \top_I.branch[16].block[8].um_I.iw[3] ;
 wire \top_I.branch[16].block[8].um_I.iw[4] ;
 wire \top_I.branch[16].block[8].um_I.iw[5] ;
 wire \top_I.branch[16].block[8].um_I.iw[6] ;
 wire \top_I.branch[16].block[8].um_I.iw[7] ;
 wire \top_I.branch[16].block[8].um_I.iw[8] ;
 wire \top_I.branch[16].block[8].um_I.iw[9] ;
 wire \top_I.branch[16].block[8].um_I.k_zero ;
 wire \top_I.branch[16].block[8].um_I.pg_vdd ;
 wire \top_I.branch[16].block[9].um_I.ana[2] ;
 wire \top_I.branch[16].block[9].um_I.ana[3] ;
 wire \top_I.branch[16].block[9].um_I.ana[4] ;
 wire \top_I.branch[16].block[9].um_I.ana[5] ;
 wire \top_I.branch[16].block[9].um_I.ana[6] ;
 wire \top_I.branch[16].block[9].um_I.ana[7] ;
 wire \top_I.branch[16].block[9].um_I.clk ;
 wire \top_I.branch[16].block[9].um_I.ena ;
 wire \top_I.branch[16].block[9].um_I.iw[10] ;
 wire \top_I.branch[16].block[9].um_I.iw[11] ;
 wire \top_I.branch[16].block[9].um_I.iw[12] ;
 wire \top_I.branch[16].block[9].um_I.iw[13] ;
 wire \top_I.branch[16].block[9].um_I.iw[14] ;
 wire \top_I.branch[16].block[9].um_I.iw[15] ;
 wire \top_I.branch[16].block[9].um_I.iw[16] ;
 wire \top_I.branch[16].block[9].um_I.iw[17] ;
 wire \top_I.branch[16].block[9].um_I.iw[1] ;
 wire \top_I.branch[16].block[9].um_I.iw[2] ;
 wire \top_I.branch[16].block[9].um_I.iw[3] ;
 wire \top_I.branch[16].block[9].um_I.iw[4] ;
 wire \top_I.branch[16].block[9].um_I.iw[5] ;
 wire \top_I.branch[16].block[9].um_I.iw[6] ;
 wire \top_I.branch[16].block[9].um_I.iw[7] ;
 wire \top_I.branch[16].block[9].um_I.iw[8] ;
 wire \top_I.branch[16].block[9].um_I.iw[9] ;
 wire \top_I.branch[16].block[9].um_I.k_zero ;
 wire \top_I.branch[16].block[9].um_I.pg_vdd ;
 wire \top_I.branch[16].l_addr[0] ;
 wire \top_I.branch[16].l_addr[3] ;
 wire \top_I.branch[17].block[0].um_I.ana[2] ;
 wire \top_I.branch[17].block[0].um_I.ana[3] ;
 wire \top_I.branch[17].block[0].um_I.ana[4] ;
 wire \top_I.branch[17].block[0].um_I.ana[5] ;
 wire \top_I.branch[17].block[0].um_I.ana[6] ;
 wire \top_I.branch[17].block[0].um_I.ana[7] ;
 wire \top_I.branch[17].block[0].um_I.clk ;
 wire \top_I.branch[17].block[0].um_I.ena ;
 wire \top_I.branch[17].block[0].um_I.iw[10] ;
 wire \top_I.branch[17].block[0].um_I.iw[11] ;
 wire \top_I.branch[17].block[0].um_I.iw[12] ;
 wire \top_I.branch[17].block[0].um_I.iw[13] ;
 wire \top_I.branch[17].block[0].um_I.iw[14] ;
 wire \top_I.branch[17].block[0].um_I.iw[15] ;
 wire \top_I.branch[17].block[0].um_I.iw[16] ;
 wire \top_I.branch[17].block[0].um_I.iw[17] ;
 wire \top_I.branch[17].block[0].um_I.iw[1] ;
 wire \top_I.branch[17].block[0].um_I.iw[2] ;
 wire \top_I.branch[17].block[0].um_I.iw[3] ;
 wire \top_I.branch[17].block[0].um_I.iw[4] ;
 wire \top_I.branch[17].block[0].um_I.iw[5] ;
 wire \top_I.branch[17].block[0].um_I.iw[6] ;
 wire \top_I.branch[17].block[0].um_I.iw[7] ;
 wire \top_I.branch[17].block[0].um_I.iw[8] ;
 wire \top_I.branch[17].block[0].um_I.iw[9] ;
 wire \top_I.branch[17].block[0].um_I.k_zero ;
 wire \top_I.branch[17].block[0].um_I.pg_vdd ;
 wire \top_I.branch[17].block[10].um_I.ana[2] ;
 wire \top_I.branch[17].block[10].um_I.ana[3] ;
 wire \top_I.branch[17].block[10].um_I.ana[4] ;
 wire \top_I.branch[17].block[10].um_I.ana[5] ;
 wire \top_I.branch[17].block[10].um_I.ana[6] ;
 wire \top_I.branch[17].block[10].um_I.ana[7] ;
 wire \top_I.branch[17].block[10].um_I.clk ;
 wire \top_I.branch[17].block[10].um_I.ena ;
 wire \top_I.branch[17].block[10].um_I.iw[10] ;
 wire \top_I.branch[17].block[10].um_I.iw[11] ;
 wire \top_I.branch[17].block[10].um_I.iw[12] ;
 wire \top_I.branch[17].block[10].um_I.iw[13] ;
 wire \top_I.branch[17].block[10].um_I.iw[14] ;
 wire \top_I.branch[17].block[10].um_I.iw[15] ;
 wire \top_I.branch[17].block[10].um_I.iw[16] ;
 wire \top_I.branch[17].block[10].um_I.iw[17] ;
 wire \top_I.branch[17].block[10].um_I.iw[1] ;
 wire \top_I.branch[17].block[10].um_I.iw[2] ;
 wire \top_I.branch[17].block[10].um_I.iw[3] ;
 wire \top_I.branch[17].block[10].um_I.iw[4] ;
 wire \top_I.branch[17].block[10].um_I.iw[5] ;
 wire \top_I.branch[17].block[10].um_I.iw[6] ;
 wire \top_I.branch[17].block[10].um_I.iw[7] ;
 wire \top_I.branch[17].block[10].um_I.iw[8] ;
 wire \top_I.branch[17].block[10].um_I.iw[9] ;
 wire \top_I.branch[17].block[10].um_I.k_zero ;
 wire \top_I.branch[17].block[10].um_I.pg_vdd ;
 wire \top_I.branch[17].block[11].um_I.ana[2] ;
 wire \top_I.branch[17].block[11].um_I.ana[3] ;
 wire \top_I.branch[17].block[11].um_I.ana[4] ;
 wire \top_I.branch[17].block[11].um_I.ana[5] ;
 wire \top_I.branch[17].block[11].um_I.ana[6] ;
 wire \top_I.branch[17].block[11].um_I.ana[7] ;
 wire \top_I.branch[17].block[11].um_I.clk ;
 wire \top_I.branch[17].block[11].um_I.ena ;
 wire \top_I.branch[17].block[11].um_I.iw[10] ;
 wire \top_I.branch[17].block[11].um_I.iw[11] ;
 wire \top_I.branch[17].block[11].um_I.iw[12] ;
 wire \top_I.branch[17].block[11].um_I.iw[13] ;
 wire \top_I.branch[17].block[11].um_I.iw[14] ;
 wire \top_I.branch[17].block[11].um_I.iw[15] ;
 wire \top_I.branch[17].block[11].um_I.iw[16] ;
 wire \top_I.branch[17].block[11].um_I.iw[17] ;
 wire \top_I.branch[17].block[11].um_I.iw[1] ;
 wire \top_I.branch[17].block[11].um_I.iw[2] ;
 wire \top_I.branch[17].block[11].um_I.iw[3] ;
 wire \top_I.branch[17].block[11].um_I.iw[4] ;
 wire \top_I.branch[17].block[11].um_I.iw[5] ;
 wire \top_I.branch[17].block[11].um_I.iw[6] ;
 wire \top_I.branch[17].block[11].um_I.iw[7] ;
 wire \top_I.branch[17].block[11].um_I.iw[8] ;
 wire \top_I.branch[17].block[11].um_I.iw[9] ;
 wire \top_I.branch[17].block[11].um_I.k_zero ;
 wire \top_I.branch[17].block[11].um_I.pg_vdd ;
 wire \top_I.branch[17].block[12].um_I.ana[2] ;
 wire \top_I.branch[17].block[12].um_I.ana[3] ;
 wire \top_I.branch[17].block[12].um_I.ana[4] ;
 wire \top_I.branch[17].block[12].um_I.ana[5] ;
 wire \top_I.branch[17].block[12].um_I.ana[6] ;
 wire \top_I.branch[17].block[12].um_I.ana[7] ;
 wire \top_I.branch[17].block[12].um_I.clk ;
 wire \top_I.branch[17].block[12].um_I.ena ;
 wire \top_I.branch[17].block[12].um_I.iw[10] ;
 wire \top_I.branch[17].block[12].um_I.iw[11] ;
 wire \top_I.branch[17].block[12].um_I.iw[12] ;
 wire \top_I.branch[17].block[12].um_I.iw[13] ;
 wire \top_I.branch[17].block[12].um_I.iw[14] ;
 wire \top_I.branch[17].block[12].um_I.iw[15] ;
 wire \top_I.branch[17].block[12].um_I.iw[16] ;
 wire \top_I.branch[17].block[12].um_I.iw[17] ;
 wire \top_I.branch[17].block[12].um_I.iw[1] ;
 wire \top_I.branch[17].block[12].um_I.iw[2] ;
 wire \top_I.branch[17].block[12].um_I.iw[3] ;
 wire \top_I.branch[17].block[12].um_I.iw[4] ;
 wire \top_I.branch[17].block[12].um_I.iw[5] ;
 wire \top_I.branch[17].block[12].um_I.iw[6] ;
 wire \top_I.branch[17].block[12].um_I.iw[7] ;
 wire \top_I.branch[17].block[12].um_I.iw[8] ;
 wire \top_I.branch[17].block[12].um_I.iw[9] ;
 wire \top_I.branch[17].block[12].um_I.k_zero ;
 wire \top_I.branch[17].block[12].um_I.pg_vdd ;
 wire \top_I.branch[17].block[13].um_I.ana[2] ;
 wire \top_I.branch[17].block[13].um_I.ana[3] ;
 wire \top_I.branch[17].block[13].um_I.ana[4] ;
 wire \top_I.branch[17].block[13].um_I.ana[5] ;
 wire \top_I.branch[17].block[13].um_I.ana[6] ;
 wire \top_I.branch[17].block[13].um_I.ana[7] ;
 wire \top_I.branch[17].block[13].um_I.clk ;
 wire \top_I.branch[17].block[13].um_I.ena ;
 wire \top_I.branch[17].block[13].um_I.iw[10] ;
 wire \top_I.branch[17].block[13].um_I.iw[11] ;
 wire \top_I.branch[17].block[13].um_I.iw[12] ;
 wire \top_I.branch[17].block[13].um_I.iw[13] ;
 wire \top_I.branch[17].block[13].um_I.iw[14] ;
 wire \top_I.branch[17].block[13].um_I.iw[15] ;
 wire \top_I.branch[17].block[13].um_I.iw[16] ;
 wire \top_I.branch[17].block[13].um_I.iw[17] ;
 wire \top_I.branch[17].block[13].um_I.iw[1] ;
 wire \top_I.branch[17].block[13].um_I.iw[2] ;
 wire \top_I.branch[17].block[13].um_I.iw[3] ;
 wire \top_I.branch[17].block[13].um_I.iw[4] ;
 wire \top_I.branch[17].block[13].um_I.iw[5] ;
 wire \top_I.branch[17].block[13].um_I.iw[6] ;
 wire \top_I.branch[17].block[13].um_I.iw[7] ;
 wire \top_I.branch[17].block[13].um_I.iw[8] ;
 wire \top_I.branch[17].block[13].um_I.iw[9] ;
 wire \top_I.branch[17].block[13].um_I.k_zero ;
 wire \top_I.branch[17].block[13].um_I.pg_vdd ;
 wire \top_I.branch[17].block[14].um_I.ana[2] ;
 wire \top_I.branch[17].block[14].um_I.ana[3] ;
 wire \top_I.branch[17].block[14].um_I.ana[4] ;
 wire \top_I.branch[17].block[14].um_I.ana[5] ;
 wire \top_I.branch[17].block[14].um_I.ana[6] ;
 wire \top_I.branch[17].block[14].um_I.ana[7] ;
 wire \top_I.branch[17].block[14].um_I.clk ;
 wire \top_I.branch[17].block[14].um_I.ena ;
 wire \top_I.branch[17].block[14].um_I.iw[10] ;
 wire \top_I.branch[17].block[14].um_I.iw[11] ;
 wire \top_I.branch[17].block[14].um_I.iw[12] ;
 wire \top_I.branch[17].block[14].um_I.iw[13] ;
 wire \top_I.branch[17].block[14].um_I.iw[14] ;
 wire \top_I.branch[17].block[14].um_I.iw[15] ;
 wire \top_I.branch[17].block[14].um_I.iw[16] ;
 wire \top_I.branch[17].block[14].um_I.iw[17] ;
 wire \top_I.branch[17].block[14].um_I.iw[1] ;
 wire \top_I.branch[17].block[14].um_I.iw[2] ;
 wire \top_I.branch[17].block[14].um_I.iw[3] ;
 wire \top_I.branch[17].block[14].um_I.iw[4] ;
 wire \top_I.branch[17].block[14].um_I.iw[5] ;
 wire \top_I.branch[17].block[14].um_I.iw[6] ;
 wire \top_I.branch[17].block[14].um_I.iw[7] ;
 wire \top_I.branch[17].block[14].um_I.iw[8] ;
 wire \top_I.branch[17].block[14].um_I.iw[9] ;
 wire \top_I.branch[17].block[14].um_I.k_zero ;
 wire \top_I.branch[17].block[14].um_I.pg_vdd ;
 wire \top_I.branch[17].block[15].um_I.ana[2] ;
 wire \top_I.branch[17].block[15].um_I.ana[3] ;
 wire \top_I.branch[17].block[15].um_I.ana[4] ;
 wire \top_I.branch[17].block[15].um_I.ana[5] ;
 wire \top_I.branch[17].block[15].um_I.ana[6] ;
 wire \top_I.branch[17].block[15].um_I.ana[7] ;
 wire \top_I.branch[17].block[15].um_I.clk ;
 wire \top_I.branch[17].block[15].um_I.ena ;
 wire \top_I.branch[17].block[15].um_I.iw[10] ;
 wire \top_I.branch[17].block[15].um_I.iw[11] ;
 wire \top_I.branch[17].block[15].um_I.iw[12] ;
 wire \top_I.branch[17].block[15].um_I.iw[13] ;
 wire \top_I.branch[17].block[15].um_I.iw[14] ;
 wire \top_I.branch[17].block[15].um_I.iw[15] ;
 wire \top_I.branch[17].block[15].um_I.iw[16] ;
 wire \top_I.branch[17].block[15].um_I.iw[17] ;
 wire \top_I.branch[17].block[15].um_I.iw[1] ;
 wire \top_I.branch[17].block[15].um_I.iw[2] ;
 wire \top_I.branch[17].block[15].um_I.iw[3] ;
 wire \top_I.branch[17].block[15].um_I.iw[4] ;
 wire \top_I.branch[17].block[15].um_I.iw[5] ;
 wire \top_I.branch[17].block[15].um_I.iw[6] ;
 wire \top_I.branch[17].block[15].um_I.iw[7] ;
 wire \top_I.branch[17].block[15].um_I.iw[8] ;
 wire \top_I.branch[17].block[15].um_I.iw[9] ;
 wire \top_I.branch[17].block[15].um_I.k_zero ;
 wire \top_I.branch[17].block[15].um_I.pg_vdd ;
 wire \top_I.branch[17].block[1].um_I.ana[2] ;
 wire \top_I.branch[17].block[1].um_I.ana[3] ;
 wire \top_I.branch[17].block[1].um_I.ana[4] ;
 wire \top_I.branch[17].block[1].um_I.ana[5] ;
 wire \top_I.branch[17].block[1].um_I.ana[6] ;
 wire \top_I.branch[17].block[1].um_I.ana[7] ;
 wire \top_I.branch[17].block[1].um_I.clk ;
 wire \top_I.branch[17].block[1].um_I.ena ;
 wire \top_I.branch[17].block[1].um_I.iw[10] ;
 wire \top_I.branch[17].block[1].um_I.iw[11] ;
 wire \top_I.branch[17].block[1].um_I.iw[12] ;
 wire \top_I.branch[17].block[1].um_I.iw[13] ;
 wire \top_I.branch[17].block[1].um_I.iw[14] ;
 wire \top_I.branch[17].block[1].um_I.iw[15] ;
 wire \top_I.branch[17].block[1].um_I.iw[16] ;
 wire \top_I.branch[17].block[1].um_I.iw[17] ;
 wire \top_I.branch[17].block[1].um_I.iw[1] ;
 wire \top_I.branch[17].block[1].um_I.iw[2] ;
 wire \top_I.branch[17].block[1].um_I.iw[3] ;
 wire \top_I.branch[17].block[1].um_I.iw[4] ;
 wire \top_I.branch[17].block[1].um_I.iw[5] ;
 wire \top_I.branch[17].block[1].um_I.iw[6] ;
 wire \top_I.branch[17].block[1].um_I.iw[7] ;
 wire \top_I.branch[17].block[1].um_I.iw[8] ;
 wire \top_I.branch[17].block[1].um_I.iw[9] ;
 wire \top_I.branch[17].block[1].um_I.k_zero ;
 wire \top_I.branch[17].block[1].um_I.pg_vdd ;
 wire \top_I.branch[17].block[2].um_I.ana[2] ;
 wire \top_I.branch[17].block[2].um_I.ana[3] ;
 wire \top_I.branch[17].block[2].um_I.ana[4] ;
 wire \top_I.branch[17].block[2].um_I.ana[5] ;
 wire \top_I.branch[17].block[2].um_I.ana[6] ;
 wire \top_I.branch[17].block[2].um_I.ana[7] ;
 wire \top_I.branch[17].block[2].um_I.clk ;
 wire \top_I.branch[17].block[2].um_I.ena ;
 wire \top_I.branch[17].block[2].um_I.iw[10] ;
 wire \top_I.branch[17].block[2].um_I.iw[11] ;
 wire \top_I.branch[17].block[2].um_I.iw[12] ;
 wire \top_I.branch[17].block[2].um_I.iw[13] ;
 wire \top_I.branch[17].block[2].um_I.iw[14] ;
 wire \top_I.branch[17].block[2].um_I.iw[15] ;
 wire \top_I.branch[17].block[2].um_I.iw[16] ;
 wire \top_I.branch[17].block[2].um_I.iw[17] ;
 wire \top_I.branch[17].block[2].um_I.iw[1] ;
 wire \top_I.branch[17].block[2].um_I.iw[2] ;
 wire \top_I.branch[17].block[2].um_I.iw[3] ;
 wire \top_I.branch[17].block[2].um_I.iw[4] ;
 wire \top_I.branch[17].block[2].um_I.iw[5] ;
 wire \top_I.branch[17].block[2].um_I.iw[6] ;
 wire \top_I.branch[17].block[2].um_I.iw[7] ;
 wire \top_I.branch[17].block[2].um_I.iw[8] ;
 wire \top_I.branch[17].block[2].um_I.iw[9] ;
 wire \top_I.branch[17].block[2].um_I.k_zero ;
 wire \top_I.branch[17].block[2].um_I.pg_vdd ;
 wire \top_I.branch[17].block[3].um_I.ana[2] ;
 wire \top_I.branch[17].block[3].um_I.ana[3] ;
 wire \top_I.branch[17].block[3].um_I.ana[4] ;
 wire \top_I.branch[17].block[3].um_I.ana[5] ;
 wire \top_I.branch[17].block[3].um_I.ana[6] ;
 wire \top_I.branch[17].block[3].um_I.ana[7] ;
 wire \top_I.branch[17].block[3].um_I.clk ;
 wire \top_I.branch[17].block[3].um_I.ena ;
 wire \top_I.branch[17].block[3].um_I.iw[10] ;
 wire \top_I.branch[17].block[3].um_I.iw[11] ;
 wire \top_I.branch[17].block[3].um_I.iw[12] ;
 wire \top_I.branch[17].block[3].um_I.iw[13] ;
 wire \top_I.branch[17].block[3].um_I.iw[14] ;
 wire \top_I.branch[17].block[3].um_I.iw[15] ;
 wire \top_I.branch[17].block[3].um_I.iw[16] ;
 wire \top_I.branch[17].block[3].um_I.iw[17] ;
 wire \top_I.branch[17].block[3].um_I.iw[1] ;
 wire \top_I.branch[17].block[3].um_I.iw[2] ;
 wire \top_I.branch[17].block[3].um_I.iw[3] ;
 wire \top_I.branch[17].block[3].um_I.iw[4] ;
 wire \top_I.branch[17].block[3].um_I.iw[5] ;
 wire \top_I.branch[17].block[3].um_I.iw[6] ;
 wire \top_I.branch[17].block[3].um_I.iw[7] ;
 wire \top_I.branch[17].block[3].um_I.iw[8] ;
 wire \top_I.branch[17].block[3].um_I.iw[9] ;
 wire \top_I.branch[17].block[3].um_I.k_zero ;
 wire \top_I.branch[17].block[3].um_I.pg_vdd ;
 wire \top_I.branch[17].block[4].um_I.ana[2] ;
 wire \top_I.branch[17].block[4].um_I.ana[3] ;
 wire \top_I.branch[17].block[4].um_I.ana[4] ;
 wire \top_I.branch[17].block[4].um_I.ana[5] ;
 wire \top_I.branch[17].block[4].um_I.ana[6] ;
 wire \top_I.branch[17].block[4].um_I.ana[7] ;
 wire \top_I.branch[17].block[4].um_I.clk ;
 wire \top_I.branch[17].block[4].um_I.ena ;
 wire \top_I.branch[17].block[4].um_I.iw[10] ;
 wire \top_I.branch[17].block[4].um_I.iw[11] ;
 wire \top_I.branch[17].block[4].um_I.iw[12] ;
 wire \top_I.branch[17].block[4].um_I.iw[13] ;
 wire \top_I.branch[17].block[4].um_I.iw[14] ;
 wire \top_I.branch[17].block[4].um_I.iw[15] ;
 wire \top_I.branch[17].block[4].um_I.iw[16] ;
 wire \top_I.branch[17].block[4].um_I.iw[17] ;
 wire \top_I.branch[17].block[4].um_I.iw[1] ;
 wire \top_I.branch[17].block[4].um_I.iw[2] ;
 wire \top_I.branch[17].block[4].um_I.iw[3] ;
 wire \top_I.branch[17].block[4].um_I.iw[4] ;
 wire \top_I.branch[17].block[4].um_I.iw[5] ;
 wire \top_I.branch[17].block[4].um_I.iw[6] ;
 wire \top_I.branch[17].block[4].um_I.iw[7] ;
 wire \top_I.branch[17].block[4].um_I.iw[8] ;
 wire \top_I.branch[17].block[4].um_I.iw[9] ;
 wire \top_I.branch[17].block[4].um_I.k_zero ;
 wire \top_I.branch[17].block[4].um_I.pg_vdd ;
 wire \top_I.branch[17].block[5].um_I.ana[2] ;
 wire \top_I.branch[17].block[5].um_I.ana[3] ;
 wire \top_I.branch[17].block[5].um_I.ana[4] ;
 wire \top_I.branch[17].block[5].um_I.ana[5] ;
 wire \top_I.branch[17].block[5].um_I.ana[6] ;
 wire \top_I.branch[17].block[5].um_I.ana[7] ;
 wire \top_I.branch[17].block[5].um_I.clk ;
 wire \top_I.branch[17].block[5].um_I.ena ;
 wire \top_I.branch[17].block[5].um_I.iw[10] ;
 wire \top_I.branch[17].block[5].um_I.iw[11] ;
 wire \top_I.branch[17].block[5].um_I.iw[12] ;
 wire \top_I.branch[17].block[5].um_I.iw[13] ;
 wire \top_I.branch[17].block[5].um_I.iw[14] ;
 wire \top_I.branch[17].block[5].um_I.iw[15] ;
 wire \top_I.branch[17].block[5].um_I.iw[16] ;
 wire \top_I.branch[17].block[5].um_I.iw[17] ;
 wire \top_I.branch[17].block[5].um_I.iw[1] ;
 wire \top_I.branch[17].block[5].um_I.iw[2] ;
 wire \top_I.branch[17].block[5].um_I.iw[3] ;
 wire \top_I.branch[17].block[5].um_I.iw[4] ;
 wire \top_I.branch[17].block[5].um_I.iw[5] ;
 wire \top_I.branch[17].block[5].um_I.iw[6] ;
 wire \top_I.branch[17].block[5].um_I.iw[7] ;
 wire \top_I.branch[17].block[5].um_I.iw[8] ;
 wire \top_I.branch[17].block[5].um_I.iw[9] ;
 wire \top_I.branch[17].block[5].um_I.k_zero ;
 wire \top_I.branch[17].block[5].um_I.pg_vdd ;
 wire \top_I.branch[17].block[6].um_I.ana[2] ;
 wire \top_I.branch[17].block[6].um_I.ana[3] ;
 wire \top_I.branch[17].block[6].um_I.ana[4] ;
 wire \top_I.branch[17].block[6].um_I.ana[5] ;
 wire \top_I.branch[17].block[6].um_I.ana[6] ;
 wire \top_I.branch[17].block[6].um_I.ana[7] ;
 wire \top_I.branch[17].block[6].um_I.clk ;
 wire \top_I.branch[17].block[6].um_I.ena ;
 wire \top_I.branch[17].block[6].um_I.iw[10] ;
 wire \top_I.branch[17].block[6].um_I.iw[11] ;
 wire \top_I.branch[17].block[6].um_I.iw[12] ;
 wire \top_I.branch[17].block[6].um_I.iw[13] ;
 wire \top_I.branch[17].block[6].um_I.iw[14] ;
 wire \top_I.branch[17].block[6].um_I.iw[15] ;
 wire \top_I.branch[17].block[6].um_I.iw[16] ;
 wire \top_I.branch[17].block[6].um_I.iw[17] ;
 wire \top_I.branch[17].block[6].um_I.iw[1] ;
 wire \top_I.branch[17].block[6].um_I.iw[2] ;
 wire \top_I.branch[17].block[6].um_I.iw[3] ;
 wire \top_I.branch[17].block[6].um_I.iw[4] ;
 wire \top_I.branch[17].block[6].um_I.iw[5] ;
 wire \top_I.branch[17].block[6].um_I.iw[6] ;
 wire \top_I.branch[17].block[6].um_I.iw[7] ;
 wire \top_I.branch[17].block[6].um_I.iw[8] ;
 wire \top_I.branch[17].block[6].um_I.iw[9] ;
 wire \top_I.branch[17].block[6].um_I.k_zero ;
 wire \top_I.branch[17].block[6].um_I.pg_vdd ;
 wire \top_I.branch[17].block[7].um_I.ana[2] ;
 wire \top_I.branch[17].block[7].um_I.ana[3] ;
 wire \top_I.branch[17].block[7].um_I.ana[4] ;
 wire \top_I.branch[17].block[7].um_I.ana[5] ;
 wire \top_I.branch[17].block[7].um_I.ana[6] ;
 wire \top_I.branch[17].block[7].um_I.ana[7] ;
 wire \top_I.branch[17].block[7].um_I.clk ;
 wire \top_I.branch[17].block[7].um_I.ena ;
 wire \top_I.branch[17].block[7].um_I.iw[10] ;
 wire \top_I.branch[17].block[7].um_I.iw[11] ;
 wire \top_I.branch[17].block[7].um_I.iw[12] ;
 wire \top_I.branch[17].block[7].um_I.iw[13] ;
 wire \top_I.branch[17].block[7].um_I.iw[14] ;
 wire \top_I.branch[17].block[7].um_I.iw[15] ;
 wire \top_I.branch[17].block[7].um_I.iw[16] ;
 wire \top_I.branch[17].block[7].um_I.iw[17] ;
 wire \top_I.branch[17].block[7].um_I.iw[1] ;
 wire \top_I.branch[17].block[7].um_I.iw[2] ;
 wire \top_I.branch[17].block[7].um_I.iw[3] ;
 wire \top_I.branch[17].block[7].um_I.iw[4] ;
 wire \top_I.branch[17].block[7].um_I.iw[5] ;
 wire \top_I.branch[17].block[7].um_I.iw[6] ;
 wire \top_I.branch[17].block[7].um_I.iw[7] ;
 wire \top_I.branch[17].block[7].um_I.iw[8] ;
 wire \top_I.branch[17].block[7].um_I.iw[9] ;
 wire \top_I.branch[17].block[7].um_I.k_zero ;
 wire \top_I.branch[17].block[7].um_I.pg_vdd ;
 wire \top_I.branch[17].block[8].um_I.ana[2] ;
 wire \top_I.branch[17].block[8].um_I.ana[3] ;
 wire \top_I.branch[17].block[8].um_I.ana[4] ;
 wire \top_I.branch[17].block[8].um_I.ana[5] ;
 wire \top_I.branch[17].block[8].um_I.ana[6] ;
 wire \top_I.branch[17].block[8].um_I.ana[7] ;
 wire \top_I.branch[17].block[8].um_I.clk ;
 wire \top_I.branch[17].block[8].um_I.ena ;
 wire \top_I.branch[17].block[8].um_I.iw[10] ;
 wire \top_I.branch[17].block[8].um_I.iw[11] ;
 wire \top_I.branch[17].block[8].um_I.iw[12] ;
 wire \top_I.branch[17].block[8].um_I.iw[13] ;
 wire \top_I.branch[17].block[8].um_I.iw[14] ;
 wire \top_I.branch[17].block[8].um_I.iw[15] ;
 wire \top_I.branch[17].block[8].um_I.iw[16] ;
 wire \top_I.branch[17].block[8].um_I.iw[17] ;
 wire \top_I.branch[17].block[8].um_I.iw[1] ;
 wire \top_I.branch[17].block[8].um_I.iw[2] ;
 wire \top_I.branch[17].block[8].um_I.iw[3] ;
 wire \top_I.branch[17].block[8].um_I.iw[4] ;
 wire \top_I.branch[17].block[8].um_I.iw[5] ;
 wire \top_I.branch[17].block[8].um_I.iw[6] ;
 wire \top_I.branch[17].block[8].um_I.iw[7] ;
 wire \top_I.branch[17].block[8].um_I.iw[8] ;
 wire \top_I.branch[17].block[8].um_I.iw[9] ;
 wire \top_I.branch[17].block[8].um_I.k_zero ;
 wire \top_I.branch[17].block[8].um_I.pg_vdd ;
 wire \top_I.branch[17].block[9].um_I.ana[2] ;
 wire \top_I.branch[17].block[9].um_I.ana[3] ;
 wire \top_I.branch[17].block[9].um_I.ana[4] ;
 wire \top_I.branch[17].block[9].um_I.ana[5] ;
 wire \top_I.branch[17].block[9].um_I.ana[6] ;
 wire \top_I.branch[17].block[9].um_I.ana[7] ;
 wire \top_I.branch[17].block[9].um_I.clk ;
 wire \top_I.branch[17].block[9].um_I.ena ;
 wire \top_I.branch[17].block[9].um_I.iw[10] ;
 wire \top_I.branch[17].block[9].um_I.iw[11] ;
 wire \top_I.branch[17].block[9].um_I.iw[12] ;
 wire \top_I.branch[17].block[9].um_I.iw[13] ;
 wire \top_I.branch[17].block[9].um_I.iw[14] ;
 wire \top_I.branch[17].block[9].um_I.iw[15] ;
 wire \top_I.branch[17].block[9].um_I.iw[16] ;
 wire \top_I.branch[17].block[9].um_I.iw[17] ;
 wire \top_I.branch[17].block[9].um_I.iw[1] ;
 wire \top_I.branch[17].block[9].um_I.iw[2] ;
 wire \top_I.branch[17].block[9].um_I.iw[3] ;
 wire \top_I.branch[17].block[9].um_I.iw[4] ;
 wire \top_I.branch[17].block[9].um_I.iw[5] ;
 wire \top_I.branch[17].block[9].um_I.iw[6] ;
 wire \top_I.branch[17].block[9].um_I.iw[7] ;
 wire \top_I.branch[17].block[9].um_I.iw[8] ;
 wire \top_I.branch[17].block[9].um_I.iw[9] ;
 wire \top_I.branch[17].block[9].um_I.k_zero ;
 wire \top_I.branch[17].block[9].um_I.pg_vdd ;
 wire \top_I.branch[17].l_addr[0] ;
 wire \top_I.branch[17].l_addr[3] ;
 wire \top_I.branch[18].block[0].um_I.ana[2] ;
 wire \top_I.branch[18].block[0].um_I.ana[3] ;
 wire \top_I.branch[18].block[0].um_I.ana[4] ;
 wire \top_I.branch[18].block[0].um_I.ana[5] ;
 wire \top_I.branch[18].block[0].um_I.ana[6] ;
 wire \top_I.branch[18].block[0].um_I.ana[7] ;
 wire \top_I.branch[18].block[0].um_I.clk ;
 wire \top_I.branch[18].block[0].um_I.ena ;
 wire \top_I.branch[18].block[0].um_I.iw[10] ;
 wire \top_I.branch[18].block[0].um_I.iw[11] ;
 wire \top_I.branch[18].block[0].um_I.iw[12] ;
 wire \top_I.branch[18].block[0].um_I.iw[13] ;
 wire \top_I.branch[18].block[0].um_I.iw[14] ;
 wire \top_I.branch[18].block[0].um_I.iw[15] ;
 wire \top_I.branch[18].block[0].um_I.iw[16] ;
 wire \top_I.branch[18].block[0].um_I.iw[17] ;
 wire \top_I.branch[18].block[0].um_I.iw[1] ;
 wire \top_I.branch[18].block[0].um_I.iw[2] ;
 wire \top_I.branch[18].block[0].um_I.iw[3] ;
 wire \top_I.branch[18].block[0].um_I.iw[4] ;
 wire \top_I.branch[18].block[0].um_I.iw[5] ;
 wire \top_I.branch[18].block[0].um_I.iw[6] ;
 wire \top_I.branch[18].block[0].um_I.iw[7] ;
 wire \top_I.branch[18].block[0].um_I.iw[8] ;
 wire \top_I.branch[18].block[0].um_I.iw[9] ;
 wire \top_I.branch[18].block[0].um_I.k_zero ;
 wire \top_I.branch[18].block[0].um_I.pg_vdd ;
 wire \top_I.branch[18].block[10].um_I.ana[2] ;
 wire \top_I.branch[18].block[10].um_I.ana[3] ;
 wire \top_I.branch[18].block[10].um_I.ana[4] ;
 wire \top_I.branch[18].block[10].um_I.ana[5] ;
 wire \top_I.branch[18].block[10].um_I.ana[6] ;
 wire \top_I.branch[18].block[10].um_I.ana[7] ;
 wire \top_I.branch[18].block[10].um_I.clk ;
 wire \top_I.branch[18].block[10].um_I.ena ;
 wire \top_I.branch[18].block[10].um_I.iw[10] ;
 wire \top_I.branch[18].block[10].um_I.iw[11] ;
 wire \top_I.branch[18].block[10].um_I.iw[12] ;
 wire \top_I.branch[18].block[10].um_I.iw[13] ;
 wire \top_I.branch[18].block[10].um_I.iw[14] ;
 wire \top_I.branch[18].block[10].um_I.iw[15] ;
 wire \top_I.branch[18].block[10].um_I.iw[16] ;
 wire \top_I.branch[18].block[10].um_I.iw[17] ;
 wire \top_I.branch[18].block[10].um_I.iw[1] ;
 wire \top_I.branch[18].block[10].um_I.iw[2] ;
 wire \top_I.branch[18].block[10].um_I.iw[3] ;
 wire \top_I.branch[18].block[10].um_I.iw[4] ;
 wire \top_I.branch[18].block[10].um_I.iw[5] ;
 wire \top_I.branch[18].block[10].um_I.iw[6] ;
 wire \top_I.branch[18].block[10].um_I.iw[7] ;
 wire \top_I.branch[18].block[10].um_I.iw[8] ;
 wire \top_I.branch[18].block[10].um_I.iw[9] ;
 wire \top_I.branch[18].block[10].um_I.k_zero ;
 wire \top_I.branch[18].block[10].um_I.pg_vdd ;
 wire \top_I.branch[18].block[11].um_I.ana[2] ;
 wire \top_I.branch[18].block[11].um_I.ana[3] ;
 wire \top_I.branch[18].block[11].um_I.ana[4] ;
 wire \top_I.branch[18].block[11].um_I.ana[5] ;
 wire \top_I.branch[18].block[11].um_I.ana[6] ;
 wire \top_I.branch[18].block[11].um_I.ana[7] ;
 wire \top_I.branch[18].block[11].um_I.clk ;
 wire \top_I.branch[18].block[11].um_I.ena ;
 wire \top_I.branch[18].block[11].um_I.iw[10] ;
 wire \top_I.branch[18].block[11].um_I.iw[11] ;
 wire \top_I.branch[18].block[11].um_I.iw[12] ;
 wire \top_I.branch[18].block[11].um_I.iw[13] ;
 wire \top_I.branch[18].block[11].um_I.iw[14] ;
 wire \top_I.branch[18].block[11].um_I.iw[15] ;
 wire \top_I.branch[18].block[11].um_I.iw[16] ;
 wire \top_I.branch[18].block[11].um_I.iw[17] ;
 wire \top_I.branch[18].block[11].um_I.iw[1] ;
 wire \top_I.branch[18].block[11].um_I.iw[2] ;
 wire \top_I.branch[18].block[11].um_I.iw[3] ;
 wire \top_I.branch[18].block[11].um_I.iw[4] ;
 wire \top_I.branch[18].block[11].um_I.iw[5] ;
 wire \top_I.branch[18].block[11].um_I.iw[6] ;
 wire \top_I.branch[18].block[11].um_I.iw[7] ;
 wire \top_I.branch[18].block[11].um_I.iw[8] ;
 wire \top_I.branch[18].block[11].um_I.iw[9] ;
 wire \top_I.branch[18].block[11].um_I.k_zero ;
 wire \top_I.branch[18].block[11].um_I.pg_vdd ;
 wire \top_I.branch[18].block[12].um_I.ana[2] ;
 wire \top_I.branch[18].block[12].um_I.ana[3] ;
 wire \top_I.branch[18].block[12].um_I.ana[4] ;
 wire \top_I.branch[18].block[12].um_I.ana[5] ;
 wire \top_I.branch[18].block[12].um_I.ana[6] ;
 wire \top_I.branch[18].block[12].um_I.ana[7] ;
 wire \top_I.branch[18].block[12].um_I.clk ;
 wire \top_I.branch[18].block[12].um_I.ena ;
 wire \top_I.branch[18].block[12].um_I.iw[10] ;
 wire \top_I.branch[18].block[12].um_I.iw[11] ;
 wire \top_I.branch[18].block[12].um_I.iw[12] ;
 wire \top_I.branch[18].block[12].um_I.iw[13] ;
 wire \top_I.branch[18].block[12].um_I.iw[14] ;
 wire \top_I.branch[18].block[12].um_I.iw[15] ;
 wire \top_I.branch[18].block[12].um_I.iw[16] ;
 wire \top_I.branch[18].block[12].um_I.iw[17] ;
 wire \top_I.branch[18].block[12].um_I.iw[1] ;
 wire \top_I.branch[18].block[12].um_I.iw[2] ;
 wire \top_I.branch[18].block[12].um_I.iw[3] ;
 wire \top_I.branch[18].block[12].um_I.iw[4] ;
 wire \top_I.branch[18].block[12].um_I.iw[5] ;
 wire \top_I.branch[18].block[12].um_I.iw[6] ;
 wire \top_I.branch[18].block[12].um_I.iw[7] ;
 wire \top_I.branch[18].block[12].um_I.iw[8] ;
 wire \top_I.branch[18].block[12].um_I.iw[9] ;
 wire \top_I.branch[18].block[12].um_I.k_zero ;
 wire \top_I.branch[18].block[12].um_I.pg_vdd ;
 wire \top_I.branch[18].block[13].um_I.ana[2] ;
 wire \top_I.branch[18].block[13].um_I.ana[3] ;
 wire \top_I.branch[18].block[13].um_I.ana[4] ;
 wire \top_I.branch[18].block[13].um_I.ana[5] ;
 wire \top_I.branch[18].block[13].um_I.ana[6] ;
 wire \top_I.branch[18].block[13].um_I.ana[7] ;
 wire \top_I.branch[18].block[13].um_I.clk ;
 wire \top_I.branch[18].block[13].um_I.ena ;
 wire \top_I.branch[18].block[13].um_I.iw[10] ;
 wire \top_I.branch[18].block[13].um_I.iw[11] ;
 wire \top_I.branch[18].block[13].um_I.iw[12] ;
 wire \top_I.branch[18].block[13].um_I.iw[13] ;
 wire \top_I.branch[18].block[13].um_I.iw[14] ;
 wire \top_I.branch[18].block[13].um_I.iw[15] ;
 wire \top_I.branch[18].block[13].um_I.iw[16] ;
 wire \top_I.branch[18].block[13].um_I.iw[17] ;
 wire \top_I.branch[18].block[13].um_I.iw[1] ;
 wire \top_I.branch[18].block[13].um_I.iw[2] ;
 wire \top_I.branch[18].block[13].um_I.iw[3] ;
 wire \top_I.branch[18].block[13].um_I.iw[4] ;
 wire \top_I.branch[18].block[13].um_I.iw[5] ;
 wire \top_I.branch[18].block[13].um_I.iw[6] ;
 wire \top_I.branch[18].block[13].um_I.iw[7] ;
 wire \top_I.branch[18].block[13].um_I.iw[8] ;
 wire \top_I.branch[18].block[13].um_I.iw[9] ;
 wire \top_I.branch[18].block[13].um_I.k_zero ;
 wire \top_I.branch[18].block[13].um_I.pg_vdd ;
 wire \top_I.branch[18].block[14].um_I.ana[2] ;
 wire \top_I.branch[18].block[14].um_I.ana[3] ;
 wire \top_I.branch[18].block[14].um_I.ana[4] ;
 wire \top_I.branch[18].block[14].um_I.ana[5] ;
 wire \top_I.branch[18].block[14].um_I.ana[6] ;
 wire \top_I.branch[18].block[14].um_I.ana[7] ;
 wire \top_I.branch[18].block[14].um_I.clk ;
 wire \top_I.branch[18].block[14].um_I.ena ;
 wire \top_I.branch[18].block[14].um_I.iw[10] ;
 wire \top_I.branch[18].block[14].um_I.iw[11] ;
 wire \top_I.branch[18].block[14].um_I.iw[12] ;
 wire \top_I.branch[18].block[14].um_I.iw[13] ;
 wire \top_I.branch[18].block[14].um_I.iw[14] ;
 wire \top_I.branch[18].block[14].um_I.iw[15] ;
 wire \top_I.branch[18].block[14].um_I.iw[16] ;
 wire \top_I.branch[18].block[14].um_I.iw[17] ;
 wire \top_I.branch[18].block[14].um_I.iw[1] ;
 wire \top_I.branch[18].block[14].um_I.iw[2] ;
 wire \top_I.branch[18].block[14].um_I.iw[3] ;
 wire \top_I.branch[18].block[14].um_I.iw[4] ;
 wire \top_I.branch[18].block[14].um_I.iw[5] ;
 wire \top_I.branch[18].block[14].um_I.iw[6] ;
 wire \top_I.branch[18].block[14].um_I.iw[7] ;
 wire \top_I.branch[18].block[14].um_I.iw[8] ;
 wire \top_I.branch[18].block[14].um_I.iw[9] ;
 wire \top_I.branch[18].block[14].um_I.k_zero ;
 wire \top_I.branch[18].block[14].um_I.pg_vdd ;
 wire \top_I.branch[18].block[15].um_I.ana[2] ;
 wire \top_I.branch[18].block[15].um_I.ana[3] ;
 wire \top_I.branch[18].block[15].um_I.ana[4] ;
 wire \top_I.branch[18].block[15].um_I.ana[5] ;
 wire \top_I.branch[18].block[15].um_I.ana[6] ;
 wire \top_I.branch[18].block[15].um_I.ana[7] ;
 wire \top_I.branch[18].block[15].um_I.clk ;
 wire \top_I.branch[18].block[15].um_I.ena ;
 wire \top_I.branch[18].block[15].um_I.iw[10] ;
 wire \top_I.branch[18].block[15].um_I.iw[11] ;
 wire \top_I.branch[18].block[15].um_I.iw[12] ;
 wire \top_I.branch[18].block[15].um_I.iw[13] ;
 wire \top_I.branch[18].block[15].um_I.iw[14] ;
 wire \top_I.branch[18].block[15].um_I.iw[15] ;
 wire \top_I.branch[18].block[15].um_I.iw[16] ;
 wire \top_I.branch[18].block[15].um_I.iw[17] ;
 wire \top_I.branch[18].block[15].um_I.iw[1] ;
 wire \top_I.branch[18].block[15].um_I.iw[2] ;
 wire \top_I.branch[18].block[15].um_I.iw[3] ;
 wire \top_I.branch[18].block[15].um_I.iw[4] ;
 wire \top_I.branch[18].block[15].um_I.iw[5] ;
 wire \top_I.branch[18].block[15].um_I.iw[6] ;
 wire \top_I.branch[18].block[15].um_I.iw[7] ;
 wire \top_I.branch[18].block[15].um_I.iw[8] ;
 wire \top_I.branch[18].block[15].um_I.iw[9] ;
 wire \top_I.branch[18].block[15].um_I.k_zero ;
 wire \top_I.branch[18].block[15].um_I.pg_vdd ;
 wire \top_I.branch[18].block[1].um_I.ana[2] ;
 wire \top_I.branch[18].block[1].um_I.ana[3] ;
 wire \top_I.branch[18].block[1].um_I.ana[4] ;
 wire \top_I.branch[18].block[1].um_I.ana[5] ;
 wire \top_I.branch[18].block[1].um_I.ana[6] ;
 wire \top_I.branch[18].block[1].um_I.ana[7] ;
 wire \top_I.branch[18].block[1].um_I.clk ;
 wire \top_I.branch[18].block[1].um_I.ena ;
 wire \top_I.branch[18].block[1].um_I.iw[10] ;
 wire \top_I.branch[18].block[1].um_I.iw[11] ;
 wire \top_I.branch[18].block[1].um_I.iw[12] ;
 wire \top_I.branch[18].block[1].um_I.iw[13] ;
 wire \top_I.branch[18].block[1].um_I.iw[14] ;
 wire \top_I.branch[18].block[1].um_I.iw[15] ;
 wire \top_I.branch[18].block[1].um_I.iw[16] ;
 wire \top_I.branch[18].block[1].um_I.iw[17] ;
 wire \top_I.branch[18].block[1].um_I.iw[1] ;
 wire \top_I.branch[18].block[1].um_I.iw[2] ;
 wire \top_I.branch[18].block[1].um_I.iw[3] ;
 wire \top_I.branch[18].block[1].um_I.iw[4] ;
 wire \top_I.branch[18].block[1].um_I.iw[5] ;
 wire \top_I.branch[18].block[1].um_I.iw[6] ;
 wire \top_I.branch[18].block[1].um_I.iw[7] ;
 wire \top_I.branch[18].block[1].um_I.iw[8] ;
 wire \top_I.branch[18].block[1].um_I.iw[9] ;
 wire \top_I.branch[18].block[1].um_I.k_zero ;
 wire \top_I.branch[18].block[1].um_I.pg_vdd ;
 wire \top_I.branch[18].block[2].um_I.ana[2] ;
 wire \top_I.branch[18].block[2].um_I.ana[3] ;
 wire \top_I.branch[18].block[2].um_I.ana[4] ;
 wire \top_I.branch[18].block[2].um_I.ana[5] ;
 wire \top_I.branch[18].block[2].um_I.ana[6] ;
 wire \top_I.branch[18].block[2].um_I.ana[7] ;
 wire \top_I.branch[18].block[2].um_I.clk ;
 wire \top_I.branch[18].block[2].um_I.ena ;
 wire \top_I.branch[18].block[2].um_I.iw[10] ;
 wire \top_I.branch[18].block[2].um_I.iw[11] ;
 wire \top_I.branch[18].block[2].um_I.iw[12] ;
 wire \top_I.branch[18].block[2].um_I.iw[13] ;
 wire \top_I.branch[18].block[2].um_I.iw[14] ;
 wire \top_I.branch[18].block[2].um_I.iw[15] ;
 wire \top_I.branch[18].block[2].um_I.iw[16] ;
 wire \top_I.branch[18].block[2].um_I.iw[17] ;
 wire \top_I.branch[18].block[2].um_I.iw[1] ;
 wire \top_I.branch[18].block[2].um_I.iw[2] ;
 wire \top_I.branch[18].block[2].um_I.iw[3] ;
 wire \top_I.branch[18].block[2].um_I.iw[4] ;
 wire \top_I.branch[18].block[2].um_I.iw[5] ;
 wire \top_I.branch[18].block[2].um_I.iw[6] ;
 wire \top_I.branch[18].block[2].um_I.iw[7] ;
 wire \top_I.branch[18].block[2].um_I.iw[8] ;
 wire \top_I.branch[18].block[2].um_I.iw[9] ;
 wire \top_I.branch[18].block[2].um_I.k_zero ;
 wire \top_I.branch[18].block[2].um_I.pg_vdd ;
 wire \top_I.branch[18].block[3].um_I.ana[2] ;
 wire \top_I.branch[18].block[3].um_I.ana[3] ;
 wire \top_I.branch[18].block[3].um_I.ana[4] ;
 wire \top_I.branch[18].block[3].um_I.ana[5] ;
 wire \top_I.branch[18].block[3].um_I.ana[6] ;
 wire \top_I.branch[18].block[3].um_I.ana[7] ;
 wire \top_I.branch[18].block[3].um_I.clk ;
 wire \top_I.branch[18].block[3].um_I.ena ;
 wire \top_I.branch[18].block[3].um_I.iw[10] ;
 wire \top_I.branch[18].block[3].um_I.iw[11] ;
 wire \top_I.branch[18].block[3].um_I.iw[12] ;
 wire \top_I.branch[18].block[3].um_I.iw[13] ;
 wire \top_I.branch[18].block[3].um_I.iw[14] ;
 wire \top_I.branch[18].block[3].um_I.iw[15] ;
 wire \top_I.branch[18].block[3].um_I.iw[16] ;
 wire \top_I.branch[18].block[3].um_I.iw[17] ;
 wire \top_I.branch[18].block[3].um_I.iw[1] ;
 wire \top_I.branch[18].block[3].um_I.iw[2] ;
 wire \top_I.branch[18].block[3].um_I.iw[3] ;
 wire \top_I.branch[18].block[3].um_I.iw[4] ;
 wire \top_I.branch[18].block[3].um_I.iw[5] ;
 wire \top_I.branch[18].block[3].um_I.iw[6] ;
 wire \top_I.branch[18].block[3].um_I.iw[7] ;
 wire \top_I.branch[18].block[3].um_I.iw[8] ;
 wire \top_I.branch[18].block[3].um_I.iw[9] ;
 wire \top_I.branch[18].block[3].um_I.k_zero ;
 wire \top_I.branch[18].block[3].um_I.pg_vdd ;
 wire \top_I.branch[18].block[4].um_I.ana[2] ;
 wire \top_I.branch[18].block[4].um_I.ana[3] ;
 wire \top_I.branch[18].block[4].um_I.ana[4] ;
 wire \top_I.branch[18].block[4].um_I.ana[5] ;
 wire \top_I.branch[18].block[4].um_I.ana[6] ;
 wire \top_I.branch[18].block[4].um_I.ana[7] ;
 wire \top_I.branch[18].block[4].um_I.clk ;
 wire \top_I.branch[18].block[4].um_I.ena ;
 wire \top_I.branch[18].block[4].um_I.iw[10] ;
 wire \top_I.branch[18].block[4].um_I.iw[11] ;
 wire \top_I.branch[18].block[4].um_I.iw[12] ;
 wire \top_I.branch[18].block[4].um_I.iw[13] ;
 wire \top_I.branch[18].block[4].um_I.iw[14] ;
 wire \top_I.branch[18].block[4].um_I.iw[15] ;
 wire \top_I.branch[18].block[4].um_I.iw[16] ;
 wire \top_I.branch[18].block[4].um_I.iw[17] ;
 wire \top_I.branch[18].block[4].um_I.iw[1] ;
 wire \top_I.branch[18].block[4].um_I.iw[2] ;
 wire \top_I.branch[18].block[4].um_I.iw[3] ;
 wire \top_I.branch[18].block[4].um_I.iw[4] ;
 wire \top_I.branch[18].block[4].um_I.iw[5] ;
 wire \top_I.branch[18].block[4].um_I.iw[6] ;
 wire \top_I.branch[18].block[4].um_I.iw[7] ;
 wire \top_I.branch[18].block[4].um_I.iw[8] ;
 wire \top_I.branch[18].block[4].um_I.iw[9] ;
 wire \top_I.branch[18].block[4].um_I.k_zero ;
 wire \top_I.branch[18].block[4].um_I.pg_vdd ;
 wire \top_I.branch[18].block[5].um_I.ana[2] ;
 wire \top_I.branch[18].block[5].um_I.ana[3] ;
 wire \top_I.branch[18].block[5].um_I.ana[4] ;
 wire \top_I.branch[18].block[5].um_I.ana[5] ;
 wire \top_I.branch[18].block[5].um_I.ana[6] ;
 wire \top_I.branch[18].block[5].um_I.ana[7] ;
 wire \top_I.branch[18].block[5].um_I.clk ;
 wire \top_I.branch[18].block[5].um_I.ena ;
 wire \top_I.branch[18].block[5].um_I.iw[10] ;
 wire \top_I.branch[18].block[5].um_I.iw[11] ;
 wire \top_I.branch[18].block[5].um_I.iw[12] ;
 wire \top_I.branch[18].block[5].um_I.iw[13] ;
 wire \top_I.branch[18].block[5].um_I.iw[14] ;
 wire \top_I.branch[18].block[5].um_I.iw[15] ;
 wire \top_I.branch[18].block[5].um_I.iw[16] ;
 wire \top_I.branch[18].block[5].um_I.iw[17] ;
 wire \top_I.branch[18].block[5].um_I.iw[1] ;
 wire \top_I.branch[18].block[5].um_I.iw[2] ;
 wire \top_I.branch[18].block[5].um_I.iw[3] ;
 wire \top_I.branch[18].block[5].um_I.iw[4] ;
 wire \top_I.branch[18].block[5].um_I.iw[5] ;
 wire \top_I.branch[18].block[5].um_I.iw[6] ;
 wire \top_I.branch[18].block[5].um_I.iw[7] ;
 wire \top_I.branch[18].block[5].um_I.iw[8] ;
 wire \top_I.branch[18].block[5].um_I.iw[9] ;
 wire \top_I.branch[18].block[5].um_I.k_zero ;
 wire \top_I.branch[18].block[5].um_I.pg_vdd ;
 wire \top_I.branch[18].block[6].um_I.ana[2] ;
 wire \top_I.branch[18].block[6].um_I.ana[3] ;
 wire \top_I.branch[18].block[6].um_I.ana[4] ;
 wire \top_I.branch[18].block[6].um_I.ana[5] ;
 wire \top_I.branch[18].block[6].um_I.ana[6] ;
 wire \top_I.branch[18].block[6].um_I.ana[7] ;
 wire \top_I.branch[18].block[6].um_I.clk ;
 wire \top_I.branch[18].block[6].um_I.ena ;
 wire \top_I.branch[18].block[6].um_I.iw[10] ;
 wire \top_I.branch[18].block[6].um_I.iw[11] ;
 wire \top_I.branch[18].block[6].um_I.iw[12] ;
 wire \top_I.branch[18].block[6].um_I.iw[13] ;
 wire \top_I.branch[18].block[6].um_I.iw[14] ;
 wire \top_I.branch[18].block[6].um_I.iw[15] ;
 wire \top_I.branch[18].block[6].um_I.iw[16] ;
 wire \top_I.branch[18].block[6].um_I.iw[17] ;
 wire \top_I.branch[18].block[6].um_I.iw[1] ;
 wire \top_I.branch[18].block[6].um_I.iw[2] ;
 wire \top_I.branch[18].block[6].um_I.iw[3] ;
 wire \top_I.branch[18].block[6].um_I.iw[4] ;
 wire \top_I.branch[18].block[6].um_I.iw[5] ;
 wire \top_I.branch[18].block[6].um_I.iw[6] ;
 wire \top_I.branch[18].block[6].um_I.iw[7] ;
 wire \top_I.branch[18].block[6].um_I.iw[8] ;
 wire \top_I.branch[18].block[6].um_I.iw[9] ;
 wire \top_I.branch[18].block[6].um_I.k_zero ;
 wire \top_I.branch[18].block[6].um_I.pg_vdd ;
 wire \top_I.branch[18].block[7].um_I.ana[2] ;
 wire \top_I.branch[18].block[7].um_I.ana[3] ;
 wire \top_I.branch[18].block[7].um_I.ana[4] ;
 wire \top_I.branch[18].block[7].um_I.ana[5] ;
 wire \top_I.branch[18].block[7].um_I.ana[6] ;
 wire \top_I.branch[18].block[7].um_I.ana[7] ;
 wire \top_I.branch[18].block[7].um_I.clk ;
 wire \top_I.branch[18].block[7].um_I.ena ;
 wire \top_I.branch[18].block[7].um_I.iw[10] ;
 wire \top_I.branch[18].block[7].um_I.iw[11] ;
 wire \top_I.branch[18].block[7].um_I.iw[12] ;
 wire \top_I.branch[18].block[7].um_I.iw[13] ;
 wire \top_I.branch[18].block[7].um_I.iw[14] ;
 wire \top_I.branch[18].block[7].um_I.iw[15] ;
 wire \top_I.branch[18].block[7].um_I.iw[16] ;
 wire \top_I.branch[18].block[7].um_I.iw[17] ;
 wire \top_I.branch[18].block[7].um_I.iw[1] ;
 wire \top_I.branch[18].block[7].um_I.iw[2] ;
 wire \top_I.branch[18].block[7].um_I.iw[3] ;
 wire \top_I.branch[18].block[7].um_I.iw[4] ;
 wire \top_I.branch[18].block[7].um_I.iw[5] ;
 wire \top_I.branch[18].block[7].um_I.iw[6] ;
 wire \top_I.branch[18].block[7].um_I.iw[7] ;
 wire \top_I.branch[18].block[7].um_I.iw[8] ;
 wire \top_I.branch[18].block[7].um_I.iw[9] ;
 wire \top_I.branch[18].block[7].um_I.k_zero ;
 wire \top_I.branch[18].block[7].um_I.pg_vdd ;
 wire \top_I.branch[18].block[8].um_I.ana[2] ;
 wire \top_I.branch[18].block[8].um_I.ana[3] ;
 wire \top_I.branch[18].block[8].um_I.ana[4] ;
 wire \top_I.branch[18].block[8].um_I.ana[5] ;
 wire \top_I.branch[18].block[8].um_I.ana[6] ;
 wire \top_I.branch[18].block[8].um_I.ana[7] ;
 wire \top_I.branch[18].block[8].um_I.clk ;
 wire \top_I.branch[18].block[8].um_I.ena ;
 wire \top_I.branch[18].block[8].um_I.iw[10] ;
 wire \top_I.branch[18].block[8].um_I.iw[11] ;
 wire \top_I.branch[18].block[8].um_I.iw[12] ;
 wire \top_I.branch[18].block[8].um_I.iw[13] ;
 wire \top_I.branch[18].block[8].um_I.iw[14] ;
 wire \top_I.branch[18].block[8].um_I.iw[15] ;
 wire \top_I.branch[18].block[8].um_I.iw[16] ;
 wire \top_I.branch[18].block[8].um_I.iw[17] ;
 wire \top_I.branch[18].block[8].um_I.iw[1] ;
 wire \top_I.branch[18].block[8].um_I.iw[2] ;
 wire \top_I.branch[18].block[8].um_I.iw[3] ;
 wire \top_I.branch[18].block[8].um_I.iw[4] ;
 wire \top_I.branch[18].block[8].um_I.iw[5] ;
 wire \top_I.branch[18].block[8].um_I.iw[6] ;
 wire \top_I.branch[18].block[8].um_I.iw[7] ;
 wire \top_I.branch[18].block[8].um_I.iw[8] ;
 wire \top_I.branch[18].block[8].um_I.iw[9] ;
 wire \top_I.branch[18].block[8].um_I.k_zero ;
 wire \top_I.branch[18].block[8].um_I.pg_vdd ;
 wire \top_I.branch[18].block[9].um_I.ana[2] ;
 wire \top_I.branch[18].block[9].um_I.ana[3] ;
 wire \top_I.branch[18].block[9].um_I.ana[4] ;
 wire \top_I.branch[18].block[9].um_I.ana[5] ;
 wire \top_I.branch[18].block[9].um_I.ana[6] ;
 wire \top_I.branch[18].block[9].um_I.ana[7] ;
 wire \top_I.branch[18].block[9].um_I.clk ;
 wire \top_I.branch[18].block[9].um_I.ena ;
 wire \top_I.branch[18].block[9].um_I.iw[10] ;
 wire \top_I.branch[18].block[9].um_I.iw[11] ;
 wire \top_I.branch[18].block[9].um_I.iw[12] ;
 wire \top_I.branch[18].block[9].um_I.iw[13] ;
 wire \top_I.branch[18].block[9].um_I.iw[14] ;
 wire \top_I.branch[18].block[9].um_I.iw[15] ;
 wire \top_I.branch[18].block[9].um_I.iw[16] ;
 wire \top_I.branch[18].block[9].um_I.iw[17] ;
 wire \top_I.branch[18].block[9].um_I.iw[1] ;
 wire \top_I.branch[18].block[9].um_I.iw[2] ;
 wire \top_I.branch[18].block[9].um_I.iw[3] ;
 wire \top_I.branch[18].block[9].um_I.iw[4] ;
 wire \top_I.branch[18].block[9].um_I.iw[5] ;
 wire \top_I.branch[18].block[9].um_I.iw[6] ;
 wire \top_I.branch[18].block[9].um_I.iw[7] ;
 wire \top_I.branch[18].block[9].um_I.iw[8] ;
 wire \top_I.branch[18].block[9].um_I.iw[9] ;
 wire \top_I.branch[18].block[9].um_I.k_zero ;
 wire \top_I.branch[18].block[9].um_I.pg_vdd ;
 wire \top_I.branch[18].l_addr[0] ;
 wire \top_I.branch[18].l_addr[1] ;
 wire \top_I.branch[19].block[0].um_I.ana[2] ;
 wire \top_I.branch[19].block[0].um_I.ana[3] ;
 wire \top_I.branch[19].block[0].um_I.ana[4] ;
 wire \top_I.branch[19].block[0].um_I.ana[5] ;
 wire \top_I.branch[19].block[0].um_I.ana[6] ;
 wire \top_I.branch[19].block[0].um_I.ana[7] ;
 wire \top_I.branch[19].block[0].um_I.clk ;
 wire \top_I.branch[19].block[0].um_I.ena ;
 wire \top_I.branch[19].block[0].um_I.iw[10] ;
 wire \top_I.branch[19].block[0].um_I.iw[11] ;
 wire \top_I.branch[19].block[0].um_I.iw[12] ;
 wire \top_I.branch[19].block[0].um_I.iw[13] ;
 wire \top_I.branch[19].block[0].um_I.iw[14] ;
 wire \top_I.branch[19].block[0].um_I.iw[15] ;
 wire \top_I.branch[19].block[0].um_I.iw[16] ;
 wire \top_I.branch[19].block[0].um_I.iw[17] ;
 wire \top_I.branch[19].block[0].um_I.iw[1] ;
 wire \top_I.branch[19].block[0].um_I.iw[2] ;
 wire \top_I.branch[19].block[0].um_I.iw[3] ;
 wire \top_I.branch[19].block[0].um_I.iw[4] ;
 wire \top_I.branch[19].block[0].um_I.iw[5] ;
 wire \top_I.branch[19].block[0].um_I.iw[6] ;
 wire \top_I.branch[19].block[0].um_I.iw[7] ;
 wire \top_I.branch[19].block[0].um_I.iw[8] ;
 wire \top_I.branch[19].block[0].um_I.iw[9] ;
 wire \top_I.branch[19].block[0].um_I.k_zero ;
 wire \top_I.branch[19].block[0].um_I.pg_vdd ;
 wire \top_I.branch[19].block[10].um_I.ana[2] ;
 wire \top_I.branch[19].block[10].um_I.ana[3] ;
 wire \top_I.branch[19].block[10].um_I.ana[4] ;
 wire \top_I.branch[19].block[10].um_I.ana[5] ;
 wire \top_I.branch[19].block[10].um_I.ana[6] ;
 wire \top_I.branch[19].block[10].um_I.ana[7] ;
 wire \top_I.branch[19].block[10].um_I.clk ;
 wire \top_I.branch[19].block[10].um_I.ena ;
 wire \top_I.branch[19].block[10].um_I.iw[10] ;
 wire \top_I.branch[19].block[10].um_I.iw[11] ;
 wire \top_I.branch[19].block[10].um_I.iw[12] ;
 wire \top_I.branch[19].block[10].um_I.iw[13] ;
 wire \top_I.branch[19].block[10].um_I.iw[14] ;
 wire \top_I.branch[19].block[10].um_I.iw[15] ;
 wire \top_I.branch[19].block[10].um_I.iw[16] ;
 wire \top_I.branch[19].block[10].um_I.iw[17] ;
 wire \top_I.branch[19].block[10].um_I.iw[1] ;
 wire \top_I.branch[19].block[10].um_I.iw[2] ;
 wire \top_I.branch[19].block[10].um_I.iw[3] ;
 wire \top_I.branch[19].block[10].um_I.iw[4] ;
 wire \top_I.branch[19].block[10].um_I.iw[5] ;
 wire \top_I.branch[19].block[10].um_I.iw[6] ;
 wire \top_I.branch[19].block[10].um_I.iw[7] ;
 wire \top_I.branch[19].block[10].um_I.iw[8] ;
 wire \top_I.branch[19].block[10].um_I.iw[9] ;
 wire \top_I.branch[19].block[10].um_I.k_zero ;
 wire \top_I.branch[19].block[10].um_I.pg_vdd ;
 wire \top_I.branch[19].block[11].um_I.ana[2] ;
 wire \top_I.branch[19].block[11].um_I.ana[3] ;
 wire \top_I.branch[19].block[11].um_I.ana[4] ;
 wire \top_I.branch[19].block[11].um_I.ana[5] ;
 wire \top_I.branch[19].block[11].um_I.ana[6] ;
 wire \top_I.branch[19].block[11].um_I.ana[7] ;
 wire \top_I.branch[19].block[11].um_I.clk ;
 wire \top_I.branch[19].block[11].um_I.ena ;
 wire \top_I.branch[19].block[11].um_I.iw[10] ;
 wire \top_I.branch[19].block[11].um_I.iw[11] ;
 wire \top_I.branch[19].block[11].um_I.iw[12] ;
 wire \top_I.branch[19].block[11].um_I.iw[13] ;
 wire \top_I.branch[19].block[11].um_I.iw[14] ;
 wire \top_I.branch[19].block[11].um_I.iw[15] ;
 wire \top_I.branch[19].block[11].um_I.iw[16] ;
 wire \top_I.branch[19].block[11].um_I.iw[17] ;
 wire \top_I.branch[19].block[11].um_I.iw[1] ;
 wire \top_I.branch[19].block[11].um_I.iw[2] ;
 wire \top_I.branch[19].block[11].um_I.iw[3] ;
 wire \top_I.branch[19].block[11].um_I.iw[4] ;
 wire \top_I.branch[19].block[11].um_I.iw[5] ;
 wire \top_I.branch[19].block[11].um_I.iw[6] ;
 wire \top_I.branch[19].block[11].um_I.iw[7] ;
 wire \top_I.branch[19].block[11].um_I.iw[8] ;
 wire \top_I.branch[19].block[11].um_I.iw[9] ;
 wire \top_I.branch[19].block[11].um_I.k_zero ;
 wire \top_I.branch[19].block[11].um_I.pg_vdd ;
 wire \top_I.branch[19].block[12].um_I.ana[2] ;
 wire \top_I.branch[19].block[12].um_I.ana[3] ;
 wire \top_I.branch[19].block[12].um_I.ana[4] ;
 wire \top_I.branch[19].block[12].um_I.ana[5] ;
 wire \top_I.branch[19].block[12].um_I.ana[6] ;
 wire \top_I.branch[19].block[12].um_I.ana[7] ;
 wire \top_I.branch[19].block[12].um_I.clk ;
 wire \top_I.branch[19].block[12].um_I.ena ;
 wire \top_I.branch[19].block[12].um_I.iw[10] ;
 wire \top_I.branch[19].block[12].um_I.iw[11] ;
 wire \top_I.branch[19].block[12].um_I.iw[12] ;
 wire \top_I.branch[19].block[12].um_I.iw[13] ;
 wire \top_I.branch[19].block[12].um_I.iw[14] ;
 wire \top_I.branch[19].block[12].um_I.iw[15] ;
 wire \top_I.branch[19].block[12].um_I.iw[16] ;
 wire \top_I.branch[19].block[12].um_I.iw[17] ;
 wire \top_I.branch[19].block[12].um_I.iw[1] ;
 wire \top_I.branch[19].block[12].um_I.iw[2] ;
 wire \top_I.branch[19].block[12].um_I.iw[3] ;
 wire \top_I.branch[19].block[12].um_I.iw[4] ;
 wire \top_I.branch[19].block[12].um_I.iw[5] ;
 wire \top_I.branch[19].block[12].um_I.iw[6] ;
 wire \top_I.branch[19].block[12].um_I.iw[7] ;
 wire \top_I.branch[19].block[12].um_I.iw[8] ;
 wire \top_I.branch[19].block[12].um_I.iw[9] ;
 wire \top_I.branch[19].block[12].um_I.k_zero ;
 wire \top_I.branch[19].block[12].um_I.pg_vdd ;
 wire \top_I.branch[19].block[13].um_I.ana[2] ;
 wire \top_I.branch[19].block[13].um_I.ana[3] ;
 wire \top_I.branch[19].block[13].um_I.ana[4] ;
 wire \top_I.branch[19].block[13].um_I.ana[5] ;
 wire \top_I.branch[19].block[13].um_I.ana[6] ;
 wire \top_I.branch[19].block[13].um_I.ana[7] ;
 wire \top_I.branch[19].block[13].um_I.clk ;
 wire \top_I.branch[19].block[13].um_I.ena ;
 wire \top_I.branch[19].block[13].um_I.iw[10] ;
 wire \top_I.branch[19].block[13].um_I.iw[11] ;
 wire \top_I.branch[19].block[13].um_I.iw[12] ;
 wire \top_I.branch[19].block[13].um_I.iw[13] ;
 wire \top_I.branch[19].block[13].um_I.iw[14] ;
 wire \top_I.branch[19].block[13].um_I.iw[15] ;
 wire \top_I.branch[19].block[13].um_I.iw[16] ;
 wire \top_I.branch[19].block[13].um_I.iw[17] ;
 wire \top_I.branch[19].block[13].um_I.iw[1] ;
 wire \top_I.branch[19].block[13].um_I.iw[2] ;
 wire \top_I.branch[19].block[13].um_I.iw[3] ;
 wire \top_I.branch[19].block[13].um_I.iw[4] ;
 wire \top_I.branch[19].block[13].um_I.iw[5] ;
 wire \top_I.branch[19].block[13].um_I.iw[6] ;
 wire \top_I.branch[19].block[13].um_I.iw[7] ;
 wire \top_I.branch[19].block[13].um_I.iw[8] ;
 wire \top_I.branch[19].block[13].um_I.iw[9] ;
 wire \top_I.branch[19].block[13].um_I.k_zero ;
 wire \top_I.branch[19].block[13].um_I.pg_vdd ;
 wire \top_I.branch[19].block[14].um_I.ana[2] ;
 wire \top_I.branch[19].block[14].um_I.ana[3] ;
 wire \top_I.branch[19].block[14].um_I.ana[4] ;
 wire \top_I.branch[19].block[14].um_I.ana[5] ;
 wire \top_I.branch[19].block[14].um_I.ana[6] ;
 wire \top_I.branch[19].block[14].um_I.ana[7] ;
 wire \top_I.branch[19].block[14].um_I.clk ;
 wire \top_I.branch[19].block[14].um_I.ena ;
 wire \top_I.branch[19].block[14].um_I.iw[10] ;
 wire \top_I.branch[19].block[14].um_I.iw[11] ;
 wire \top_I.branch[19].block[14].um_I.iw[12] ;
 wire \top_I.branch[19].block[14].um_I.iw[13] ;
 wire \top_I.branch[19].block[14].um_I.iw[14] ;
 wire \top_I.branch[19].block[14].um_I.iw[15] ;
 wire \top_I.branch[19].block[14].um_I.iw[16] ;
 wire \top_I.branch[19].block[14].um_I.iw[17] ;
 wire \top_I.branch[19].block[14].um_I.iw[1] ;
 wire \top_I.branch[19].block[14].um_I.iw[2] ;
 wire \top_I.branch[19].block[14].um_I.iw[3] ;
 wire \top_I.branch[19].block[14].um_I.iw[4] ;
 wire \top_I.branch[19].block[14].um_I.iw[5] ;
 wire \top_I.branch[19].block[14].um_I.iw[6] ;
 wire \top_I.branch[19].block[14].um_I.iw[7] ;
 wire \top_I.branch[19].block[14].um_I.iw[8] ;
 wire \top_I.branch[19].block[14].um_I.iw[9] ;
 wire \top_I.branch[19].block[14].um_I.k_zero ;
 wire \top_I.branch[19].block[14].um_I.pg_vdd ;
 wire \top_I.branch[19].block[15].um_I.ana[2] ;
 wire \top_I.branch[19].block[15].um_I.ana[3] ;
 wire \top_I.branch[19].block[15].um_I.ana[4] ;
 wire \top_I.branch[19].block[15].um_I.ana[5] ;
 wire \top_I.branch[19].block[15].um_I.ana[6] ;
 wire \top_I.branch[19].block[15].um_I.ana[7] ;
 wire \top_I.branch[19].block[15].um_I.clk ;
 wire \top_I.branch[19].block[15].um_I.ena ;
 wire \top_I.branch[19].block[15].um_I.iw[10] ;
 wire \top_I.branch[19].block[15].um_I.iw[11] ;
 wire \top_I.branch[19].block[15].um_I.iw[12] ;
 wire \top_I.branch[19].block[15].um_I.iw[13] ;
 wire \top_I.branch[19].block[15].um_I.iw[14] ;
 wire \top_I.branch[19].block[15].um_I.iw[15] ;
 wire \top_I.branch[19].block[15].um_I.iw[16] ;
 wire \top_I.branch[19].block[15].um_I.iw[17] ;
 wire \top_I.branch[19].block[15].um_I.iw[1] ;
 wire \top_I.branch[19].block[15].um_I.iw[2] ;
 wire \top_I.branch[19].block[15].um_I.iw[3] ;
 wire \top_I.branch[19].block[15].um_I.iw[4] ;
 wire \top_I.branch[19].block[15].um_I.iw[5] ;
 wire \top_I.branch[19].block[15].um_I.iw[6] ;
 wire \top_I.branch[19].block[15].um_I.iw[7] ;
 wire \top_I.branch[19].block[15].um_I.iw[8] ;
 wire \top_I.branch[19].block[15].um_I.iw[9] ;
 wire \top_I.branch[19].block[15].um_I.k_zero ;
 wire \top_I.branch[19].block[15].um_I.pg_vdd ;
 wire \top_I.branch[19].block[1].um_I.ana[2] ;
 wire \top_I.branch[19].block[1].um_I.ana[3] ;
 wire \top_I.branch[19].block[1].um_I.ana[4] ;
 wire \top_I.branch[19].block[1].um_I.ana[5] ;
 wire \top_I.branch[19].block[1].um_I.ana[6] ;
 wire \top_I.branch[19].block[1].um_I.ana[7] ;
 wire \top_I.branch[19].block[1].um_I.clk ;
 wire \top_I.branch[19].block[1].um_I.ena ;
 wire \top_I.branch[19].block[1].um_I.iw[10] ;
 wire \top_I.branch[19].block[1].um_I.iw[11] ;
 wire \top_I.branch[19].block[1].um_I.iw[12] ;
 wire \top_I.branch[19].block[1].um_I.iw[13] ;
 wire \top_I.branch[19].block[1].um_I.iw[14] ;
 wire \top_I.branch[19].block[1].um_I.iw[15] ;
 wire \top_I.branch[19].block[1].um_I.iw[16] ;
 wire \top_I.branch[19].block[1].um_I.iw[17] ;
 wire \top_I.branch[19].block[1].um_I.iw[1] ;
 wire \top_I.branch[19].block[1].um_I.iw[2] ;
 wire \top_I.branch[19].block[1].um_I.iw[3] ;
 wire \top_I.branch[19].block[1].um_I.iw[4] ;
 wire \top_I.branch[19].block[1].um_I.iw[5] ;
 wire \top_I.branch[19].block[1].um_I.iw[6] ;
 wire \top_I.branch[19].block[1].um_I.iw[7] ;
 wire \top_I.branch[19].block[1].um_I.iw[8] ;
 wire \top_I.branch[19].block[1].um_I.iw[9] ;
 wire \top_I.branch[19].block[1].um_I.k_zero ;
 wire \top_I.branch[19].block[1].um_I.pg_vdd ;
 wire \top_I.branch[19].block[2].um_I.ana[2] ;
 wire \top_I.branch[19].block[2].um_I.ana[3] ;
 wire \top_I.branch[19].block[2].um_I.ana[4] ;
 wire \top_I.branch[19].block[2].um_I.ana[5] ;
 wire \top_I.branch[19].block[2].um_I.ana[6] ;
 wire \top_I.branch[19].block[2].um_I.ana[7] ;
 wire \top_I.branch[19].block[2].um_I.clk ;
 wire \top_I.branch[19].block[2].um_I.ena ;
 wire \top_I.branch[19].block[2].um_I.iw[10] ;
 wire \top_I.branch[19].block[2].um_I.iw[11] ;
 wire \top_I.branch[19].block[2].um_I.iw[12] ;
 wire \top_I.branch[19].block[2].um_I.iw[13] ;
 wire \top_I.branch[19].block[2].um_I.iw[14] ;
 wire \top_I.branch[19].block[2].um_I.iw[15] ;
 wire \top_I.branch[19].block[2].um_I.iw[16] ;
 wire \top_I.branch[19].block[2].um_I.iw[17] ;
 wire \top_I.branch[19].block[2].um_I.iw[1] ;
 wire \top_I.branch[19].block[2].um_I.iw[2] ;
 wire \top_I.branch[19].block[2].um_I.iw[3] ;
 wire \top_I.branch[19].block[2].um_I.iw[4] ;
 wire \top_I.branch[19].block[2].um_I.iw[5] ;
 wire \top_I.branch[19].block[2].um_I.iw[6] ;
 wire \top_I.branch[19].block[2].um_I.iw[7] ;
 wire \top_I.branch[19].block[2].um_I.iw[8] ;
 wire \top_I.branch[19].block[2].um_I.iw[9] ;
 wire \top_I.branch[19].block[2].um_I.k_zero ;
 wire \top_I.branch[19].block[2].um_I.pg_vdd ;
 wire \top_I.branch[19].block[3].um_I.ana[2] ;
 wire \top_I.branch[19].block[3].um_I.ana[3] ;
 wire \top_I.branch[19].block[3].um_I.ana[4] ;
 wire \top_I.branch[19].block[3].um_I.ana[5] ;
 wire \top_I.branch[19].block[3].um_I.ana[6] ;
 wire \top_I.branch[19].block[3].um_I.ana[7] ;
 wire \top_I.branch[19].block[3].um_I.clk ;
 wire \top_I.branch[19].block[3].um_I.ena ;
 wire \top_I.branch[19].block[3].um_I.iw[10] ;
 wire \top_I.branch[19].block[3].um_I.iw[11] ;
 wire \top_I.branch[19].block[3].um_I.iw[12] ;
 wire \top_I.branch[19].block[3].um_I.iw[13] ;
 wire \top_I.branch[19].block[3].um_I.iw[14] ;
 wire \top_I.branch[19].block[3].um_I.iw[15] ;
 wire \top_I.branch[19].block[3].um_I.iw[16] ;
 wire \top_I.branch[19].block[3].um_I.iw[17] ;
 wire \top_I.branch[19].block[3].um_I.iw[1] ;
 wire \top_I.branch[19].block[3].um_I.iw[2] ;
 wire \top_I.branch[19].block[3].um_I.iw[3] ;
 wire \top_I.branch[19].block[3].um_I.iw[4] ;
 wire \top_I.branch[19].block[3].um_I.iw[5] ;
 wire \top_I.branch[19].block[3].um_I.iw[6] ;
 wire \top_I.branch[19].block[3].um_I.iw[7] ;
 wire \top_I.branch[19].block[3].um_I.iw[8] ;
 wire \top_I.branch[19].block[3].um_I.iw[9] ;
 wire \top_I.branch[19].block[3].um_I.k_zero ;
 wire \top_I.branch[19].block[3].um_I.pg_vdd ;
 wire \top_I.branch[19].block[4].um_I.ana[2] ;
 wire \top_I.branch[19].block[4].um_I.ana[3] ;
 wire \top_I.branch[19].block[4].um_I.ana[4] ;
 wire \top_I.branch[19].block[4].um_I.ana[5] ;
 wire \top_I.branch[19].block[4].um_I.ana[6] ;
 wire \top_I.branch[19].block[4].um_I.ana[7] ;
 wire \top_I.branch[19].block[4].um_I.clk ;
 wire \top_I.branch[19].block[4].um_I.ena ;
 wire \top_I.branch[19].block[4].um_I.iw[10] ;
 wire \top_I.branch[19].block[4].um_I.iw[11] ;
 wire \top_I.branch[19].block[4].um_I.iw[12] ;
 wire \top_I.branch[19].block[4].um_I.iw[13] ;
 wire \top_I.branch[19].block[4].um_I.iw[14] ;
 wire \top_I.branch[19].block[4].um_I.iw[15] ;
 wire \top_I.branch[19].block[4].um_I.iw[16] ;
 wire \top_I.branch[19].block[4].um_I.iw[17] ;
 wire \top_I.branch[19].block[4].um_I.iw[1] ;
 wire \top_I.branch[19].block[4].um_I.iw[2] ;
 wire \top_I.branch[19].block[4].um_I.iw[3] ;
 wire \top_I.branch[19].block[4].um_I.iw[4] ;
 wire \top_I.branch[19].block[4].um_I.iw[5] ;
 wire \top_I.branch[19].block[4].um_I.iw[6] ;
 wire \top_I.branch[19].block[4].um_I.iw[7] ;
 wire \top_I.branch[19].block[4].um_I.iw[8] ;
 wire \top_I.branch[19].block[4].um_I.iw[9] ;
 wire \top_I.branch[19].block[4].um_I.k_zero ;
 wire \top_I.branch[19].block[4].um_I.pg_vdd ;
 wire \top_I.branch[19].block[5].um_I.ana[2] ;
 wire \top_I.branch[19].block[5].um_I.ana[3] ;
 wire \top_I.branch[19].block[5].um_I.ana[4] ;
 wire \top_I.branch[19].block[5].um_I.ana[5] ;
 wire \top_I.branch[19].block[5].um_I.ana[6] ;
 wire \top_I.branch[19].block[5].um_I.ana[7] ;
 wire \top_I.branch[19].block[5].um_I.clk ;
 wire \top_I.branch[19].block[5].um_I.ena ;
 wire \top_I.branch[19].block[5].um_I.iw[10] ;
 wire \top_I.branch[19].block[5].um_I.iw[11] ;
 wire \top_I.branch[19].block[5].um_I.iw[12] ;
 wire \top_I.branch[19].block[5].um_I.iw[13] ;
 wire \top_I.branch[19].block[5].um_I.iw[14] ;
 wire \top_I.branch[19].block[5].um_I.iw[15] ;
 wire \top_I.branch[19].block[5].um_I.iw[16] ;
 wire \top_I.branch[19].block[5].um_I.iw[17] ;
 wire \top_I.branch[19].block[5].um_I.iw[1] ;
 wire \top_I.branch[19].block[5].um_I.iw[2] ;
 wire \top_I.branch[19].block[5].um_I.iw[3] ;
 wire \top_I.branch[19].block[5].um_I.iw[4] ;
 wire \top_I.branch[19].block[5].um_I.iw[5] ;
 wire \top_I.branch[19].block[5].um_I.iw[6] ;
 wire \top_I.branch[19].block[5].um_I.iw[7] ;
 wire \top_I.branch[19].block[5].um_I.iw[8] ;
 wire \top_I.branch[19].block[5].um_I.iw[9] ;
 wire \top_I.branch[19].block[5].um_I.k_zero ;
 wire \top_I.branch[19].block[5].um_I.pg_vdd ;
 wire \top_I.branch[19].block[6].um_I.ana[2] ;
 wire \top_I.branch[19].block[6].um_I.ana[3] ;
 wire \top_I.branch[19].block[6].um_I.ana[4] ;
 wire \top_I.branch[19].block[6].um_I.ana[5] ;
 wire \top_I.branch[19].block[6].um_I.ana[6] ;
 wire \top_I.branch[19].block[6].um_I.ana[7] ;
 wire \top_I.branch[19].block[6].um_I.clk ;
 wire \top_I.branch[19].block[6].um_I.ena ;
 wire \top_I.branch[19].block[6].um_I.iw[10] ;
 wire \top_I.branch[19].block[6].um_I.iw[11] ;
 wire \top_I.branch[19].block[6].um_I.iw[12] ;
 wire \top_I.branch[19].block[6].um_I.iw[13] ;
 wire \top_I.branch[19].block[6].um_I.iw[14] ;
 wire \top_I.branch[19].block[6].um_I.iw[15] ;
 wire \top_I.branch[19].block[6].um_I.iw[16] ;
 wire \top_I.branch[19].block[6].um_I.iw[17] ;
 wire \top_I.branch[19].block[6].um_I.iw[1] ;
 wire \top_I.branch[19].block[6].um_I.iw[2] ;
 wire \top_I.branch[19].block[6].um_I.iw[3] ;
 wire \top_I.branch[19].block[6].um_I.iw[4] ;
 wire \top_I.branch[19].block[6].um_I.iw[5] ;
 wire \top_I.branch[19].block[6].um_I.iw[6] ;
 wire \top_I.branch[19].block[6].um_I.iw[7] ;
 wire \top_I.branch[19].block[6].um_I.iw[8] ;
 wire \top_I.branch[19].block[6].um_I.iw[9] ;
 wire \top_I.branch[19].block[6].um_I.k_zero ;
 wire \top_I.branch[19].block[6].um_I.pg_vdd ;
 wire \top_I.branch[19].block[7].um_I.ana[2] ;
 wire \top_I.branch[19].block[7].um_I.ana[3] ;
 wire \top_I.branch[19].block[7].um_I.ana[4] ;
 wire \top_I.branch[19].block[7].um_I.ana[5] ;
 wire \top_I.branch[19].block[7].um_I.ana[6] ;
 wire \top_I.branch[19].block[7].um_I.ana[7] ;
 wire \top_I.branch[19].block[7].um_I.clk ;
 wire \top_I.branch[19].block[7].um_I.ena ;
 wire \top_I.branch[19].block[7].um_I.iw[10] ;
 wire \top_I.branch[19].block[7].um_I.iw[11] ;
 wire \top_I.branch[19].block[7].um_I.iw[12] ;
 wire \top_I.branch[19].block[7].um_I.iw[13] ;
 wire \top_I.branch[19].block[7].um_I.iw[14] ;
 wire \top_I.branch[19].block[7].um_I.iw[15] ;
 wire \top_I.branch[19].block[7].um_I.iw[16] ;
 wire \top_I.branch[19].block[7].um_I.iw[17] ;
 wire \top_I.branch[19].block[7].um_I.iw[1] ;
 wire \top_I.branch[19].block[7].um_I.iw[2] ;
 wire \top_I.branch[19].block[7].um_I.iw[3] ;
 wire \top_I.branch[19].block[7].um_I.iw[4] ;
 wire \top_I.branch[19].block[7].um_I.iw[5] ;
 wire \top_I.branch[19].block[7].um_I.iw[6] ;
 wire \top_I.branch[19].block[7].um_I.iw[7] ;
 wire \top_I.branch[19].block[7].um_I.iw[8] ;
 wire \top_I.branch[19].block[7].um_I.iw[9] ;
 wire \top_I.branch[19].block[7].um_I.k_zero ;
 wire \top_I.branch[19].block[7].um_I.pg_vdd ;
 wire \top_I.branch[19].block[8].um_I.ana[2] ;
 wire \top_I.branch[19].block[8].um_I.ana[3] ;
 wire \top_I.branch[19].block[8].um_I.ana[4] ;
 wire \top_I.branch[19].block[8].um_I.ana[5] ;
 wire \top_I.branch[19].block[8].um_I.ana[6] ;
 wire \top_I.branch[19].block[8].um_I.ana[7] ;
 wire \top_I.branch[19].block[8].um_I.clk ;
 wire \top_I.branch[19].block[8].um_I.ena ;
 wire \top_I.branch[19].block[8].um_I.iw[10] ;
 wire \top_I.branch[19].block[8].um_I.iw[11] ;
 wire \top_I.branch[19].block[8].um_I.iw[12] ;
 wire \top_I.branch[19].block[8].um_I.iw[13] ;
 wire \top_I.branch[19].block[8].um_I.iw[14] ;
 wire \top_I.branch[19].block[8].um_I.iw[15] ;
 wire \top_I.branch[19].block[8].um_I.iw[16] ;
 wire \top_I.branch[19].block[8].um_I.iw[17] ;
 wire \top_I.branch[19].block[8].um_I.iw[1] ;
 wire \top_I.branch[19].block[8].um_I.iw[2] ;
 wire \top_I.branch[19].block[8].um_I.iw[3] ;
 wire \top_I.branch[19].block[8].um_I.iw[4] ;
 wire \top_I.branch[19].block[8].um_I.iw[5] ;
 wire \top_I.branch[19].block[8].um_I.iw[6] ;
 wire \top_I.branch[19].block[8].um_I.iw[7] ;
 wire \top_I.branch[19].block[8].um_I.iw[8] ;
 wire \top_I.branch[19].block[8].um_I.iw[9] ;
 wire \top_I.branch[19].block[8].um_I.k_zero ;
 wire \top_I.branch[19].block[8].um_I.pg_vdd ;
 wire \top_I.branch[19].block[9].um_I.ana[2] ;
 wire \top_I.branch[19].block[9].um_I.ana[3] ;
 wire \top_I.branch[19].block[9].um_I.ana[4] ;
 wire \top_I.branch[19].block[9].um_I.ana[5] ;
 wire \top_I.branch[19].block[9].um_I.ana[6] ;
 wire \top_I.branch[19].block[9].um_I.ana[7] ;
 wire \top_I.branch[19].block[9].um_I.clk ;
 wire \top_I.branch[19].block[9].um_I.ena ;
 wire \top_I.branch[19].block[9].um_I.iw[10] ;
 wire \top_I.branch[19].block[9].um_I.iw[11] ;
 wire \top_I.branch[19].block[9].um_I.iw[12] ;
 wire \top_I.branch[19].block[9].um_I.iw[13] ;
 wire \top_I.branch[19].block[9].um_I.iw[14] ;
 wire \top_I.branch[19].block[9].um_I.iw[15] ;
 wire \top_I.branch[19].block[9].um_I.iw[16] ;
 wire \top_I.branch[19].block[9].um_I.iw[17] ;
 wire \top_I.branch[19].block[9].um_I.iw[1] ;
 wire \top_I.branch[19].block[9].um_I.iw[2] ;
 wire \top_I.branch[19].block[9].um_I.iw[3] ;
 wire \top_I.branch[19].block[9].um_I.iw[4] ;
 wire \top_I.branch[19].block[9].um_I.iw[5] ;
 wire \top_I.branch[19].block[9].um_I.iw[6] ;
 wire \top_I.branch[19].block[9].um_I.iw[7] ;
 wire \top_I.branch[19].block[9].um_I.iw[8] ;
 wire \top_I.branch[19].block[9].um_I.iw[9] ;
 wire \top_I.branch[19].block[9].um_I.k_zero ;
 wire \top_I.branch[19].block[9].um_I.pg_vdd ;
 wire \top_I.branch[19].l_addr[0] ;
 wire \top_I.branch[19].l_addr[1] ;
 wire \top_I.branch[1].block[0].um_I.ana[2] ;
 wire \top_I.branch[1].block[0].um_I.ana[3] ;
 wire \top_I.branch[1].block[0].um_I.ana[4] ;
 wire \top_I.branch[1].block[0].um_I.ana[5] ;
 wire \top_I.branch[1].block[0].um_I.ana[6] ;
 wire \top_I.branch[1].block[0].um_I.ana[7] ;
 wire \top_I.branch[1].block[0].um_I.clk ;
 wire \top_I.branch[1].block[0].um_I.ena ;
 wire \top_I.branch[1].block[0].um_I.iw[10] ;
 wire \top_I.branch[1].block[0].um_I.iw[11] ;
 wire \top_I.branch[1].block[0].um_I.iw[12] ;
 wire \top_I.branch[1].block[0].um_I.iw[13] ;
 wire \top_I.branch[1].block[0].um_I.iw[14] ;
 wire \top_I.branch[1].block[0].um_I.iw[15] ;
 wire \top_I.branch[1].block[0].um_I.iw[16] ;
 wire \top_I.branch[1].block[0].um_I.iw[17] ;
 wire \top_I.branch[1].block[0].um_I.iw[1] ;
 wire \top_I.branch[1].block[0].um_I.iw[2] ;
 wire \top_I.branch[1].block[0].um_I.iw[3] ;
 wire \top_I.branch[1].block[0].um_I.iw[4] ;
 wire \top_I.branch[1].block[0].um_I.iw[5] ;
 wire \top_I.branch[1].block[0].um_I.iw[6] ;
 wire \top_I.branch[1].block[0].um_I.iw[7] ;
 wire \top_I.branch[1].block[0].um_I.iw[8] ;
 wire \top_I.branch[1].block[0].um_I.iw[9] ;
 wire \top_I.branch[1].block[0].um_I.k_zero ;
 wire \top_I.branch[1].block[0].um_I.pg_vdd ;
 wire \top_I.branch[1].block[10].um_I.ana[2] ;
 wire \top_I.branch[1].block[10].um_I.ana[3] ;
 wire \top_I.branch[1].block[10].um_I.ana[4] ;
 wire \top_I.branch[1].block[10].um_I.ana[5] ;
 wire \top_I.branch[1].block[10].um_I.ana[6] ;
 wire \top_I.branch[1].block[10].um_I.ana[7] ;
 wire \top_I.branch[1].block[10].um_I.clk ;
 wire \top_I.branch[1].block[10].um_I.ena ;
 wire \top_I.branch[1].block[10].um_I.iw[10] ;
 wire \top_I.branch[1].block[10].um_I.iw[11] ;
 wire \top_I.branch[1].block[10].um_I.iw[12] ;
 wire \top_I.branch[1].block[10].um_I.iw[13] ;
 wire \top_I.branch[1].block[10].um_I.iw[14] ;
 wire \top_I.branch[1].block[10].um_I.iw[15] ;
 wire \top_I.branch[1].block[10].um_I.iw[16] ;
 wire \top_I.branch[1].block[10].um_I.iw[17] ;
 wire \top_I.branch[1].block[10].um_I.iw[1] ;
 wire \top_I.branch[1].block[10].um_I.iw[2] ;
 wire \top_I.branch[1].block[10].um_I.iw[3] ;
 wire \top_I.branch[1].block[10].um_I.iw[4] ;
 wire \top_I.branch[1].block[10].um_I.iw[5] ;
 wire \top_I.branch[1].block[10].um_I.iw[6] ;
 wire \top_I.branch[1].block[10].um_I.iw[7] ;
 wire \top_I.branch[1].block[10].um_I.iw[8] ;
 wire \top_I.branch[1].block[10].um_I.iw[9] ;
 wire \top_I.branch[1].block[10].um_I.k_zero ;
 wire \top_I.branch[1].block[10].um_I.pg_vdd ;
 wire \top_I.branch[1].block[11].um_I.ana[2] ;
 wire \top_I.branch[1].block[11].um_I.ana[3] ;
 wire \top_I.branch[1].block[11].um_I.ana[4] ;
 wire \top_I.branch[1].block[11].um_I.ana[5] ;
 wire \top_I.branch[1].block[11].um_I.ana[6] ;
 wire \top_I.branch[1].block[11].um_I.ana[7] ;
 wire \top_I.branch[1].block[11].um_I.clk ;
 wire \top_I.branch[1].block[11].um_I.ena ;
 wire \top_I.branch[1].block[11].um_I.iw[10] ;
 wire \top_I.branch[1].block[11].um_I.iw[11] ;
 wire \top_I.branch[1].block[11].um_I.iw[12] ;
 wire \top_I.branch[1].block[11].um_I.iw[13] ;
 wire \top_I.branch[1].block[11].um_I.iw[14] ;
 wire \top_I.branch[1].block[11].um_I.iw[15] ;
 wire \top_I.branch[1].block[11].um_I.iw[16] ;
 wire \top_I.branch[1].block[11].um_I.iw[17] ;
 wire \top_I.branch[1].block[11].um_I.iw[1] ;
 wire \top_I.branch[1].block[11].um_I.iw[2] ;
 wire \top_I.branch[1].block[11].um_I.iw[3] ;
 wire \top_I.branch[1].block[11].um_I.iw[4] ;
 wire \top_I.branch[1].block[11].um_I.iw[5] ;
 wire \top_I.branch[1].block[11].um_I.iw[6] ;
 wire \top_I.branch[1].block[11].um_I.iw[7] ;
 wire \top_I.branch[1].block[11].um_I.iw[8] ;
 wire \top_I.branch[1].block[11].um_I.iw[9] ;
 wire \top_I.branch[1].block[11].um_I.k_zero ;
 wire \top_I.branch[1].block[11].um_I.pg_vdd ;
 wire \top_I.branch[1].block[12].um_I.ana[2] ;
 wire \top_I.branch[1].block[12].um_I.ana[3] ;
 wire \top_I.branch[1].block[12].um_I.ana[4] ;
 wire \top_I.branch[1].block[12].um_I.ana[5] ;
 wire \top_I.branch[1].block[12].um_I.ana[6] ;
 wire \top_I.branch[1].block[12].um_I.ana[7] ;
 wire \top_I.branch[1].block[12].um_I.clk ;
 wire \top_I.branch[1].block[12].um_I.ena ;
 wire \top_I.branch[1].block[12].um_I.iw[10] ;
 wire \top_I.branch[1].block[12].um_I.iw[11] ;
 wire \top_I.branch[1].block[12].um_I.iw[12] ;
 wire \top_I.branch[1].block[12].um_I.iw[13] ;
 wire \top_I.branch[1].block[12].um_I.iw[14] ;
 wire \top_I.branch[1].block[12].um_I.iw[15] ;
 wire \top_I.branch[1].block[12].um_I.iw[16] ;
 wire \top_I.branch[1].block[12].um_I.iw[17] ;
 wire \top_I.branch[1].block[12].um_I.iw[1] ;
 wire \top_I.branch[1].block[12].um_I.iw[2] ;
 wire \top_I.branch[1].block[12].um_I.iw[3] ;
 wire \top_I.branch[1].block[12].um_I.iw[4] ;
 wire \top_I.branch[1].block[12].um_I.iw[5] ;
 wire \top_I.branch[1].block[12].um_I.iw[6] ;
 wire \top_I.branch[1].block[12].um_I.iw[7] ;
 wire \top_I.branch[1].block[12].um_I.iw[8] ;
 wire \top_I.branch[1].block[12].um_I.iw[9] ;
 wire \top_I.branch[1].block[12].um_I.k_zero ;
 wire \top_I.branch[1].block[12].um_I.pg_vdd ;
 wire \top_I.branch[1].block[13].um_I.ana[2] ;
 wire \top_I.branch[1].block[13].um_I.ana[3] ;
 wire \top_I.branch[1].block[13].um_I.ana[4] ;
 wire \top_I.branch[1].block[13].um_I.ana[5] ;
 wire \top_I.branch[1].block[13].um_I.ana[6] ;
 wire \top_I.branch[1].block[13].um_I.ana[7] ;
 wire \top_I.branch[1].block[13].um_I.clk ;
 wire \top_I.branch[1].block[13].um_I.ena ;
 wire \top_I.branch[1].block[13].um_I.iw[10] ;
 wire \top_I.branch[1].block[13].um_I.iw[11] ;
 wire \top_I.branch[1].block[13].um_I.iw[12] ;
 wire \top_I.branch[1].block[13].um_I.iw[13] ;
 wire \top_I.branch[1].block[13].um_I.iw[14] ;
 wire \top_I.branch[1].block[13].um_I.iw[15] ;
 wire \top_I.branch[1].block[13].um_I.iw[16] ;
 wire \top_I.branch[1].block[13].um_I.iw[17] ;
 wire \top_I.branch[1].block[13].um_I.iw[1] ;
 wire \top_I.branch[1].block[13].um_I.iw[2] ;
 wire \top_I.branch[1].block[13].um_I.iw[3] ;
 wire \top_I.branch[1].block[13].um_I.iw[4] ;
 wire \top_I.branch[1].block[13].um_I.iw[5] ;
 wire \top_I.branch[1].block[13].um_I.iw[6] ;
 wire \top_I.branch[1].block[13].um_I.iw[7] ;
 wire \top_I.branch[1].block[13].um_I.iw[8] ;
 wire \top_I.branch[1].block[13].um_I.iw[9] ;
 wire \top_I.branch[1].block[13].um_I.k_zero ;
 wire \top_I.branch[1].block[13].um_I.pg_vdd ;
 wire \top_I.branch[1].block[14].um_I.ana[2] ;
 wire \top_I.branch[1].block[14].um_I.ana[3] ;
 wire \top_I.branch[1].block[14].um_I.ana[4] ;
 wire \top_I.branch[1].block[14].um_I.ana[5] ;
 wire \top_I.branch[1].block[14].um_I.ana[6] ;
 wire \top_I.branch[1].block[14].um_I.ana[7] ;
 wire \top_I.branch[1].block[14].um_I.clk ;
 wire \top_I.branch[1].block[14].um_I.ena ;
 wire \top_I.branch[1].block[14].um_I.iw[10] ;
 wire \top_I.branch[1].block[14].um_I.iw[11] ;
 wire \top_I.branch[1].block[14].um_I.iw[12] ;
 wire \top_I.branch[1].block[14].um_I.iw[13] ;
 wire \top_I.branch[1].block[14].um_I.iw[14] ;
 wire \top_I.branch[1].block[14].um_I.iw[15] ;
 wire \top_I.branch[1].block[14].um_I.iw[16] ;
 wire \top_I.branch[1].block[14].um_I.iw[17] ;
 wire \top_I.branch[1].block[14].um_I.iw[1] ;
 wire \top_I.branch[1].block[14].um_I.iw[2] ;
 wire \top_I.branch[1].block[14].um_I.iw[3] ;
 wire \top_I.branch[1].block[14].um_I.iw[4] ;
 wire \top_I.branch[1].block[14].um_I.iw[5] ;
 wire \top_I.branch[1].block[14].um_I.iw[6] ;
 wire \top_I.branch[1].block[14].um_I.iw[7] ;
 wire \top_I.branch[1].block[14].um_I.iw[8] ;
 wire \top_I.branch[1].block[14].um_I.iw[9] ;
 wire \top_I.branch[1].block[14].um_I.k_zero ;
 wire \top_I.branch[1].block[14].um_I.pg_vdd ;
 wire \top_I.branch[1].block[15].um_I.ana[2] ;
 wire \top_I.branch[1].block[15].um_I.ana[3] ;
 wire \top_I.branch[1].block[15].um_I.ana[4] ;
 wire \top_I.branch[1].block[15].um_I.ana[5] ;
 wire \top_I.branch[1].block[15].um_I.ana[6] ;
 wire \top_I.branch[1].block[15].um_I.ana[7] ;
 wire \top_I.branch[1].block[15].um_I.clk ;
 wire \top_I.branch[1].block[15].um_I.ena ;
 wire \top_I.branch[1].block[15].um_I.iw[10] ;
 wire \top_I.branch[1].block[15].um_I.iw[11] ;
 wire \top_I.branch[1].block[15].um_I.iw[12] ;
 wire \top_I.branch[1].block[15].um_I.iw[13] ;
 wire \top_I.branch[1].block[15].um_I.iw[14] ;
 wire \top_I.branch[1].block[15].um_I.iw[15] ;
 wire \top_I.branch[1].block[15].um_I.iw[16] ;
 wire \top_I.branch[1].block[15].um_I.iw[17] ;
 wire \top_I.branch[1].block[15].um_I.iw[1] ;
 wire \top_I.branch[1].block[15].um_I.iw[2] ;
 wire \top_I.branch[1].block[15].um_I.iw[3] ;
 wire \top_I.branch[1].block[15].um_I.iw[4] ;
 wire \top_I.branch[1].block[15].um_I.iw[5] ;
 wire \top_I.branch[1].block[15].um_I.iw[6] ;
 wire \top_I.branch[1].block[15].um_I.iw[7] ;
 wire \top_I.branch[1].block[15].um_I.iw[8] ;
 wire \top_I.branch[1].block[15].um_I.iw[9] ;
 wire \top_I.branch[1].block[15].um_I.k_zero ;
 wire \top_I.branch[1].block[15].um_I.pg_vdd ;
 wire \top_I.branch[1].block[1].um_I.ana[2] ;
 wire \top_I.branch[1].block[1].um_I.ana[3] ;
 wire \top_I.branch[1].block[1].um_I.ana[4] ;
 wire \top_I.branch[1].block[1].um_I.ana[5] ;
 wire \top_I.branch[1].block[1].um_I.ana[6] ;
 wire \top_I.branch[1].block[1].um_I.ana[7] ;
 wire \top_I.branch[1].block[1].um_I.clk ;
 wire \top_I.branch[1].block[1].um_I.ena ;
 wire \top_I.branch[1].block[1].um_I.iw[10] ;
 wire \top_I.branch[1].block[1].um_I.iw[11] ;
 wire \top_I.branch[1].block[1].um_I.iw[12] ;
 wire \top_I.branch[1].block[1].um_I.iw[13] ;
 wire \top_I.branch[1].block[1].um_I.iw[14] ;
 wire \top_I.branch[1].block[1].um_I.iw[15] ;
 wire \top_I.branch[1].block[1].um_I.iw[16] ;
 wire \top_I.branch[1].block[1].um_I.iw[17] ;
 wire \top_I.branch[1].block[1].um_I.iw[1] ;
 wire \top_I.branch[1].block[1].um_I.iw[2] ;
 wire \top_I.branch[1].block[1].um_I.iw[3] ;
 wire \top_I.branch[1].block[1].um_I.iw[4] ;
 wire \top_I.branch[1].block[1].um_I.iw[5] ;
 wire \top_I.branch[1].block[1].um_I.iw[6] ;
 wire \top_I.branch[1].block[1].um_I.iw[7] ;
 wire \top_I.branch[1].block[1].um_I.iw[8] ;
 wire \top_I.branch[1].block[1].um_I.iw[9] ;
 wire \top_I.branch[1].block[1].um_I.k_zero ;
 wire \top_I.branch[1].block[1].um_I.pg_vdd ;
 wire \top_I.branch[1].block[2].um_I.ana[2] ;
 wire \top_I.branch[1].block[2].um_I.ana[3] ;
 wire \top_I.branch[1].block[2].um_I.ana[4] ;
 wire \top_I.branch[1].block[2].um_I.ana[5] ;
 wire \top_I.branch[1].block[2].um_I.ana[6] ;
 wire \top_I.branch[1].block[2].um_I.ana[7] ;
 wire \top_I.branch[1].block[2].um_I.clk ;
 wire \top_I.branch[1].block[2].um_I.ena ;
 wire \top_I.branch[1].block[2].um_I.iw[10] ;
 wire \top_I.branch[1].block[2].um_I.iw[11] ;
 wire \top_I.branch[1].block[2].um_I.iw[12] ;
 wire \top_I.branch[1].block[2].um_I.iw[13] ;
 wire \top_I.branch[1].block[2].um_I.iw[14] ;
 wire \top_I.branch[1].block[2].um_I.iw[15] ;
 wire \top_I.branch[1].block[2].um_I.iw[16] ;
 wire \top_I.branch[1].block[2].um_I.iw[17] ;
 wire \top_I.branch[1].block[2].um_I.iw[1] ;
 wire \top_I.branch[1].block[2].um_I.iw[2] ;
 wire \top_I.branch[1].block[2].um_I.iw[3] ;
 wire \top_I.branch[1].block[2].um_I.iw[4] ;
 wire \top_I.branch[1].block[2].um_I.iw[5] ;
 wire \top_I.branch[1].block[2].um_I.iw[6] ;
 wire \top_I.branch[1].block[2].um_I.iw[7] ;
 wire \top_I.branch[1].block[2].um_I.iw[8] ;
 wire \top_I.branch[1].block[2].um_I.iw[9] ;
 wire \top_I.branch[1].block[2].um_I.k_zero ;
 wire \top_I.branch[1].block[2].um_I.pg_vdd ;
 wire \top_I.branch[1].block[3].um_I.ana[2] ;
 wire \top_I.branch[1].block[3].um_I.ana[3] ;
 wire \top_I.branch[1].block[3].um_I.ana[4] ;
 wire \top_I.branch[1].block[3].um_I.ana[5] ;
 wire \top_I.branch[1].block[3].um_I.ana[6] ;
 wire \top_I.branch[1].block[3].um_I.ana[7] ;
 wire \top_I.branch[1].block[3].um_I.clk ;
 wire \top_I.branch[1].block[3].um_I.ena ;
 wire \top_I.branch[1].block[3].um_I.iw[10] ;
 wire \top_I.branch[1].block[3].um_I.iw[11] ;
 wire \top_I.branch[1].block[3].um_I.iw[12] ;
 wire \top_I.branch[1].block[3].um_I.iw[13] ;
 wire \top_I.branch[1].block[3].um_I.iw[14] ;
 wire \top_I.branch[1].block[3].um_I.iw[15] ;
 wire \top_I.branch[1].block[3].um_I.iw[16] ;
 wire \top_I.branch[1].block[3].um_I.iw[17] ;
 wire \top_I.branch[1].block[3].um_I.iw[1] ;
 wire \top_I.branch[1].block[3].um_I.iw[2] ;
 wire \top_I.branch[1].block[3].um_I.iw[3] ;
 wire \top_I.branch[1].block[3].um_I.iw[4] ;
 wire \top_I.branch[1].block[3].um_I.iw[5] ;
 wire \top_I.branch[1].block[3].um_I.iw[6] ;
 wire \top_I.branch[1].block[3].um_I.iw[7] ;
 wire \top_I.branch[1].block[3].um_I.iw[8] ;
 wire \top_I.branch[1].block[3].um_I.iw[9] ;
 wire \top_I.branch[1].block[3].um_I.k_zero ;
 wire \top_I.branch[1].block[3].um_I.pg_vdd ;
 wire \top_I.branch[1].block[4].um_I.ana[2] ;
 wire \top_I.branch[1].block[4].um_I.ana[3] ;
 wire \top_I.branch[1].block[4].um_I.ana[4] ;
 wire \top_I.branch[1].block[4].um_I.ana[5] ;
 wire \top_I.branch[1].block[4].um_I.ana[6] ;
 wire \top_I.branch[1].block[4].um_I.ana[7] ;
 wire \top_I.branch[1].block[4].um_I.clk ;
 wire \top_I.branch[1].block[4].um_I.ena ;
 wire \top_I.branch[1].block[4].um_I.iw[10] ;
 wire \top_I.branch[1].block[4].um_I.iw[11] ;
 wire \top_I.branch[1].block[4].um_I.iw[12] ;
 wire \top_I.branch[1].block[4].um_I.iw[13] ;
 wire \top_I.branch[1].block[4].um_I.iw[14] ;
 wire \top_I.branch[1].block[4].um_I.iw[15] ;
 wire \top_I.branch[1].block[4].um_I.iw[16] ;
 wire \top_I.branch[1].block[4].um_I.iw[17] ;
 wire \top_I.branch[1].block[4].um_I.iw[1] ;
 wire \top_I.branch[1].block[4].um_I.iw[2] ;
 wire \top_I.branch[1].block[4].um_I.iw[3] ;
 wire \top_I.branch[1].block[4].um_I.iw[4] ;
 wire \top_I.branch[1].block[4].um_I.iw[5] ;
 wire \top_I.branch[1].block[4].um_I.iw[6] ;
 wire \top_I.branch[1].block[4].um_I.iw[7] ;
 wire \top_I.branch[1].block[4].um_I.iw[8] ;
 wire \top_I.branch[1].block[4].um_I.iw[9] ;
 wire \top_I.branch[1].block[4].um_I.k_zero ;
 wire \top_I.branch[1].block[4].um_I.pg_vdd ;
 wire \top_I.branch[1].block[5].um_I.ana[2] ;
 wire \top_I.branch[1].block[5].um_I.ana[3] ;
 wire \top_I.branch[1].block[5].um_I.ana[4] ;
 wire \top_I.branch[1].block[5].um_I.ana[5] ;
 wire \top_I.branch[1].block[5].um_I.ana[6] ;
 wire \top_I.branch[1].block[5].um_I.ana[7] ;
 wire \top_I.branch[1].block[5].um_I.clk ;
 wire \top_I.branch[1].block[5].um_I.ena ;
 wire \top_I.branch[1].block[5].um_I.iw[10] ;
 wire \top_I.branch[1].block[5].um_I.iw[11] ;
 wire \top_I.branch[1].block[5].um_I.iw[12] ;
 wire \top_I.branch[1].block[5].um_I.iw[13] ;
 wire \top_I.branch[1].block[5].um_I.iw[14] ;
 wire \top_I.branch[1].block[5].um_I.iw[15] ;
 wire \top_I.branch[1].block[5].um_I.iw[16] ;
 wire \top_I.branch[1].block[5].um_I.iw[17] ;
 wire \top_I.branch[1].block[5].um_I.iw[1] ;
 wire \top_I.branch[1].block[5].um_I.iw[2] ;
 wire \top_I.branch[1].block[5].um_I.iw[3] ;
 wire \top_I.branch[1].block[5].um_I.iw[4] ;
 wire \top_I.branch[1].block[5].um_I.iw[5] ;
 wire \top_I.branch[1].block[5].um_I.iw[6] ;
 wire \top_I.branch[1].block[5].um_I.iw[7] ;
 wire \top_I.branch[1].block[5].um_I.iw[8] ;
 wire \top_I.branch[1].block[5].um_I.iw[9] ;
 wire \top_I.branch[1].block[5].um_I.k_zero ;
 wire \top_I.branch[1].block[5].um_I.pg_vdd ;
 wire \top_I.branch[1].block[6].um_I.ana[2] ;
 wire \top_I.branch[1].block[6].um_I.ana[3] ;
 wire \top_I.branch[1].block[6].um_I.ana[4] ;
 wire \top_I.branch[1].block[6].um_I.ana[5] ;
 wire \top_I.branch[1].block[6].um_I.ana[6] ;
 wire \top_I.branch[1].block[6].um_I.ana[7] ;
 wire \top_I.branch[1].block[6].um_I.clk ;
 wire \top_I.branch[1].block[6].um_I.ena ;
 wire \top_I.branch[1].block[6].um_I.iw[10] ;
 wire \top_I.branch[1].block[6].um_I.iw[11] ;
 wire \top_I.branch[1].block[6].um_I.iw[12] ;
 wire \top_I.branch[1].block[6].um_I.iw[13] ;
 wire \top_I.branch[1].block[6].um_I.iw[14] ;
 wire \top_I.branch[1].block[6].um_I.iw[15] ;
 wire \top_I.branch[1].block[6].um_I.iw[16] ;
 wire \top_I.branch[1].block[6].um_I.iw[17] ;
 wire \top_I.branch[1].block[6].um_I.iw[1] ;
 wire \top_I.branch[1].block[6].um_I.iw[2] ;
 wire \top_I.branch[1].block[6].um_I.iw[3] ;
 wire \top_I.branch[1].block[6].um_I.iw[4] ;
 wire \top_I.branch[1].block[6].um_I.iw[5] ;
 wire \top_I.branch[1].block[6].um_I.iw[6] ;
 wire \top_I.branch[1].block[6].um_I.iw[7] ;
 wire \top_I.branch[1].block[6].um_I.iw[8] ;
 wire \top_I.branch[1].block[6].um_I.iw[9] ;
 wire \top_I.branch[1].block[6].um_I.k_zero ;
 wire \top_I.branch[1].block[6].um_I.pg_vdd ;
 wire \top_I.branch[1].block[7].um_I.ana[2] ;
 wire \top_I.branch[1].block[7].um_I.ana[3] ;
 wire \top_I.branch[1].block[7].um_I.ana[4] ;
 wire \top_I.branch[1].block[7].um_I.ana[5] ;
 wire \top_I.branch[1].block[7].um_I.ana[6] ;
 wire \top_I.branch[1].block[7].um_I.ana[7] ;
 wire \top_I.branch[1].block[7].um_I.clk ;
 wire \top_I.branch[1].block[7].um_I.ena ;
 wire \top_I.branch[1].block[7].um_I.iw[10] ;
 wire \top_I.branch[1].block[7].um_I.iw[11] ;
 wire \top_I.branch[1].block[7].um_I.iw[12] ;
 wire \top_I.branch[1].block[7].um_I.iw[13] ;
 wire \top_I.branch[1].block[7].um_I.iw[14] ;
 wire \top_I.branch[1].block[7].um_I.iw[15] ;
 wire \top_I.branch[1].block[7].um_I.iw[16] ;
 wire \top_I.branch[1].block[7].um_I.iw[17] ;
 wire \top_I.branch[1].block[7].um_I.iw[1] ;
 wire \top_I.branch[1].block[7].um_I.iw[2] ;
 wire \top_I.branch[1].block[7].um_I.iw[3] ;
 wire \top_I.branch[1].block[7].um_I.iw[4] ;
 wire \top_I.branch[1].block[7].um_I.iw[5] ;
 wire \top_I.branch[1].block[7].um_I.iw[6] ;
 wire \top_I.branch[1].block[7].um_I.iw[7] ;
 wire \top_I.branch[1].block[7].um_I.iw[8] ;
 wire \top_I.branch[1].block[7].um_I.iw[9] ;
 wire \top_I.branch[1].block[7].um_I.k_zero ;
 wire \top_I.branch[1].block[7].um_I.pg_vdd ;
 wire \top_I.branch[1].block[8].um_I.ana[2] ;
 wire \top_I.branch[1].block[8].um_I.ana[3] ;
 wire \top_I.branch[1].block[8].um_I.ana[4] ;
 wire \top_I.branch[1].block[8].um_I.ana[5] ;
 wire \top_I.branch[1].block[8].um_I.ana[6] ;
 wire \top_I.branch[1].block[8].um_I.ana[7] ;
 wire \top_I.branch[1].block[8].um_I.clk ;
 wire \top_I.branch[1].block[8].um_I.ena ;
 wire \top_I.branch[1].block[8].um_I.iw[10] ;
 wire \top_I.branch[1].block[8].um_I.iw[11] ;
 wire \top_I.branch[1].block[8].um_I.iw[12] ;
 wire \top_I.branch[1].block[8].um_I.iw[13] ;
 wire \top_I.branch[1].block[8].um_I.iw[14] ;
 wire \top_I.branch[1].block[8].um_I.iw[15] ;
 wire \top_I.branch[1].block[8].um_I.iw[16] ;
 wire \top_I.branch[1].block[8].um_I.iw[17] ;
 wire \top_I.branch[1].block[8].um_I.iw[1] ;
 wire \top_I.branch[1].block[8].um_I.iw[2] ;
 wire \top_I.branch[1].block[8].um_I.iw[3] ;
 wire \top_I.branch[1].block[8].um_I.iw[4] ;
 wire \top_I.branch[1].block[8].um_I.iw[5] ;
 wire \top_I.branch[1].block[8].um_I.iw[6] ;
 wire \top_I.branch[1].block[8].um_I.iw[7] ;
 wire \top_I.branch[1].block[8].um_I.iw[8] ;
 wire \top_I.branch[1].block[8].um_I.iw[9] ;
 wire \top_I.branch[1].block[8].um_I.k_zero ;
 wire \top_I.branch[1].block[8].um_I.pg_vdd ;
 wire \top_I.branch[1].block[9].um_I.ana[2] ;
 wire \top_I.branch[1].block[9].um_I.ana[3] ;
 wire \top_I.branch[1].block[9].um_I.ana[4] ;
 wire \top_I.branch[1].block[9].um_I.ana[5] ;
 wire \top_I.branch[1].block[9].um_I.ana[6] ;
 wire \top_I.branch[1].block[9].um_I.ana[7] ;
 wire \top_I.branch[1].block[9].um_I.clk ;
 wire \top_I.branch[1].block[9].um_I.ena ;
 wire \top_I.branch[1].block[9].um_I.iw[10] ;
 wire \top_I.branch[1].block[9].um_I.iw[11] ;
 wire \top_I.branch[1].block[9].um_I.iw[12] ;
 wire \top_I.branch[1].block[9].um_I.iw[13] ;
 wire \top_I.branch[1].block[9].um_I.iw[14] ;
 wire \top_I.branch[1].block[9].um_I.iw[15] ;
 wire \top_I.branch[1].block[9].um_I.iw[16] ;
 wire \top_I.branch[1].block[9].um_I.iw[17] ;
 wire \top_I.branch[1].block[9].um_I.iw[1] ;
 wire \top_I.branch[1].block[9].um_I.iw[2] ;
 wire \top_I.branch[1].block[9].um_I.iw[3] ;
 wire \top_I.branch[1].block[9].um_I.iw[4] ;
 wire \top_I.branch[1].block[9].um_I.iw[5] ;
 wire \top_I.branch[1].block[9].um_I.iw[6] ;
 wire \top_I.branch[1].block[9].um_I.iw[7] ;
 wire \top_I.branch[1].block[9].um_I.iw[8] ;
 wire \top_I.branch[1].block[9].um_I.iw[9] ;
 wire \top_I.branch[1].block[9].um_I.k_zero ;
 wire \top_I.branch[1].block[9].um_I.pg_vdd ;
 wire \top_I.branch[1].l_addr[0] ;
 wire \top_I.branch[1].l_k_one ;
 wire \top_I.branch[20].block[0].um_I.ana[2] ;
 wire \top_I.branch[20].block[0].um_I.ana[3] ;
 wire \top_I.branch[20].block[0].um_I.ana[4] ;
 wire \top_I.branch[20].block[0].um_I.ana[5] ;
 wire \top_I.branch[20].block[0].um_I.ana[6] ;
 wire \top_I.branch[20].block[0].um_I.ana[7] ;
 wire \top_I.branch[20].block[0].um_I.clk ;
 wire \top_I.branch[20].block[0].um_I.ena ;
 wire \top_I.branch[20].block[0].um_I.iw[10] ;
 wire \top_I.branch[20].block[0].um_I.iw[11] ;
 wire \top_I.branch[20].block[0].um_I.iw[12] ;
 wire \top_I.branch[20].block[0].um_I.iw[13] ;
 wire \top_I.branch[20].block[0].um_I.iw[14] ;
 wire \top_I.branch[20].block[0].um_I.iw[15] ;
 wire \top_I.branch[20].block[0].um_I.iw[16] ;
 wire \top_I.branch[20].block[0].um_I.iw[17] ;
 wire \top_I.branch[20].block[0].um_I.iw[1] ;
 wire \top_I.branch[20].block[0].um_I.iw[2] ;
 wire \top_I.branch[20].block[0].um_I.iw[3] ;
 wire \top_I.branch[20].block[0].um_I.iw[4] ;
 wire \top_I.branch[20].block[0].um_I.iw[5] ;
 wire \top_I.branch[20].block[0].um_I.iw[6] ;
 wire \top_I.branch[20].block[0].um_I.iw[7] ;
 wire \top_I.branch[20].block[0].um_I.iw[8] ;
 wire \top_I.branch[20].block[0].um_I.iw[9] ;
 wire \top_I.branch[20].block[0].um_I.k_zero ;
 wire \top_I.branch[20].block[0].um_I.pg_vdd ;
 wire \top_I.branch[20].block[10].um_I.ana[2] ;
 wire \top_I.branch[20].block[10].um_I.ana[3] ;
 wire \top_I.branch[20].block[10].um_I.ana[4] ;
 wire \top_I.branch[20].block[10].um_I.ana[5] ;
 wire \top_I.branch[20].block[10].um_I.ana[6] ;
 wire \top_I.branch[20].block[10].um_I.ana[7] ;
 wire \top_I.branch[20].block[10].um_I.clk ;
 wire \top_I.branch[20].block[10].um_I.ena ;
 wire \top_I.branch[20].block[10].um_I.iw[10] ;
 wire \top_I.branch[20].block[10].um_I.iw[11] ;
 wire \top_I.branch[20].block[10].um_I.iw[12] ;
 wire \top_I.branch[20].block[10].um_I.iw[13] ;
 wire \top_I.branch[20].block[10].um_I.iw[14] ;
 wire \top_I.branch[20].block[10].um_I.iw[15] ;
 wire \top_I.branch[20].block[10].um_I.iw[16] ;
 wire \top_I.branch[20].block[10].um_I.iw[17] ;
 wire \top_I.branch[20].block[10].um_I.iw[1] ;
 wire \top_I.branch[20].block[10].um_I.iw[2] ;
 wire \top_I.branch[20].block[10].um_I.iw[3] ;
 wire \top_I.branch[20].block[10].um_I.iw[4] ;
 wire \top_I.branch[20].block[10].um_I.iw[5] ;
 wire \top_I.branch[20].block[10].um_I.iw[6] ;
 wire \top_I.branch[20].block[10].um_I.iw[7] ;
 wire \top_I.branch[20].block[10].um_I.iw[8] ;
 wire \top_I.branch[20].block[10].um_I.iw[9] ;
 wire \top_I.branch[20].block[10].um_I.k_zero ;
 wire \top_I.branch[20].block[10].um_I.pg_vdd ;
 wire \top_I.branch[20].block[11].um_I.ana[2] ;
 wire \top_I.branch[20].block[11].um_I.ana[3] ;
 wire \top_I.branch[20].block[11].um_I.ana[4] ;
 wire \top_I.branch[20].block[11].um_I.ana[5] ;
 wire \top_I.branch[20].block[11].um_I.ana[6] ;
 wire \top_I.branch[20].block[11].um_I.ana[7] ;
 wire \top_I.branch[20].block[11].um_I.clk ;
 wire \top_I.branch[20].block[11].um_I.ena ;
 wire \top_I.branch[20].block[11].um_I.iw[10] ;
 wire \top_I.branch[20].block[11].um_I.iw[11] ;
 wire \top_I.branch[20].block[11].um_I.iw[12] ;
 wire \top_I.branch[20].block[11].um_I.iw[13] ;
 wire \top_I.branch[20].block[11].um_I.iw[14] ;
 wire \top_I.branch[20].block[11].um_I.iw[15] ;
 wire \top_I.branch[20].block[11].um_I.iw[16] ;
 wire \top_I.branch[20].block[11].um_I.iw[17] ;
 wire \top_I.branch[20].block[11].um_I.iw[1] ;
 wire \top_I.branch[20].block[11].um_I.iw[2] ;
 wire \top_I.branch[20].block[11].um_I.iw[3] ;
 wire \top_I.branch[20].block[11].um_I.iw[4] ;
 wire \top_I.branch[20].block[11].um_I.iw[5] ;
 wire \top_I.branch[20].block[11].um_I.iw[6] ;
 wire \top_I.branch[20].block[11].um_I.iw[7] ;
 wire \top_I.branch[20].block[11].um_I.iw[8] ;
 wire \top_I.branch[20].block[11].um_I.iw[9] ;
 wire \top_I.branch[20].block[11].um_I.k_zero ;
 wire \top_I.branch[20].block[11].um_I.pg_vdd ;
 wire \top_I.branch[20].block[12].um_I.ana[2] ;
 wire \top_I.branch[20].block[12].um_I.ana[3] ;
 wire \top_I.branch[20].block[12].um_I.ana[4] ;
 wire \top_I.branch[20].block[12].um_I.ana[5] ;
 wire \top_I.branch[20].block[12].um_I.ana[6] ;
 wire \top_I.branch[20].block[12].um_I.ana[7] ;
 wire \top_I.branch[20].block[12].um_I.clk ;
 wire \top_I.branch[20].block[12].um_I.ena ;
 wire \top_I.branch[20].block[12].um_I.iw[10] ;
 wire \top_I.branch[20].block[12].um_I.iw[11] ;
 wire \top_I.branch[20].block[12].um_I.iw[12] ;
 wire \top_I.branch[20].block[12].um_I.iw[13] ;
 wire \top_I.branch[20].block[12].um_I.iw[14] ;
 wire \top_I.branch[20].block[12].um_I.iw[15] ;
 wire \top_I.branch[20].block[12].um_I.iw[16] ;
 wire \top_I.branch[20].block[12].um_I.iw[17] ;
 wire \top_I.branch[20].block[12].um_I.iw[1] ;
 wire \top_I.branch[20].block[12].um_I.iw[2] ;
 wire \top_I.branch[20].block[12].um_I.iw[3] ;
 wire \top_I.branch[20].block[12].um_I.iw[4] ;
 wire \top_I.branch[20].block[12].um_I.iw[5] ;
 wire \top_I.branch[20].block[12].um_I.iw[6] ;
 wire \top_I.branch[20].block[12].um_I.iw[7] ;
 wire \top_I.branch[20].block[12].um_I.iw[8] ;
 wire \top_I.branch[20].block[12].um_I.iw[9] ;
 wire \top_I.branch[20].block[12].um_I.k_zero ;
 wire \top_I.branch[20].block[12].um_I.pg_vdd ;
 wire \top_I.branch[20].block[13].um_I.ana[2] ;
 wire \top_I.branch[20].block[13].um_I.ana[3] ;
 wire \top_I.branch[20].block[13].um_I.ana[4] ;
 wire \top_I.branch[20].block[13].um_I.ana[5] ;
 wire \top_I.branch[20].block[13].um_I.ana[6] ;
 wire \top_I.branch[20].block[13].um_I.ana[7] ;
 wire \top_I.branch[20].block[13].um_I.clk ;
 wire \top_I.branch[20].block[13].um_I.ena ;
 wire \top_I.branch[20].block[13].um_I.iw[10] ;
 wire \top_I.branch[20].block[13].um_I.iw[11] ;
 wire \top_I.branch[20].block[13].um_I.iw[12] ;
 wire \top_I.branch[20].block[13].um_I.iw[13] ;
 wire \top_I.branch[20].block[13].um_I.iw[14] ;
 wire \top_I.branch[20].block[13].um_I.iw[15] ;
 wire \top_I.branch[20].block[13].um_I.iw[16] ;
 wire \top_I.branch[20].block[13].um_I.iw[17] ;
 wire \top_I.branch[20].block[13].um_I.iw[1] ;
 wire \top_I.branch[20].block[13].um_I.iw[2] ;
 wire \top_I.branch[20].block[13].um_I.iw[3] ;
 wire \top_I.branch[20].block[13].um_I.iw[4] ;
 wire \top_I.branch[20].block[13].um_I.iw[5] ;
 wire \top_I.branch[20].block[13].um_I.iw[6] ;
 wire \top_I.branch[20].block[13].um_I.iw[7] ;
 wire \top_I.branch[20].block[13].um_I.iw[8] ;
 wire \top_I.branch[20].block[13].um_I.iw[9] ;
 wire \top_I.branch[20].block[13].um_I.k_zero ;
 wire \top_I.branch[20].block[13].um_I.pg_vdd ;
 wire \top_I.branch[20].block[14].um_I.ana[2] ;
 wire \top_I.branch[20].block[14].um_I.ana[3] ;
 wire \top_I.branch[20].block[14].um_I.ana[4] ;
 wire \top_I.branch[20].block[14].um_I.ana[5] ;
 wire \top_I.branch[20].block[14].um_I.ana[6] ;
 wire \top_I.branch[20].block[14].um_I.ana[7] ;
 wire \top_I.branch[20].block[14].um_I.clk ;
 wire \top_I.branch[20].block[14].um_I.ena ;
 wire \top_I.branch[20].block[14].um_I.iw[10] ;
 wire \top_I.branch[20].block[14].um_I.iw[11] ;
 wire \top_I.branch[20].block[14].um_I.iw[12] ;
 wire \top_I.branch[20].block[14].um_I.iw[13] ;
 wire \top_I.branch[20].block[14].um_I.iw[14] ;
 wire \top_I.branch[20].block[14].um_I.iw[15] ;
 wire \top_I.branch[20].block[14].um_I.iw[16] ;
 wire \top_I.branch[20].block[14].um_I.iw[17] ;
 wire \top_I.branch[20].block[14].um_I.iw[1] ;
 wire \top_I.branch[20].block[14].um_I.iw[2] ;
 wire \top_I.branch[20].block[14].um_I.iw[3] ;
 wire \top_I.branch[20].block[14].um_I.iw[4] ;
 wire \top_I.branch[20].block[14].um_I.iw[5] ;
 wire \top_I.branch[20].block[14].um_I.iw[6] ;
 wire \top_I.branch[20].block[14].um_I.iw[7] ;
 wire \top_I.branch[20].block[14].um_I.iw[8] ;
 wire \top_I.branch[20].block[14].um_I.iw[9] ;
 wire \top_I.branch[20].block[14].um_I.k_zero ;
 wire \top_I.branch[20].block[14].um_I.ow[0] ;
 wire \top_I.branch[20].block[14].um_I.ow[10] ;
 wire \top_I.branch[20].block[14].um_I.ow[11] ;
 wire \top_I.branch[20].block[14].um_I.ow[12] ;
 wire \top_I.branch[20].block[14].um_I.ow[13] ;
 wire \top_I.branch[20].block[14].um_I.ow[14] ;
 wire \top_I.branch[20].block[14].um_I.ow[15] ;
 wire \top_I.branch[20].block[14].um_I.ow[16] ;
 wire \top_I.branch[20].block[14].um_I.ow[17] ;
 wire \top_I.branch[20].block[14].um_I.ow[18] ;
 wire \top_I.branch[20].block[14].um_I.ow[19] ;
 wire \top_I.branch[20].block[14].um_I.ow[1] ;
 wire \top_I.branch[20].block[14].um_I.ow[20] ;
 wire \top_I.branch[20].block[14].um_I.ow[21] ;
 wire \top_I.branch[20].block[14].um_I.ow[22] ;
 wire \top_I.branch[20].block[14].um_I.ow[23] ;
 wire \top_I.branch[20].block[14].um_I.ow[2] ;
 wire \top_I.branch[20].block[14].um_I.ow[3] ;
 wire \top_I.branch[20].block[14].um_I.ow[4] ;
 wire \top_I.branch[20].block[14].um_I.ow[5] ;
 wire \top_I.branch[20].block[14].um_I.ow[6] ;
 wire \top_I.branch[20].block[14].um_I.ow[7] ;
 wire \top_I.branch[20].block[14].um_I.ow[8] ;
 wire \top_I.branch[20].block[14].um_I.ow[9] ;
 wire \top_I.branch[20].block[14].um_I.pg_vdd ;
 wire \top_I.branch[20].block[15].um_I.ana[2] ;
 wire \top_I.branch[20].block[15].um_I.ana[3] ;
 wire \top_I.branch[20].block[15].um_I.ana[4] ;
 wire \top_I.branch[20].block[15].um_I.ana[5] ;
 wire \top_I.branch[20].block[15].um_I.ana[6] ;
 wire \top_I.branch[20].block[15].um_I.ana[7] ;
 wire \top_I.branch[20].block[15].um_I.clk ;
 wire \top_I.branch[20].block[15].um_I.ena ;
 wire \top_I.branch[20].block[15].um_I.iw[10] ;
 wire \top_I.branch[20].block[15].um_I.iw[11] ;
 wire \top_I.branch[20].block[15].um_I.iw[12] ;
 wire \top_I.branch[20].block[15].um_I.iw[13] ;
 wire \top_I.branch[20].block[15].um_I.iw[14] ;
 wire \top_I.branch[20].block[15].um_I.iw[15] ;
 wire \top_I.branch[20].block[15].um_I.iw[16] ;
 wire \top_I.branch[20].block[15].um_I.iw[17] ;
 wire \top_I.branch[20].block[15].um_I.iw[1] ;
 wire \top_I.branch[20].block[15].um_I.iw[2] ;
 wire \top_I.branch[20].block[15].um_I.iw[3] ;
 wire \top_I.branch[20].block[15].um_I.iw[4] ;
 wire \top_I.branch[20].block[15].um_I.iw[5] ;
 wire \top_I.branch[20].block[15].um_I.iw[6] ;
 wire \top_I.branch[20].block[15].um_I.iw[7] ;
 wire \top_I.branch[20].block[15].um_I.iw[8] ;
 wire \top_I.branch[20].block[15].um_I.iw[9] ;
 wire \top_I.branch[20].block[15].um_I.k_zero ;
 wire \top_I.branch[20].block[15].um_I.pg_vdd ;
 wire \top_I.branch[20].block[1].um_I.ana[2] ;
 wire \top_I.branch[20].block[1].um_I.ana[3] ;
 wire \top_I.branch[20].block[1].um_I.ana[4] ;
 wire \top_I.branch[20].block[1].um_I.ana[5] ;
 wire \top_I.branch[20].block[1].um_I.ana[6] ;
 wire \top_I.branch[20].block[1].um_I.ana[7] ;
 wire \top_I.branch[20].block[1].um_I.clk ;
 wire \top_I.branch[20].block[1].um_I.ena ;
 wire \top_I.branch[20].block[1].um_I.iw[10] ;
 wire \top_I.branch[20].block[1].um_I.iw[11] ;
 wire \top_I.branch[20].block[1].um_I.iw[12] ;
 wire \top_I.branch[20].block[1].um_I.iw[13] ;
 wire \top_I.branch[20].block[1].um_I.iw[14] ;
 wire \top_I.branch[20].block[1].um_I.iw[15] ;
 wire \top_I.branch[20].block[1].um_I.iw[16] ;
 wire \top_I.branch[20].block[1].um_I.iw[17] ;
 wire \top_I.branch[20].block[1].um_I.iw[1] ;
 wire \top_I.branch[20].block[1].um_I.iw[2] ;
 wire \top_I.branch[20].block[1].um_I.iw[3] ;
 wire \top_I.branch[20].block[1].um_I.iw[4] ;
 wire \top_I.branch[20].block[1].um_I.iw[5] ;
 wire \top_I.branch[20].block[1].um_I.iw[6] ;
 wire \top_I.branch[20].block[1].um_I.iw[7] ;
 wire \top_I.branch[20].block[1].um_I.iw[8] ;
 wire \top_I.branch[20].block[1].um_I.iw[9] ;
 wire \top_I.branch[20].block[1].um_I.k_zero ;
 wire \top_I.branch[20].block[1].um_I.pg_vdd ;
 wire \top_I.branch[20].block[2].um_I.ana[2] ;
 wire \top_I.branch[20].block[2].um_I.ana[3] ;
 wire \top_I.branch[20].block[2].um_I.ana[4] ;
 wire \top_I.branch[20].block[2].um_I.ana[5] ;
 wire \top_I.branch[20].block[2].um_I.ana[6] ;
 wire \top_I.branch[20].block[2].um_I.ana[7] ;
 wire \top_I.branch[20].block[2].um_I.clk ;
 wire \top_I.branch[20].block[2].um_I.ena ;
 wire \top_I.branch[20].block[2].um_I.iw[10] ;
 wire \top_I.branch[20].block[2].um_I.iw[11] ;
 wire \top_I.branch[20].block[2].um_I.iw[12] ;
 wire \top_I.branch[20].block[2].um_I.iw[13] ;
 wire \top_I.branch[20].block[2].um_I.iw[14] ;
 wire \top_I.branch[20].block[2].um_I.iw[15] ;
 wire \top_I.branch[20].block[2].um_I.iw[16] ;
 wire \top_I.branch[20].block[2].um_I.iw[17] ;
 wire \top_I.branch[20].block[2].um_I.iw[1] ;
 wire \top_I.branch[20].block[2].um_I.iw[2] ;
 wire \top_I.branch[20].block[2].um_I.iw[3] ;
 wire \top_I.branch[20].block[2].um_I.iw[4] ;
 wire \top_I.branch[20].block[2].um_I.iw[5] ;
 wire \top_I.branch[20].block[2].um_I.iw[6] ;
 wire \top_I.branch[20].block[2].um_I.iw[7] ;
 wire \top_I.branch[20].block[2].um_I.iw[8] ;
 wire \top_I.branch[20].block[2].um_I.iw[9] ;
 wire \top_I.branch[20].block[2].um_I.k_zero ;
 wire \top_I.branch[20].block[2].um_I.pg_vdd ;
 wire \top_I.branch[20].block[3].um_I.ana[2] ;
 wire \top_I.branch[20].block[3].um_I.ana[3] ;
 wire \top_I.branch[20].block[3].um_I.ana[4] ;
 wire \top_I.branch[20].block[3].um_I.ana[5] ;
 wire \top_I.branch[20].block[3].um_I.ana[6] ;
 wire \top_I.branch[20].block[3].um_I.ana[7] ;
 wire \top_I.branch[20].block[3].um_I.clk ;
 wire \top_I.branch[20].block[3].um_I.ena ;
 wire \top_I.branch[20].block[3].um_I.iw[10] ;
 wire \top_I.branch[20].block[3].um_I.iw[11] ;
 wire \top_I.branch[20].block[3].um_I.iw[12] ;
 wire \top_I.branch[20].block[3].um_I.iw[13] ;
 wire \top_I.branch[20].block[3].um_I.iw[14] ;
 wire \top_I.branch[20].block[3].um_I.iw[15] ;
 wire \top_I.branch[20].block[3].um_I.iw[16] ;
 wire \top_I.branch[20].block[3].um_I.iw[17] ;
 wire \top_I.branch[20].block[3].um_I.iw[1] ;
 wire \top_I.branch[20].block[3].um_I.iw[2] ;
 wire \top_I.branch[20].block[3].um_I.iw[3] ;
 wire \top_I.branch[20].block[3].um_I.iw[4] ;
 wire \top_I.branch[20].block[3].um_I.iw[5] ;
 wire \top_I.branch[20].block[3].um_I.iw[6] ;
 wire \top_I.branch[20].block[3].um_I.iw[7] ;
 wire \top_I.branch[20].block[3].um_I.iw[8] ;
 wire \top_I.branch[20].block[3].um_I.iw[9] ;
 wire \top_I.branch[20].block[3].um_I.k_zero ;
 wire \top_I.branch[20].block[3].um_I.pg_vdd ;
 wire \top_I.branch[20].block[4].um_I.ana[2] ;
 wire \top_I.branch[20].block[4].um_I.ana[3] ;
 wire \top_I.branch[20].block[4].um_I.ana[4] ;
 wire \top_I.branch[20].block[4].um_I.ana[5] ;
 wire \top_I.branch[20].block[4].um_I.ana[6] ;
 wire \top_I.branch[20].block[4].um_I.ana[7] ;
 wire \top_I.branch[20].block[4].um_I.clk ;
 wire \top_I.branch[20].block[4].um_I.ena ;
 wire \top_I.branch[20].block[4].um_I.iw[10] ;
 wire \top_I.branch[20].block[4].um_I.iw[11] ;
 wire \top_I.branch[20].block[4].um_I.iw[12] ;
 wire \top_I.branch[20].block[4].um_I.iw[13] ;
 wire \top_I.branch[20].block[4].um_I.iw[14] ;
 wire \top_I.branch[20].block[4].um_I.iw[15] ;
 wire \top_I.branch[20].block[4].um_I.iw[16] ;
 wire \top_I.branch[20].block[4].um_I.iw[17] ;
 wire \top_I.branch[20].block[4].um_I.iw[1] ;
 wire \top_I.branch[20].block[4].um_I.iw[2] ;
 wire \top_I.branch[20].block[4].um_I.iw[3] ;
 wire \top_I.branch[20].block[4].um_I.iw[4] ;
 wire \top_I.branch[20].block[4].um_I.iw[5] ;
 wire \top_I.branch[20].block[4].um_I.iw[6] ;
 wire \top_I.branch[20].block[4].um_I.iw[7] ;
 wire \top_I.branch[20].block[4].um_I.iw[8] ;
 wire \top_I.branch[20].block[4].um_I.iw[9] ;
 wire \top_I.branch[20].block[4].um_I.k_zero ;
 wire \top_I.branch[20].block[4].um_I.pg_vdd ;
 wire \top_I.branch[20].block[5].um_I.ana[2] ;
 wire \top_I.branch[20].block[5].um_I.ana[3] ;
 wire \top_I.branch[20].block[5].um_I.ana[4] ;
 wire \top_I.branch[20].block[5].um_I.ana[5] ;
 wire \top_I.branch[20].block[5].um_I.ana[6] ;
 wire \top_I.branch[20].block[5].um_I.ana[7] ;
 wire \top_I.branch[20].block[5].um_I.clk ;
 wire \top_I.branch[20].block[5].um_I.ena ;
 wire \top_I.branch[20].block[5].um_I.iw[10] ;
 wire \top_I.branch[20].block[5].um_I.iw[11] ;
 wire \top_I.branch[20].block[5].um_I.iw[12] ;
 wire \top_I.branch[20].block[5].um_I.iw[13] ;
 wire \top_I.branch[20].block[5].um_I.iw[14] ;
 wire \top_I.branch[20].block[5].um_I.iw[15] ;
 wire \top_I.branch[20].block[5].um_I.iw[16] ;
 wire \top_I.branch[20].block[5].um_I.iw[17] ;
 wire \top_I.branch[20].block[5].um_I.iw[1] ;
 wire \top_I.branch[20].block[5].um_I.iw[2] ;
 wire \top_I.branch[20].block[5].um_I.iw[3] ;
 wire \top_I.branch[20].block[5].um_I.iw[4] ;
 wire \top_I.branch[20].block[5].um_I.iw[5] ;
 wire \top_I.branch[20].block[5].um_I.iw[6] ;
 wire \top_I.branch[20].block[5].um_I.iw[7] ;
 wire \top_I.branch[20].block[5].um_I.iw[8] ;
 wire \top_I.branch[20].block[5].um_I.iw[9] ;
 wire \top_I.branch[20].block[5].um_I.k_zero ;
 wire \top_I.branch[20].block[5].um_I.pg_vdd ;
 wire \top_I.branch[20].block[6].um_I.ana[2] ;
 wire \top_I.branch[20].block[6].um_I.ana[3] ;
 wire \top_I.branch[20].block[6].um_I.ana[4] ;
 wire \top_I.branch[20].block[6].um_I.ana[5] ;
 wire \top_I.branch[20].block[6].um_I.ana[6] ;
 wire \top_I.branch[20].block[6].um_I.ana[7] ;
 wire \top_I.branch[20].block[6].um_I.clk ;
 wire \top_I.branch[20].block[6].um_I.ena ;
 wire \top_I.branch[20].block[6].um_I.iw[10] ;
 wire \top_I.branch[20].block[6].um_I.iw[11] ;
 wire \top_I.branch[20].block[6].um_I.iw[12] ;
 wire \top_I.branch[20].block[6].um_I.iw[13] ;
 wire \top_I.branch[20].block[6].um_I.iw[14] ;
 wire \top_I.branch[20].block[6].um_I.iw[15] ;
 wire \top_I.branch[20].block[6].um_I.iw[16] ;
 wire \top_I.branch[20].block[6].um_I.iw[17] ;
 wire \top_I.branch[20].block[6].um_I.iw[1] ;
 wire \top_I.branch[20].block[6].um_I.iw[2] ;
 wire \top_I.branch[20].block[6].um_I.iw[3] ;
 wire \top_I.branch[20].block[6].um_I.iw[4] ;
 wire \top_I.branch[20].block[6].um_I.iw[5] ;
 wire \top_I.branch[20].block[6].um_I.iw[6] ;
 wire \top_I.branch[20].block[6].um_I.iw[7] ;
 wire \top_I.branch[20].block[6].um_I.iw[8] ;
 wire \top_I.branch[20].block[6].um_I.iw[9] ;
 wire \top_I.branch[20].block[6].um_I.k_zero ;
 wire \top_I.branch[20].block[6].um_I.pg_vdd ;
 wire \top_I.branch[20].block[7].um_I.ana[2] ;
 wire \top_I.branch[20].block[7].um_I.ana[3] ;
 wire \top_I.branch[20].block[7].um_I.ana[4] ;
 wire \top_I.branch[20].block[7].um_I.ana[5] ;
 wire \top_I.branch[20].block[7].um_I.ana[6] ;
 wire \top_I.branch[20].block[7].um_I.ana[7] ;
 wire \top_I.branch[20].block[7].um_I.clk ;
 wire \top_I.branch[20].block[7].um_I.ena ;
 wire \top_I.branch[20].block[7].um_I.iw[10] ;
 wire \top_I.branch[20].block[7].um_I.iw[11] ;
 wire \top_I.branch[20].block[7].um_I.iw[12] ;
 wire \top_I.branch[20].block[7].um_I.iw[13] ;
 wire \top_I.branch[20].block[7].um_I.iw[14] ;
 wire \top_I.branch[20].block[7].um_I.iw[15] ;
 wire \top_I.branch[20].block[7].um_I.iw[16] ;
 wire \top_I.branch[20].block[7].um_I.iw[17] ;
 wire \top_I.branch[20].block[7].um_I.iw[1] ;
 wire \top_I.branch[20].block[7].um_I.iw[2] ;
 wire \top_I.branch[20].block[7].um_I.iw[3] ;
 wire \top_I.branch[20].block[7].um_I.iw[4] ;
 wire \top_I.branch[20].block[7].um_I.iw[5] ;
 wire \top_I.branch[20].block[7].um_I.iw[6] ;
 wire \top_I.branch[20].block[7].um_I.iw[7] ;
 wire \top_I.branch[20].block[7].um_I.iw[8] ;
 wire \top_I.branch[20].block[7].um_I.iw[9] ;
 wire \top_I.branch[20].block[7].um_I.k_zero ;
 wire \top_I.branch[20].block[7].um_I.pg_vdd ;
 wire \top_I.branch[20].block[8].um_I.ana[2] ;
 wire \top_I.branch[20].block[8].um_I.ana[3] ;
 wire \top_I.branch[20].block[8].um_I.ana[4] ;
 wire \top_I.branch[20].block[8].um_I.ana[5] ;
 wire \top_I.branch[20].block[8].um_I.ana[6] ;
 wire \top_I.branch[20].block[8].um_I.ana[7] ;
 wire \top_I.branch[20].block[8].um_I.clk ;
 wire \top_I.branch[20].block[8].um_I.ena ;
 wire \top_I.branch[20].block[8].um_I.iw[10] ;
 wire \top_I.branch[20].block[8].um_I.iw[11] ;
 wire \top_I.branch[20].block[8].um_I.iw[12] ;
 wire \top_I.branch[20].block[8].um_I.iw[13] ;
 wire \top_I.branch[20].block[8].um_I.iw[14] ;
 wire \top_I.branch[20].block[8].um_I.iw[15] ;
 wire \top_I.branch[20].block[8].um_I.iw[16] ;
 wire \top_I.branch[20].block[8].um_I.iw[17] ;
 wire \top_I.branch[20].block[8].um_I.iw[1] ;
 wire \top_I.branch[20].block[8].um_I.iw[2] ;
 wire \top_I.branch[20].block[8].um_I.iw[3] ;
 wire \top_I.branch[20].block[8].um_I.iw[4] ;
 wire \top_I.branch[20].block[8].um_I.iw[5] ;
 wire \top_I.branch[20].block[8].um_I.iw[6] ;
 wire \top_I.branch[20].block[8].um_I.iw[7] ;
 wire \top_I.branch[20].block[8].um_I.iw[8] ;
 wire \top_I.branch[20].block[8].um_I.iw[9] ;
 wire \top_I.branch[20].block[8].um_I.k_zero ;
 wire \top_I.branch[20].block[8].um_I.pg_vdd ;
 wire \top_I.branch[20].block[9].um_I.ana[2] ;
 wire \top_I.branch[20].block[9].um_I.ana[3] ;
 wire \top_I.branch[20].block[9].um_I.ana[4] ;
 wire \top_I.branch[20].block[9].um_I.ana[5] ;
 wire \top_I.branch[20].block[9].um_I.ana[6] ;
 wire \top_I.branch[20].block[9].um_I.ana[7] ;
 wire \top_I.branch[20].block[9].um_I.clk ;
 wire \top_I.branch[20].block[9].um_I.ena ;
 wire \top_I.branch[20].block[9].um_I.iw[10] ;
 wire \top_I.branch[20].block[9].um_I.iw[11] ;
 wire \top_I.branch[20].block[9].um_I.iw[12] ;
 wire \top_I.branch[20].block[9].um_I.iw[13] ;
 wire \top_I.branch[20].block[9].um_I.iw[14] ;
 wire \top_I.branch[20].block[9].um_I.iw[15] ;
 wire \top_I.branch[20].block[9].um_I.iw[16] ;
 wire \top_I.branch[20].block[9].um_I.iw[17] ;
 wire \top_I.branch[20].block[9].um_I.iw[1] ;
 wire \top_I.branch[20].block[9].um_I.iw[2] ;
 wire \top_I.branch[20].block[9].um_I.iw[3] ;
 wire \top_I.branch[20].block[9].um_I.iw[4] ;
 wire \top_I.branch[20].block[9].um_I.iw[5] ;
 wire \top_I.branch[20].block[9].um_I.iw[6] ;
 wire \top_I.branch[20].block[9].um_I.iw[7] ;
 wire \top_I.branch[20].block[9].um_I.iw[8] ;
 wire \top_I.branch[20].block[9].um_I.iw[9] ;
 wire \top_I.branch[20].block[9].um_I.k_zero ;
 wire \top_I.branch[20].block[9].um_I.pg_vdd ;
 wire \top_I.branch[20].l_addr[0] ;
 wire \top_I.branch[20].l_addr[1] ;
 wire \top_I.branch[21].block[0].um_I.ana[2] ;
 wire \top_I.branch[21].block[0].um_I.ana[3] ;
 wire \top_I.branch[21].block[0].um_I.ana[4] ;
 wire \top_I.branch[21].block[0].um_I.ana[5] ;
 wire \top_I.branch[21].block[0].um_I.ana[6] ;
 wire \top_I.branch[21].block[0].um_I.ana[7] ;
 wire \top_I.branch[21].block[0].um_I.clk ;
 wire \top_I.branch[21].block[0].um_I.ena ;
 wire \top_I.branch[21].block[0].um_I.iw[10] ;
 wire \top_I.branch[21].block[0].um_I.iw[11] ;
 wire \top_I.branch[21].block[0].um_I.iw[12] ;
 wire \top_I.branch[21].block[0].um_I.iw[13] ;
 wire \top_I.branch[21].block[0].um_I.iw[14] ;
 wire \top_I.branch[21].block[0].um_I.iw[15] ;
 wire \top_I.branch[21].block[0].um_I.iw[16] ;
 wire \top_I.branch[21].block[0].um_I.iw[17] ;
 wire \top_I.branch[21].block[0].um_I.iw[1] ;
 wire \top_I.branch[21].block[0].um_I.iw[2] ;
 wire \top_I.branch[21].block[0].um_I.iw[3] ;
 wire \top_I.branch[21].block[0].um_I.iw[4] ;
 wire \top_I.branch[21].block[0].um_I.iw[5] ;
 wire \top_I.branch[21].block[0].um_I.iw[6] ;
 wire \top_I.branch[21].block[0].um_I.iw[7] ;
 wire \top_I.branch[21].block[0].um_I.iw[8] ;
 wire \top_I.branch[21].block[0].um_I.iw[9] ;
 wire \top_I.branch[21].block[0].um_I.k_zero ;
 wire \top_I.branch[21].block[0].um_I.pg_vdd ;
 wire \top_I.branch[21].block[10].um_I.ana[2] ;
 wire \top_I.branch[21].block[10].um_I.ana[3] ;
 wire \top_I.branch[21].block[10].um_I.ana[4] ;
 wire \top_I.branch[21].block[10].um_I.ana[5] ;
 wire \top_I.branch[21].block[10].um_I.ana[6] ;
 wire \top_I.branch[21].block[10].um_I.ana[7] ;
 wire \top_I.branch[21].block[10].um_I.clk ;
 wire \top_I.branch[21].block[10].um_I.ena ;
 wire \top_I.branch[21].block[10].um_I.iw[10] ;
 wire \top_I.branch[21].block[10].um_I.iw[11] ;
 wire \top_I.branch[21].block[10].um_I.iw[12] ;
 wire \top_I.branch[21].block[10].um_I.iw[13] ;
 wire \top_I.branch[21].block[10].um_I.iw[14] ;
 wire \top_I.branch[21].block[10].um_I.iw[15] ;
 wire \top_I.branch[21].block[10].um_I.iw[16] ;
 wire \top_I.branch[21].block[10].um_I.iw[17] ;
 wire \top_I.branch[21].block[10].um_I.iw[1] ;
 wire \top_I.branch[21].block[10].um_I.iw[2] ;
 wire \top_I.branch[21].block[10].um_I.iw[3] ;
 wire \top_I.branch[21].block[10].um_I.iw[4] ;
 wire \top_I.branch[21].block[10].um_I.iw[5] ;
 wire \top_I.branch[21].block[10].um_I.iw[6] ;
 wire \top_I.branch[21].block[10].um_I.iw[7] ;
 wire \top_I.branch[21].block[10].um_I.iw[8] ;
 wire \top_I.branch[21].block[10].um_I.iw[9] ;
 wire \top_I.branch[21].block[10].um_I.k_zero ;
 wire \top_I.branch[21].block[10].um_I.pg_vdd ;
 wire \top_I.branch[21].block[11].um_I.ana[2] ;
 wire \top_I.branch[21].block[11].um_I.ana[3] ;
 wire \top_I.branch[21].block[11].um_I.ana[4] ;
 wire \top_I.branch[21].block[11].um_I.ana[5] ;
 wire \top_I.branch[21].block[11].um_I.ana[6] ;
 wire \top_I.branch[21].block[11].um_I.ana[7] ;
 wire \top_I.branch[21].block[11].um_I.clk ;
 wire \top_I.branch[21].block[11].um_I.ena ;
 wire \top_I.branch[21].block[11].um_I.iw[10] ;
 wire \top_I.branch[21].block[11].um_I.iw[11] ;
 wire \top_I.branch[21].block[11].um_I.iw[12] ;
 wire \top_I.branch[21].block[11].um_I.iw[13] ;
 wire \top_I.branch[21].block[11].um_I.iw[14] ;
 wire \top_I.branch[21].block[11].um_I.iw[15] ;
 wire \top_I.branch[21].block[11].um_I.iw[16] ;
 wire \top_I.branch[21].block[11].um_I.iw[17] ;
 wire \top_I.branch[21].block[11].um_I.iw[1] ;
 wire \top_I.branch[21].block[11].um_I.iw[2] ;
 wire \top_I.branch[21].block[11].um_I.iw[3] ;
 wire \top_I.branch[21].block[11].um_I.iw[4] ;
 wire \top_I.branch[21].block[11].um_I.iw[5] ;
 wire \top_I.branch[21].block[11].um_I.iw[6] ;
 wire \top_I.branch[21].block[11].um_I.iw[7] ;
 wire \top_I.branch[21].block[11].um_I.iw[8] ;
 wire \top_I.branch[21].block[11].um_I.iw[9] ;
 wire \top_I.branch[21].block[11].um_I.k_zero ;
 wire \top_I.branch[21].block[11].um_I.pg_vdd ;
 wire \top_I.branch[21].block[12].um_I.ana[2] ;
 wire \top_I.branch[21].block[12].um_I.ana[3] ;
 wire \top_I.branch[21].block[12].um_I.ana[4] ;
 wire \top_I.branch[21].block[12].um_I.ana[5] ;
 wire \top_I.branch[21].block[12].um_I.ana[6] ;
 wire \top_I.branch[21].block[12].um_I.ana[7] ;
 wire \top_I.branch[21].block[12].um_I.clk ;
 wire \top_I.branch[21].block[12].um_I.ena ;
 wire \top_I.branch[21].block[12].um_I.iw[10] ;
 wire \top_I.branch[21].block[12].um_I.iw[11] ;
 wire \top_I.branch[21].block[12].um_I.iw[12] ;
 wire \top_I.branch[21].block[12].um_I.iw[13] ;
 wire \top_I.branch[21].block[12].um_I.iw[14] ;
 wire \top_I.branch[21].block[12].um_I.iw[15] ;
 wire \top_I.branch[21].block[12].um_I.iw[16] ;
 wire \top_I.branch[21].block[12].um_I.iw[17] ;
 wire \top_I.branch[21].block[12].um_I.iw[1] ;
 wire \top_I.branch[21].block[12].um_I.iw[2] ;
 wire \top_I.branch[21].block[12].um_I.iw[3] ;
 wire \top_I.branch[21].block[12].um_I.iw[4] ;
 wire \top_I.branch[21].block[12].um_I.iw[5] ;
 wire \top_I.branch[21].block[12].um_I.iw[6] ;
 wire \top_I.branch[21].block[12].um_I.iw[7] ;
 wire \top_I.branch[21].block[12].um_I.iw[8] ;
 wire \top_I.branch[21].block[12].um_I.iw[9] ;
 wire \top_I.branch[21].block[12].um_I.k_zero ;
 wire \top_I.branch[21].block[12].um_I.pg_vdd ;
 wire \top_I.branch[21].block[13].um_I.ana[2] ;
 wire \top_I.branch[21].block[13].um_I.ana[3] ;
 wire \top_I.branch[21].block[13].um_I.ana[4] ;
 wire \top_I.branch[21].block[13].um_I.ana[5] ;
 wire \top_I.branch[21].block[13].um_I.ana[6] ;
 wire \top_I.branch[21].block[13].um_I.ana[7] ;
 wire \top_I.branch[21].block[13].um_I.clk ;
 wire \top_I.branch[21].block[13].um_I.ena ;
 wire \top_I.branch[21].block[13].um_I.iw[10] ;
 wire \top_I.branch[21].block[13].um_I.iw[11] ;
 wire \top_I.branch[21].block[13].um_I.iw[12] ;
 wire \top_I.branch[21].block[13].um_I.iw[13] ;
 wire \top_I.branch[21].block[13].um_I.iw[14] ;
 wire \top_I.branch[21].block[13].um_I.iw[15] ;
 wire \top_I.branch[21].block[13].um_I.iw[16] ;
 wire \top_I.branch[21].block[13].um_I.iw[17] ;
 wire \top_I.branch[21].block[13].um_I.iw[1] ;
 wire \top_I.branch[21].block[13].um_I.iw[2] ;
 wire \top_I.branch[21].block[13].um_I.iw[3] ;
 wire \top_I.branch[21].block[13].um_I.iw[4] ;
 wire \top_I.branch[21].block[13].um_I.iw[5] ;
 wire \top_I.branch[21].block[13].um_I.iw[6] ;
 wire \top_I.branch[21].block[13].um_I.iw[7] ;
 wire \top_I.branch[21].block[13].um_I.iw[8] ;
 wire \top_I.branch[21].block[13].um_I.iw[9] ;
 wire \top_I.branch[21].block[13].um_I.k_zero ;
 wire \top_I.branch[21].block[13].um_I.pg_vdd ;
 wire \top_I.branch[21].block[14].um_I.ana[2] ;
 wire \top_I.branch[21].block[14].um_I.ana[3] ;
 wire \top_I.branch[21].block[14].um_I.ana[4] ;
 wire \top_I.branch[21].block[14].um_I.ana[5] ;
 wire \top_I.branch[21].block[14].um_I.ana[6] ;
 wire \top_I.branch[21].block[14].um_I.ana[7] ;
 wire \top_I.branch[21].block[14].um_I.clk ;
 wire \top_I.branch[21].block[14].um_I.ena ;
 wire \top_I.branch[21].block[14].um_I.iw[10] ;
 wire \top_I.branch[21].block[14].um_I.iw[11] ;
 wire \top_I.branch[21].block[14].um_I.iw[12] ;
 wire \top_I.branch[21].block[14].um_I.iw[13] ;
 wire \top_I.branch[21].block[14].um_I.iw[14] ;
 wire \top_I.branch[21].block[14].um_I.iw[15] ;
 wire \top_I.branch[21].block[14].um_I.iw[16] ;
 wire \top_I.branch[21].block[14].um_I.iw[17] ;
 wire \top_I.branch[21].block[14].um_I.iw[1] ;
 wire \top_I.branch[21].block[14].um_I.iw[2] ;
 wire \top_I.branch[21].block[14].um_I.iw[3] ;
 wire \top_I.branch[21].block[14].um_I.iw[4] ;
 wire \top_I.branch[21].block[14].um_I.iw[5] ;
 wire \top_I.branch[21].block[14].um_I.iw[6] ;
 wire \top_I.branch[21].block[14].um_I.iw[7] ;
 wire \top_I.branch[21].block[14].um_I.iw[8] ;
 wire \top_I.branch[21].block[14].um_I.iw[9] ;
 wire \top_I.branch[21].block[14].um_I.k_zero ;
 wire \top_I.branch[21].block[14].um_I.pg_vdd ;
 wire \top_I.branch[21].block[15].um_I.ana[2] ;
 wire \top_I.branch[21].block[15].um_I.ana[3] ;
 wire \top_I.branch[21].block[15].um_I.ana[4] ;
 wire \top_I.branch[21].block[15].um_I.ana[5] ;
 wire \top_I.branch[21].block[15].um_I.ana[6] ;
 wire \top_I.branch[21].block[15].um_I.ana[7] ;
 wire \top_I.branch[21].block[15].um_I.clk ;
 wire \top_I.branch[21].block[15].um_I.ena ;
 wire \top_I.branch[21].block[15].um_I.iw[10] ;
 wire \top_I.branch[21].block[15].um_I.iw[11] ;
 wire \top_I.branch[21].block[15].um_I.iw[12] ;
 wire \top_I.branch[21].block[15].um_I.iw[13] ;
 wire \top_I.branch[21].block[15].um_I.iw[14] ;
 wire \top_I.branch[21].block[15].um_I.iw[15] ;
 wire \top_I.branch[21].block[15].um_I.iw[16] ;
 wire \top_I.branch[21].block[15].um_I.iw[17] ;
 wire \top_I.branch[21].block[15].um_I.iw[1] ;
 wire \top_I.branch[21].block[15].um_I.iw[2] ;
 wire \top_I.branch[21].block[15].um_I.iw[3] ;
 wire \top_I.branch[21].block[15].um_I.iw[4] ;
 wire \top_I.branch[21].block[15].um_I.iw[5] ;
 wire \top_I.branch[21].block[15].um_I.iw[6] ;
 wire \top_I.branch[21].block[15].um_I.iw[7] ;
 wire \top_I.branch[21].block[15].um_I.iw[8] ;
 wire \top_I.branch[21].block[15].um_I.iw[9] ;
 wire \top_I.branch[21].block[15].um_I.k_zero ;
 wire \top_I.branch[21].block[15].um_I.pg_vdd ;
 wire \top_I.branch[21].block[1].um_I.ana[2] ;
 wire \top_I.branch[21].block[1].um_I.ana[3] ;
 wire \top_I.branch[21].block[1].um_I.ana[4] ;
 wire \top_I.branch[21].block[1].um_I.ana[5] ;
 wire \top_I.branch[21].block[1].um_I.ana[6] ;
 wire \top_I.branch[21].block[1].um_I.ana[7] ;
 wire \top_I.branch[21].block[1].um_I.clk ;
 wire \top_I.branch[21].block[1].um_I.ena ;
 wire \top_I.branch[21].block[1].um_I.iw[10] ;
 wire \top_I.branch[21].block[1].um_I.iw[11] ;
 wire \top_I.branch[21].block[1].um_I.iw[12] ;
 wire \top_I.branch[21].block[1].um_I.iw[13] ;
 wire \top_I.branch[21].block[1].um_I.iw[14] ;
 wire \top_I.branch[21].block[1].um_I.iw[15] ;
 wire \top_I.branch[21].block[1].um_I.iw[16] ;
 wire \top_I.branch[21].block[1].um_I.iw[17] ;
 wire \top_I.branch[21].block[1].um_I.iw[1] ;
 wire \top_I.branch[21].block[1].um_I.iw[2] ;
 wire \top_I.branch[21].block[1].um_I.iw[3] ;
 wire \top_I.branch[21].block[1].um_I.iw[4] ;
 wire \top_I.branch[21].block[1].um_I.iw[5] ;
 wire \top_I.branch[21].block[1].um_I.iw[6] ;
 wire \top_I.branch[21].block[1].um_I.iw[7] ;
 wire \top_I.branch[21].block[1].um_I.iw[8] ;
 wire \top_I.branch[21].block[1].um_I.iw[9] ;
 wire \top_I.branch[21].block[1].um_I.k_zero ;
 wire \top_I.branch[21].block[1].um_I.pg_vdd ;
 wire \top_I.branch[21].block[2].um_I.ana[2] ;
 wire \top_I.branch[21].block[2].um_I.ana[3] ;
 wire \top_I.branch[21].block[2].um_I.ana[4] ;
 wire \top_I.branch[21].block[2].um_I.ana[5] ;
 wire \top_I.branch[21].block[2].um_I.ana[6] ;
 wire \top_I.branch[21].block[2].um_I.ana[7] ;
 wire \top_I.branch[21].block[2].um_I.clk ;
 wire \top_I.branch[21].block[2].um_I.ena ;
 wire \top_I.branch[21].block[2].um_I.iw[10] ;
 wire \top_I.branch[21].block[2].um_I.iw[11] ;
 wire \top_I.branch[21].block[2].um_I.iw[12] ;
 wire \top_I.branch[21].block[2].um_I.iw[13] ;
 wire \top_I.branch[21].block[2].um_I.iw[14] ;
 wire \top_I.branch[21].block[2].um_I.iw[15] ;
 wire \top_I.branch[21].block[2].um_I.iw[16] ;
 wire \top_I.branch[21].block[2].um_I.iw[17] ;
 wire \top_I.branch[21].block[2].um_I.iw[1] ;
 wire \top_I.branch[21].block[2].um_I.iw[2] ;
 wire \top_I.branch[21].block[2].um_I.iw[3] ;
 wire \top_I.branch[21].block[2].um_I.iw[4] ;
 wire \top_I.branch[21].block[2].um_I.iw[5] ;
 wire \top_I.branch[21].block[2].um_I.iw[6] ;
 wire \top_I.branch[21].block[2].um_I.iw[7] ;
 wire \top_I.branch[21].block[2].um_I.iw[8] ;
 wire \top_I.branch[21].block[2].um_I.iw[9] ;
 wire \top_I.branch[21].block[2].um_I.k_zero ;
 wire \top_I.branch[21].block[2].um_I.pg_vdd ;
 wire \top_I.branch[21].block[3].um_I.ana[2] ;
 wire \top_I.branch[21].block[3].um_I.ana[3] ;
 wire \top_I.branch[21].block[3].um_I.ana[4] ;
 wire \top_I.branch[21].block[3].um_I.ana[5] ;
 wire \top_I.branch[21].block[3].um_I.ana[6] ;
 wire \top_I.branch[21].block[3].um_I.ana[7] ;
 wire \top_I.branch[21].block[3].um_I.clk ;
 wire \top_I.branch[21].block[3].um_I.ena ;
 wire \top_I.branch[21].block[3].um_I.iw[10] ;
 wire \top_I.branch[21].block[3].um_I.iw[11] ;
 wire \top_I.branch[21].block[3].um_I.iw[12] ;
 wire \top_I.branch[21].block[3].um_I.iw[13] ;
 wire \top_I.branch[21].block[3].um_I.iw[14] ;
 wire \top_I.branch[21].block[3].um_I.iw[15] ;
 wire \top_I.branch[21].block[3].um_I.iw[16] ;
 wire \top_I.branch[21].block[3].um_I.iw[17] ;
 wire \top_I.branch[21].block[3].um_I.iw[1] ;
 wire \top_I.branch[21].block[3].um_I.iw[2] ;
 wire \top_I.branch[21].block[3].um_I.iw[3] ;
 wire \top_I.branch[21].block[3].um_I.iw[4] ;
 wire \top_I.branch[21].block[3].um_I.iw[5] ;
 wire \top_I.branch[21].block[3].um_I.iw[6] ;
 wire \top_I.branch[21].block[3].um_I.iw[7] ;
 wire \top_I.branch[21].block[3].um_I.iw[8] ;
 wire \top_I.branch[21].block[3].um_I.iw[9] ;
 wire \top_I.branch[21].block[3].um_I.k_zero ;
 wire \top_I.branch[21].block[3].um_I.pg_vdd ;
 wire \top_I.branch[21].block[4].um_I.ana[2] ;
 wire \top_I.branch[21].block[4].um_I.ana[3] ;
 wire \top_I.branch[21].block[4].um_I.ana[4] ;
 wire \top_I.branch[21].block[4].um_I.ana[5] ;
 wire \top_I.branch[21].block[4].um_I.ana[6] ;
 wire \top_I.branch[21].block[4].um_I.ana[7] ;
 wire \top_I.branch[21].block[4].um_I.clk ;
 wire \top_I.branch[21].block[4].um_I.ena ;
 wire \top_I.branch[21].block[4].um_I.iw[10] ;
 wire \top_I.branch[21].block[4].um_I.iw[11] ;
 wire \top_I.branch[21].block[4].um_I.iw[12] ;
 wire \top_I.branch[21].block[4].um_I.iw[13] ;
 wire \top_I.branch[21].block[4].um_I.iw[14] ;
 wire \top_I.branch[21].block[4].um_I.iw[15] ;
 wire \top_I.branch[21].block[4].um_I.iw[16] ;
 wire \top_I.branch[21].block[4].um_I.iw[17] ;
 wire \top_I.branch[21].block[4].um_I.iw[1] ;
 wire \top_I.branch[21].block[4].um_I.iw[2] ;
 wire \top_I.branch[21].block[4].um_I.iw[3] ;
 wire \top_I.branch[21].block[4].um_I.iw[4] ;
 wire \top_I.branch[21].block[4].um_I.iw[5] ;
 wire \top_I.branch[21].block[4].um_I.iw[6] ;
 wire \top_I.branch[21].block[4].um_I.iw[7] ;
 wire \top_I.branch[21].block[4].um_I.iw[8] ;
 wire \top_I.branch[21].block[4].um_I.iw[9] ;
 wire \top_I.branch[21].block[4].um_I.k_zero ;
 wire \top_I.branch[21].block[4].um_I.pg_vdd ;
 wire \top_I.branch[21].block[5].um_I.ana[2] ;
 wire \top_I.branch[21].block[5].um_I.ana[3] ;
 wire \top_I.branch[21].block[5].um_I.ana[4] ;
 wire \top_I.branch[21].block[5].um_I.ana[5] ;
 wire \top_I.branch[21].block[5].um_I.ana[6] ;
 wire \top_I.branch[21].block[5].um_I.ana[7] ;
 wire \top_I.branch[21].block[5].um_I.clk ;
 wire \top_I.branch[21].block[5].um_I.ena ;
 wire \top_I.branch[21].block[5].um_I.iw[10] ;
 wire \top_I.branch[21].block[5].um_I.iw[11] ;
 wire \top_I.branch[21].block[5].um_I.iw[12] ;
 wire \top_I.branch[21].block[5].um_I.iw[13] ;
 wire \top_I.branch[21].block[5].um_I.iw[14] ;
 wire \top_I.branch[21].block[5].um_I.iw[15] ;
 wire \top_I.branch[21].block[5].um_I.iw[16] ;
 wire \top_I.branch[21].block[5].um_I.iw[17] ;
 wire \top_I.branch[21].block[5].um_I.iw[1] ;
 wire \top_I.branch[21].block[5].um_I.iw[2] ;
 wire \top_I.branch[21].block[5].um_I.iw[3] ;
 wire \top_I.branch[21].block[5].um_I.iw[4] ;
 wire \top_I.branch[21].block[5].um_I.iw[5] ;
 wire \top_I.branch[21].block[5].um_I.iw[6] ;
 wire \top_I.branch[21].block[5].um_I.iw[7] ;
 wire \top_I.branch[21].block[5].um_I.iw[8] ;
 wire \top_I.branch[21].block[5].um_I.iw[9] ;
 wire \top_I.branch[21].block[5].um_I.k_zero ;
 wire \top_I.branch[21].block[5].um_I.pg_vdd ;
 wire \top_I.branch[21].block[6].um_I.ana[2] ;
 wire \top_I.branch[21].block[6].um_I.ana[3] ;
 wire \top_I.branch[21].block[6].um_I.ana[4] ;
 wire \top_I.branch[21].block[6].um_I.ana[5] ;
 wire \top_I.branch[21].block[6].um_I.ana[6] ;
 wire \top_I.branch[21].block[6].um_I.ana[7] ;
 wire \top_I.branch[21].block[6].um_I.clk ;
 wire \top_I.branch[21].block[6].um_I.ena ;
 wire \top_I.branch[21].block[6].um_I.iw[10] ;
 wire \top_I.branch[21].block[6].um_I.iw[11] ;
 wire \top_I.branch[21].block[6].um_I.iw[12] ;
 wire \top_I.branch[21].block[6].um_I.iw[13] ;
 wire \top_I.branch[21].block[6].um_I.iw[14] ;
 wire \top_I.branch[21].block[6].um_I.iw[15] ;
 wire \top_I.branch[21].block[6].um_I.iw[16] ;
 wire \top_I.branch[21].block[6].um_I.iw[17] ;
 wire \top_I.branch[21].block[6].um_I.iw[1] ;
 wire \top_I.branch[21].block[6].um_I.iw[2] ;
 wire \top_I.branch[21].block[6].um_I.iw[3] ;
 wire \top_I.branch[21].block[6].um_I.iw[4] ;
 wire \top_I.branch[21].block[6].um_I.iw[5] ;
 wire \top_I.branch[21].block[6].um_I.iw[6] ;
 wire \top_I.branch[21].block[6].um_I.iw[7] ;
 wire \top_I.branch[21].block[6].um_I.iw[8] ;
 wire \top_I.branch[21].block[6].um_I.iw[9] ;
 wire \top_I.branch[21].block[6].um_I.k_zero ;
 wire \top_I.branch[21].block[6].um_I.pg_vdd ;
 wire \top_I.branch[21].block[7].um_I.ana[2] ;
 wire \top_I.branch[21].block[7].um_I.ana[3] ;
 wire \top_I.branch[21].block[7].um_I.ana[4] ;
 wire \top_I.branch[21].block[7].um_I.ana[5] ;
 wire \top_I.branch[21].block[7].um_I.ana[6] ;
 wire \top_I.branch[21].block[7].um_I.ana[7] ;
 wire \top_I.branch[21].block[7].um_I.clk ;
 wire \top_I.branch[21].block[7].um_I.ena ;
 wire \top_I.branch[21].block[7].um_I.iw[10] ;
 wire \top_I.branch[21].block[7].um_I.iw[11] ;
 wire \top_I.branch[21].block[7].um_I.iw[12] ;
 wire \top_I.branch[21].block[7].um_I.iw[13] ;
 wire \top_I.branch[21].block[7].um_I.iw[14] ;
 wire \top_I.branch[21].block[7].um_I.iw[15] ;
 wire \top_I.branch[21].block[7].um_I.iw[16] ;
 wire \top_I.branch[21].block[7].um_I.iw[17] ;
 wire \top_I.branch[21].block[7].um_I.iw[1] ;
 wire \top_I.branch[21].block[7].um_I.iw[2] ;
 wire \top_I.branch[21].block[7].um_I.iw[3] ;
 wire \top_I.branch[21].block[7].um_I.iw[4] ;
 wire \top_I.branch[21].block[7].um_I.iw[5] ;
 wire \top_I.branch[21].block[7].um_I.iw[6] ;
 wire \top_I.branch[21].block[7].um_I.iw[7] ;
 wire \top_I.branch[21].block[7].um_I.iw[8] ;
 wire \top_I.branch[21].block[7].um_I.iw[9] ;
 wire \top_I.branch[21].block[7].um_I.k_zero ;
 wire \top_I.branch[21].block[7].um_I.pg_vdd ;
 wire \top_I.branch[21].block[8].um_I.ana[2] ;
 wire \top_I.branch[21].block[8].um_I.ana[3] ;
 wire \top_I.branch[21].block[8].um_I.ana[4] ;
 wire \top_I.branch[21].block[8].um_I.ana[5] ;
 wire \top_I.branch[21].block[8].um_I.ana[6] ;
 wire \top_I.branch[21].block[8].um_I.ana[7] ;
 wire \top_I.branch[21].block[8].um_I.clk ;
 wire \top_I.branch[21].block[8].um_I.ena ;
 wire \top_I.branch[21].block[8].um_I.iw[10] ;
 wire \top_I.branch[21].block[8].um_I.iw[11] ;
 wire \top_I.branch[21].block[8].um_I.iw[12] ;
 wire \top_I.branch[21].block[8].um_I.iw[13] ;
 wire \top_I.branch[21].block[8].um_I.iw[14] ;
 wire \top_I.branch[21].block[8].um_I.iw[15] ;
 wire \top_I.branch[21].block[8].um_I.iw[16] ;
 wire \top_I.branch[21].block[8].um_I.iw[17] ;
 wire \top_I.branch[21].block[8].um_I.iw[1] ;
 wire \top_I.branch[21].block[8].um_I.iw[2] ;
 wire \top_I.branch[21].block[8].um_I.iw[3] ;
 wire \top_I.branch[21].block[8].um_I.iw[4] ;
 wire \top_I.branch[21].block[8].um_I.iw[5] ;
 wire \top_I.branch[21].block[8].um_I.iw[6] ;
 wire \top_I.branch[21].block[8].um_I.iw[7] ;
 wire \top_I.branch[21].block[8].um_I.iw[8] ;
 wire \top_I.branch[21].block[8].um_I.iw[9] ;
 wire \top_I.branch[21].block[8].um_I.k_zero ;
 wire \top_I.branch[21].block[8].um_I.pg_vdd ;
 wire \top_I.branch[21].block[9].um_I.ana[2] ;
 wire \top_I.branch[21].block[9].um_I.ana[3] ;
 wire \top_I.branch[21].block[9].um_I.ana[4] ;
 wire \top_I.branch[21].block[9].um_I.ana[5] ;
 wire \top_I.branch[21].block[9].um_I.ana[6] ;
 wire \top_I.branch[21].block[9].um_I.ana[7] ;
 wire \top_I.branch[21].block[9].um_I.clk ;
 wire \top_I.branch[21].block[9].um_I.ena ;
 wire \top_I.branch[21].block[9].um_I.iw[10] ;
 wire \top_I.branch[21].block[9].um_I.iw[11] ;
 wire \top_I.branch[21].block[9].um_I.iw[12] ;
 wire \top_I.branch[21].block[9].um_I.iw[13] ;
 wire \top_I.branch[21].block[9].um_I.iw[14] ;
 wire \top_I.branch[21].block[9].um_I.iw[15] ;
 wire \top_I.branch[21].block[9].um_I.iw[16] ;
 wire \top_I.branch[21].block[9].um_I.iw[17] ;
 wire \top_I.branch[21].block[9].um_I.iw[1] ;
 wire \top_I.branch[21].block[9].um_I.iw[2] ;
 wire \top_I.branch[21].block[9].um_I.iw[3] ;
 wire \top_I.branch[21].block[9].um_I.iw[4] ;
 wire \top_I.branch[21].block[9].um_I.iw[5] ;
 wire \top_I.branch[21].block[9].um_I.iw[6] ;
 wire \top_I.branch[21].block[9].um_I.iw[7] ;
 wire \top_I.branch[21].block[9].um_I.iw[8] ;
 wire \top_I.branch[21].block[9].um_I.iw[9] ;
 wire \top_I.branch[21].block[9].um_I.k_zero ;
 wire \top_I.branch[21].block[9].um_I.pg_vdd ;
 wire \top_I.branch[21].l_addr[0] ;
 wire \top_I.branch[21].l_addr[1] ;
 wire \top_I.branch[22].block[0].um_I.ana[2] ;
 wire \top_I.branch[22].block[0].um_I.ana[3] ;
 wire \top_I.branch[22].block[0].um_I.ana[4] ;
 wire \top_I.branch[22].block[0].um_I.ana[5] ;
 wire \top_I.branch[22].block[0].um_I.ana[6] ;
 wire \top_I.branch[22].block[0].um_I.ana[7] ;
 wire \top_I.branch[22].block[0].um_I.clk ;
 wire \top_I.branch[22].block[0].um_I.ena ;
 wire \top_I.branch[22].block[0].um_I.iw[10] ;
 wire \top_I.branch[22].block[0].um_I.iw[11] ;
 wire \top_I.branch[22].block[0].um_I.iw[12] ;
 wire \top_I.branch[22].block[0].um_I.iw[13] ;
 wire \top_I.branch[22].block[0].um_I.iw[14] ;
 wire \top_I.branch[22].block[0].um_I.iw[15] ;
 wire \top_I.branch[22].block[0].um_I.iw[16] ;
 wire \top_I.branch[22].block[0].um_I.iw[17] ;
 wire \top_I.branch[22].block[0].um_I.iw[1] ;
 wire \top_I.branch[22].block[0].um_I.iw[2] ;
 wire \top_I.branch[22].block[0].um_I.iw[3] ;
 wire \top_I.branch[22].block[0].um_I.iw[4] ;
 wire \top_I.branch[22].block[0].um_I.iw[5] ;
 wire \top_I.branch[22].block[0].um_I.iw[6] ;
 wire \top_I.branch[22].block[0].um_I.iw[7] ;
 wire \top_I.branch[22].block[0].um_I.iw[8] ;
 wire \top_I.branch[22].block[0].um_I.iw[9] ;
 wire \top_I.branch[22].block[0].um_I.k_zero ;
 wire \top_I.branch[22].block[0].um_I.pg_vdd ;
 wire \top_I.branch[22].block[10].um_I.ana[2] ;
 wire \top_I.branch[22].block[10].um_I.ana[3] ;
 wire \top_I.branch[22].block[10].um_I.ana[4] ;
 wire \top_I.branch[22].block[10].um_I.ana[5] ;
 wire \top_I.branch[22].block[10].um_I.ana[6] ;
 wire \top_I.branch[22].block[10].um_I.ana[7] ;
 wire \top_I.branch[22].block[10].um_I.clk ;
 wire \top_I.branch[22].block[10].um_I.ena ;
 wire \top_I.branch[22].block[10].um_I.iw[10] ;
 wire \top_I.branch[22].block[10].um_I.iw[11] ;
 wire \top_I.branch[22].block[10].um_I.iw[12] ;
 wire \top_I.branch[22].block[10].um_I.iw[13] ;
 wire \top_I.branch[22].block[10].um_I.iw[14] ;
 wire \top_I.branch[22].block[10].um_I.iw[15] ;
 wire \top_I.branch[22].block[10].um_I.iw[16] ;
 wire \top_I.branch[22].block[10].um_I.iw[17] ;
 wire \top_I.branch[22].block[10].um_I.iw[1] ;
 wire \top_I.branch[22].block[10].um_I.iw[2] ;
 wire \top_I.branch[22].block[10].um_I.iw[3] ;
 wire \top_I.branch[22].block[10].um_I.iw[4] ;
 wire \top_I.branch[22].block[10].um_I.iw[5] ;
 wire \top_I.branch[22].block[10].um_I.iw[6] ;
 wire \top_I.branch[22].block[10].um_I.iw[7] ;
 wire \top_I.branch[22].block[10].um_I.iw[8] ;
 wire \top_I.branch[22].block[10].um_I.iw[9] ;
 wire \top_I.branch[22].block[10].um_I.k_zero ;
 wire \top_I.branch[22].block[10].um_I.pg_vdd ;
 wire \top_I.branch[22].block[11].um_I.ana[2] ;
 wire \top_I.branch[22].block[11].um_I.ana[3] ;
 wire \top_I.branch[22].block[11].um_I.ana[4] ;
 wire \top_I.branch[22].block[11].um_I.ana[5] ;
 wire \top_I.branch[22].block[11].um_I.ana[6] ;
 wire \top_I.branch[22].block[11].um_I.ana[7] ;
 wire \top_I.branch[22].block[11].um_I.clk ;
 wire \top_I.branch[22].block[11].um_I.ena ;
 wire \top_I.branch[22].block[11].um_I.iw[10] ;
 wire \top_I.branch[22].block[11].um_I.iw[11] ;
 wire \top_I.branch[22].block[11].um_I.iw[12] ;
 wire \top_I.branch[22].block[11].um_I.iw[13] ;
 wire \top_I.branch[22].block[11].um_I.iw[14] ;
 wire \top_I.branch[22].block[11].um_I.iw[15] ;
 wire \top_I.branch[22].block[11].um_I.iw[16] ;
 wire \top_I.branch[22].block[11].um_I.iw[17] ;
 wire \top_I.branch[22].block[11].um_I.iw[1] ;
 wire \top_I.branch[22].block[11].um_I.iw[2] ;
 wire \top_I.branch[22].block[11].um_I.iw[3] ;
 wire \top_I.branch[22].block[11].um_I.iw[4] ;
 wire \top_I.branch[22].block[11].um_I.iw[5] ;
 wire \top_I.branch[22].block[11].um_I.iw[6] ;
 wire \top_I.branch[22].block[11].um_I.iw[7] ;
 wire \top_I.branch[22].block[11].um_I.iw[8] ;
 wire \top_I.branch[22].block[11].um_I.iw[9] ;
 wire \top_I.branch[22].block[11].um_I.k_zero ;
 wire \top_I.branch[22].block[11].um_I.pg_vdd ;
 wire \top_I.branch[22].block[12].um_I.ana[2] ;
 wire \top_I.branch[22].block[12].um_I.ana[3] ;
 wire \top_I.branch[22].block[12].um_I.ana[4] ;
 wire \top_I.branch[22].block[12].um_I.ana[5] ;
 wire \top_I.branch[22].block[12].um_I.ana[6] ;
 wire \top_I.branch[22].block[12].um_I.ana[7] ;
 wire \top_I.branch[22].block[12].um_I.clk ;
 wire \top_I.branch[22].block[12].um_I.ena ;
 wire \top_I.branch[22].block[12].um_I.iw[10] ;
 wire \top_I.branch[22].block[12].um_I.iw[11] ;
 wire \top_I.branch[22].block[12].um_I.iw[12] ;
 wire \top_I.branch[22].block[12].um_I.iw[13] ;
 wire \top_I.branch[22].block[12].um_I.iw[14] ;
 wire \top_I.branch[22].block[12].um_I.iw[15] ;
 wire \top_I.branch[22].block[12].um_I.iw[16] ;
 wire \top_I.branch[22].block[12].um_I.iw[17] ;
 wire \top_I.branch[22].block[12].um_I.iw[1] ;
 wire \top_I.branch[22].block[12].um_I.iw[2] ;
 wire \top_I.branch[22].block[12].um_I.iw[3] ;
 wire \top_I.branch[22].block[12].um_I.iw[4] ;
 wire \top_I.branch[22].block[12].um_I.iw[5] ;
 wire \top_I.branch[22].block[12].um_I.iw[6] ;
 wire \top_I.branch[22].block[12].um_I.iw[7] ;
 wire \top_I.branch[22].block[12].um_I.iw[8] ;
 wire \top_I.branch[22].block[12].um_I.iw[9] ;
 wire \top_I.branch[22].block[12].um_I.k_zero ;
 wire \top_I.branch[22].block[12].um_I.pg_vdd ;
 wire \top_I.branch[22].block[13].um_I.ana[2] ;
 wire \top_I.branch[22].block[13].um_I.ana[3] ;
 wire \top_I.branch[22].block[13].um_I.ana[4] ;
 wire \top_I.branch[22].block[13].um_I.ana[5] ;
 wire \top_I.branch[22].block[13].um_I.ana[6] ;
 wire \top_I.branch[22].block[13].um_I.ana[7] ;
 wire \top_I.branch[22].block[13].um_I.clk ;
 wire \top_I.branch[22].block[13].um_I.ena ;
 wire \top_I.branch[22].block[13].um_I.iw[10] ;
 wire \top_I.branch[22].block[13].um_I.iw[11] ;
 wire \top_I.branch[22].block[13].um_I.iw[12] ;
 wire \top_I.branch[22].block[13].um_I.iw[13] ;
 wire \top_I.branch[22].block[13].um_I.iw[14] ;
 wire \top_I.branch[22].block[13].um_I.iw[15] ;
 wire \top_I.branch[22].block[13].um_I.iw[16] ;
 wire \top_I.branch[22].block[13].um_I.iw[17] ;
 wire \top_I.branch[22].block[13].um_I.iw[1] ;
 wire \top_I.branch[22].block[13].um_I.iw[2] ;
 wire \top_I.branch[22].block[13].um_I.iw[3] ;
 wire \top_I.branch[22].block[13].um_I.iw[4] ;
 wire \top_I.branch[22].block[13].um_I.iw[5] ;
 wire \top_I.branch[22].block[13].um_I.iw[6] ;
 wire \top_I.branch[22].block[13].um_I.iw[7] ;
 wire \top_I.branch[22].block[13].um_I.iw[8] ;
 wire \top_I.branch[22].block[13].um_I.iw[9] ;
 wire \top_I.branch[22].block[13].um_I.k_zero ;
 wire \top_I.branch[22].block[13].um_I.pg_vdd ;
 wire \top_I.branch[22].block[14].um_I.ana[2] ;
 wire \top_I.branch[22].block[14].um_I.ana[3] ;
 wire \top_I.branch[22].block[14].um_I.ana[4] ;
 wire \top_I.branch[22].block[14].um_I.ana[5] ;
 wire \top_I.branch[22].block[14].um_I.ana[6] ;
 wire \top_I.branch[22].block[14].um_I.ana[7] ;
 wire \top_I.branch[22].block[14].um_I.clk ;
 wire \top_I.branch[22].block[14].um_I.ena ;
 wire \top_I.branch[22].block[14].um_I.iw[10] ;
 wire \top_I.branch[22].block[14].um_I.iw[11] ;
 wire \top_I.branch[22].block[14].um_I.iw[12] ;
 wire \top_I.branch[22].block[14].um_I.iw[13] ;
 wire \top_I.branch[22].block[14].um_I.iw[14] ;
 wire \top_I.branch[22].block[14].um_I.iw[15] ;
 wire \top_I.branch[22].block[14].um_I.iw[16] ;
 wire \top_I.branch[22].block[14].um_I.iw[17] ;
 wire \top_I.branch[22].block[14].um_I.iw[1] ;
 wire \top_I.branch[22].block[14].um_I.iw[2] ;
 wire \top_I.branch[22].block[14].um_I.iw[3] ;
 wire \top_I.branch[22].block[14].um_I.iw[4] ;
 wire \top_I.branch[22].block[14].um_I.iw[5] ;
 wire \top_I.branch[22].block[14].um_I.iw[6] ;
 wire \top_I.branch[22].block[14].um_I.iw[7] ;
 wire \top_I.branch[22].block[14].um_I.iw[8] ;
 wire \top_I.branch[22].block[14].um_I.iw[9] ;
 wire \top_I.branch[22].block[14].um_I.k_zero ;
 wire \top_I.branch[22].block[14].um_I.pg_vdd ;
 wire \top_I.branch[22].block[15].um_I.ana[2] ;
 wire \top_I.branch[22].block[15].um_I.ana[3] ;
 wire \top_I.branch[22].block[15].um_I.ana[4] ;
 wire \top_I.branch[22].block[15].um_I.ana[5] ;
 wire \top_I.branch[22].block[15].um_I.ana[6] ;
 wire \top_I.branch[22].block[15].um_I.ana[7] ;
 wire \top_I.branch[22].block[15].um_I.clk ;
 wire \top_I.branch[22].block[15].um_I.ena ;
 wire \top_I.branch[22].block[15].um_I.iw[10] ;
 wire \top_I.branch[22].block[15].um_I.iw[11] ;
 wire \top_I.branch[22].block[15].um_I.iw[12] ;
 wire \top_I.branch[22].block[15].um_I.iw[13] ;
 wire \top_I.branch[22].block[15].um_I.iw[14] ;
 wire \top_I.branch[22].block[15].um_I.iw[15] ;
 wire \top_I.branch[22].block[15].um_I.iw[16] ;
 wire \top_I.branch[22].block[15].um_I.iw[17] ;
 wire \top_I.branch[22].block[15].um_I.iw[1] ;
 wire \top_I.branch[22].block[15].um_I.iw[2] ;
 wire \top_I.branch[22].block[15].um_I.iw[3] ;
 wire \top_I.branch[22].block[15].um_I.iw[4] ;
 wire \top_I.branch[22].block[15].um_I.iw[5] ;
 wire \top_I.branch[22].block[15].um_I.iw[6] ;
 wire \top_I.branch[22].block[15].um_I.iw[7] ;
 wire \top_I.branch[22].block[15].um_I.iw[8] ;
 wire \top_I.branch[22].block[15].um_I.iw[9] ;
 wire \top_I.branch[22].block[15].um_I.k_zero ;
 wire \top_I.branch[22].block[15].um_I.pg_vdd ;
 wire \top_I.branch[22].block[1].um_I.ana[2] ;
 wire \top_I.branch[22].block[1].um_I.ana[3] ;
 wire \top_I.branch[22].block[1].um_I.ana[4] ;
 wire \top_I.branch[22].block[1].um_I.ana[5] ;
 wire \top_I.branch[22].block[1].um_I.ana[6] ;
 wire \top_I.branch[22].block[1].um_I.ana[7] ;
 wire \top_I.branch[22].block[1].um_I.clk ;
 wire \top_I.branch[22].block[1].um_I.ena ;
 wire \top_I.branch[22].block[1].um_I.iw[10] ;
 wire \top_I.branch[22].block[1].um_I.iw[11] ;
 wire \top_I.branch[22].block[1].um_I.iw[12] ;
 wire \top_I.branch[22].block[1].um_I.iw[13] ;
 wire \top_I.branch[22].block[1].um_I.iw[14] ;
 wire \top_I.branch[22].block[1].um_I.iw[15] ;
 wire \top_I.branch[22].block[1].um_I.iw[16] ;
 wire \top_I.branch[22].block[1].um_I.iw[17] ;
 wire \top_I.branch[22].block[1].um_I.iw[1] ;
 wire \top_I.branch[22].block[1].um_I.iw[2] ;
 wire \top_I.branch[22].block[1].um_I.iw[3] ;
 wire \top_I.branch[22].block[1].um_I.iw[4] ;
 wire \top_I.branch[22].block[1].um_I.iw[5] ;
 wire \top_I.branch[22].block[1].um_I.iw[6] ;
 wire \top_I.branch[22].block[1].um_I.iw[7] ;
 wire \top_I.branch[22].block[1].um_I.iw[8] ;
 wire \top_I.branch[22].block[1].um_I.iw[9] ;
 wire \top_I.branch[22].block[1].um_I.k_zero ;
 wire \top_I.branch[22].block[1].um_I.pg_vdd ;
 wire \top_I.branch[22].block[2].um_I.ana[2] ;
 wire \top_I.branch[22].block[2].um_I.ana[3] ;
 wire \top_I.branch[22].block[2].um_I.ana[4] ;
 wire \top_I.branch[22].block[2].um_I.ana[5] ;
 wire \top_I.branch[22].block[2].um_I.ana[6] ;
 wire \top_I.branch[22].block[2].um_I.ana[7] ;
 wire \top_I.branch[22].block[2].um_I.clk ;
 wire \top_I.branch[22].block[2].um_I.ena ;
 wire \top_I.branch[22].block[2].um_I.iw[10] ;
 wire \top_I.branch[22].block[2].um_I.iw[11] ;
 wire \top_I.branch[22].block[2].um_I.iw[12] ;
 wire \top_I.branch[22].block[2].um_I.iw[13] ;
 wire \top_I.branch[22].block[2].um_I.iw[14] ;
 wire \top_I.branch[22].block[2].um_I.iw[15] ;
 wire \top_I.branch[22].block[2].um_I.iw[16] ;
 wire \top_I.branch[22].block[2].um_I.iw[17] ;
 wire \top_I.branch[22].block[2].um_I.iw[1] ;
 wire \top_I.branch[22].block[2].um_I.iw[2] ;
 wire \top_I.branch[22].block[2].um_I.iw[3] ;
 wire \top_I.branch[22].block[2].um_I.iw[4] ;
 wire \top_I.branch[22].block[2].um_I.iw[5] ;
 wire \top_I.branch[22].block[2].um_I.iw[6] ;
 wire \top_I.branch[22].block[2].um_I.iw[7] ;
 wire \top_I.branch[22].block[2].um_I.iw[8] ;
 wire \top_I.branch[22].block[2].um_I.iw[9] ;
 wire \top_I.branch[22].block[2].um_I.k_zero ;
 wire \top_I.branch[22].block[2].um_I.pg_vdd ;
 wire \top_I.branch[22].block[3].um_I.ana[2] ;
 wire \top_I.branch[22].block[3].um_I.ana[3] ;
 wire \top_I.branch[22].block[3].um_I.ana[4] ;
 wire \top_I.branch[22].block[3].um_I.ana[5] ;
 wire \top_I.branch[22].block[3].um_I.ana[6] ;
 wire \top_I.branch[22].block[3].um_I.ana[7] ;
 wire \top_I.branch[22].block[3].um_I.clk ;
 wire \top_I.branch[22].block[3].um_I.ena ;
 wire \top_I.branch[22].block[3].um_I.iw[10] ;
 wire \top_I.branch[22].block[3].um_I.iw[11] ;
 wire \top_I.branch[22].block[3].um_I.iw[12] ;
 wire \top_I.branch[22].block[3].um_I.iw[13] ;
 wire \top_I.branch[22].block[3].um_I.iw[14] ;
 wire \top_I.branch[22].block[3].um_I.iw[15] ;
 wire \top_I.branch[22].block[3].um_I.iw[16] ;
 wire \top_I.branch[22].block[3].um_I.iw[17] ;
 wire \top_I.branch[22].block[3].um_I.iw[1] ;
 wire \top_I.branch[22].block[3].um_I.iw[2] ;
 wire \top_I.branch[22].block[3].um_I.iw[3] ;
 wire \top_I.branch[22].block[3].um_I.iw[4] ;
 wire \top_I.branch[22].block[3].um_I.iw[5] ;
 wire \top_I.branch[22].block[3].um_I.iw[6] ;
 wire \top_I.branch[22].block[3].um_I.iw[7] ;
 wire \top_I.branch[22].block[3].um_I.iw[8] ;
 wire \top_I.branch[22].block[3].um_I.iw[9] ;
 wire \top_I.branch[22].block[3].um_I.k_zero ;
 wire \top_I.branch[22].block[3].um_I.pg_vdd ;
 wire \top_I.branch[22].block[4].um_I.ana[2] ;
 wire \top_I.branch[22].block[4].um_I.ana[3] ;
 wire \top_I.branch[22].block[4].um_I.ana[4] ;
 wire \top_I.branch[22].block[4].um_I.ana[5] ;
 wire \top_I.branch[22].block[4].um_I.ana[6] ;
 wire \top_I.branch[22].block[4].um_I.ana[7] ;
 wire \top_I.branch[22].block[4].um_I.clk ;
 wire \top_I.branch[22].block[4].um_I.ena ;
 wire \top_I.branch[22].block[4].um_I.iw[10] ;
 wire \top_I.branch[22].block[4].um_I.iw[11] ;
 wire \top_I.branch[22].block[4].um_I.iw[12] ;
 wire \top_I.branch[22].block[4].um_I.iw[13] ;
 wire \top_I.branch[22].block[4].um_I.iw[14] ;
 wire \top_I.branch[22].block[4].um_I.iw[15] ;
 wire \top_I.branch[22].block[4].um_I.iw[16] ;
 wire \top_I.branch[22].block[4].um_I.iw[17] ;
 wire \top_I.branch[22].block[4].um_I.iw[1] ;
 wire \top_I.branch[22].block[4].um_I.iw[2] ;
 wire \top_I.branch[22].block[4].um_I.iw[3] ;
 wire \top_I.branch[22].block[4].um_I.iw[4] ;
 wire \top_I.branch[22].block[4].um_I.iw[5] ;
 wire \top_I.branch[22].block[4].um_I.iw[6] ;
 wire \top_I.branch[22].block[4].um_I.iw[7] ;
 wire \top_I.branch[22].block[4].um_I.iw[8] ;
 wire \top_I.branch[22].block[4].um_I.iw[9] ;
 wire \top_I.branch[22].block[4].um_I.k_zero ;
 wire \top_I.branch[22].block[4].um_I.pg_vdd ;
 wire \top_I.branch[22].block[5].um_I.ana[2] ;
 wire \top_I.branch[22].block[5].um_I.ana[3] ;
 wire \top_I.branch[22].block[5].um_I.ana[4] ;
 wire \top_I.branch[22].block[5].um_I.ana[5] ;
 wire \top_I.branch[22].block[5].um_I.ana[6] ;
 wire \top_I.branch[22].block[5].um_I.ana[7] ;
 wire \top_I.branch[22].block[5].um_I.clk ;
 wire \top_I.branch[22].block[5].um_I.ena ;
 wire \top_I.branch[22].block[5].um_I.iw[10] ;
 wire \top_I.branch[22].block[5].um_I.iw[11] ;
 wire \top_I.branch[22].block[5].um_I.iw[12] ;
 wire \top_I.branch[22].block[5].um_I.iw[13] ;
 wire \top_I.branch[22].block[5].um_I.iw[14] ;
 wire \top_I.branch[22].block[5].um_I.iw[15] ;
 wire \top_I.branch[22].block[5].um_I.iw[16] ;
 wire \top_I.branch[22].block[5].um_I.iw[17] ;
 wire \top_I.branch[22].block[5].um_I.iw[1] ;
 wire \top_I.branch[22].block[5].um_I.iw[2] ;
 wire \top_I.branch[22].block[5].um_I.iw[3] ;
 wire \top_I.branch[22].block[5].um_I.iw[4] ;
 wire \top_I.branch[22].block[5].um_I.iw[5] ;
 wire \top_I.branch[22].block[5].um_I.iw[6] ;
 wire \top_I.branch[22].block[5].um_I.iw[7] ;
 wire \top_I.branch[22].block[5].um_I.iw[8] ;
 wire \top_I.branch[22].block[5].um_I.iw[9] ;
 wire \top_I.branch[22].block[5].um_I.k_zero ;
 wire \top_I.branch[22].block[5].um_I.pg_vdd ;
 wire \top_I.branch[22].block[6].um_I.ana[2] ;
 wire \top_I.branch[22].block[6].um_I.ana[3] ;
 wire \top_I.branch[22].block[6].um_I.ana[4] ;
 wire \top_I.branch[22].block[6].um_I.ana[5] ;
 wire \top_I.branch[22].block[6].um_I.ana[6] ;
 wire \top_I.branch[22].block[6].um_I.ana[7] ;
 wire \top_I.branch[22].block[6].um_I.clk ;
 wire \top_I.branch[22].block[6].um_I.ena ;
 wire \top_I.branch[22].block[6].um_I.iw[10] ;
 wire \top_I.branch[22].block[6].um_I.iw[11] ;
 wire \top_I.branch[22].block[6].um_I.iw[12] ;
 wire \top_I.branch[22].block[6].um_I.iw[13] ;
 wire \top_I.branch[22].block[6].um_I.iw[14] ;
 wire \top_I.branch[22].block[6].um_I.iw[15] ;
 wire \top_I.branch[22].block[6].um_I.iw[16] ;
 wire \top_I.branch[22].block[6].um_I.iw[17] ;
 wire \top_I.branch[22].block[6].um_I.iw[1] ;
 wire \top_I.branch[22].block[6].um_I.iw[2] ;
 wire \top_I.branch[22].block[6].um_I.iw[3] ;
 wire \top_I.branch[22].block[6].um_I.iw[4] ;
 wire \top_I.branch[22].block[6].um_I.iw[5] ;
 wire \top_I.branch[22].block[6].um_I.iw[6] ;
 wire \top_I.branch[22].block[6].um_I.iw[7] ;
 wire \top_I.branch[22].block[6].um_I.iw[8] ;
 wire \top_I.branch[22].block[6].um_I.iw[9] ;
 wire \top_I.branch[22].block[6].um_I.k_zero ;
 wire \top_I.branch[22].block[6].um_I.pg_vdd ;
 wire \top_I.branch[22].block[7].um_I.ana[2] ;
 wire \top_I.branch[22].block[7].um_I.ana[3] ;
 wire \top_I.branch[22].block[7].um_I.ana[4] ;
 wire \top_I.branch[22].block[7].um_I.ana[5] ;
 wire \top_I.branch[22].block[7].um_I.ana[6] ;
 wire \top_I.branch[22].block[7].um_I.ana[7] ;
 wire \top_I.branch[22].block[7].um_I.clk ;
 wire \top_I.branch[22].block[7].um_I.ena ;
 wire \top_I.branch[22].block[7].um_I.iw[10] ;
 wire \top_I.branch[22].block[7].um_I.iw[11] ;
 wire \top_I.branch[22].block[7].um_I.iw[12] ;
 wire \top_I.branch[22].block[7].um_I.iw[13] ;
 wire \top_I.branch[22].block[7].um_I.iw[14] ;
 wire \top_I.branch[22].block[7].um_I.iw[15] ;
 wire \top_I.branch[22].block[7].um_I.iw[16] ;
 wire \top_I.branch[22].block[7].um_I.iw[17] ;
 wire \top_I.branch[22].block[7].um_I.iw[1] ;
 wire \top_I.branch[22].block[7].um_I.iw[2] ;
 wire \top_I.branch[22].block[7].um_I.iw[3] ;
 wire \top_I.branch[22].block[7].um_I.iw[4] ;
 wire \top_I.branch[22].block[7].um_I.iw[5] ;
 wire \top_I.branch[22].block[7].um_I.iw[6] ;
 wire \top_I.branch[22].block[7].um_I.iw[7] ;
 wire \top_I.branch[22].block[7].um_I.iw[8] ;
 wire \top_I.branch[22].block[7].um_I.iw[9] ;
 wire \top_I.branch[22].block[7].um_I.k_zero ;
 wire \top_I.branch[22].block[7].um_I.pg_vdd ;
 wire \top_I.branch[22].block[8].um_I.ana[2] ;
 wire \top_I.branch[22].block[8].um_I.ana[3] ;
 wire \top_I.branch[22].block[8].um_I.ana[4] ;
 wire \top_I.branch[22].block[8].um_I.ana[5] ;
 wire \top_I.branch[22].block[8].um_I.ana[6] ;
 wire \top_I.branch[22].block[8].um_I.ana[7] ;
 wire \top_I.branch[22].block[8].um_I.clk ;
 wire \top_I.branch[22].block[8].um_I.ena ;
 wire \top_I.branch[22].block[8].um_I.iw[10] ;
 wire \top_I.branch[22].block[8].um_I.iw[11] ;
 wire \top_I.branch[22].block[8].um_I.iw[12] ;
 wire \top_I.branch[22].block[8].um_I.iw[13] ;
 wire \top_I.branch[22].block[8].um_I.iw[14] ;
 wire \top_I.branch[22].block[8].um_I.iw[15] ;
 wire \top_I.branch[22].block[8].um_I.iw[16] ;
 wire \top_I.branch[22].block[8].um_I.iw[17] ;
 wire \top_I.branch[22].block[8].um_I.iw[1] ;
 wire \top_I.branch[22].block[8].um_I.iw[2] ;
 wire \top_I.branch[22].block[8].um_I.iw[3] ;
 wire \top_I.branch[22].block[8].um_I.iw[4] ;
 wire \top_I.branch[22].block[8].um_I.iw[5] ;
 wire \top_I.branch[22].block[8].um_I.iw[6] ;
 wire \top_I.branch[22].block[8].um_I.iw[7] ;
 wire \top_I.branch[22].block[8].um_I.iw[8] ;
 wire \top_I.branch[22].block[8].um_I.iw[9] ;
 wire \top_I.branch[22].block[8].um_I.k_zero ;
 wire \top_I.branch[22].block[8].um_I.pg_vdd ;
 wire \top_I.branch[22].block[9].um_I.ana[2] ;
 wire \top_I.branch[22].block[9].um_I.ana[3] ;
 wire \top_I.branch[22].block[9].um_I.ana[4] ;
 wire \top_I.branch[22].block[9].um_I.ana[5] ;
 wire \top_I.branch[22].block[9].um_I.ana[6] ;
 wire \top_I.branch[22].block[9].um_I.ana[7] ;
 wire \top_I.branch[22].block[9].um_I.clk ;
 wire \top_I.branch[22].block[9].um_I.ena ;
 wire \top_I.branch[22].block[9].um_I.iw[10] ;
 wire \top_I.branch[22].block[9].um_I.iw[11] ;
 wire \top_I.branch[22].block[9].um_I.iw[12] ;
 wire \top_I.branch[22].block[9].um_I.iw[13] ;
 wire \top_I.branch[22].block[9].um_I.iw[14] ;
 wire \top_I.branch[22].block[9].um_I.iw[15] ;
 wire \top_I.branch[22].block[9].um_I.iw[16] ;
 wire \top_I.branch[22].block[9].um_I.iw[17] ;
 wire \top_I.branch[22].block[9].um_I.iw[1] ;
 wire \top_I.branch[22].block[9].um_I.iw[2] ;
 wire \top_I.branch[22].block[9].um_I.iw[3] ;
 wire \top_I.branch[22].block[9].um_I.iw[4] ;
 wire \top_I.branch[22].block[9].um_I.iw[5] ;
 wire \top_I.branch[22].block[9].um_I.iw[6] ;
 wire \top_I.branch[22].block[9].um_I.iw[7] ;
 wire \top_I.branch[22].block[9].um_I.iw[8] ;
 wire \top_I.branch[22].block[9].um_I.iw[9] ;
 wire \top_I.branch[22].block[9].um_I.k_zero ;
 wire \top_I.branch[22].block[9].um_I.pg_vdd ;
 wire \top_I.branch[22].l_addr[0] ;
 wire \top_I.branch[22].l_addr[2] ;
 wire \top_I.branch[23].block[0].um_I.ana[2] ;
 wire \top_I.branch[23].block[0].um_I.ana[3] ;
 wire \top_I.branch[23].block[0].um_I.ana[4] ;
 wire \top_I.branch[23].block[0].um_I.ana[5] ;
 wire \top_I.branch[23].block[0].um_I.ana[6] ;
 wire \top_I.branch[23].block[0].um_I.ana[7] ;
 wire \top_I.branch[23].block[0].um_I.clk ;
 wire \top_I.branch[23].block[0].um_I.ena ;
 wire \top_I.branch[23].block[0].um_I.iw[10] ;
 wire \top_I.branch[23].block[0].um_I.iw[11] ;
 wire \top_I.branch[23].block[0].um_I.iw[12] ;
 wire \top_I.branch[23].block[0].um_I.iw[13] ;
 wire \top_I.branch[23].block[0].um_I.iw[14] ;
 wire \top_I.branch[23].block[0].um_I.iw[15] ;
 wire \top_I.branch[23].block[0].um_I.iw[16] ;
 wire \top_I.branch[23].block[0].um_I.iw[17] ;
 wire \top_I.branch[23].block[0].um_I.iw[1] ;
 wire \top_I.branch[23].block[0].um_I.iw[2] ;
 wire \top_I.branch[23].block[0].um_I.iw[3] ;
 wire \top_I.branch[23].block[0].um_I.iw[4] ;
 wire \top_I.branch[23].block[0].um_I.iw[5] ;
 wire \top_I.branch[23].block[0].um_I.iw[6] ;
 wire \top_I.branch[23].block[0].um_I.iw[7] ;
 wire \top_I.branch[23].block[0].um_I.iw[8] ;
 wire \top_I.branch[23].block[0].um_I.iw[9] ;
 wire \top_I.branch[23].block[0].um_I.k_zero ;
 wire \top_I.branch[23].block[0].um_I.pg_vdd ;
 wire \top_I.branch[23].block[10].um_I.ana[2] ;
 wire \top_I.branch[23].block[10].um_I.ana[3] ;
 wire \top_I.branch[23].block[10].um_I.ana[4] ;
 wire \top_I.branch[23].block[10].um_I.ana[5] ;
 wire \top_I.branch[23].block[10].um_I.ana[6] ;
 wire \top_I.branch[23].block[10].um_I.ana[7] ;
 wire \top_I.branch[23].block[10].um_I.clk ;
 wire \top_I.branch[23].block[10].um_I.ena ;
 wire \top_I.branch[23].block[10].um_I.iw[10] ;
 wire \top_I.branch[23].block[10].um_I.iw[11] ;
 wire \top_I.branch[23].block[10].um_I.iw[12] ;
 wire \top_I.branch[23].block[10].um_I.iw[13] ;
 wire \top_I.branch[23].block[10].um_I.iw[14] ;
 wire \top_I.branch[23].block[10].um_I.iw[15] ;
 wire \top_I.branch[23].block[10].um_I.iw[16] ;
 wire \top_I.branch[23].block[10].um_I.iw[17] ;
 wire \top_I.branch[23].block[10].um_I.iw[1] ;
 wire \top_I.branch[23].block[10].um_I.iw[2] ;
 wire \top_I.branch[23].block[10].um_I.iw[3] ;
 wire \top_I.branch[23].block[10].um_I.iw[4] ;
 wire \top_I.branch[23].block[10].um_I.iw[5] ;
 wire \top_I.branch[23].block[10].um_I.iw[6] ;
 wire \top_I.branch[23].block[10].um_I.iw[7] ;
 wire \top_I.branch[23].block[10].um_I.iw[8] ;
 wire \top_I.branch[23].block[10].um_I.iw[9] ;
 wire \top_I.branch[23].block[10].um_I.k_zero ;
 wire \top_I.branch[23].block[10].um_I.pg_vdd ;
 wire \top_I.branch[23].block[11].um_I.ana[2] ;
 wire \top_I.branch[23].block[11].um_I.ana[3] ;
 wire \top_I.branch[23].block[11].um_I.ana[4] ;
 wire \top_I.branch[23].block[11].um_I.ana[5] ;
 wire \top_I.branch[23].block[11].um_I.ana[6] ;
 wire \top_I.branch[23].block[11].um_I.ana[7] ;
 wire \top_I.branch[23].block[11].um_I.clk ;
 wire \top_I.branch[23].block[11].um_I.ena ;
 wire \top_I.branch[23].block[11].um_I.iw[10] ;
 wire \top_I.branch[23].block[11].um_I.iw[11] ;
 wire \top_I.branch[23].block[11].um_I.iw[12] ;
 wire \top_I.branch[23].block[11].um_I.iw[13] ;
 wire \top_I.branch[23].block[11].um_I.iw[14] ;
 wire \top_I.branch[23].block[11].um_I.iw[15] ;
 wire \top_I.branch[23].block[11].um_I.iw[16] ;
 wire \top_I.branch[23].block[11].um_I.iw[17] ;
 wire \top_I.branch[23].block[11].um_I.iw[1] ;
 wire \top_I.branch[23].block[11].um_I.iw[2] ;
 wire \top_I.branch[23].block[11].um_I.iw[3] ;
 wire \top_I.branch[23].block[11].um_I.iw[4] ;
 wire \top_I.branch[23].block[11].um_I.iw[5] ;
 wire \top_I.branch[23].block[11].um_I.iw[6] ;
 wire \top_I.branch[23].block[11].um_I.iw[7] ;
 wire \top_I.branch[23].block[11].um_I.iw[8] ;
 wire \top_I.branch[23].block[11].um_I.iw[9] ;
 wire \top_I.branch[23].block[11].um_I.k_zero ;
 wire \top_I.branch[23].block[11].um_I.pg_vdd ;
 wire \top_I.branch[23].block[12].um_I.ana[2] ;
 wire \top_I.branch[23].block[12].um_I.ana[3] ;
 wire \top_I.branch[23].block[12].um_I.ana[4] ;
 wire \top_I.branch[23].block[12].um_I.ana[5] ;
 wire \top_I.branch[23].block[12].um_I.ana[6] ;
 wire \top_I.branch[23].block[12].um_I.ana[7] ;
 wire \top_I.branch[23].block[12].um_I.clk ;
 wire \top_I.branch[23].block[12].um_I.ena ;
 wire \top_I.branch[23].block[12].um_I.iw[10] ;
 wire \top_I.branch[23].block[12].um_I.iw[11] ;
 wire \top_I.branch[23].block[12].um_I.iw[12] ;
 wire \top_I.branch[23].block[12].um_I.iw[13] ;
 wire \top_I.branch[23].block[12].um_I.iw[14] ;
 wire \top_I.branch[23].block[12].um_I.iw[15] ;
 wire \top_I.branch[23].block[12].um_I.iw[16] ;
 wire \top_I.branch[23].block[12].um_I.iw[17] ;
 wire \top_I.branch[23].block[12].um_I.iw[1] ;
 wire \top_I.branch[23].block[12].um_I.iw[2] ;
 wire \top_I.branch[23].block[12].um_I.iw[3] ;
 wire \top_I.branch[23].block[12].um_I.iw[4] ;
 wire \top_I.branch[23].block[12].um_I.iw[5] ;
 wire \top_I.branch[23].block[12].um_I.iw[6] ;
 wire \top_I.branch[23].block[12].um_I.iw[7] ;
 wire \top_I.branch[23].block[12].um_I.iw[8] ;
 wire \top_I.branch[23].block[12].um_I.iw[9] ;
 wire \top_I.branch[23].block[12].um_I.k_zero ;
 wire \top_I.branch[23].block[12].um_I.pg_vdd ;
 wire \top_I.branch[23].block[13].um_I.ana[2] ;
 wire \top_I.branch[23].block[13].um_I.ana[3] ;
 wire \top_I.branch[23].block[13].um_I.ana[4] ;
 wire \top_I.branch[23].block[13].um_I.ana[5] ;
 wire \top_I.branch[23].block[13].um_I.ana[6] ;
 wire \top_I.branch[23].block[13].um_I.ana[7] ;
 wire \top_I.branch[23].block[13].um_I.clk ;
 wire \top_I.branch[23].block[13].um_I.ena ;
 wire \top_I.branch[23].block[13].um_I.iw[10] ;
 wire \top_I.branch[23].block[13].um_I.iw[11] ;
 wire \top_I.branch[23].block[13].um_I.iw[12] ;
 wire \top_I.branch[23].block[13].um_I.iw[13] ;
 wire \top_I.branch[23].block[13].um_I.iw[14] ;
 wire \top_I.branch[23].block[13].um_I.iw[15] ;
 wire \top_I.branch[23].block[13].um_I.iw[16] ;
 wire \top_I.branch[23].block[13].um_I.iw[17] ;
 wire \top_I.branch[23].block[13].um_I.iw[1] ;
 wire \top_I.branch[23].block[13].um_I.iw[2] ;
 wire \top_I.branch[23].block[13].um_I.iw[3] ;
 wire \top_I.branch[23].block[13].um_I.iw[4] ;
 wire \top_I.branch[23].block[13].um_I.iw[5] ;
 wire \top_I.branch[23].block[13].um_I.iw[6] ;
 wire \top_I.branch[23].block[13].um_I.iw[7] ;
 wire \top_I.branch[23].block[13].um_I.iw[8] ;
 wire \top_I.branch[23].block[13].um_I.iw[9] ;
 wire \top_I.branch[23].block[13].um_I.k_zero ;
 wire \top_I.branch[23].block[13].um_I.pg_vdd ;
 wire \top_I.branch[23].block[14].um_I.ana[2] ;
 wire \top_I.branch[23].block[14].um_I.ana[3] ;
 wire \top_I.branch[23].block[14].um_I.ana[4] ;
 wire \top_I.branch[23].block[14].um_I.ana[5] ;
 wire \top_I.branch[23].block[14].um_I.ana[6] ;
 wire \top_I.branch[23].block[14].um_I.ana[7] ;
 wire \top_I.branch[23].block[14].um_I.clk ;
 wire \top_I.branch[23].block[14].um_I.ena ;
 wire \top_I.branch[23].block[14].um_I.iw[10] ;
 wire \top_I.branch[23].block[14].um_I.iw[11] ;
 wire \top_I.branch[23].block[14].um_I.iw[12] ;
 wire \top_I.branch[23].block[14].um_I.iw[13] ;
 wire \top_I.branch[23].block[14].um_I.iw[14] ;
 wire \top_I.branch[23].block[14].um_I.iw[15] ;
 wire \top_I.branch[23].block[14].um_I.iw[16] ;
 wire \top_I.branch[23].block[14].um_I.iw[17] ;
 wire \top_I.branch[23].block[14].um_I.iw[1] ;
 wire \top_I.branch[23].block[14].um_I.iw[2] ;
 wire \top_I.branch[23].block[14].um_I.iw[3] ;
 wire \top_I.branch[23].block[14].um_I.iw[4] ;
 wire \top_I.branch[23].block[14].um_I.iw[5] ;
 wire \top_I.branch[23].block[14].um_I.iw[6] ;
 wire \top_I.branch[23].block[14].um_I.iw[7] ;
 wire \top_I.branch[23].block[14].um_I.iw[8] ;
 wire \top_I.branch[23].block[14].um_I.iw[9] ;
 wire \top_I.branch[23].block[14].um_I.k_zero ;
 wire \top_I.branch[23].block[14].um_I.pg_vdd ;
 wire \top_I.branch[23].block[15].um_I.ana[2] ;
 wire \top_I.branch[23].block[15].um_I.ana[3] ;
 wire \top_I.branch[23].block[15].um_I.ana[4] ;
 wire \top_I.branch[23].block[15].um_I.ana[5] ;
 wire \top_I.branch[23].block[15].um_I.ana[6] ;
 wire \top_I.branch[23].block[15].um_I.ana[7] ;
 wire \top_I.branch[23].block[15].um_I.clk ;
 wire \top_I.branch[23].block[15].um_I.ena ;
 wire \top_I.branch[23].block[15].um_I.iw[10] ;
 wire \top_I.branch[23].block[15].um_I.iw[11] ;
 wire \top_I.branch[23].block[15].um_I.iw[12] ;
 wire \top_I.branch[23].block[15].um_I.iw[13] ;
 wire \top_I.branch[23].block[15].um_I.iw[14] ;
 wire \top_I.branch[23].block[15].um_I.iw[15] ;
 wire \top_I.branch[23].block[15].um_I.iw[16] ;
 wire \top_I.branch[23].block[15].um_I.iw[17] ;
 wire \top_I.branch[23].block[15].um_I.iw[1] ;
 wire \top_I.branch[23].block[15].um_I.iw[2] ;
 wire \top_I.branch[23].block[15].um_I.iw[3] ;
 wire \top_I.branch[23].block[15].um_I.iw[4] ;
 wire \top_I.branch[23].block[15].um_I.iw[5] ;
 wire \top_I.branch[23].block[15].um_I.iw[6] ;
 wire \top_I.branch[23].block[15].um_I.iw[7] ;
 wire \top_I.branch[23].block[15].um_I.iw[8] ;
 wire \top_I.branch[23].block[15].um_I.iw[9] ;
 wire \top_I.branch[23].block[15].um_I.k_zero ;
 wire \top_I.branch[23].block[15].um_I.pg_vdd ;
 wire \top_I.branch[23].block[1].um_I.ana[2] ;
 wire \top_I.branch[23].block[1].um_I.ana[3] ;
 wire \top_I.branch[23].block[1].um_I.ana[4] ;
 wire \top_I.branch[23].block[1].um_I.ana[5] ;
 wire \top_I.branch[23].block[1].um_I.ana[6] ;
 wire \top_I.branch[23].block[1].um_I.ana[7] ;
 wire \top_I.branch[23].block[1].um_I.clk ;
 wire \top_I.branch[23].block[1].um_I.ena ;
 wire \top_I.branch[23].block[1].um_I.iw[10] ;
 wire \top_I.branch[23].block[1].um_I.iw[11] ;
 wire \top_I.branch[23].block[1].um_I.iw[12] ;
 wire \top_I.branch[23].block[1].um_I.iw[13] ;
 wire \top_I.branch[23].block[1].um_I.iw[14] ;
 wire \top_I.branch[23].block[1].um_I.iw[15] ;
 wire \top_I.branch[23].block[1].um_I.iw[16] ;
 wire \top_I.branch[23].block[1].um_I.iw[17] ;
 wire \top_I.branch[23].block[1].um_I.iw[1] ;
 wire \top_I.branch[23].block[1].um_I.iw[2] ;
 wire \top_I.branch[23].block[1].um_I.iw[3] ;
 wire \top_I.branch[23].block[1].um_I.iw[4] ;
 wire \top_I.branch[23].block[1].um_I.iw[5] ;
 wire \top_I.branch[23].block[1].um_I.iw[6] ;
 wire \top_I.branch[23].block[1].um_I.iw[7] ;
 wire \top_I.branch[23].block[1].um_I.iw[8] ;
 wire \top_I.branch[23].block[1].um_I.iw[9] ;
 wire \top_I.branch[23].block[1].um_I.k_zero ;
 wire \top_I.branch[23].block[1].um_I.pg_vdd ;
 wire \top_I.branch[23].block[2].um_I.ana[2] ;
 wire \top_I.branch[23].block[2].um_I.ana[3] ;
 wire \top_I.branch[23].block[2].um_I.ana[4] ;
 wire \top_I.branch[23].block[2].um_I.ana[5] ;
 wire \top_I.branch[23].block[2].um_I.ana[6] ;
 wire \top_I.branch[23].block[2].um_I.ana[7] ;
 wire \top_I.branch[23].block[2].um_I.clk ;
 wire \top_I.branch[23].block[2].um_I.ena ;
 wire \top_I.branch[23].block[2].um_I.iw[10] ;
 wire \top_I.branch[23].block[2].um_I.iw[11] ;
 wire \top_I.branch[23].block[2].um_I.iw[12] ;
 wire \top_I.branch[23].block[2].um_I.iw[13] ;
 wire \top_I.branch[23].block[2].um_I.iw[14] ;
 wire \top_I.branch[23].block[2].um_I.iw[15] ;
 wire \top_I.branch[23].block[2].um_I.iw[16] ;
 wire \top_I.branch[23].block[2].um_I.iw[17] ;
 wire \top_I.branch[23].block[2].um_I.iw[1] ;
 wire \top_I.branch[23].block[2].um_I.iw[2] ;
 wire \top_I.branch[23].block[2].um_I.iw[3] ;
 wire \top_I.branch[23].block[2].um_I.iw[4] ;
 wire \top_I.branch[23].block[2].um_I.iw[5] ;
 wire \top_I.branch[23].block[2].um_I.iw[6] ;
 wire \top_I.branch[23].block[2].um_I.iw[7] ;
 wire \top_I.branch[23].block[2].um_I.iw[8] ;
 wire \top_I.branch[23].block[2].um_I.iw[9] ;
 wire \top_I.branch[23].block[2].um_I.k_zero ;
 wire \top_I.branch[23].block[2].um_I.pg_vdd ;
 wire \top_I.branch[23].block[3].um_I.ana[2] ;
 wire \top_I.branch[23].block[3].um_I.ana[3] ;
 wire \top_I.branch[23].block[3].um_I.ana[4] ;
 wire \top_I.branch[23].block[3].um_I.ana[5] ;
 wire \top_I.branch[23].block[3].um_I.ana[6] ;
 wire \top_I.branch[23].block[3].um_I.ana[7] ;
 wire \top_I.branch[23].block[3].um_I.clk ;
 wire \top_I.branch[23].block[3].um_I.ena ;
 wire \top_I.branch[23].block[3].um_I.iw[10] ;
 wire \top_I.branch[23].block[3].um_I.iw[11] ;
 wire \top_I.branch[23].block[3].um_I.iw[12] ;
 wire \top_I.branch[23].block[3].um_I.iw[13] ;
 wire \top_I.branch[23].block[3].um_I.iw[14] ;
 wire \top_I.branch[23].block[3].um_I.iw[15] ;
 wire \top_I.branch[23].block[3].um_I.iw[16] ;
 wire \top_I.branch[23].block[3].um_I.iw[17] ;
 wire \top_I.branch[23].block[3].um_I.iw[1] ;
 wire \top_I.branch[23].block[3].um_I.iw[2] ;
 wire \top_I.branch[23].block[3].um_I.iw[3] ;
 wire \top_I.branch[23].block[3].um_I.iw[4] ;
 wire \top_I.branch[23].block[3].um_I.iw[5] ;
 wire \top_I.branch[23].block[3].um_I.iw[6] ;
 wire \top_I.branch[23].block[3].um_I.iw[7] ;
 wire \top_I.branch[23].block[3].um_I.iw[8] ;
 wire \top_I.branch[23].block[3].um_I.iw[9] ;
 wire \top_I.branch[23].block[3].um_I.k_zero ;
 wire \top_I.branch[23].block[3].um_I.pg_vdd ;
 wire \top_I.branch[23].block[4].um_I.ana[2] ;
 wire \top_I.branch[23].block[4].um_I.ana[3] ;
 wire \top_I.branch[23].block[4].um_I.ana[4] ;
 wire \top_I.branch[23].block[4].um_I.ana[5] ;
 wire \top_I.branch[23].block[4].um_I.ana[6] ;
 wire \top_I.branch[23].block[4].um_I.ana[7] ;
 wire \top_I.branch[23].block[4].um_I.clk ;
 wire \top_I.branch[23].block[4].um_I.ena ;
 wire \top_I.branch[23].block[4].um_I.iw[10] ;
 wire \top_I.branch[23].block[4].um_I.iw[11] ;
 wire \top_I.branch[23].block[4].um_I.iw[12] ;
 wire \top_I.branch[23].block[4].um_I.iw[13] ;
 wire \top_I.branch[23].block[4].um_I.iw[14] ;
 wire \top_I.branch[23].block[4].um_I.iw[15] ;
 wire \top_I.branch[23].block[4].um_I.iw[16] ;
 wire \top_I.branch[23].block[4].um_I.iw[17] ;
 wire \top_I.branch[23].block[4].um_I.iw[1] ;
 wire \top_I.branch[23].block[4].um_I.iw[2] ;
 wire \top_I.branch[23].block[4].um_I.iw[3] ;
 wire \top_I.branch[23].block[4].um_I.iw[4] ;
 wire \top_I.branch[23].block[4].um_I.iw[5] ;
 wire \top_I.branch[23].block[4].um_I.iw[6] ;
 wire \top_I.branch[23].block[4].um_I.iw[7] ;
 wire \top_I.branch[23].block[4].um_I.iw[8] ;
 wire \top_I.branch[23].block[4].um_I.iw[9] ;
 wire \top_I.branch[23].block[4].um_I.k_zero ;
 wire \top_I.branch[23].block[4].um_I.pg_vdd ;
 wire \top_I.branch[23].block[5].um_I.ana[2] ;
 wire \top_I.branch[23].block[5].um_I.ana[3] ;
 wire \top_I.branch[23].block[5].um_I.ana[4] ;
 wire \top_I.branch[23].block[5].um_I.ana[5] ;
 wire \top_I.branch[23].block[5].um_I.ana[6] ;
 wire \top_I.branch[23].block[5].um_I.ana[7] ;
 wire \top_I.branch[23].block[5].um_I.clk ;
 wire \top_I.branch[23].block[5].um_I.ena ;
 wire \top_I.branch[23].block[5].um_I.iw[10] ;
 wire \top_I.branch[23].block[5].um_I.iw[11] ;
 wire \top_I.branch[23].block[5].um_I.iw[12] ;
 wire \top_I.branch[23].block[5].um_I.iw[13] ;
 wire \top_I.branch[23].block[5].um_I.iw[14] ;
 wire \top_I.branch[23].block[5].um_I.iw[15] ;
 wire \top_I.branch[23].block[5].um_I.iw[16] ;
 wire \top_I.branch[23].block[5].um_I.iw[17] ;
 wire \top_I.branch[23].block[5].um_I.iw[1] ;
 wire \top_I.branch[23].block[5].um_I.iw[2] ;
 wire \top_I.branch[23].block[5].um_I.iw[3] ;
 wire \top_I.branch[23].block[5].um_I.iw[4] ;
 wire \top_I.branch[23].block[5].um_I.iw[5] ;
 wire \top_I.branch[23].block[5].um_I.iw[6] ;
 wire \top_I.branch[23].block[5].um_I.iw[7] ;
 wire \top_I.branch[23].block[5].um_I.iw[8] ;
 wire \top_I.branch[23].block[5].um_I.iw[9] ;
 wire \top_I.branch[23].block[5].um_I.k_zero ;
 wire \top_I.branch[23].block[5].um_I.pg_vdd ;
 wire \top_I.branch[23].block[6].um_I.ana[2] ;
 wire \top_I.branch[23].block[6].um_I.ana[3] ;
 wire \top_I.branch[23].block[6].um_I.ana[4] ;
 wire \top_I.branch[23].block[6].um_I.ana[5] ;
 wire \top_I.branch[23].block[6].um_I.ana[6] ;
 wire \top_I.branch[23].block[6].um_I.ana[7] ;
 wire \top_I.branch[23].block[6].um_I.clk ;
 wire \top_I.branch[23].block[6].um_I.ena ;
 wire \top_I.branch[23].block[6].um_I.iw[10] ;
 wire \top_I.branch[23].block[6].um_I.iw[11] ;
 wire \top_I.branch[23].block[6].um_I.iw[12] ;
 wire \top_I.branch[23].block[6].um_I.iw[13] ;
 wire \top_I.branch[23].block[6].um_I.iw[14] ;
 wire \top_I.branch[23].block[6].um_I.iw[15] ;
 wire \top_I.branch[23].block[6].um_I.iw[16] ;
 wire \top_I.branch[23].block[6].um_I.iw[17] ;
 wire \top_I.branch[23].block[6].um_I.iw[1] ;
 wire \top_I.branch[23].block[6].um_I.iw[2] ;
 wire \top_I.branch[23].block[6].um_I.iw[3] ;
 wire \top_I.branch[23].block[6].um_I.iw[4] ;
 wire \top_I.branch[23].block[6].um_I.iw[5] ;
 wire \top_I.branch[23].block[6].um_I.iw[6] ;
 wire \top_I.branch[23].block[6].um_I.iw[7] ;
 wire \top_I.branch[23].block[6].um_I.iw[8] ;
 wire \top_I.branch[23].block[6].um_I.iw[9] ;
 wire \top_I.branch[23].block[6].um_I.k_zero ;
 wire \top_I.branch[23].block[6].um_I.pg_vdd ;
 wire \top_I.branch[23].block[7].um_I.ana[2] ;
 wire \top_I.branch[23].block[7].um_I.ana[3] ;
 wire \top_I.branch[23].block[7].um_I.ana[4] ;
 wire \top_I.branch[23].block[7].um_I.ana[5] ;
 wire \top_I.branch[23].block[7].um_I.ana[6] ;
 wire \top_I.branch[23].block[7].um_I.ana[7] ;
 wire \top_I.branch[23].block[7].um_I.clk ;
 wire \top_I.branch[23].block[7].um_I.ena ;
 wire \top_I.branch[23].block[7].um_I.iw[10] ;
 wire \top_I.branch[23].block[7].um_I.iw[11] ;
 wire \top_I.branch[23].block[7].um_I.iw[12] ;
 wire \top_I.branch[23].block[7].um_I.iw[13] ;
 wire \top_I.branch[23].block[7].um_I.iw[14] ;
 wire \top_I.branch[23].block[7].um_I.iw[15] ;
 wire \top_I.branch[23].block[7].um_I.iw[16] ;
 wire \top_I.branch[23].block[7].um_I.iw[17] ;
 wire \top_I.branch[23].block[7].um_I.iw[1] ;
 wire \top_I.branch[23].block[7].um_I.iw[2] ;
 wire \top_I.branch[23].block[7].um_I.iw[3] ;
 wire \top_I.branch[23].block[7].um_I.iw[4] ;
 wire \top_I.branch[23].block[7].um_I.iw[5] ;
 wire \top_I.branch[23].block[7].um_I.iw[6] ;
 wire \top_I.branch[23].block[7].um_I.iw[7] ;
 wire \top_I.branch[23].block[7].um_I.iw[8] ;
 wire \top_I.branch[23].block[7].um_I.iw[9] ;
 wire \top_I.branch[23].block[7].um_I.k_zero ;
 wire \top_I.branch[23].block[7].um_I.pg_vdd ;
 wire \top_I.branch[23].block[8].um_I.ana[2] ;
 wire \top_I.branch[23].block[8].um_I.ana[3] ;
 wire \top_I.branch[23].block[8].um_I.ana[4] ;
 wire \top_I.branch[23].block[8].um_I.ana[5] ;
 wire \top_I.branch[23].block[8].um_I.ana[6] ;
 wire \top_I.branch[23].block[8].um_I.ana[7] ;
 wire \top_I.branch[23].block[8].um_I.clk ;
 wire \top_I.branch[23].block[8].um_I.ena ;
 wire \top_I.branch[23].block[8].um_I.iw[10] ;
 wire \top_I.branch[23].block[8].um_I.iw[11] ;
 wire \top_I.branch[23].block[8].um_I.iw[12] ;
 wire \top_I.branch[23].block[8].um_I.iw[13] ;
 wire \top_I.branch[23].block[8].um_I.iw[14] ;
 wire \top_I.branch[23].block[8].um_I.iw[15] ;
 wire \top_I.branch[23].block[8].um_I.iw[16] ;
 wire \top_I.branch[23].block[8].um_I.iw[17] ;
 wire \top_I.branch[23].block[8].um_I.iw[1] ;
 wire \top_I.branch[23].block[8].um_I.iw[2] ;
 wire \top_I.branch[23].block[8].um_I.iw[3] ;
 wire \top_I.branch[23].block[8].um_I.iw[4] ;
 wire \top_I.branch[23].block[8].um_I.iw[5] ;
 wire \top_I.branch[23].block[8].um_I.iw[6] ;
 wire \top_I.branch[23].block[8].um_I.iw[7] ;
 wire \top_I.branch[23].block[8].um_I.iw[8] ;
 wire \top_I.branch[23].block[8].um_I.iw[9] ;
 wire \top_I.branch[23].block[8].um_I.k_zero ;
 wire \top_I.branch[23].block[8].um_I.pg_vdd ;
 wire \top_I.branch[23].block[9].um_I.ana[2] ;
 wire \top_I.branch[23].block[9].um_I.ana[3] ;
 wire \top_I.branch[23].block[9].um_I.ana[4] ;
 wire \top_I.branch[23].block[9].um_I.ana[5] ;
 wire \top_I.branch[23].block[9].um_I.ana[6] ;
 wire \top_I.branch[23].block[9].um_I.ana[7] ;
 wire \top_I.branch[23].block[9].um_I.clk ;
 wire \top_I.branch[23].block[9].um_I.ena ;
 wire \top_I.branch[23].block[9].um_I.iw[10] ;
 wire \top_I.branch[23].block[9].um_I.iw[11] ;
 wire \top_I.branch[23].block[9].um_I.iw[12] ;
 wire \top_I.branch[23].block[9].um_I.iw[13] ;
 wire \top_I.branch[23].block[9].um_I.iw[14] ;
 wire \top_I.branch[23].block[9].um_I.iw[15] ;
 wire \top_I.branch[23].block[9].um_I.iw[16] ;
 wire \top_I.branch[23].block[9].um_I.iw[17] ;
 wire \top_I.branch[23].block[9].um_I.iw[1] ;
 wire \top_I.branch[23].block[9].um_I.iw[2] ;
 wire \top_I.branch[23].block[9].um_I.iw[3] ;
 wire \top_I.branch[23].block[9].um_I.iw[4] ;
 wire \top_I.branch[23].block[9].um_I.iw[5] ;
 wire \top_I.branch[23].block[9].um_I.iw[6] ;
 wire \top_I.branch[23].block[9].um_I.iw[7] ;
 wire \top_I.branch[23].block[9].um_I.iw[8] ;
 wire \top_I.branch[23].block[9].um_I.iw[9] ;
 wire \top_I.branch[23].block[9].um_I.k_zero ;
 wire \top_I.branch[23].block[9].um_I.pg_vdd ;
 wire \top_I.branch[23].l_addr[0] ;
 wire \top_I.branch[23].l_addr[2] ;
 wire \top_I.branch[2].block[0].um_I.ana[2] ;
 wire \top_I.branch[2].block[0].um_I.ana[3] ;
 wire \top_I.branch[2].block[0].um_I.ana[4] ;
 wire \top_I.branch[2].block[0].um_I.ana[5] ;
 wire \top_I.branch[2].block[0].um_I.ana[6] ;
 wire \top_I.branch[2].block[0].um_I.ana[7] ;
 wire \top_I.branch[2].block[0].um_I.clk ;
 wire \top_I.branch[2].block[0].um_I.ena ;
 wire \top_I.branch[2].block[0].um_I.iw[10] ;
 wire \top_I.branch[2].block[0].um_I.iw[11] ;
 wire \top_I.branch[2].block[0].um_I.iw[12] ;
 wire \top_I.branch[2].block[0].um_I.iw[13] ;
 wire \top_I.branch[2].block[0].um_I.iw[14] ;
 wire \top_I.branch[2].block[0].um_I.iw[15] ;
 wire \top_I.branch[2].block[0].um_I.iw[16] ;
 wire \top_I.branch[2].block[0].um_I.iw[17] ;
 wire \top_I.branch[2].block[0].um_I.iw[1] ;
 wire \top_I.branch[2].block[0].um_I.iw[2] ;
 wire \top_I.branch[2].block[0].um_I.iw[3] ;
 wire \top_I.branch[2].block[0].um_I.iw[4] ;
 wire \top_I.branch[2].block[0].um_I.iw[5] ;
 wire \top_I.branch[2].block[0].um_I.iw[6] ;
 wire \top_I.branch[2].block[0].um_I.iw[7] ;
 wire \top_I.branch[2].block[0].um_I.iw[8] ;
 wire \top_I.branch[2].block[0].um_I.iw[9] ;
 wire \top_I.branch[2].block[0].um_I.k_zero ;
 wire \top_I.branch[2].block[0].um_I.pg_vdd ;
 wire \top_I.branch[2].block[10].um_I.ana[2] ;
 wire \top_I.branch[2].block[10].um_I.ana[3] ;
 wire \top_I.branch[2].block[10].um_I.ana[4] ;
 wire \top_I.branch[2].block[10].um_I.ana[5] ;
 wire \top_I.branch[2].block[10].um_I.ana[6] ;
 wire \top_I.branch[2].block[10].um_I.ana[7] ;
 wire \top_I.branch[2].block[10].um_I.clk ;
 wire \top_I.branch[2].block[10].um_I.ena ;
 wire \top_I.branch[2].block[10].um_I.iw[10] ;
 wire \top_I.branch[2].block[10].um_I.iw[11] ;
 wire \top_I.branch[2].block[10].um_I.iw[12] ;
 wire \top_I.branch[2].block[10].um_I.iw[13] ;
 wire \top_I.branch[2].block[10].um_I.iw[14] ;
 wire \top_I.branch[2].block[10].um_I.iw[15] ;
 wire \top_I.branch[2].block[10].um_I.iw[16] ;
 wire \top_I.branch[2].block[10].um_I.iw[17] ;
 wire \top_I.branch[2].block[10].um_I.iw[1] ;
 wire \top_I.branch[2].block[10].um_I.iw[2] ;
 wire \top_I.branch[2].block[10].um_I.iw[3] ;
 wire \top_I.branch[2].block[10].um_I.iw[4] ;
 wire \top_I.branch[2].block[10].um_I.iw[5] ;
 wire \top_I.branch[2].block[10].um_I.iw[6] ;
 wire \top_I.branch[2].block[10].um_I.iw[7] ;
 wire \top_I.branch[2].block[10].um_I.iw[8] ;
 wire \top_I.branch[2].block[10].um_I.iw[9] ;
 wire \top_I.branch[2].block[10].um_I.k_zero ;
 wire \top_I.branch[2].block[10].um_I.pg_vdd ;
 wire \top_I.branch[2].block[11].um_I.ana[2] ;
 wire \top_I.branch[2].block[11].um_I.ana[3] ;
 wire \top_I.branch[2].block[11].um_I.ana[4] ;
 wire \top_I.branch[2].block[11].um_I.ana[5] ;
 wire \top_I.branch[2].block[11].um_I.ana[6] ;
 wire \top_I.branch[2].block[11].um_I.ana[7] ;
 wire \top_I.branch[2].block[11].um_I.clk ;
 wire \top_I.branch[2].block[11].um_I.ena ;
 wire \top_I.branch[2].block[11].um_I.iw[10] ;
 wire \top_I.branch[2].block[11].um_I.iw[11] ;
 wire \top_I.branch[2].block[11].um_I.iw[12] ;
 wire \top_I.branch[2].block[11].um_I.iw[13] ;
 wire \top_I.branch[2].block[11].um_I.iw[14] ;
 wire \top_I.branch[2].block[11].um_I.iw[15] ;
 wire \top_I.branch[2].block[11].um_I.iw[16] ;
 wire \top_I.branch[2].block[11].um_I.iw[17] ;
 wire \top_I.branch[2].block[11].um_I.iw[1] ;
 wire \top_I.branch[2].block[11].um_I.iw[2] ;
 wire \top_I.branch[2].block[11].um_I.iw[3] ;
 wire \top_I.branch[2].block[11].um_I.iw[4] ;
 wire \top_I.branch[2].block[11].um_I.iw[5] ;
 wire \top_I.branch[2].block[11].um_I.iw[6] ;
 wire \top_I.branch[2].block[11].um_I.iw[7] ;
 wire \top_I.branch[2].block[11].um_I.iw[8] ;
 wire \top_I.branch[2].block[11].um_I.iw[9] ;
 wire \top_I.branch[2].block[11].um_I.k_zero ;
 wire \top_I.branch[2].block[11].um_I.pg_vdd ;
 wire \top_I.branch[2].block[12].um_I.ana[2] ;
 wire \top_I.branch[2].block[12].um_I.ana[3] ;
 wire \top_I.branch[2].block[12].um_I.ana[4] ;
 wire \top_I.branch[2].block[12].um_I.ana[5] ;
 wire \top_I.branch[2].block[12].um_I.ana[6] ;
 wire \top_I.branch[2].block[12].um_I.ana[7] ;
 wire \top_I.branch[2].block[12].um_I.clk ;
 wire \top_I.branch[2].block[12].um_I.ena ;
 wire \top_I.branch[2].block[12].um_I.iw[10] ;
 wire \top_I.branch[2].block[12].um_I.iw[11] ;
 wire \top_I.branch[2].block[12].um_I.iw[12] ;
 wire \top_I.branch[2].block[12].um_I.iw[13] ;
 wire \top_I.branch[2].block[12].um_I.iw[14] ;
 wire \top_I.branch[2].block[12].um_I.iw[15] ;
 wire \top_I.branch[2].block[12].um_I.iw[16] ;
 wire \top_I.branch[2].block[12].um_I.iw[17] ;
 wire \top_I.branch[2].block[12].um_I.iw[1] ;
 wire \top_I.branch[2].block[12].um_I.iw[2] ;
 wire \top_I.branch[2].block[12].um_I.iw[3] ;
 wire \top_I.branch[2].block[12].um_I.iw[4] ;
 wire \top_I.branch[2].block[12].um_I.iw[5] ;
 wire \top_I.branch[2].block[12].um_I.iw[6] ;
 wire \top_I.branch[2].block[12].um_I.iw[7] ;
 wire \top_I.branch[2].block[12].um_I.iw[8] ;
 wire \top_I.branch[2].block[12].um_I.iw[9] ;
 wire \top_I.branch[2].block[12].um_I.k_zero ;
 wire \top_I.branch[2].block[12].um_I.pg_vdd ;
 wire \top_I.branch[2].block[13].um_I.ana[2] ;
 wire \top_I.branch[2].block[13].um_I.ana[3] ;
 wire \top_I.branch[2].block[13].um_I.ana[4] ;
 wire \top_I.branch[2].block[13].um_I.ana[5] ;
 wire \top_I.branch[2].block[13].um_I.ana[6] ;
 wire \top_I.branch[2].block[13].um_I.ana[7] ;
 wire \top_I.branch[2].block[13].um_I.clk ;
 wire \top_I.branch[2].block[13].um_I.ena ;
 wire \top_I.branch[2].block[13].um_I.iw[10] ;
 wire \top_I.branch[2].block[13].um_I.iw[11] ;
 wire \top_I.branch[2].block[13].um_I.iw[12] ;
 wire \top_I.branch[2].block[13].um_I.iw[13] ;
 wire \top_I.branch[2].block[13].um_I.iw[14] ;
 wire \top_I.branch[2].block[13].um_I.iw[15] ;
 wire \top_I.branch[2].block[13].um_I.iw[16] ;
 wire \top_I.branch[2].block[13].um_I.iw[17] ;
 wire \top_I.branch[2].block[13].um_I.iw[1] ;
 wire \top_I.branch[2].block[13].um_I.iw[2] ;
 wire \top_I.branch[2].block[13].um_I.iw[3] ;
 wire \top_I.branch[2].block[13].um_I.iw[4] ;
 wire \top_I.branch[2].block[13].um_I.iw[5] ;
 wire \top_I.branch[2].block[13].um_I.iw[6] ;
 wire \top_I.branch[2].block[13].um_I.iw[7] ;
 wire \top_I.branch[2].block[13].um_I.iw[8] ;
 wire \top_I.branch[2].block[13].um_I.iw[9] ;
 wire \top_I.branch[2].block[13].um_I.k_zero ;
 wire \top_I.branch[2].block[13].um_I.pg_vdd ;
 wire \top_I.branch[2].block[14].um_I.ana[2] ;
 wire \top_I.branch[2].block[14].um_I.ana[3] ;
 wire \top_I.branch[2].block[14].um_I.ana[4] ;
 wire \top_I.branch[2].block[14].um_I.ana[5] ;
 wire \top_I.branch[2].block[14].um_I.ana[6] ;
 wire \top_I.branch[2].block[14].um_I.ana[7] ;
 wire \top_I.branch[2].block[14].um_I.clk ;
 wire \top_I.branch[2].block[14].um_I.ena ;
 wire \top_I.branch[2].block[14].um_I.iw[10] ;
 wire \top_I.branch[2].block[14].um_I.iw[11] ;
 wire \top_I.branch[2].block[14].um_I.iw[12] ;
 wire \top_I.branch[2].block[14].um_I.iw[13] ;
 wire \top_I.branch[2].block[14].um_I.iw[14] ;
 wire \top_I.branch[2].block[14].um_I.iw[15] ;
 wire \top_I.branch[2].block[14].um_I.iw[16] ;
 wire \top_I.branch[2].block[14].um_I.iw[17] ;
 wire \top_I.branch[2].block[14].um_I.iw[1] ;
 wire \top_I.branch[2].block[14].um_I.iw[2] ;
 wire \top_I.branch[2].block[14].um_I.iw[3] ;
 wire \top_I.branch[2].block[14].um_I.iw[4] ;
 wire \top_I.branch[2].block[14].um_I.iw[5] ;
 wire \top_I.branch[2].block[14].um_I.iw[6] ;
 wire \top_I.branch[2].block[14].um_I.iw[7] ;
 wire \top_I.branch[2].block[14].um_I.iw[8] ;
 wire \top_I.branch[2].block[14].um_I.iw[9] ;
 wire \top_I.branch[2].block[14].um_I.k_zero ;
 wire \top_I.branch[2].block[14].um_I.pg_vdd ;
 wire \top_I.branch[2].block[15].um_I.ana[2] ;
 wire \top_I.branch[2].block[15].um_I.ana[3] ;
 wire \top_I.branch[2].block[15].um_I.ana[4] ;
 wire \top_I.branch[2].block[15].um_I.ana[5] ;
 wire \top_I.branch[2].block[15].um_I.ana[6] ;
 wire \top_I.branch[2].block[15].um_I.ana[7] ;
 wire \top_I.branch[2].block[15].um_I.clk ;
 wire \top_I.branch[2].block[15].um_I.ena ;
 wire \top_I.branch[2].block[15].um_I.iw[10] ;
 wire \top_I.branch[2].block[15].um_I.iw[11] ;
 wire \top_I.branch[2].block[15].um_I.iw[12] ;
 wire \top_I.branch[2].block[15].um_I.iw[13] ;
 wire \top_I.branch[2].block[15].um_I.iw[14] ;
 wire \top_I.branch[2].block[15].um_I.iw[15] ;
 wire \top_I.branch[2].block[15].um_I.iw[16] ;
 wire \top_I.branch[2].block[15].um_I.iw[17] ;
 wire \top_I.branch[2].block[15].um_I.iw[1] ;
 wire \top_I.branch[2].block[15].um_I.iw[2] ;
 wire \top_I.branch[2].block[15].um_I.iw[3] ;
 wire \top_I.branch[2].block[15].um_I.iw[4] ;
 wire \top_I.branch[2].block[15].um_I.iw[5] ;
 wire \top_I.branch[2].block[15].um_I.iw[6] ;
 wire \top_I.branch[2].block[15].um_I.iw[7] ;
 wire \top_I.branch[2].block[15].um_I.iw[8] ;
 wire \top_I.branch[2].block[15].um_I.iw[9] ;
 wire \top_I.branch[2].block[15].um_I.k_zero ;
 wire \top_I.branch[2].block[15].um_I.pg_vdd ;
 wire \top_I.branch[2].block[1].um_I.ana[2] ;
 wire \top_I.branch[2].block[1].um_I.ana[3] ;
 wire \top_I.branch[2].block[1].um_I.ana[4] ;
 wire \top_I.branch[2].block[1].um_I.ana[5] ;
 wire \top_I.branch[2].block[1].um_I.ana[6] ;
 wire \top_I.branch[2].block[1].um_I.ana[7] ;
 wire \top_I.branch[2].block[1].um_I.clk ;
 wire \top_I.branch[2].block[1].um_I.ena ;
 wire \top_I.branch[2].block[1].um_I.iw[10] ;
 wire \top_I.branch[2].block[1].um_I.iw[11] ;
 wire \top_I.branch[2].block[1].um_I.iw[12] ;
 wire \top_I.branch[2].block[1].um_I.iw[13] ;
 wire \top_I.branch[2].block[1].um_I.iw[14] ;
 wire \top_I.branch[2].block[1].um_I.iw[15] ;
 wire \top_I.branch[2].block[1].um_I.iw[16] ;
 wire \top_I.branch[2].block[1].um_I.iw[17] ;
 wire \top_I.branch[2].block[1].um_I.iw[1] ;
 wire \top_I.branch[2].block[1].um_I.iw[2] ;
 wire \top_I.branch[2].block[1].um_I.iw[3] ;
 wire \top_I.branch[2].block[1].um_I.iw[4] ;
 wire \top_I.branch[2].block[1].um_I.iw[5] ;
 wire \top_I.branch[2].block[1].um_I.iw[6] ;
 wire \top_I.branch[2].block[1].um_I.iw[7] ;
 wire \top_I.branch[2].block[1].um_I.iw[8] ;
 wire \top_I.branch[2].block[1].um_I.iw[9] ;
 wire \top_I.branch[2].block[1].um_I.k_zero ;
 wire \top_I.branch[2].block[1].um_I.pg_vdd ;
 wire \top_I.branch[2].block[2].um_I.ana[2] ;
 wire \top_I.branch[2].block[2].um_I.ana[3] ;
 wire \top_I.branch[2].block[2].um_I.ana[4] ;
 wire \top_I.branch[2].block[2].um_I.ana[5] ;
 wire \top_I.branch[2].block[2].um_I.ana[6] ;
 wire \top_I.branch[2].block[2].um_I.ana[7] ;
 wire \top_I.branch[2].block[2].um_I.clk ;
 wire \top_I.branch[2].block[2].um_I.ena ;
 wire \top_I.branch[2].block[2].um_I.iw[10] ;
 wire \top_I.branch[2].block[2].um_I.iw[11] ;
 wire \top_I.branch[2].block[2].um_I.iw[12] ;
 wire \top_I.branch[2].block[2].um_I.iw[13] ;
 wire \top_I.branch[2].block[2].um_I.iw[14] ;
 wire \top_I.branch[2].block[2].um_I.iw[15] ;
 wire \top_I.branch[2].block[2].um_I.iw[16] ;
 wire \top_I.branch[2].block[2].um_I.iw[17] ;
 wire \top_I.branch[2].block[2].um_I.iw[1] ;
 wire \top_I.branch[2].block[2].um_I.iw[2] ;
 wire \top_I.branch[2].block[2].um_I.iw[3] ;
 wire \top_I.branch[2].block[2].um_I.iw[4] ;
 wire \top_I.branch[2].block[2].um_I.iw[5] ;
 wire \top_I.branch[2].block[2].um_I.iw[6] ;
 wire \top_I.branch[2].block[2].um_I.iw[7] ;
 wire \top_I.branch[2].block[2].um_I.iw[8] ;
 wire \top_I.branch[2].block[2].um_I.iw[9] ;
 wire \top_I.branch[2].block[2].um_I.k_zero ;
 wire \top_I.branch[2].block[2].um_I.pg_vdd ;
 wire \top_I.branch[2].block[3].um_I.ana[2] ;
 wire \top_I.branch[2].block[3].um_I.ana[3] ;
 wire \top_I.branch[2].block[3].um_I.ana[4] ;
 wire \top_I.branch[2].block[3].um_I.ana[5] ;
 wire \top_I.branch[2].block[3].um_I.ana[6] ;
 wire \top_I.branch[2].block[3].um_I.ana[7] ;
 wire \top_I.branch[2].block[3].um_I.clk ;
 wire \top_I.branch[2].block[3].um_I.ena ;
 wire \top_I.branch[2].block[3].um_I.iw[10] ;
 wire \top_I.branch[2].block[3].um_I.iw[11] ;
 wire \top_I.branch[2].block[3].um_I.iw[12] ;
 wire \top_I.branch[2].block[3].um_I.iw[13] ;
 wire \top_I.branch[2].block[3].um_I.iw[14] ;
 wire \top_I.branch[2].block[3].um_I.iw[15] ;
 wire \top_I.branch[2].block[3].um_I.iw[16] ;
 wire \top_I.branch[2].block[3].um_I.iw[17] ;
 wire \top_I.branch[2].block[3].um_I.iw[1] ;
 wire \top_I.branch[2].block[3].um_I.iw[2] ;
 wire \top_I.branch[2].block[3].um_I.iw[3] ;
 wire \top_I.branch[2].block[3].um_I.iw[4] ;
 wire \top_I.branch[2].block[3].um_I.iw[5] ;
 wire \top_I.branch[2].block[3].um_I.iw[6] ;
 wire \top_I.branch[2].block[3].um_I.iw[7] ;
 wire \top_I.branch[2].block[3].um_I.iw[8] ;
 wire \top_I.branch[2].block[3].um_I.iw[9] ;
 wire \top_I.branch[2].block[3].um_I.k_zero ;
 wire \top_I.branch[2].block[3].um_I.pg_vdd ;
 wire \top_I.branch[2].block[4].um_I.ana[2] ;
 wire \top_I.branch[2].block[4].um_I.ana[3] ;
 wire \top_I.branch[2].block[4].um_I.ana[4] ;
 wire \top_I.branch[2].block[4].um_I.ana[5] ;
 wire \top_I.branch[2].block[4].um_I.ana[6] ;
 wire \top_I.branch[2].block[4].um_I.ana[7] ;
 wire \top_I.branch[2].block[4].um_I.clk ;
 wire \top_I.branch[2].block[4].um_I.ena ;
 wire \top_I.branch[2].block[4].um_I.iw[10] ;
 wire \top_I.branch[2].block[4].um_I.iw[11] ;
 wire \top_I.branch[2].block[4].um_I.iw[12] ;
 wire \top_I.branch[2].block[4].um_I.iw[13] ;
 wire \top_I.branch[2].block[4].um_I.iw[14] ;
 wire \top_I.branch[2].block[4].um_I.iw[15] ;
 wire \top_I.branch[2].block[4].um_I.iw[16] ;
 wire \top_I.branch[2].block[4].um_I.iw[17] ;
 wire \top_I.branch[2].block[4].um_I.iw[1] ;
 wire \top_I.branch[2].block[4].um_I.iw[2] ;
 wire \top_I.branch[2].block[4].um_I.iw[3] ;
 wire \top_I.branch[2].block[4].um_I.iw[4] ;
 wire \top_I.branch[2].block[4].um_I.iw[5] ;
 wire \top_I.branch[2].block[4].um_I.iw[6] ;
 wire \top_I.branch[2].block[4].um_I.iw[7] ;
 wire \top_I.branch[2].block[4].um_I.iw[8] ;
 wire \top_I.branch[2].block[4].um_I.iw[9] ;
 wire \top_I.branch[2].block[4].um_I.k_zero ;
 wire \top_I.branch[2].block[4].um_I.pg_vdd ;
 wire \top_I.branch[2].block[5].um_I.ana[2] ;
 wire \top_I.branch[2].block[5].um_I.ana[3] ;
 wire \top_I.branch[2].block[5].um_I.ana[4] ;
 wire \top_I.branch[2].block[5].um_I.ana[5] ;
 wire \top_I.branch[2].block[5].um_I.ana[6] ;
 wire \top_I.branch[2].block[5].um_I.ana[7] ;
 wire \top_I.branch[2].block[5].um_I.clk ;
 wire \top_I.branch[2].block[5].um_I.ena ;
 wire \top_I.branch[2].block[5].um_I.iw[10] ;
 wire \top_I.branch[2].block[5].um_I.iw[11] ;
 wire \top_I.branch[2].block[5].um_I.iw[12] ;
 wire \top_I.branch[2].block[5].um_I.iw[13] ;
 wire \top_I.branch[2].block[5].um_I.iw[14] ;
 wire \top_I.branch[2].block[5].um_I.iw[15] ;
 wire \top_I.branch[2].block[5].um_I.iw[16] ;
 wire \top_I.branch[2].block[5].um_I.iw[17] ;
 wire \top_I.branch[2].block[5].um_I.iw[1] ;
 wire \top_I.branch[2].block[5].um_I.iw[2] ;
 wire \top_I.branch[2].block[5].um_I.iw[3] ;
 wire \top_I.branch[2].block[5].um_I.iw[4] ;
 wire \top_I.branch[2].block[5].um_I.iw[5] ;
 wire \top_I.branch[2].block[5].um_I.iw[6] ;
 wire \top_I.branch[2].block[5].um_I.iw[7] ;
 wire \top_I.branch[2].block[5].um_I.iw[8] ;
 wire \top_I.branch[2].block[5].um_I.iw[9] ;
 wire \top_I.branch[2].block[5].um_I.k_zero ;
 wire \top_I.branch[2].block[5].um_I.pg_vdd ;
 wire \top_I.branch[2].block[6].um_I.ana[2] ;
 wire \top_I.branch[2].block[6].um_I.ana[3] ;
 wire \top_I.branch[2].block[6].um_I.ana[4] ;
 wire \top_I.branch[2].block[6].um_I.ana[5] ;
 wire \top_I.branch[2].block[6].um_I.ana[6] ;
 wire \top_I.branch[2].block[6].um_I.ana[7] ;
 wire \top_I.branch[2].block[6].um_I.clk ;
 wire \top_I.branch[2].block[6].um_I.ena ;
 wire \top_I.branch[2].block[6].um_I.iw[10] ;
 wire \top_I.branch[2].block[6].um_I.iw[11] ;
 wire \top_I.branch[2].block[6].um_I.iw[12] ;
 wire \top_I.branch[2].block[6].um_I.iw[13] ;
 wire \top_I.branch[2].block[6].um_I.iw[14] ;
 wire \top_I.branch[2].block[6].um_I.iw[15] ;
 wire \top_I.branch[2].block[6].um_I.iw[16] ;
 wire \top_I.branch[2].block[6].um_I.iw[17] ;
 wire \top_I.branch[2].block[6].um_I.iw[1] ;
 wire \top_I.branch[2].block[6].um_I.iw[2] ;
 wire \top_I.branch[2].block[6].um_I.iw[3] ;
 wire \top_I.branch[2].block[6].um_I.iw[4] ;
 wire \top_I.branch[2].block[6].um_I.iw[5] ;
 wire \top_I.branch[2].block[6].um_I.iw[6] ;
 wire \top_I.branch[2].block[6].um_I.iw[7] ;
 wire \top_I.branch[2].block[6].um_I.iw[8] ;
 wire \top_I.branch[2].block[6].um_I.iw[9] ;
 wire \top_I.branch[2].block[6].um_I.k_zero ;
 wire \top_I.branch[2].block[6].um_I.pg_vdd ;
 wire \top_I.branch[2].block[7].um_I.ana[2] ;
 wire \top_I.branch[2].block[7].um_I.ana[3] ;
 wire \top_I.branch[2].block[7].um_I.ana[4] ;
 wire \top_I.branch[2].block[7].um_I.ana[5] ;
 wire \top_I.branch[2].block[7].um_I.ana[6] ;
 wire \top_I.branch[2].block[7].um_I.ana[7] ;
 wire \top_I.branch[2].block[7].um_I.clk ;
 wire \top_I.branch[2].block[7].um_I.ena ;
 wire \top_I.branch[2].block[7].um_I.iw[10] ;
 wire \top_I.branch[2].block[7].um_I.iw[11] ;
 wire \top_I.branch[2].block[7].um_I.iw[12] ;
 wire \top_I.branch[2].block[7].um_I.iw[13] ;
 wire \top_I.branch[2].block[7].um_I.iw[14] ;
 wire \top_I.branch[2].block[7].um_I.iw[15] ;
 wire \top_I.branch[2].block[7].um_I.iw[16] ;
 wire \top_I.branch[2].block[7].um_I.iw[17] ;
 wire \top_I.branch[2].block[7].um_I.iw[1] ;
 wire \top_I.branch[2].block[7].um_I.iw[2] ;
 wire \top_I.branch[2].block[7].um_I.iw[3] ;
 wire \top_I.branch[2].block[7].um_I.iw[4] ;
 wire \top_I.branch[2].block[7].um_I.iw[5] ;
 wire \top_I.branch[2].block[7].um_I.iw[6] ;
 wire \top_I.branch[2].block[7].um_I.iw[7] ;
 wire \top_I.branch[2].block[7].um_I.iw[8] ;
 wire \top_I.branch[2].block[7].um_I.iw[9] ;
 wire \top_I.branch[2].block[7].um_I.k_zero ;
 wire \top_I.branch[2].block[7].um_I.pg_vdd ;
 wire \top_I.branch[2].block[8].um_I.ana[2] ;
 wire \top_I.branch[2].block[8].um_I.ana[3] ;
 wire \top_I.branch[2].block[8].um_I.ana[4] ;
 wire \top_I.branch[2].block[8].um_I.ana[5] ;
 wire \top_I.branch[2].block[8].um_I.ana[6] ;
 wire \top_I.branch[2].block[8].um_I.ana[7] ;
 wire \top_I.branch[2].block[8].um_I.clk ;
 wire \top_I.branch[2].block[8].um_I.ena ;
 wire \top_I.branch[2].block[8].um_I.iw[10] ;
 wire \top_I.branch[2].block[8].um_I.iw[11] ;
 wire \top_I.branch[2].block[8].um_I.iw[12] ;
 wire \top_I.branch[2].block[8].um_I.iw[13] ;
 wire \top_I.branch[2].block[8].um_I.iw[14] ;
 wire \top_I.branch[2].block[8].um_I.iw[15] ;
 wire \top_I.branch[2].block[8].um_I.iw[16] ;
 wire \top_I.branch[2].block[8].um_I.iw[17] ;
 wire \top_I.branch[2].block[8].um_I.iw[1] ;
 wire \top_I.branch[2].block[8].um_I.iw[2] ;
 wire \top_I.branch[2].block[8].um_I.iw[3] ;
 wire \top_I.branch[2].block[8].um_I.iw[4] ;
 wire \top_I.branch[2].block[8].um_I.iw[5] ;
 wire \top_I.branch[2].block[8].um_I.iw[6] ;
 wire \top_I.branch[2].block[8].um_I.iw[7] ;
 wire \top_I.branch[2].block[8].um_I.iw[8] ;
 wire \top_I.branch[2].block[8].um_I.iw[9] ;
 wire \top_I.branch[2].block[8].um_I.k_zero ;
 wire \top_I.branch[2].block[8].um_I.pg_vdd ;
 wire \top_I.branch[2].block[9].um_I.ana[2] ;
 wire \top_I.branch[2].block[9].um_I.ana[3] ;
 wire \top_I.branch[2].block[9].um_I.ana[4] ;
 wire \top_I.branch[2].block[9].um_I.ana[5] ;
 wire \top_I.branch[2].block[9].um_I.ana[6] ;
 wire \top_I.branch[2].block[9].um_I.ana[7] ;
 wire \top_I.branch[2].block[9].um_I.clk ;
 wire \top_I.branch[2].block[9].um_I.ena ;
 wire \top_I.branch[2].block[9].um_I.iw[10] ;
 wire \top_I.branch[2].block[9].um_I.iw[11] ;
 wire \top_I.branch[2].block[9].um_I.iw[12] ;
 wire \top_I.branch[2].block[9].um_I.iw[13] ;
 wire \top_I.branch[2].block[9].um_I.iw[14] ;
 wire \top_I.branch[2].block[9].um_I.iw[15] ;
 wire \top_I.branch[2].block[9].um_I.iw[16] ;
 wire \top_I.branch[2].block[9].um_I.iw[17] ;
 wire \top_I.branch[2].block[9].um_I.iw[1] ;
 wire \top_I.branch[2].block[9].um_I.iw[2] ;
 wire \top_I.branch[2].block[9].um_I.iw[3] ;
 wire \top_I.branch[2].block[9].um_I.iw[4] ;
 wire \top_I.branch[2].block[9].um_I.iw[5] ;
 wire \top_I.branch[2].block[9].um_I.iw[6] ;
 wire \top_I.branch[2].block[9].um_I.iw[7] ;
 wire \top_I.branch[2].block[9].um_I.iw[8] ;
 wire \top_I.branch[2].block[9].um_I.iw[9] ;
 wire \top_I.branch[2].block[9].um_I.k_zero ;
 wire \top_I.branch[2].block[9].um_I.pg_vdd ;
 wire \top_I.branch[2].l_addr[0] ;
 wire \top_I.branch[2].l_addr[1] ;
 wire \top_I.branch[3].block[0].um_I.ana[2] ;
 wire \top_I.branch[3].block[0].um_I.ana[3] ;
 wire \top_I.branch[3].block[0].um_I.ana[4] ;
 wire \top_I.branch[3].block[0].um_I.ana[5] ;
 wire \top_I.branch[3].block[0].um_I.ana[6] ;
 wire \top_I.branch[3].block[0].um_I.ana[7] ;
 wire \top_I.branch[3].block[0].um_I.clk ;
 wire \top_I.branch[3].block[0].um_I.ena ;
 wire \top_I.branch[3].block[0].um_I.iw[10] ;
 wire \top_I.branch[3].block[0].um_I.iw[11] ;
 wire \top_I.branch[3].block[0].um_I.iw[12] ;
 wire \top_I.branch[3].block[0].um_I.iw[13] ;
 wire \top_I.branch[3].block[0].um_I.iw[14] ;
 wire \top_I.branch[3].block[0].um_I.iw[15] ;
 wire \top_I.branch[3].block[0].um_I.iw[16] ;
 wire \top_I.branch[3].block[0].um_I.iw[17] ;
 wire \top_I.branch[3].block[0].um_I.iw[1] ;
 wire \top_I.branch[3].block[0].um_I.iw[2] ;
 wire \top_I.branch[3].block[0].um_I.iw[3] ;
 wire \top_I.branch[3].block[0].um_I.iw[4] ;
 wire \top_I.branch[3].block[0].um_I.iw[5] ;
 wire \top_I.branch[3].block[0].um_I.iw[6] ;
 wire \top_I.branch[3].block[0].um_I.iw[7] ;
 wire \top_I.branch[3].block[0].um_I.iw[8] ;
 wire \top_I.branch[3].block[0].um_I.iw[9] ;
 wire \top_I.branch[3].block[0].um_I.k_zero ;
 wire \top_I.branch[3].block[0].um_I.pg_vdd ;
 wire \top_I.branch[3].block[10].um_I.ana[2] ;
 wire \top_I.branch[3].block[10].um_I.ana[3] ;
 wire \top_I.branch[3].block[10].um_I.ana[4] ;
 wire \top_I.branch[3].block[10].um_I.ana[5] ;
 wire \top_I.branch[3].block[10].um_I.ana[6] ;
 wire \top_I.branch[3].block[10].um_I.ana[7] ;
 wire \top_I.branch[3].block[10].um_I.clk ;
 wire \top_I.branch[3].block[10].um_I.ena ;
 wire \top_I.branch[3].block[10].um_I.iw[10] ;
 wire \top_I.branch[3].block[10].um_I.iw[11] ;
 wire \top_I.branch[3].block[10].um_I.iw[12] ;
 wire \top_I.branch[3].block[10].um_I.iw[13] ;
 wire \top_I.branch[3].block[10].um_I.iw[14] ;
 wire \top_I.branch[3].block[10].um_I.iw[15] ;
 wire \top_I.branch[3].block[10].um_I.iw[16] ;
 wire \top_I.branch[3].block[10].um_I.iw[17] ;
 wire \top_I.branch[3].block[10].um_I.iw[1] ;
 wire \top_I.branch[3].block[10].um_I.iw[2] ;
 wire \top_I.branch[3].block[10].um_I.iw[3] ;
 wire \top_I.branch[3].block[10].um_I.iw[4] ;
 wire \top_I.branch[3].block[10].um_I.iw[5] ;
 wire \top_I.branch[3].block[10].um_I.iw[6] ;
 wire \top_I.branch[3].block[10].um_I.iw[7] ;
 wire \top_I.branch[3].block[10].um_I.iw[8] ;
 wire \top_I.branch[3].block[10].um_I.iw[9] ;
 wire \top_I.branch[3].block[10].um_I.k_zero ;
 wire \top_I.branch[3].block[10].um_I.pg_vdd ;
 wire \top_I.branch[3].block[11].um_I.ana[2] ;
 wire \top_I.branch[3].block[11].um_I.ana[3] ;
 wire \top_I.branch[3].block[11].um_I.ana[4] ;
 wire \top_I.branch[3].block[11].um_I.ana[5] ;
 wire \top_I.branch[3].block[11].um_I.ana[6] ;
 wire \top_I.branch[3].block[11].um_I.ana[7] ;
 wire \top_I.branch[3].block[11].um_I.clk ;
 wire \top_I.branch[3].block[11].um_I.ena ;
 wire \top_I.branch[3].block[11].um_I.iw[10] ;
 wire \top_I.branch[3].block[11].um_I.iw[11] ;
 wire \top_I.branch[3].block[11].um_I.iw[12] ;
 wire \top_I.branch[3].block[11].um_I.iw[13] ;
 wire \top_I.branch[3].block[11].um_I.iw[14] ;
 wire \top_I.branch[3].block[11].um_I.iw[15] ;
 wire \top_I.branch[3].block[11].um_I.iw[16] ;
 wire \top_I.branch[3].block[11].um_I.iw[17] ;
 wire \top_I.branch[3].block[11].um_I.iw[1] ;
 wire \top_I.branch[3].block[11].um_I.iw[2] ;
 wire \top_I.branch[3].block[11].um_I.iw[3] ;
 wire \top_I.branch[3].block[11].um_I.iw[4] ;
 wire \top_I.branch[3].block[11].um_I.iw[5] ;
 wire \top_I.branch[3].block[11].um_I.iw[6] ;
 wire \top_I.branch[3].block[11].um_I.iw[7] ;
 wire \top_I.branch[3].block[11].um_I.iw[8] ;
 wire \top_I.branch[3].block[11].um_I.iw[9] ;
 wire \top_I.branch[3].block[11].um_I.k_zero ;
 wire \top_I.branch[3].block[11].um_I.pg_vdd ;
 wire \top_I.branch[3].block[12].um_I.ana[2] ;
 wire \top_I.branch[3].block[12].um_I.ana[3] ;
 wire \top_I.branch[3].block[12].um_I.ana[4] ;
 wire \top_I.branch[3].block[12].um_I.ana[5] ;
 wire \top_I.branch[3].block[12].um_I.ana[6] ;
 wire \top_I.branch[3].block[12].um_I.ana[7] ;
 wire \top_I.branch[3].block[12].um_I.clk ;
 wire \top_I.branch[3].block[12].um_I.ena ;
 wire \top_I.branch[3].block[12].um_I.iw[10] ;
 wire \top_I.branch[3].block[12].um_I.iw[11] ;
 wire \top_I.branch[3].block[12].um_I.iw[12] ;
 wire \top_I.branch[3].block[12].um_I.iw[13] ;
 wire \top_I.branch[3].block[12].um_I.iw[14] ;
 wire \top_I.branch[3].block[12].um_I.iw[15] ;
 wire \top_I.branch[3].block[12].um_I.iw[16] ;
 wire \top_I.branch[3].block[12].um_I.iw[17] ;
 wire \top_I.branch[3].block[12].um_I.iw[1] ;
 wire \top_I.branch[3].block[12].um_I.iw[2] ;
 wire \top_I.branch[3].block[12].um_I.iw[3] ;
 wire \top_I.branch[3].block[12].um_I.iw[4] ;
 wire \top_I.branch[3].block[12].um_I.iw[5] ;
 wire \top_I.branch[3].block[12].um_I.iw[6] ;
 wire \top_I.branch[3].block[12].um_I.iw[7] ;
 wire \top_I.branch[3].block[12].um_I.iw[8] ;
 wire \top_I.branch[3].block[12].um_I.iw[9] ;
 wire \top_I.branch[3].block[12].um_I.k_zero ;
 wire \top_I.branch[3].block[12].um_I.pg_vdd ;
 wire \top_I.branch[3].block[13].um_I.ana[2] ;
 wire \top_I.branch[3].block[13].um_I.ana[3] ;
 wire \top_I.branch[3].block[13].um_I.ana[4] ;
 wire \top_I.branch[3].block[13].um_I.ana[5] ;
 wire \top_I.branch[3].block[13].um_I.ana[6] ;
 wire \top_I.branch[3].block[13].um_I.ana[7] ;
 wire \top_I.branch[3].block[13].um_I.clk ;
 wire \top_I.branch[3].block[13].um_I.ena ;
 wire \top_I.branch[3].block[13].um_I.iw[10] ;
 wire \top_I.branch[3].block[13].um_I.iw[11] ;
 wire \top_I.branch[3].block[13].um_I.iw[12] ;
 wire \top_I.branch[3].block[13].um_I.iw[13] ;
 wire \top_I.branch[3].block[13].um_I.iw[14] ;
 wire \top_I.branch[3].block[13].um_I.iw[15] ;
 wire \top_I.branch[3].block[13].um_I.iw[16] ;
 wire \top_I.branch[3].block[13].um_I.iw[17] ;
 wire \top_I.branch[3].block[13].um_I.iw[1] ;
 wire \top_I.branch[3].block[13].um_I.iw[2] ;
 wire \top_I.branch[3].block[13].um_I.iw[3] ;
 wire \top_I.branch[3].block[13].um_I.iw[4] ;
 wire \top_I.branch[3].block[13].um_I.iw[5] ;
 wire \top_I.branch[3].block[13].um_I.iw[6] ;
 wire \top_I.branch[3].block[13].um_I.iw[7] ;
 wire \top_I.branch[3].block[13].um_I.iw[8] ;
 wire \top_I.branch[3].block[13].um_I.iw[9] ;
 wire \top_I.branch[3].block[13].um_I.k_zero ;
 wire \top_I.branch[3].block[13].um_I.pg_vdd ;
 wire \top_I.branch[3].block[14].um_I.ana[2] ;
 wire \top_I.branch[3].block[14].um_I.ana[3] ;
 wire \top_I.branch[3].block[14].um_I.ana[4] ;
 wire \top_I.branch[3].block[14].um_I.ana[5] ;
 wire \top_I.branch[3].block[14].um_I.ana[6] ;
 wire \top_I.branch[3].block[14].um_I.ana[7] ;
 wire \top_I.branch[3].block[14].um_I.clk ;
 wire \top_I.branch[3].block[14].um_I.ena ;
 wire \top_I.branch[3].block[14].um_I.iw[10] ;
 wire \top_I.branch[3].block[14].um_I.iw[11] ;
 wire \top_I.branch[3].block[14].um_I.iw[12] ;
 wire \top_I.branch[3].block[14].um_I.iw[13] ;
 wire \top_I.branch[3].block[14].um_I.iw[14] ;
 wire \top_I.branch[3].block[14].um_I.iw[15] ;
 wire \top_I.branch[3].block[14].um_I.iw[16] ;
 wire \top_I.branch[3].block[14].um_I.iw[17] ;
 wire \top_I.branch[3].block[14].um_I.iw[1] ;
 wire \top_I.branch[3].block[14].um_I.iw[2] ;
 wire \top_I.branch[3].block[14].um_I.iw[3] ;
 wire \top_I.branch[3].block[14].um_I.iw[4] ;
 wire \top_I.branch[3].block[14].um_I.iw[5] ;
 wire \top_I.branch[3].block[14].um_I.iw[6] ;
 wire \top_I.branch[3].block[14].um_I.iw[7] ;
 wire \top_I.branch[3].block[14].um_I.iw[8] ;
 wire \top_I.branch[3].block[14].um_I.iw[9] ;
 wire \top_I.branch[3].block[14].um_I.k_zero ;
 wire \top_I.branch[3].block[14].um_I.pg_vdd ;
 wire \top_I.branch[3].block[15].um_I.ana[2] ;
 wire \top_I.branch[3].block[15].um_I.ana[3] ;
 wire \top_I.branch[3].block[15].um_I.ana[4] ;
 wire \top_I.branch[3].block[15].um_I.ana[5] ;
 wire \top_I.branch[3].block[15].um_I.ana[6] ;
 wire \top_I.branch[3].block[15].um_I.ana[7] ;
 wire \top_I.branch[3].block[15].um_I.clk ;
 wire \top_I.branch[3].block[15].um_I.ena ;
 wire \top_I.branch[3].block[15].um_I.iw[10] ;
 wire \top_I.branch[3].block[15].um_I.iw[11] ;
 wire \top_I.branch[3].block[15].um_I.iw[12] ;
 wire \top_I.branch[3].block[15].um_I.iw[13] ;
 wire \top_I.branch[3].block[15].um_I.iw[14] ;
 wire \top_I.branch[3].block[15].um_I.iw[15] ;
 wire \top_I.branch[3].block[15].um_I.iw[16] ;
 wire \top_I.branch[3].block[15].um_I.iw[17] ;
 wire \top_I.branch[3].block[15].um_I.iw[1] ;
 wire \top_I.branch[3].block[15].um_I.iw[2] ;
 wire \top_I.branch[3].block[15].um_I.iw[3] ;
 wire \top_I.branch[3].block[15].um_I.iw[4] ;
 wire \top_I.branch[3].block[15].um_I.iw[5] ;
 wire \top_I.branch[3].block[15].um_I.iw[6] ;
 wire \top_I.branch[3].block[15].um_I.iw[7] ;
 wire \top_I.branch[3].block[15].um_I.iw[8] ;
 wire \top_I.branch[3].block[15].um_I.iw[9] ;
 wire \top_I.branch[3].block[15].um_I.k_zero ;
 wire \top_I.branch[3].block[15].um_I.pg_vdd ;
 wire \top_I.branch[3].block[1].um_I.ana[2] ;
 wire \top_I.branch[3].block[1].um_I.ana[3] ;
 wire \top_I.branch[3].block[1].um_I.ana[4] ;
 wire \top_I.branch[3].block[1].um_I.ana[5] ;
 wire \top_I.branch[3].block[1].um_I.ana[6] ;
 wire \top_I.branch[3].block[1].um_I.ana[7] ;
 wire \top_I.branch[3].block[1].um_I.clk ;
 wire \top_I.branch[3].block[1].um_I.ena ;
 wire \top_I.branch[3].block[1].um_I.iw[10] ;
 wire \top_I.branch[3].block[1].um_I.iw[11] ;
 wire \top_I.branch[3].block[1].um_I.iw[12] ;
 wire \top_I.branch[3].block[1].um_I.iw[13] ;
 wire \top_I.branch[3].block[1].um_I.iw[14] ;
 wire \top_I.branch[3].block[1].um_I.iw[15] ;
 wire \top_I.branch[3].block[1].um_I.iw[16] ;
 wire \top_I.branch[3].block[1].um_I.iw[17] ;
 wire \top_I.branch[3].block[1].um_I.iw[1] ;
 wire \top_I.branch[3].block[1].um_I.iw[2] ;
 wire \top_I.branch[3].block[1].um_I.iw[3] ;
 wire \top_I.branch[3].block[1].um_I.iw[4] ;
 wire \top_I.branch[3].block[1].um_I.iw[5] ;
 wire \top_I.branch[3].block[1].um_I.iw[6] ;
 wire \top_I.branch[3].block[1].um_I.iw[7] ;
 wire \top_I.branch[3].block[1].um_I.iw[8] ;
 wire \top_I.branch[3].block[1].um_I.iw[9] ;
 wire \top_I.branch[3].block[1].um_I.k_zero ;
 wire \top_I.branch[3].block[1].um_I.pg_vdd ;
 wire \top_I.branch[3].block[2].um_I.ana[2] ;
 wire \top_I.branch[3].block[2].um_I.ana[3] ;
 wire \top_I.branch[3].block[2].um_I.ana[4] ;
 wire \top_I.branch[3].block[2].um_I.ana[5] ;
 wire \top_I.branch[3].block[2].um_I.ana[6] ;
 wire \top_I.branch[3].block[2].um_I.ana[7] ;
 wire \top_I.branch[3].block[2].um_I.clk ;
 wire \top_I.branch[3].block[2].um_I.ena ;
 wire \top_I.branch[3].block[2].um_I.iw[10] ;
 wire \top_I.branch[3].block[2].um_I.iw[11] ;
 wire \top_I.branch[3].block[2].um_I.iw[12] ;
 wire \top_I.branch[3].block[2].um_I.iw[13] ;
 wire \top_I.branch[3].block[2].um_I.iw[14] ;
 wire \top_I.branch[3].block[2].um_I.iw[15] ;
 wire \top_I.branch[3].block[2].um_I.iw[16] ;
 wire \top_I.branch[3].block[2].um_I.iw[17] ;
 wire \top_I.branch[3].block[2].um_I.iw[1] ;
 wire \top_I.branch[3].block[2].um_I.iw[2] ;
 wire \top_I.branch[3].block[2].um_I.iw[3] ;
 wire \top_I.branch[3].block[2].um_I.iw[4] ;
 wire \top_I.branch[3].block[2].um_I.iw[5] ;
 wire \top_I.branch[3].block[2].um_I.iw[6] ;
 wire \top_I.branch[3].block[2].um_I.iw[7] ;
 wire \top_I.branch[3].block[2].um_I.iw[8] ;
 wire \top_I.branch[3].block[2].um_I.iw[9] ;
 wire \top_I.branch[3].block[2].um_I.k_zero ;
 wire \top_I.branch[3].block[2].um_I.pg_vdd ;
 wire \top_I.branch[3].block[3].um_I.ana[2] ;
 wire \top_I.branch[3].block[3].um_I.ana[3] ;
 wire \top_I.branch[3].block[3].um_I.ana[4] ;
 wire \top_I.branch[3].block[3].um_I.ana[5] ;
 wire \top_I.branch[3].block[3].um_I.ana[6] ;
 wire \top_I.branch[3].block[3].um_I.ana[7] ;
 wire \top_I.branch[3].block[3].um_I.clk ;
 wire \top_I.branch[3].block[3].um_I.ena ;
 wire \top_I.branch[3].block[3].um_I.iw[10] ;
 wire \top_I.branch[3].block[3].um_I.iw[11] ;
 wire \top_I.branch[3].block[3].um_I.iw[12] ;
 wire \top_I.branch[3].block[3].um_I.iw[13] ;
 wire \top_I.branch[3].block[3].um_I.iw[14] ;
 wire \top_I.branch[3].block[3].um_I.iw[15] ;
 wire \top_I.branch[3].block[3].um_I.iw[16] ;
 wire \top_I.branch[3].block[3].um_I.iw[17] ;
 wire \top_I.branch[3].block[3].um_I.iw[1] ;
 wire \top_I.branch[3].block[3].um_I.iw[2] ;
 wire \top_I.branch[3].block[3].um_I.iw[3] ;
 wire \top_I.branch[3].block[3].um_I.iw[4] ;
 wire \top_I.branch[3].block[3].um_I.iw[5] ;
 wire \top_I.branch[3].block[3].um_I.iw[6] ;
 wire \top_I.branch[3].block[3].um_I.iw[7] ;
 wire \top_I.branch[3].block[3].um_I.iw[8] ;
 wire \top_I.branch[3].block[3].um_I.iw[9] ;
 wire \top_I.branch[3].block[3].um_I.k_zero ;
 wire \top_I.branch[3].block[3].um_I.pg_vdd ;
 wire \top_I.branch[3].block[4].um_I.ana[2] ;
 wire \top_I.branch[3].block[4].um_I.ana[3] ;
 wire \top_I.branch[3].block[4].um_I.ana[4] ;
 wire \top_I.branch[3].block[4].um_I.ana[5] ;
 wire \top_I.branch[3].block[4].um_I.ana[6] ;
 wire \top_I.branch[3].block[4].um_I.ana[7] ;
 wire \top_I.branch[3].block[4].um_I.clk ;
 wire \top_I.branch[3].block[4].um_I.ena ;
 wire \top_I.branch[3].block[4].um_I.iw[10] ;
 wire \top_I.branch[3].block[4].um_I.iw[11] ;
 wire \top_I.branch[3].block[4].um_I.iw[12] ;
 wire \top_I.branch[3].block[4].um_I.iw[13] ;
 wire \top_I.branch[3].block[4].um_I.iw[14] ;
 wire \top_I.branch[3].block[4].um_I.iw[15] ;
 wire \top_I.branch[3].block[4].um_I.iw[16] ;
 wire \top_I.branch[3].block[4].um_I.iw[17] ;
 wire \top_I.branch[3].block[4].um_I.iw[1] ;
 wire \top_I.branch[3].block[4].um_I.iw[2] ;
 wire \top_I.branch[3].block[4].um_I.iw[3] ;
 wire \top_I.branch[3].block[4].um_I.iw[4] ;
 wire \top_I.branch[3].block[4].um_I.iw[5] ;
 wire \top_I.branch[3].block[4].um_I.iw[6] ;
 wire \top_I.branch[3].block[4].um_I.iw[7] ;
 wire \top_I.branch[3].block[4].um_I.iw[8] ;
 wire \top_I.branch[3].block[4].um_I.iw[9] ;
 wire \top_I.branch[3].block[4].um_I.k_zero ;
 wire \top_I.branch[3].block[4].um_I.pg_vdd ;
 wire \top_I.branch[3].block[5].um_I.ana[2] ;
 wire \top_I.branch[3].block[5].um_I.ana[3] ;
 wire \top_I.branch[3].block[5].um_I.ana[4] ;
 wire \top_I.branch[3].block[5].um_I.ana[5] ;
 wire \top_I.branch[3].block[5].um_I.ana[6] ;
 wire \top_I.branch[3].block[5].um_I.ana[7] ;
 wire \top_I.branch[3].block[5].um_I.clk ;
 wire \top_I.branch[3].block[5].um_I.ena ;
 wire \top_I.branch[3].block[5].um_I.iw[10] ;
 wire \top_I.branch[3].block[5].um_I.iw[11] ;
 wire \top_I.branch[3].block[5].um_I.iw[12] ;
 wire \top_I.branch[3].block[5].um_I.iw[13] ;
 wire \top_I.branch[3].block[5].um_I.iw[14] ;
 wire \top_I.branch[3].block[5].um_I.iw[15] ;
 wire \top_I.branch[3].block[5].um_I.iw[16] ;
 wire \top_I.branch[3].block[5].um_I.iw[17] ;
 wire \top_I.branch[3].block[5].um_I.iw[1] ;
 wire \top_I.branch[3].block[5].um_I.iw[2] ;
 wire \top_I.branch[3].block[5].um_I.iw[3] ;
 wire \top_I.branch[3].block[5].um_I.iw[4] ;
 wire \top_I.branch[3].block[5].um_I.iw[5] ;
 wire \top_I.branch[3].block[5].um_I.iw[6] ;
 wire \top_I.branch[3].block[5].um_I.iw[7] ;
 wire \top_I.branch[3].block[5].um_I.iw[8] ;
 wire \top_I.branch[3].block[5].um_I.iw[9] ;
 wire \top_I.branch[3].block[5].um_I.k_zero ;
 wire \top_I.branch[3].block[5].um_I.pg_vdd ;
 wire \top_I.branch[3].block[6].um_I.ana[2] ;
 wire \top_I.branch[3].block[6].um_I.ana[3] ;
 wire \top_I.branch[3].block[6].um_I.ana[4] ;
 wire \top_I.branch[3].block[6].um_I.ana[5] ;
 wire \top_I.branch[3].block[6].um_I.ana[6] ;
 wire \top_I.branch[3].block[6].um_I.ana[7] ;
 wire \top_I.branch[3].block[6].um_I.clk ;
 wire \top_I.branch[3].block[6].um_I.ena ;
 wire \top_I.branch[3].block[6].um_I.iw[10] ;
 wire \top_I.branch[3].block[6].um_I.iw[11] ;
 wire \top_I.branch[3].block[6].um_I.iw[12] ;
 wire \top_I.branch[3].block[6].um_I.iw[13] ;
 wire \top_I.branch[3].block[6].um_I.iw[14] ;
 wire \top_I.branch[3].block[6].um_I.iw[15] ;
 wire \top_I.branch[3].block[6].um_I.iw[16] ;
 wire \top_I.branch[3].block[6].um_I.iw[17] ;
 wire \top_I.branch[3].block[6].um_I.iw[1] ;
 wire \top_I.branch[3].block[6].um_I.iw[2] ;
 wire \top_I.branch[3].block[6].um_I.iw[3] ;
 wire \top_I.branch[3].block[6].um_I.iw[4] ;
 wire \top_I.branch[3].block[6].um_I.iw[5] ;
 wire \top_I.branch[3].block[6].um_I.iw[6] ;
 wire \top_I.branch[3].block[6].um_I.iw[7] ;
 wire \top_I.branch[3].block[6].um_I.iw[8] ;
 wire \top_I.branch[3].block[6].um_I.iw[9] ;
 wire \top_I.branch[3].block[6].um_I.k_zero ;
 wire \top_I.branch[3].block[6].um_I.pg_vdd ;
 wire \top_I.branch[3].block[7].um_I.ana[2] ;
 wire \top_I.branch[3].block[7].um_I.ana[3] ;
 wire \top_I.branch[3].block[7].um_I.ana[4] ;
 wire \top_I.branch[3].block[7].um_I.ana[5] ;
 wire \top_I.branch[3].block[7].um_I.ana[6] ;
 wire \top_I.branch[3].block[7].um_I.ana[7] ;
 wire \top_I.branch[3].block[7].um_I.clk ;
 wire \top_I.branch[3].block[7].um_I.ena ;
 wire \top_I.branch[3].block[7].um_I.iw[10] ;
 wire \top_I.branch[3].block[7].um_I.iw[11] ;
 wire \top_I.branch[3].block[7].um_I.iw[12] ;
 wire \top_I.branch[3].block[7].um_I.iw[13] ;
 wire \top_I.branch[3].block[7].um_I.iw[14] ;
 wire \top_I.branch[3].block[7].um_I.iw[15] ;
 wire \top_I.branch[3].block[7].um_I.iw[16] ;
 wire \top_I.branch[3].block[7].um_I.iw[17] ;
 wire \top_I.branch[3].block[7].um_I.iw[1] ;
 wire \top_I.branch[3].block[7].um_I.iw[2] ;
 wire \top_I.branch[3].block[7].um_I.iw[3] ;
 wire \top_I.branch[3].block[7].um_I.iw[4] ;
 wire \top_I.branch[3].block[7].um_I.iw[5] ;
 wire \top_I.branch[3].block[7].um_I.iw[6] ;
 wire \top_I.branch[3].block[7].um_I.iw[7] ;
 wire \top_I.branch[3].block[7].um_I.iw[8] ;
 wire \top_I.branch[3].block[7].um_I.iw[9] ;
 wire \top_I.branch[3].block[7].um_I.k_zero ;
 wire \top_I.branch[3].block[7].um_I.pg_vdd ;
 wire \top_I.branch[3].block[8].um_I.ana[2] ;
 wire \top_I.branch[3].block[8].um_I.ana[3] ;
 wire \top_I.branch[3].block[8].um_I.ana[4] ;
 wire \top_I.branch[3].block[8].um_I.ana[5] ;
 wire \top_I.branch[3].block[8].um_I.ana[6] ;
 wire \top_I.branch[3].block[8].um_I.ana[7] ;
 wire \top_I.branch[3].block[8].um_I.clk ;
 wire \top_I.branch[3].block[8].um_I.ena ;
 wire \top_I.branch[3].block[8].um_I.iw[10] ;
 wire \top_I.branch[3].block[8].um_I.iw[11] ;
 wire \top_I.branch[3].block[8].um_I.iw[12] ;
 wire \top_I.branch[3].block[8].um_I.iw[13] ;
 wire \top_I.branch[3].block[8].um_I.iw[14] ;
 wire \top_I.branch[3].block[8].um_I.iw[15] ;
 wire \top_I.branch[3].block[8].um_I.iw[16] ;
 wire \top_I.branch[3].block[8].um_I.iw[17] ;
 wire \top_I.branch[3].block[8].um_I.iw[1] ;
 wire \top_I.branch[3].block[8].um_I.iw[2] ;
 wire \top_I.branch[3].block[8].um_I.iw[3] ;
 wire \top_I.branch[3].block[8].um_I.iw[4] ;
 wire \top_I.branch[3].block[8].um_I.iw[5] ;
 wire \top_I.branch[3].block[8].um_I.iw[6] ;
 wire \top_I.branch[3].block[8].um_I.iw[7] ;
 wire \top_I.branch[3].block[8].um_I.iw[8] ;
 wire \top_I.branch[3].block[8].um_I.iw[9] ;
 wire \top_I.branch[3].block[8].um_I.k_zero ;
 wire \top_I.branch[3].block[8].um_I.pg_vdd ;
 wire \top_I.branch[3].block[9].um_I.ana[2] ;
 wire \top_I.branch[3].block[9].um_I.ana[3] ;
 wire \top_I.branch[3].block[9].um_I.ana[4] ;
 wire \top_I.branch[3].block[9].um_I.ana[5] ;
 wire \top_I.branch[3].block[9].um_I.ana[6] ;
 wire \top_I.branch[3].block[9].um_I.ana[7] ;
 wire \top_I.branch[3].block[9].um_I.clk ;
 wire \top_I.branch[3].block[9].um_I.ena ;
 wire \top_I.branch[3].block[9].um_I.iw[10] ;
 wire \top_I.branch[3].block[9].um_I.iw[11] ;
 wire \top_I.branch[3].block[9].um_I.iw[12] ;
 wire \top_I.branch[3].block[9].um_I.iw[13] ;
 wire \top_I.branch[3].block[9].um_I.iw[14] ;
 wire \top_I.branch[3].block[9].um_I.iw[15] ;
 wire \top_I.branch[3].block[9].um_I.iw[16] ;
 wire \top_I.branch[3].block[9].um_I.iw[17] ;
 wire \top_I.branch[3].block[9].um_I.iw[1] ;
 wire \top_I.branch[3].block[9].um_I.iw[2] ;
 wire \top_I.branch[3].block[9].um_I.iw[3] ;
 wire \top_I.branch[3].block[9].um_I.iw[4] ;
 wire \top_I.branch[3].block[9].um_I.iw[5] ;
 wire \top_I.branch[3].block[9].um_I.iw[6] ;
 wire \top_I.branch[3].block[9].um_I.iw[7] ;
 wire \top_I.branch[3].block[9].um_I.iw[8] ;
 wire \top_I.branch[3].block[9].um_I.iw[9] ;
 wire \top_I.branch[3].block[9].um_I.k_zero ;
 wire \top_I.branch[3].block[9].um_I.pg_vdd ;
 wire \top_I.branch[3].l_addr[0] ;
 wire \top_I.branch[3].l_addr[1] ;
 wire \top_I.branch[4].block[0].um_I.ana[2] ;
 wire \top_I.branch[4].block[0].um_I.ana[3] ;
 wire \top_I.branch[4].block[0].um_I.ana[4] ;
 wire \top_I.branch[4].block[0].um_I.ana[5] ;
 wire \top_I.branch[4].block[0].um_I.ana[6] ;
 wire \top_I.branch[4].block[0].um_I.ana[7] ;
 wire \top_I.branch[4].block[0].um_I.clk ;
 wire \top_I.branch[4].block[0].um_I.ena ;
 wire \top_I.branch[4].block[0].um_I.iw[10] ;
 wire \top_I.branch[4].block[0].um_I.iw[11] ;
 wire \top_I.branch[4].block[0].um_I.iw[12] ;
 wire \top_I.branch[4].block[0].um_I.iw[13] ;
 wire \top_I.branch[4].block[0].um_I.iw[14] ;
 wire \top_I.branch[4].block[0].um_I.iw[15] ;
 wire \top_I.branch[4].block[0].um_I.iw[16] ;
 wire \top_I.branch[4].block[0].um_I.iw[17] ;
 wire \top_I.branch[4].block[0].um_I.iw[1] ;
 wire \top_I.branch[4].block[0].um_I.iw[2] ;
 wire \top_I.branch[4].block[0].um_I.iw[3] ;
 wire \top_I.branch[4].block[0].um_I.iw[4] ;
 wire \top_I.branch[4].block[0].um_I.iw[5] ;
 wire \top_I.branch[4].block[0].um_I.iw[6] ;
 wire \top_I.branch[4].block[0].um_I.iw[7] ;
 wire \top_I.branch[4].block[0].um_I.iw[8] ;
 wire \top_I.branch[4].block[0].um_I.iw[9] ;
 wire \top_I.branch[4].block[0].um_I.k_zero ;
 wire \top_I.branch[4].block[0].um_I.pg_vdd ;
 wire \top_I.branch[4].block[10].um_I.ana[2] ;
 wire \top_I.branch[4].block[10].um_I.ana[3] ;
 wire \top_I.branch[4].block[10].um_I.ana[4] ;
 wire \top_I.branch[4].block[10].um_I.ana[5] ;
 wire \top_I.branch[4].block[10].um_I.ana[6] ;
 wire \top_I.branch[4].block[10].um_I.ana[7] ;
 wire \top_I.branch[4].block[10].um_I.clk ;
 wire \top_I.branch[4].block[10].um_I.ena ;
 wire \top_I.branch[4].block[10].um_I.iw[10] ;
 wire \top_I.branch[4].block[10].um_I.iw[11] ;
 wire \top_I.branch[4].block[10].um_I.iw[12] ;
 wire \top_I.branch[4].block[10].um_I.iw[13] ;
 wire \top_I.branch[4].block[10].um_I.iw[14] ;
 wire \top_I.branch[4].block[10].um_I.iw[15] ;
 wire \top_I.branch[4].block[10].um_I.iw[16] ;
 wire \top_I.branch[4].block[10].um_I.iw[17] ;
 wire \top_I.branch[4].block[10].um_I.iw[1] ;
 wire \top_I.branch[4].block[10].um_I.iw[2] ;
 wire \top_I.branch[4].block[10].um_I.iw[3] ;
 wire \top_I.branch[4].block[10].um_I.iw[4] ;
 wire \top_I.branch[4].block[10].um_I.iw[5] ;
 wire \top_I.branch[4].block[10].um_I.iw[6] ;
 wire \top_I.branch[4].block[10].um_I.iw[7] ;
 wire \top_I.branch[4].block[10].um_I.iw[8] ;
 wire \top_I.branch[4].block[10].um_I.iw[9] ;
 wire \top_I.branch[4].block[10].um_I.k_zero ;
 wire \top_I.branch[4].block[10].um_I.pg_vdd ;
 wire \top_I.branch[4].block[11].um_I.ana[2] ;
 wire \top_I.branch[4].block[11].um_I.ana[3] ;
 wire \top_I.branch[4].block[11].um_I.ana[4] ;
 wire \top_I.branch[4].block[11].um_I.ana[5] ;
 wire \top_I.branch[4].block[11].um_I.ana[6] ;
 wire \top_I.branch[4].block[11].um_I.ana[7] ;
 wire \top_I.branch[4].block[11].um_I.clk ;
 wire \top_I.branch[4].block[11].um_I.ena ;
 wire \top_I.branch[4].block[11].um_I.iw[10] ;
 wire \top_I.branch[4].block[11].um_I.iw[11] ;
 wire \top_I.branch[4].block[11].um_I.iw[12] ;
 wire \top_I.branch[4].block[11].um_I.iw[13] ;
 wire \top_I.branch[4].block[11].um_I.iw[14] ;
 wire \top_I.branch[4].block[11].um_I.iw[15] ;
 wire \top_I.branch[4].block[11].um_I.iw[16] ;
 wire \top_I.branch[4].block[11].um_I.iw[17] ;
 wire \top_I.branch[4].block[11].um_I.iw[1] ;
 wire \top_I.branch[4].block[11].um_I.iw[2] ;
 wire \top_I.branch[4].block[11].um_I.iw[3] ;
 wire \top_I.branch[4].block[11].um_I.iw[4] ;
 wire \top_I.branch[4].block[11].um_I.iw[5] ;
 wire \top_I.branch[4].block[11].um_I.iw[6] ;
 wire \top_I.branch[4].block[11].um_I.iw[7] ;
 wire \top_I.branch[4].block[11].um_I.iw[8] ;
 wire \top_I.branch[4].block[11].um_I.iw[9] ;
 wire \top_I.branch[4].block[11].um_I.k_zero ;
 wire \top_I.branch[4].block[11].um_I.pg_vdd ;
 wire \top_I.branch[4].block[12].um_I.ana[2] ;
 wire \top_I.branch[4].block[12].um_I.ana[3] ;
 wire \top_I.branch[4].block[12].um_I.ana[4] ;
 wire \top_I.branch[4].block[12].um_I.ana[5] ;
 wire \top_I.branch[4].block[12].um_I.ana[6] ;
 wire \top_I.branch[4].block[12].um_I.ana[7] ;
 wire \top_I.branch[4].block[12].um_I.clk ;
 wire \top_I.branch[4].block[12].um_I.ena ;
 wire \top_I.branch[4].block[12].um_I.iw[10] ;
 wire \top_I.branch[4].block[12].um_I.iw[11] ;
 wire \top_I.branch[4].block[12].um_I.iw[12] ;
 wire \top_I.branch[4].block[12].um_I.iw[13] ;
 wire \top_I.branch[4].block[12].um_I.iw[14] ;
 wire \top_I.branch[4].block[12].um_I.iw[15] ;
 wire \top_I.branch[4].block[12].um_I.iw[16] ;
 wire \top_I.branch[4].block[12].um_I.iw[17] ;
 wire \top_I.branch[4].block[12].um_I.iw[1] ;
 wire \top_I.branch[4].block[12].um_I.iw[2] ;
 wire \top_I.branch[4].block[12].um_I.iw[3] ;
 wire \top_I.branch[4].block[12].um_I.iw[4] ;
 wire \top_I.branch[4].block[12].um_I.iw[5] ;
 wire \top_I.branch[4].block[12].um_I.iw[6] ;
 wire \top_I.branch[4].block[12].um_I.iw[7] ;
 wire \top_I.branch[4].block[12].um_I.iw[8] ;
 wire \top_I.branch[4].block[12].um_I.iw[9] ;
 wire \top_I.branch[4].block[12].um_I.k_zero ;
 wire \top_I.branch[4].block[12].um_I.pg_vdd ;
 wire \top_I.branch[4].block[13].um_I.ana[2] ;
 wire \top_I.branch[4].block[13].um_I.ana[3] ;
 wire \top_I.branch[4].block[13].um_I.ana[4] ;
 wire \top_I.branch[4].block[13].um_I.ana[5] ;
 wire \top_I.branch[4].block[13].um_I.ana[6] ;
 wire \top_I.branch[4].block[13].um_I.ana[7] ;
 wire \top_I.branch[4].block[13].um_I.clk ;
 wire \top_I.branch[4].block[13].um_I.ena ;
 wire \top_I.branch[4].block[13].um_I.iw[10] ;
 wire \top_I.branch[4].block[13].um_I.iw[11] ;
 wire \top_I.branch[4].block[13].um_I.iw[12] ;
 wire \top_I.branch[4].block[13].um_I.iw[13] ;
 wire \top_I.branch[4].block[13].um_I.iw[14] ;
 wire \top_I.branch[4].block[13].um_I.iw[15] ;
 wire \top_I.branch[4].block[13].um_I.iw[16] ;
 wire \top_I.branch[4].block[13].um_I.iw[17] ;
 wire \top_I.branch[4].block[13].um_I.iw[1] ;
 wire \top_I.branch[4].block[13].um_I.iw[2] ;
 wire \top_I.branch[4].block[13].um_I.iw[3] ;
 wire \top_I.branch[4].block[13].um_I.iw[4] ;
 wire \top_I.branch[4].block[13].um_I.iw[5] ;
 wire \top_I.branch[4].block[13].um_I.iw[6] ;
 wire \top_I.branch[4].block[13].um_I.iw[7] ;
 wire \top_I.branch[4].block[13].um_I.iw[8] ;
 wire \top_I.branch[4].block[13].um_I.iw[9] ;
 wire \top_I.branch[4].block[13].um_I.k_zero ;
 wire \top_I.branch[4].block[13].um_I.pg_vdd ;
 wire \top_I.branch[4].block[14].um_I.ana[2] ;
 wire \top_I.branch[4].block[14].um_I.ana[3] ;
 wire \top_I.branch[4].block[14].um_I.ana[4] ;
 wire \top_I.branch[4].block[14].um_I.ana[5] ;
 wire \top_I.branch[4].block[14].um_I.ana[6] ;
 wire \top_I.branch[4].block[14].um_I.ana[7] ;
 wire \top_I.branch[4].block[14].um_I.clk ;
 wire \top_I.branch[4].block[14].um_I.ena ;
 wire \top_I.branch[4].block[14].um_I.iw[10] ;
 wire \top_I.branch[4].block[14].um_I.iw[11] ;
 wire \top_I.branch[4].block[14].um_I.iw[12] ;
 wire \top_I.branch[4].block[14].um_I.iw[13] ;
 wire \top_I.branch[4].block[14].um_I.iw[14] ;
 wire \top_I.branch[4].block[14].um_I.iw[15] ;
 wire \top_I.branch[4].block[14].um_I.iw[16] ;
 wire \top_I.branch[4].block[14].um_I.iw[17] ;
 wire \top_I.branch[4].block[14].um_I.iw[1] ;
 wire \top_I.branch[4].block[14].um_I.iw[2] ;
 wire \top_I.branch[4].block[14].um_I.iw[3] ;
 wire \top_I.branch[4].block[14].um_I.iw[4] ;
 wire \top_I.branch[4].block[14].um_I.iw[5] ;
 wire \top_I.branch[4].block[14].um_I.iw[6] ;
 wire \top_I.branch[4].block[14].um_I.iw[7] ;
 wire \top_I.branch[4].block[14].um_I.iw[8] ;
 wire \top_I.branch[4].block[14].um_I.iw[9] ;
 wire \top_I.branch[4].block[14].um_I.k_zero ;
 wire \top_I.branch[4].block[14].um_I.pg_vdd ;
 wire \top_I.branch[4].block[15].um_I.ana[2] ;
 wire \top_I.branch[4].block[15].um_I.ana[3] ;
 wire \top_I.branch[4].block[15].um_I.ana[4] ;
 wire \top_I.branch[4].block[15].um_I.ana[5] ;
 wire \top_I.branch[4].block[15].um_I.ana[6] ;
 wire \top_I.branch[4].block[15].um_I.ana[7] ;
 wire \top_I.branch[4].block[15].um_I.clk ;
 wire \top_I.branch[4].block[15].um_I.ena ;
 wire \top_I.branch[4].block[15].um_I.iw[10] ;
 wire \top_I.branch[4].block[15].um_I.iw[11] ;
 wire \top_I.branch[4].block[15].um_I.iw[12] ;
 wire \top_I.branch[4].block[15].um_I.iw[13] ;
 wire \top_I.branch[4].block[15].um_I.iw[14] ;
 wire \top_I.branch[4].block[15].um_I.iw[15] ;
 wire \top_I.branch[4].block[15].um_I.iw[16] ;
 wire \top_I.branch[4].block[15].um_I.iw[17] ;
 wire \top_I.branch[4].block[15].um_I.iw[1] ;
 wire \top_I.branch[4].block[15].um_I.iw[2] ;
 wire \top_I.branch[4].block[15].um_I.iw[3] ;
 wire \top_I.branch[4].block[15].um_I.iw[4] ;
 wire \top_I.branch[4].block[15].um_I.iw[5] ;
 wire \top_I.branch[4].block[15].um_I.iw[6] ;
 wire \top_I.branch[4].block[15].um_I.iw[7] ;
 wire \top_I.branch[4].block[15].um_I.iw[8] ;
 wire \top_I.branch[4].block[15].um_I.iw[9] ;
 wire \top_I.branch[4].block[15].um_I.k_zero ;
 wire \top_I.branch[4].block[15].um_I.pg_vdd ;
 wire \top_I.branch[4].block[1].um_I.ana[2] ;
 wire \top_I.branch[4].block[1].um_I.ana[3] ;
 wire \top_I.branch[4].block[1].um_I.ana[4] ;
 wire \top_I.branch[4].block[1].um_I.ana[5] ;
 wire \top_I.branch[4].block[1].um_I.ana[6] ;
 wire \top_I.branch[4].block[1].um_I.ana[7] ;
 wire \top_I.branch[4].block[1].um_I.clk ;
 wire \top_I.branch[4].block[1].um_I.ena ;
 wire \top_I.branch[4].block[1].um_I.iw[10] ;
 wire \top_I.branch[4].block[1].um_I.iw[11] ;
 wire \top_I.branch[4].block[1].um_I.iw[12] ;
 wire \top_I.branch[4].block[1].um_I.iw[13] ;
 wire \top_I.branch[4].block[1].um_I.iw[14] ;
 wire \top_I.branch[4].block[1].um_I.iw[15] ;
 wire \top_I.branch[4].block[1].um_I.iw[16] ;
 wire \top_I.branch[4].block[1].um_I.iw[17] ;
 wire \top_I.branch[4].block[1].um_I.iw[1] ;
 wire \top_I.branch[4].block[1].um_I.iw[2] ;
 wire \top_I.branch[4].block[1].um_I.iw[3] ;
 wire \top_I.branch[4].block[1].um_I.iw[4] ;
 wire \top_I.branch[4].block[1].um_I.iw[5] ;
 wire \top_I.branch[4].block[1].um_I.iw[6] ;
 wire \top_I.branch[4].block[1].um_I.iw[7] ;
 wire \top_I.branch[4].block[1].um_I.iw[8] ;
 wire \top_I.branch[4].block[1].um_I.iw[9] ;
 wire \top_I.branch[4].block[1].um_I.k_zero ;
 wire \top_I.branch[4].block[1].um_I.pg_vdd ;
 wire \top_I.branch[4].block[2].um_I.ana[2] ;
 wire \top_I.branch[4].block[2].um_I.ana[3] ;
 wire \top_I.branch[4].block[2].um_I.ana[4] ;
 wire \top_I.branch[4].block[2].um_I.ana[5] ;
 wire \top_I.branch[4].block[2].um_I.ana[6] ;
 wire \top_I.branch[4].block[2].um_I.ana[7] ;
 wire \top_I.branch[4].block[2].um_I.clk ;
 wire \top_I.branch[4].block[2].um_I.ena ;
 wire \top_I.branch[4].block[2].um_I.iw[10] ;
 wire \top_I.branch[4].block[2].um_I.iw[11] ;
 wire \top_I.branch[4].block[2].um_I.iw[12] ;
 wire \top_I.branch[4].block[2].um_I.iw[13] ;
 wire \top_I.branch[4].block[2].um_I.iw[14] ;
 wire \top_I.branch[4].block[2].um_I.iw[15] ;
 wire \top_I.branch[4].block[2].um_I.iw[16] ;
 wire \top_I.branch[4].block[2].um_I.iw[17] ;
 wire \top_I.branch[4].block[2].um_I.iw[1] ;
 wire \top_I.branch[4].block[2].um_I.iw[2] ;
 wire \top_I.branch[4].block[2].um_I.iw[3] ;
 wire \top_I.branch[4].block[2].um_I.iw[4] ;
 wire \top_I.branch[4].block[2].um_I.iw[5] ;
 wire \top_I.branch[4].block[2].um_I.iw[6] ;
 wire \top_I.branch[4].block[2].um_I.iw[7] ;
 wire \top_I.branch[4].block[2].um_I.iw[8] ;
 wire \top_I.branch[4].block[2].um_I.iw[9] ;
 wire \top_I.branch[4].block[2].um_I.k_zero ;
 wire \top_I.branch[4].block[2].um_I.pg_vdd ;
 wire \top_I.branch[4].block[3].um_I.ana[2] ;
 wire \top_I.branch[4].block[3].um_I.ana[3] ;
 wire \top_I.branch[4].block[3].um_I.ana[4] ;
 wire \top_I.branch[4].block[3].um_I.ana[5] ;
 wire \top_I.branch[4].block[3].um_I.ana[6] ;
 wire \top_I.branch[4].block[3].um_I.ana[7] ;
 wire \top_I.branch[4].block[3].um_I.clk ;
 wire \top_I.branch[4].block[3].um_I.ena ;
 wire \top_I.branch[4].block[3].um_I.iw[10] ;
 wire \top_I.branch[4].block[3].um_I.iw[11] ;
 wire \top_I.branch[4].block[3].um_I.iw[12] ;
 wire \top_I.branch[4].block[3].um_I.iw[13] ;
 wire \top_I.branch[4].block[3].um_I.iw[14] ;
 wire \top_I.branch[4].block[3].um_I.iw[15] ;
 wire \top_I.branch[4].block[3].um_I.iw[16] ;
 wire \top_I.branch[4].block[3].um_I.iw[17] ;
 wire \top_I.branch[4].block[3].um_I.iw[1] ;
 wire \top_I.branch[4].block[3].um_I.iw[2] ;
 wire \top_I.branch[4].block[3].um_I.iw[3] ;
 wire \top_I.branch[4].block[3].um_I.iw[4] ;
 wire \top_I.branch[4].block[3].um_I.iw[5] ;
 wire \top_I.branch[4].block[3].um_I.iw[6] ;
 wire \top_I.branch[4].block[3].um_I.iw[7] ;
 wire \top_I.branch[4].block[3].um_I.iw[8] ;
 wire \top_I.branch[4].block[3].um_I.iw[9] ;
 wire \top_I.branch[4].block[3].um_I.k_zero ;
 wire \top_I.branch[4].block[3].um_I.pg_vdd ;
 wire \top_I.branch[4].block[4].um_I.ana[2] ;
 wire \top_I.branch[4].block[4].um_I.ana[3] ;
 wire \top_I.branch[4].block[4].um_I.ana[4] ;
 wire \top_I.branch[4].block[4].um_I.ana[5] ;
 wire \top_I.branch[4].block[4].um_I.ana[6] ;
 wire \top_I.branch[4].block[4].um_I.ana[7] ;
 wire \top_I.branch[4].block[4].um_I.clk ;
 wire \top_I.branch[4].block[4].um_I.ena ;
 wire \top_I.branch[4].block[4].um_I.iw[10] ;
 wire \top_I.branch[4].block[4].um_I.iw[11] ;
 wire \top_I.branch[4].block[4].um_I.iw[12] ;
 wire \top_I.branch[4].block[4].um_I.iw[13] ;
 wire \top_I.branch[4].block[4].um_I.iw[14] ;
 wire \top_I.branch[4].block[4].um_I.iw[15] ;
 wire \top_I.branch[4].block[4].um_I.iw[16] ;
 wire \top_I.branch[4].block[4].um_I.iw[17] ;
 wire \top_I.branch[4].block[4].um_I.iw[1] ;
 wire \top_I.branch[4].block[4].um_I.iw[2] ;
 wire \top_I.branch[4].block[4].um_I.iw[3] ;
 wire \top_I.branch[4].block[4].um_I.iw[4] ;
 wire \top_I.branch[4].block[4].um_I.iw[5] ;
 wire \top_I.branch[4].block[4].um_I.iw[6] ;
 wire \top_I.branch[4].block[4].um_I.iw[7] ;
 wire \top_I.branch[4].block[4].um_I.iw[8] ;
 wire \top_I.branch[4].block[4].um_I.iw[9] ;
 wire \top_I.branch[4].block[4].um_I.k_zero ;
 wire \top_I.branch[4].block[4].um_I.pg_vdd ;
 wire \top_I.branch[4].block[5].um_I.ana[2] ;
 wire \top_I.branch[4].block[5].um_I.ana[3] ;
 wire \top_I.branch[4].block[5].um_I.ana[4] ;
 wire \top_I.branch[4].block[5].um_I.ana[5] ;
 wire \top_I.branch[4].block[5].um_I.ana[6] ;
 wire \top_I.branch[4].block[5].um_I.ana[7] ;
 wire \top_I.branch[4].block[5].um_I.clk ;
 wire \top_I.branch[4].block[5].um_I.ena ;
 wire \top_I.branch[4].block[5].um_I.iw[10] ;
 wire \top_I.branch[4].block[5].um_I.iw[11] ;
 wire \top_I.branch[4].block[5].um_I.iw[12] ;
 wire \top_I.branch[4].block[5].um_I.iw[13] ;
 wire \top_I.branch[4].block[5].um_I.iw[14] ;
 wire \top_I.branch[4].block[5].um_I.iw[15] ;
 wire \top_I.branch[4].block[5].um_I.iw[16] ;
 wire \top_I.branch[4].block[5].um_I.iw[17] ;
 wire \top_I.branch[4].block[5].um_I.iw[1] ;
 wire \top_I.branch[4].block[5].um_I.iw[2] ;
 wire \top_I.branch[4].block[5].um_I.iw[3] ;
 wire \top_I.branch[4].block[5].um_I.iw[4] ;
 wire \top_I.branch[4].block[5].um_I.iw[5] ;
 wire \top_I.branch[4].block[5].um_I.iw[6] ;
 wire \top_I.branch[4].block[5].um_I.iw[7] ;
 wire \top_I.branch[4].block[5].um_I.iw[8] ;
 wire \top_I.branch[4].block[5].um_I.iw[9] ;
 wire \top_I.branch[4].block[5].um_I.k_zero ;
 wire \top_I.branch[4].block[5].um_I.pg_vdd ;
 wire \top_I.branch[4].block[6].um_I.ana[2] ;
 wire \top_I.branch[4].block[6].um_I.ana[3] ;
 wire \top_I.branch[4].block[6].um_I.ana[4] ;
 wire \top_I.branch[4].block[6].um_I.ana[5] ;
 wire \top_I.branch[4].block[6].um_I.ana[6] ;
 wire \top_I.branch[4].block[6].um_I.ana[7] ;
 wire \top_I.branch[4].block[6].um_I.clk ;
 wire \top_I.branch[4].block[6].um_I.ena ;
 wire \top_I.branch[4].block[6].um_I.iw[10] ;
 wire \top_I.branch[4].block[6].um_I.iw[11] ;
 wire \top_I.branch[4].block[6].um_I.iw[12] ;
 wire \top_I.branch[4].block[6].um_I.iw[13] ;
 wire \top_I.branch[4].block[6].um_I.iw[14] ;
 wire \top_I.branch[4].block[6].um_I.iw[15] ;
 wire \top_I.branch[4].block[6].um_I.iw[16] ;
 wire \top_I.branch[4].block[6].um_I.iw[17] ;
 wire \top_I.branch[4].block[6].um_I.iw[1] ;
 wire \top_I.branch[4].block[6].um_I.iw[2] ;
 wire \top_I.branch[4].block[6].um_I.iw[3] ;
 wire \top_I.branch[4].block[6].um_I.iw[4] ;
 wire \top_I.branch[4].block[6].um_I.iw[5] ;
 wire \top_I.branch[4].block[6].um_I.iw[6] ;
 wire \top_I.branch[4].block[6].um_I.iw[7] ;
 wire \top_I.branch[4].block[6].um_I.iw[8] ;
 wire \top_I.branch[4].block[6].um_I.iw[9] ;
 wire \top_I.branch[4].block[6].um_I.k_zero ;
 wire \top_I.branch[4].block[6].um_I.pg_vdd ;
 wire \top_I.branch[4].block[7].um_I.ana[2] ;
 wire \top_I.branch[4].block[7].um_I.ana[3] ;
 wire \top_I.branch[4].block[7].um_I.ana[4] ;
 wire \top_I.branch[4].block[7].um_I.ana[5] ;
 wire \top_I.branch[4].block[7].um_I.ana[6] ;
 wire \top_I.branch[4].block[7].um_I.ana[7] ;
 wire \top_I.branch[4].block[7].um_I.clk ;
 wire \top_I.branch[4].block[7].um_I.ena ;
 wire \top_I.branch[4].block[7].um_I.iw[10] ;
 wire \top_I.branch[4].block[7].um_I.iw[11] ;
 wire \top_I.branch[4].block[7].um_I.iw[12] ;
 wire \top_I.branch[4].block[7].um_I.iw[13] ;
 wire \top_I.branch[4].block[7].um_I.iw[14] ;
 wire \top_I.branch[4].block[7].um_I.iw[15] ;
 wire \top_I.branch[4].block[7].um_I.iw[16] ;
 wire \top_I.branch[4].block[7].um_I.iw[17] ;
 wire \top_I.branch[4].block[7].um_I.iw[1] ;
 wire \top_I.branch[4].block[7].um_I.iw[2] ;
 wire \top_I.branch[4].block[7].um_I.iw[3] ;
 wire \top_I.branch[4].block[7].um_I.iw[4] ;
 wire \top_I.branch[4].block[7].um_I.iw[5] ;
 wire \top_I.branch[4].block[7].um_I.iw[6] ;
 wire \top_I.branch[4].block[7].um_I.iw[7] ;
 wire \top_I.branch[4].block[7].um_I.iw[8] ;
 wire \top_I.branch[4].block[7].um_I.iw[9] ;
 wire \top_I.branch[4].block[7].um_I.k_zero ;
 wire \top_I.branch[4].block[7].um_I.pg_vdd ;
 wire \top_I.branch[4].block[8].um_I.ana[2] ;
 wire \top_I.branch[4].block[8].um_I.ana[3] ;
 wire \top_I.branch[4].block[8].um_I.ana[4] ;
 wire \top_I.branch[4].block[8].um_I.ana[5] ;
 wire \top_I.branch[4].block[8].um_I.ana[6] ;
 wire \top_I.branch[4].block[8].um_I.ana[7] ;
 wire \top_I.branch[4].block[8].um_I.clk ;
 wire \top_I.branch[4].block[8].um_I.ena ;
 wire \top_I.branch[4].block[8].um_I.iw[10] ;
 wire \top_I.branch[4].block[8].um_I.iw[11] ;
 wire \top_I.branch[4].block[8].um_I.iw[12] ;
 wire \top_I.branch[4].block[8].um_I.iw[13] ;
 wire \top_I.branch[4].block[8].um_I.iw[14] ;
 wire \top_I.branch[4].block[8].um_I.iw[15] ;
 wire \top_I.branch[4].block[8].um_I.iw[16] ;
 wire \top_I.branch[4].block[8].um_I.iw[17] ;
 wire \top_I.branch[4].block[8].um_I.iw[1] ;
 wire \top_I.branch[4].block[8].um_I.iw[2] ;
 wire \top_I.branch[4].block[8].um_I.iw[3] ;
 wire \top_I.branch[4].block[8].um_I.iw[4] ;
 wire \top_I.branch[4].block[8].um_I.iw[5] ;
 wire \top_I.branch[4].block[8].um_I.iw[6] ;
 wire \top_I.branch[4].block[8].um_I.iw[7] ;
 wire \top_I.branch[4].block[8].um_I.iw[8] ;
 wire \top_I.branch[4].block[8].um_I.iw[9] ;
 wire \top_I.branch[4].block[8].um_I.k_zero ;
 wire \top_I.branch[4].block[8].um_I.pg_vdd ;
 wire \top_I.branch[4].block[9].um_I.ana[2] ;
 wire \top_I.branch[4].block[9].um_I.ana[3] ;
 wire \top_I.branch[4].block[9].um_I.ana[4] ;
 wire \top_I.branch[4].block[9].um_I.ana[5] ;
 wire \top_I.branch[4].block[9].um_I.ana[6] ;
 wire \top_I.branch[4].block[9].um_I.ana[7] ;
 wire \top_I.branch[4].block[9].um_I.clk ;
 wire \top_I.branch[4].block[9].um_I.ena ;
 wire \top_I.branch[4].block[9].um_I.iw[10] ;
 wire \top_I.branch[4].block[9].um_I.iw[11] ;
 wire \top_I.branch[4].block[9].um_I.iw[12] ;
 wire \top_I.branch[4].block[9].um_I.iw[13] ;
 wire \top_I.branch[4].block[9].um_I.iw[14] ;
 wire \top_I.branch[4].block[9].um_I.iw[15] ;
 wire \top_I.branch[4].block[9].um_I.iw[16] ;
 wire \top_I.branch[4].block[9].um_I.iw[17] ;
 wire \top_I.branch[4].block[9].um_I.iw[1] ;
 wire \top_I.branch[4].block[9].um_I.iw[2] ;
 wire \top_I.branch[4].block[9].um_I.iw[3] ;
 wire \top_I.branch[4].block[9].um_I.iw[4] ;
 wire \top_I.branch[4].block[9].um_I.iw[5] ;
 wire \top_I.branch[4].block[9].um_I.iw[6] ;
 wire \top_I.branch[4].block[9].um_I.iw[7] ;
 wire \top_I.branch[4].block[9].um_I.iw[8] ;
 wire \top_I.branch[4].block[9].um_I.iw[9] ;
 wire \top_I.branch[4].block[9].um_I.k_zero ;
 wire \top_I.branch[4].block[9].um_I.pg_vdd ;
 wire \top_I.branch[4].l_addr[0] ;
 wire \top_I.branch[4].l_addr[1] ;
 wire \top_I.branch[5].block[0].um_I.ana[2] ;
 wire \top_I.branch[5].block[0].um_I.ana[3] ;
 wire \top_I.branch[5].block[0].um_I.ana[4] ;
 wire \top_I.branch[5].block[0].um_I.ana[5] ;
 wire \top_I.branch[5].block[0].um_I.ana[6] ;
 wire \top_I.branch[5].block[0].um_I.ana[7] ;
 wire \top_I.branch[5].block[0].um_I.clk ;
 wire \top_I.branch[5].block[0].um_I.ena ;
 wire \top_I.branch[5].block[0].um_I.iw[10] ;
 wire \top_I.branch[5].block[0].um_I.iw[11] ;
 wire \top_I.branch[5].block[0].um_I.iw[12] ;
 wire \top_I.branch[5].block[0].um_I.iw[13] ;
 wire \top_I.branch[5].block[0].um_I.iw[14] ;
 wire \top_I.branch[5].block[0].um_I.iw[15] ;
 wire \top_I.branch[5].block[0].um_I.iw[16] ;
 wire \top_I.branch[5].block[0].um_I.iw[17] ;
 wire \top_I.branch[5].block[0].um_I.iw[1] ;
 wire \top_I.branch[5].block[0].um_I.iw[2] ;
 wire \top_I.branch[5].block[0].um_I.iw[3] ;
 wire \top_I.branch[5].block[0].um_I.iw[4] ;
 wire \top_I.branch[5].block[0].um_I.iw[5] ;
 wire \top_I.branch[5].block[0].um_I.iw[6] ;
 wire \top_I.branch[5].block[0].um_I.iw[7] ;
 wire \top_I.branch[5].block[0].um_I.iw[8] ;
 wire \top_I.branch[5].block[0].um_I.iw[9] ;
 wire \top_I.branch[5].block[0].um_I.k_zero ;
 wire \top_I.branch[5].block[0].um_I.pg_vdd ;
 wire \top_I.branch[5].block[10].um_I.ana[2] ;
 wire \top_I.branch[5].block[10].um_I.ana[3] ;
 wire \top_I.branch[5].block[10].um_I.ana[4] ;
 wire \top_I.branch[5].block[10].um_I.ana[5] ;
 wire \top_I.branch[5].block[10].um_I.ana[6] ;
 wire \top_I.branch[5].block[10].um_I.ana[7] ;
 wire \top_I.branch[5].block[10].um_I.clk ;
 wire \top_I.branch[5].block[10].um_I.ena ;
 wire \top_I.branch[5].block[10].um_I.iw[10] ;
 wire \top_I.branch[5].block[10].um_I.iw[11] ;
 wire \top_I.branch[5].block[10].um_I.iw[12] ;
 wire \top_I.branch[5].block[10].um_I.iw[13] ;
 wire \top_I.branch[5].block[10].um_I.iw[14] ;
 wire \top_I.branch[5].block[10].um_I.iw[15] ;
 wire \top_I.branch[5].block[10].um_I.iw[16] ;
 wire \top_I.branch[5].block[10].um_I.iw[17] ;
 wire \top_I.branch[5].block[10].um_I.iw[1] ;
 wire \top_I.branch[5].block[10].um_I.iw[2] ;
 wire \top_I.branch[5].block[10].um_I.iw[3] ;
 wire \top_I.branch[5].block[10].um_I.iw[4] ;
 wire \top_I.branch[5].block[10].um_I.iw[5] ;
 wire \top_I.branch[5].block[10].um_I.iw[6] ;
 wire \top_I.branch[5].block[10].um_I.iw[7] ;
 wire \top_I.branch[5].block[10].um_I.iw[8] ;
 wire \top_I.branch[5].block[10].um_I.iw[9] ;
 wire \top_I.branch[5].block[10].um_I.k_zero ;
 wire \top_I.branch[5].block[10].um_I.pg_vdd ;
 wire \top_I.branch[5].block[11].um_I.ana[2] ;
 wire \top_I.branch[5].block[11].um_I.ana[3] ;
 wire \top_I.branch[5].block[11].um_I.ana[4] ;
 wire \top_I.branch[5].block[11].um_I.ana[5] ;
 wire \top_I.branch[5].block[11].um_I.ana[6] ;
 wire \top_I.branch[5].block[11].um_I.ana[7] ;
 wire \top_I.branch[5].block[11].um_I.clk ;
 wire \top_I.branch[5].block[11].um_I.ena ;
 wire \top_I.branch[5].block[11].um_I.iw[10] ;
 wire \top_I.branch[5].block[11].um_I.iw[11] ;
 wire \top_I.branch[5].block[11].um_I.iw[12] ;
 wire \top_I.branch[5].block[11].um_I.iw[13] ;
 wire \top_I.branch[5].block[11].um_I.iw[14] ;
 wire \top_I.branch[5].block[11].um_I.iw[15] ;
 wire \top_I.branch[5].block[11].um_I.iw[16] ;
 wire \top_I.branch[5].block[11].um_I.iw[17] ;
 wire \top_I.branch[5].block[11].um_I.iw[1] ;
 wire \top_I.branch[5].block[11].um_I.iw[2] ;
 wire \top_I.branch[5].block[11].um_I.iw[3] ;
 wire \top_I.branch[5].block[11].um_I.iw[4] ;
 wire \top_I.branch[5].block[11].um_I.iw[5] ;
 wire \top_I.branch[5].block[11].um_I.iw[6] ;
 wire \top_I.branch[5].block[11].um_I.iw[7] ;
 wire \top_I.branch[5].block[11].um_I.iw[8] ;
 wire \top_I.branch[5].block[11].um_I.iw[9] ;
 wire \top_I.branch[5].block[11].um_I.k_zero ;
 wire \top_I.branch[5].block[11].um_I.pg_vdd ;
 wire \top_I.branch[5].block[12].um_I.ana[2] ;
 wire \top_I.branch[5].block[12].um_I.ana[3] ;
 wire \top_I.branch[5].block[12].um_I.ana[4] ;
 wire \top_I.branch[5].block[12].um_I.ana[5] ;
 wire \top_I.branch[5].block[12].um_I.ana[6] ;
 wire \top_I.branch[5].block[12].um_I.ana[7] ;
 wire \top_I.branch[5].block[12].um_I.clk ;
 wire \top_I.branch[5].block[12].um_I.ena ;
 wire \top_I.branch[5].block[12].um_I.iw[10] ;
 wire \top_I.branch[5].block[12].um_I.iw[11] ;
 wire \top_I.branch[5].block[12].um_I.iw[12] ;
 wire \top_I.branch[5].block[12].um_I.iw[13] ;
 wire \top_I.branch[5].block[12].um_I.iw[14] ;
 wire \top_I.branch[5].block[12].um_I.iw[15] ;
 wire \top_I.branch[5].block[12].um_I.iw[16] ;
 wire \top_I.branch[5].block[12].um_I.iw[17] ;
 wire \top_I.branch[5].block[12].um_I.iw[1] ;
 wire \top_I.branch[5].block[12].um_I.iw[2] ;
 wire \top_I.branch[5].block[12].um_I.iw[3] ;
 wire \top_I.branch[5].block[12].um_I.iw[4] ;
 wire \top_I.branch[5].block[12].um_I.iw[5] ;
 wire \top_I.branch[5].block[12].um_I.iw[6] ;
 wire \top_I.branch[5].block[12].um_I.iw[7] ;
 wire \top_I.branch[5].block[12].um_I.iw[8] ;
 wire \top_I.branch[5].block[12].um_I.iw[9] ;
 wire \top_I.branch[5].block[12].um_I.k_zero ;
 wire \top_I.branch[5].block[12].um_I.pg_vdd ;
 wire \top_I.branch[5].block[13].um_I.ana[2] ;
 wire \top_I.branch[5].block[13].um_I.ana[3] ;
 wire \top_I.branch[5].block[13].um_I.ana[4] ;
 wire \top_I.branch[5].block[13].um_I.ana[5] ;
 wire \top_I.branch[5].block[13].um_I.ana[6] ;
 wire \top_I.branch[5].block[13].um_I.ana[7] ;
 wire \top_I.branch[5].block[13].um_I.clk ;
 wire \top_I.branch[5].block[13].um_I.ena ;
 wire \top_I.branch[5].block[13].um_I.iw[10] ;
 wire \top_I.branch[5].block[13].um_I.iw[11] ;
 wire \top_I.branch[5].block[13].um_I.iw[12] ;
 wire \top_I.branch[5].block[13].um_I.iw[13] ;
 wire \top_I.branch[5].block[13].um_I.iw[14] ;
 wire \top_I.branch[5].block[13].um_I.iw[15] ;
 wire \top_I.branch[5].block[13].um_I.iw[16] ;
 wire \top_I.branch[5].block[13].um_I.iw[17] ;
 wire \top_I.branch[5].block[13].um_I.iw[1] ;
 wire \top_I.branch[5].block[13].um_I.iw[2] ;
 wire \top_I.branch[5].block[13].um_I.iw[3] ;
 wire \top_I.branch[5].block[13].um_I.iw[4] ;
 wire \top_I.branch[5].block[13].um_I.iw[5] ;
 wire \top_I.branch[5].block[13].um_I.iw[6] ;
 wire \top_I.branch[5].block[13].um_I.iw[7] ;
 wire \top_I.branch[5].block[13].um_I.iw[8] ;
 wire \top_I.branch[5].block[13].um_I.iw[9] ;
 wire \top_I.branch[5].block[13].um_I.k_zero ;
 wire \top_I.branch[5].block[13].um_I.pg_vdd ;
 wire \top_I.branch[5].block[14].um_I.ana[2] ;
 wire \top_I.branch[5].block[14].um_I.ana[3] ;
 wire \top_I.branch[5].block[14].um_I.ana[4] ;
 wire \top_I.branch[5].block[14].um_I.ana[5] ;
 wire \top_I.branch[5].block[14].um_I.ana[6] ;
 wire \top_I.branch[5].block[14].um_I.ana[7] ;
 wire \top_I.branch[5].block[14].um_I.clk ;
 wire \top_I.branch[5].block[14].um_I.ena ;
 wire \top_I.branch[5].block[14].um_I.iw[10] ;
 wire \top_I.branch[5].block[14].um_I.iw[11] ;
 wire \top_I.branch[5].block[14].um_I.iw[12] ;
 wire \top_I.branch[5].block[14].um_I.iw[13] ;
 wire \top_I.branch[5].block[14].um_I.iw[14] ;
 wire \top_I.branch[5].block[14].um_I.iw[15] ;
 wire \top_I.branch[5].block[14].um_I.iw[16] ;
 wire \top_I.branch[5].block[14].um_I.iw[17] ;
 wire \top_I.branch[5].block[14].um_I.iw[1] ;
 wire \top_I.branch[5].block[14].um_I.iw[2] ;
 wire \top_I.branch[5].block[14].um_I.iw[3] ;
 wire \top_I.branch[5].block[14].um_I.iw[4] ;
 wire \top_I.branch[5].block[14].um_I.iw[5] ;
 wire \top_I.branch[5].block[14].um_I.iw[6] ;
 wire \top_I.branch[5].block[14].um_I.iw[7] ;
 wire \top_I.branch[5].block[14].um_I.iw[8] ;
 wire \top_I.branch[5].block[14].um_I.iw[9] ;
 wire \top_I.branch[5].block[14].um_I.k_zero ;
 wire \top_I.branch[5].block[14].um_I.pg_vdd ;
 wire \top_I.branch[5].block[15].um_I.ana[2] ;
 wire \top_I.branch[5].block[15].um_I.ana[3] ;
 wire \top_I.branch[5].block[15].um_I.ana[4] ;
 wire \top_I.branch[5].block[15].um_I.ana[5] ;
 wire \top_I.branch[5].block[15].um_I.ana[6] ;
 wire \top_I.branch[5].block[15].um_I.ana[7] ;
 wire \top_I.branch[5].block[15].um_I.clk ;
 wire \top_I.branch[5].block[15].um_I.ena ;
 wire \top_I.branch[5].block[15].um_I.iw[10] ;
 wire \top_I.branch[5].block[15].um_I.iw[11] ;
 wire \top_I.branch[5].block[15].um_I.iw[12] ;
 wire \top_I.branch[5].block[15].um_I.iw[13] ;
 wire \top_I.branch[5].block[15].um_I.iw[14] ;
 wire \top_I.branch[5].block[15].um_I.iw[15] ;
 wire \top_I.branch[5].block[15].um_I.iw[16] ;
 wire \top_I.branch[5].block[15].um_I.iw[17] ;
 wire \top_I.branch[5].block[15].um_I.iw[1] ;
 wire \top_I.branch[5].block[15].um_I.iw[2] ;
 wire \top_I.branch[5].block[15].um_I.iw[3] ;
 wire \top_I.branch[5].block[15].um_I.iw[4] ;
 wire \top_I.branch[5].block[15].um_I.iw[5] ;
 wire \top_I.branch[5].block[15].um_I.iw[6] ;
 wire \top_I.branch[5].block[15].um_I.iw[7] ;
 wire \top_I.branch[5].block[15].um_I.iw[8] ;
 wire \top_I.branch[5].block[15].um_I.iw[9] ;
 wire \top_I.branch[5].block[15].um_I.k_zero ;
 wire \top_I.branch[5].block[15].um_I.pg_vdd ;
 wire \top_I.branch[5].block[1].um_I.ana[2] ;
 wire \top_I.branch[5].block[1].um_I.ana[3] ;
 wire \top_I.branch[5].block[1].um_I.ana[4] ;
 wire \top_I.branch[5].block[1].um_I.ana[5] ;
 wire \top_I.branch[5].block[1].um_I.ana[6] ;
 wire \top_I.branch[5].block[1].um_I.ana[7] ;
 wire \top_I.branch[5].block[1].um_I.clk ;
 wire \top_I.branch[5].block[1].um_I.ena ;
 wire \top_I.branch[5].block[1].um_I.iw[10] ;
 wire \top_I.branch[5].block[1].um_I.iw[11] ;
 wire \top_I.branch[5].block[1].um_I.iw[12] ;
 wire \top_I.branch[5].block[1].um_I.iw[13] ;
 wire \top_I.branch[5].block[1].um_I.iw[14] ;
 wire \top_I.branch[5].block[1].um_I.iw[15] ;
 wire \top_I.branch[5].block[1].um_I.iw[16] ;
 wire \top_I.branch[5].block[1].um_I.iw[17] ;
 wire \top_I.branch[5].block[1].um_I.iw[1] ;
 wire \top_I.branch[5].block[1].um_I.iw[2] ;
 wire \top_I.branch[5].block[1].um_I.iw[3] ;
 wire \top_I.branch[5].block[1].um_I.iw[4] ;
 wire \top_I.branch[5].block[1].um_I.iw[5] ;
 wire \top_I.branch[5].block[1].um_I.iw[6] ;
 wire \top_I.branch[5].block[1].um_I.iw[7] ;
 wire \top_I.branch[5].block[1].um_I.iw[8] ;
 wire \top_I.branch[5].block[1].um_I.iw[9] ;
 wire \top_I.branch[5].block[1].um_I.k_zero ;
 wire \top_I.branch[5].block[1].um_I.pg_vdd ;
 wire \top_I.branch[5].block[2].um_I.ana[2] ;
 wire \top_I.branch[5].block[2].um_I.ana[3] ;
 wire \top_I.branch[5].block[2].um_I.ana[4] ;
 wire \top_I.branch[5].block[2].um_I.ana[5] ;
 wire \top_I.branch[5].block[2].um_I.ana[6] ;
 wire \top_I.branch[5].block[2].um_I.ana[7] ;
 wire \top_I.branch[5].block[2].um_I.clk ;
 wire \top_I.branch[5].block[2].um_I.ena ;
 wire \top_I.branch[5].block[2].um_I.iw[10] ;
 wire \top_I.branch[5].block[2].um_I.iw[11] ;
 wire \top_I.branch[5].block[2].um_I.iw[12] ;
 wire \top_I.branch[5].block[2].um_I.iw[13] ;
 wire \top_I.branch[5].block[2].um_I.iw[14] ;
 wire \top_I.branch[5].block[2].um_I.iw[15] ;
 wire \top_I.branch[5].block[2].um_I.iw[16] ;
 wire \top_I.branch[5].block[2].um_I.iw[17] ;
 wire \top_I.branch[5].block[2].um_I.iw[1] ;
 wire \top_I.branch[5].block[2].um_I.iw[2] ;
 wire \top_I.branch[5].block[2].um_I.iw[3] ;
 wire \top_I.branch[5].block[2].um_I.iw[4] ;
 wire \top_I.branch[5].block[2].um_I.iw[5] ;
 wire \top_I.branch[5].block[2].um_I.iw[6] ;
 wire \top_I.branch[5].block[2].um_I.iw[7] ;
 wire \top_I.branch[5].block[2].um_I.iw[8] ;
 wire \top_I.branch[5].block[2].um_I.iw[9] ;
 wire \top_I.branch[5].block[2].um_I.k_zero ;
 wire \top_I.branch[5].block[2].um_I.pg_vdd ;
 wire \top_I.branch[5].block[3].um_I.ana[2] ;
 wire \top_I.branch[5].block[3].um_I.ana[3] ;
 wire \top_I.branch[5].block[3].um_I.ana[4] ;
 wire \top_I.branch[5].block[3].um_I.ana[5] ;
 wire \top_I.branch[5].block[3].um_I.ana[6] ;
 wire \top_I.branch[5].block[3].um_I.ana[7] ;
 wire \top_I.branch[5].block[3].um_I.clk ;
 wire \top_I.branch[5].block[3].um_I.ena ;
 wire \top_I.branch[5].block[3].um_I.iw[10] ;
 wire \top_I.branch[5].block[3].um_I.iw[11] ;
 wire \top_I.branch[5].block[3].um_I.iw[12] ;
 wire \top_I.branch[5].block[3].um_I.iw[13] ;
 wire \top_I.branch[5].block[3].um_I.iw[14] ;
 wire \top_I.branch[5].block[3].um_I.iw[15] ;
 wire \top_I.branch[5].block[3].um_I.iw[16] ;
 wire \top_I.branch[5].block[3].um_I.iw[17] ;
 wire \top_I.branch[5].block[3].um_I.iw[1] ;
 wire \top_I.branch[5].block[3].um_I.iw[2] ;
 wire \top_I.branch[5].block[3].um_I.iw[3] ;
 wire \top_I.branch[5].block[3].um_I.iw[4] ;
 wire \top_I.branch[5].block[3].um_I.iw[5] ;
 wire \top_I.branch[5].block[3].um_I.iw[6] ;
 wire \top_I.branch[5].block[3].um_I.iw[7] ;
 wire \top_I.branch[5].block[3].um_I.iw[8] ;
 wire \top_I.branch[5].block[3].um_I.iw[9] ;
 wire \top_I.branch[5].block[3].um_I.k_zero ;
 wire \top_I.branch[5].block[3].um_I.pg_vdd ;
 wire \top_I.branch[5].block[4].um_I.ana[2] ;
 wire \top_I.branch[5].block[4].um_I.ana[3] ;
 wire \top_I.branch[5].block[4].um_I.ana[4] ;
 wire \top_I.branch[5].block[4].um_I.ana[5] ;
 wire \top_I.branch[5].block[4].um_I.ana[6] ;
 wire \top_I.branch[5].block[4].um_I.ana[7] ;
 wire \top_I.branch[5].block[4].um_I.clk ;
 wire \top_I.branch[5].block[4].um_I.ena ;
 wire \top_I.branch[5].block[4].um_I.iw[10] ;
 wire \top_I.branch[5].block[4].um_I.iw[11] ;
 wire \top_I.branch[5].block[4].um_I.iw[12] ;
 wire \top_I.branch[5].block[4].um_I.iw[13] ;
 wire \top_I.branch[5].block[4].um_I.iw[14] ;
 wire \top_I.branch[5].block[4].um_I.iw[15] ;
 wire \top_I.branch[5].block[4].um_I.iw[16] ;
 wire \top_I.branch[5].block[4].um_I.iw[17] ;
 wire \top_I.branch[5].block[4].um_I.iw[1] ;
 wire \top_I.branch[5].block[4].um_I.iw[2] ;
 wire \top_I.branch[5].block[4].um_I.iw[3] ;
 wire \top_I.branch[5].block[4].um_I.iw[4] ;
 wire \top_I.branch[5].block[4].um_I.iw[5] ;
 wire \top_I.branch[5].block[4].um_I.iw[6] ;
 wire \top_I.branch[5].block[4].um_I.iw[7] ;
 wire \top_I.branch[5].block[4].um_I.iw[8] ;
 wire \top_I.branch[5].block[4].um_I.iw[9] ;
 wire \top_I.branch[5].block[4].um_I.k_zero ;
 wire \top_I.branch[5].block[4].um_I.pg_vdd ;
 wire \top_I.branch[5].block[5].um_I.ana[2] ;
 wire \top_I.branch[5].block[5].um_I.ana[3] ;
 wire \top_I.branch[5].block[5].um_I.ana[4] ;
 wire \top_I.branch[5].block[5].um_I.ana[5] ;
 wire \top_I.branch[5].block[5].um_I.ana[6] ;
 wire \top_I.branch[5].block[5].um_I.ana[7] ;
 wire \top_I.branch[5].block[5].um_I.clk ;
 wire \top_I.branch[5].block[5].um_I.ena ;
 wire \top_I.branch[5].block[5].um_I.iw[10] ;
 wire \top_I.branch[5].block[5].um_I.iw[11] ;
 wire \top_I.branch[5].block[5].um_I.iw[12] ;
 wire \top_I.branch[5].block[5].um_I.iw[13] ;
 wire \top_I.branch[5].block[5].um_I.iw[14] ;
 wire \top_I.branch[5].block[5].um_I.iw[15] ;
 wire \top_I.branch[5].block[5].um_I.iw[16] ;
 wire \top_I.branch[5].block[5].um_I.iw[17] ;
 wire \top_I.branch[5].block[5].um_I.iw[1] ;
 wire \top_I.branch[5].block[5].um_I.iw[2] ;
 wire \top_I.branch[5].block[5].um_I.iw[3] ;
 wire \top_I.branch[5].block[5].um_I.iw[4] ;
 wire \top_I.branch[5].block[5].um_I.iw[5] ;
 wire \top_I.branch[5].block[5].um_I.iw[6] ;
 wire \top_I.branch[5].block[5].um_I.iw[7] ;
 wire \top_I.branch[5].block[5].um_I.iw[8] ;
 wire \top_I.branch[5].block[5].um_I.iw[9] ;
 wire \top_I.branch[5].block[5].um_I.k_zero ;
 wire \top_I.branch[5].block[5].um_I.pg_vdd ;
 wire \top_I.branch[5].block[6].um_I.ana[2] ;
 wire \top_I.branch[5].block[6].um_I.ana[3] ;
 wire \top_I.branch[5].block[6].um_I.ana[4] ;
 wire \top_I.branch[5].block[6].um_I.ana[5] ;
 wire \top_I.branch[5].block[6].um_I.ana[6] ;
 wire \top_I.branch[5].block[6].um_I.ana[7] ;
 wire \top_I.branch[5].block[6].um_I.clk ;
 wire \top_I.branch[5].block[6].um_I.ena ;
 wire \top_I.branch[5].block[6].um_I.iw[10] ;
 wire \top_I.branch[5].block[6].um_I.iw[11] ;
 wire \top_I.branch[5].block[6].um_I.iw[12] ;
 wire \top_I.branch[5].block[6].um_I.iw[13] ;
 wire \top_I.branch[5].block[6].um_I.iw[14] ;
 wire \top_I.branch[5].block[6].um_I.iw[15] ;
 wire \top_I.branch[5].block[6].um_I.iw[16] ;
 wire \top_I.branch[5].block[6].um_I.iw[17] ;
 wire \top_I.branch[5].block[6].um_I.iw[1] ;
 wire \top_I.branch[5].block[6].um_I.iw[2] ;
 wire \top_I.branch[5].block[6].um_I.iw[3] ;
 wire \top_I.branch[5].block[6].um_I.iw[4] ;
 wire \top_I.branch[5].block[6].um_I.iw[5] ;
 wire \top_I.branch[5].block[6].um_I.iw[6] ;
 wire \top_I.branch[5].block[6].um_I.iw[7] ;
 wire \top_I.branch[5].block[6].um_I.iw[8] ;
 wire \top_I.branch[5].block[6].um_I.iw[9] ;
 wire \top_I.branch[5].block[6].um_I.k_zero ;
 wire \top_I.branch[5].block[6].um_I.pg_vdd ;
 wire \top_I.branch[5].block[7].um_I.ana[2] ;
 wire \top_I.branch[5].block[7].um_I.ana[3] ;
 wire \top_I.branch[5].block[7].um_I.ana[4] ;
 wire \top_I.branch[5].block[7].um_I.ana[5] ;
 wire \top_I.branch[5].block[7].um_I.ana[6] ;
 wire \top_I.branch[5].block[7].um_I.ana[7] ;
 wire \top_I.branch[5].block[7].um_I.clk ;
 wire \top_I.branch[5].block[7].um_I.ena ;
 wire \top_I.branch[5].block[7].um_I.iw[10] ;
 wire \top_I.branch[5].block[7].um_I.iw[11] ;
 wire \top_I.branch[5].block[7].um_I.iw[12] ;
 wire \top_I.branch[5].block[7].um_I.iw[13] ;
 wire \top_I.branch[5].block[7].um_I.iw[14] ;
 wire \top_I.branch[5].block[7].um_I.iw[15] ;
 wire \top_I.branch[5].block[7].um_I.iw[16] ;
 wire \top_I.branch[5].block[7].um_I.iw[17] ;
 wire \top_I.branch[5].block[7].um_I.iw[1] ;
 wire \top_I.branch[5].block[7].um_I.iw[2] ;
 wire \top_I.branch[5].block[7].um_I.iw[3] ;
 wire \top_I.branch[5].block[7].um_I.iw[4] ;
 wire \top_I.branch[5].block[7].um_I.iw[5] ;
 wire \top_I.branch[5].block[7].um_I.iw[6] ;
 wire \top_I.branch[5].block[7].um_I.iw[7] ;
 wire \top_I.branch[5].block[7].um_I.iw[8] ;
 wire \top_I.branch[5].block[7].um_I.iw[9] ;
 wire \top_I.branch[5].block[7].um_I.k_zero ;
 wire \top_I.branch[5].block[7].um_I.pg_vdd ;
 wire \top_I.branch[5].block[8].um_I.ana[2] ;
 wire \top_I.branch[5].block[8].um_I.ana[3] ;
 wire \top_I.branch[5].block[8].um_I.ana[4] ;
 wire \top_I.branch[5].block[8].um_I.ana[5] ;
 wire \top_I.branch[5].block[8].um_I.ana[6] ;
 wire \top_I.branch[5].block[8].um_I.ana[7] ;
 wire \top_I.branch[5].block[8].um_I.clk ;
 wire \top_I.branch[5].block[8].um_I.ena ;
 wire \top_I.branch[5].block[8].um_I.iw[10] ;
 wire \top_I.branch[5].block[8].um_I.iw[11] ;
 wire \top_I.branch[5].block[8].um_I.iw[12] ;
 wire \top_I.branch[5].block[8].um_I.iw[13] ;
 wire \top_I.branch[5].block[8].um_I.iw[14] ;
 wire \top_I.branch[5].block[8].um_I.iw[15] ;
 wire \top_I.branch[5].block[8].um_I.iw[16] ;
 wire \top_I.branch[5].block[8].um_I.iw[17] ;
 wire \top_I.branch[5].block[8].um_I.iw[1] ;
 wire \top_I.branch[5].block[8].um_I.iw[2] ;
 wire \top_I.branch[5].block[8].um_I.iw[3] ;
 wire \top_I.branch[5].block[8].um_I.iw[4] ;
 wire \top_I.branch[5].block[8].um_I.iw[5] ;
 wire \top_I.branch[5].block[8].um_I.iw[6] ;
 wire \top_I.branch[5].block[8].um_I.iw[7] ;
 wire \top_I.branch[5].block[8].um_I.iw[8] ;
 wire \top_I.branch[5].block[8].um_I.iw[9] ;
 wire \top_I.branch[5].block[8].um_I.k_zero ;
 wire \top_I.branch[5].block[8].um_I.pg_vdd ;
 wire \top_I.branch[5].block[9].um_I.ana[2] ;
 wire \top_I.branch[5].block[9].um_I.ana[3] ;
 wire \top_I.branch[5].block[9].um_I.ana[4] ;
 wire \top_I.branch[5].block[9].um_I.ana[5] ;
 wire \top_I.branch[5].block[9].um_I.ana[6] ;
 wire \top_I.branch[5].block[9].um_I.ana[7] ;
 wire \top_I.branch[5].block[9].um_I.clk ;
 wire \top_I.branch[5].block[9].um_I.ena ;
 wire \top_I.branch[5].block[9].um_I.iw[10] ;
 wire \top_I.branch[5].block[9].um_I.iw[11] ;
 wire \top_I.branch[5].block[9].um_I.iw[12] ;
 wire \top_I.branch[5].block[9].um_I.iw[13] ;
 wire \top_I.branch[5].block[9].um_I.iw[14] ;
 wire \top_I.branch[5].block[9].um_I.iw[15] ;
 wire \top_I.branch[5].block[9].um_I.iw[16] ;
 wire \top_I.branch[5].block[9].um_I.iw[17] ;
 wire \top_I.branch[5].block[9].um_I.iw[1] ;
 wire \top_I.branch[5].block[9].um_I.iw[2] ;
 wire \top_I.branch[5].block[9].um_I.iw[3] ;
 wire \top_I.branch[5].block[9].um_I.iw[4] ;
 wire \top_I.branch[5].block[9].um_I.iw[5] ;
 wire \top_I.branch[5].block[9].um_I.iw[6] ;
 wire \top_I.branch[5].block[9].um_I.iw[7] ;
 wire \top_I.branch[5].block[9].um_I.iw[8] ;
 wire \top_I.branch[5].block[9].um_I.iw[9] ;
 wire \top_I.branch[5].block[9].um_I.k_zero ;
 wire \top_I.branch[5].block[9].um_I.pg_vdd ;
 wire \top_I.branch[5].l_addr[0] ;
 wire \top_I.branch[5].l_addr[1] ;
 wire \top_I.branch[6].block[0].um_I.ana[2] ;
 wire \top_I.branch[6].block[0].um_I.ana[3] ;
 wire \top_I.branch[6].block[0].um_I.ana[4] ;
 wire \top_I.branch[6].block[0].um_I.ana[5] ;
 wire \top_I.branch[6].block[0].um_I.ana[6] ;
 wire \top_I.branch[6].block[0].um_I.ana[7] ;
 wire \top_I.branch[6].block[0].um_I.clk ;
 wire \top_I.branch[6].block[0].um_I.ena ;
 wire \top_I.branch[6].block[0].um_I.iw[10] ;
 wire \top_I.branch[6].block[0].um_I.iw[11] ;
 wire \top_I.branch[6].block[0].um_I.iw[12] ;
 wire \top_I.branch[6].block[0].um_I.iw[13] ;
 wire \top_I.branch[6].block[0].um_I.iw[14] ;
 wire \top_I.branch[6].block[0].um_I.iw[15] ;
 wire \top_I.branch[6].block[0].um_I.iw[16] ;
 wire \top_I.branch[6].block[0].um_I.iw[17] ;
 wire \top_I.branch[6].block[0].um_I.iw[1] ;
 wire \top_I.branch[6].block[0].um_I.iw[2] ;
 wire \top_I.branch[6].block[0].um_I.iw[3] ;
 wire \top_I.branch[6].block[0].um_I.iw[4] ;
 wire \top_I.branch[6].block[0].um_I.iw[5] ;
 wire \top_I.branch[6].block[0].um_I.iw[6] ;
 wire \top_I.branch[6].block[0].um_I.iw[7] ;
 wire \top_I.branch[6].block[0].um_I.iw[8] ;
 wire \top_I.branch[6].block[0].um_I.iw[9] ;
 wire \top_I.branch[6].block[0].um_I.k_zero ;
 wire \top_I.branch[6].block[0].um_I.pg_vdd ;
 wire \top_I.branch[6].block[10].um_I.ana[2] ;
 wire \top_I.branch[6].block[10].um_I.ana[3] ;
 wire \top_I.branch[6].block[10].um_I.ana[4] ;
 wire \top_I.branch[6].block[10].um_I.ana[5] ;
 wire \top_I.branch[6].block[10].um_I.ana[6] ;
 wire \top_I.branch[6].block[10].um_I.ana[7] ;
 wire \top_I.branch[6].block[10].um_I.clk ;
 wire \top_I.branch[6].block[10].um_I.ena ;
 wire \top_I.branch[6].block[10].um_I.iw[10] ;
 wire \top_I.branch[6].block[10].um_I.iw[11] ;
 wire \top_I.branch[6].block[10].um_I.iw[12] ;
 wire \top_I.branch[6].block[10].um_I.iw[13] ;
 wire \top_I.branch[6].block[10].um_I.iw[14] ;
 wire \top_I.branch[6].block[10].um_I.iw[15] ;
 wire \top_I.branch[6].block[10].um_I.iw[16] ;
 wire \top_I.branch[6].block[10].um_I.iw[17] ;
 wire \top_I.branch[6].block[10].um_I.iw[1] ;
 wire \top_I.branch[6].block[10].um_I.iw[2] ;
 wire \top_I.branch[6].block[10].um_I.iw[3] ;
 wire \top_I.branch[6].block[10].um_I.iw[4] ;
 wire \top_I.branch[6].block[10].um_I.iw[5] ;
 wire \top_I.branch[6].block[10].um_I.iw[6] ;
 wire \top_I.branch[6].block[10].um_I.iw[7] ;
 wire \top_I.branch[6].block[10].um_I.iw[8] ;
 wire \top_I.branch[6].block[10].um_I.iw[9] ;
 wire \top_I.branch[6].block[10].um_I.k_zero ;
 wire \top_I.branch[6].block[10].um_I.pg_vdd ;
 wire \top_I.branch[6].block[11].um_I.ana[2] ;
 wire \top_I.branch[6].block[11].um_I.ana[3] ;
 wire \top_I.branch[6].block[11].um_I.ana[4] ;
 wire \top_I.branch[6].block[11].um_I.ana[5] ;
 wire \top_I.branch[6].block[11].um_I.ana[6] ;
 wire \top_I.branch[6].block[11].um_I.ana[7] ;
 wire \top_I.branch[6].block[11].um_I.clk ;
 wire \top_I.branch[6].block[11].um_I.ena ;
 wire \top_I.branch[6].block[11].um_I.iw[10] ;
 wire \top_I.branch[6].block[11].um_I.iw[11] ;
 wire \top_I.branch[6].block[11].um_I.iw[12] ;
 wire \top_I.branch[6].block[11].um_I.iw[13] ;
 wire \top_I.branch[6].block[11].um_I.iw[14] ;
 wire \top_I.branch[6].block[11].um_I.iw[15] ;
 wire \top_I.branch[6].block[11].um_I.iw[16] ;
 wire \top_I.branch[6].block[11].um_I.iw[17] ;
 wire \top_I.branch[6].block[11].um_I.iw[1] ;
 wire \top_I.branch[6].block[11].um_I.iw[2] ;
 wire \top_I.branch[6].block[11].um_I.iw[3] ;
 wire \top_I.branch[6].block[11].um_I.iw[4] ;
 wire \top_I.branch[6].block[11].um_I.iw[5] ;
 wire \top_I.branch[6].block[11].um_I.iw[6] ;
 wire \top_I.branch[6].block[11].um_I.iw[7] ;
 wire \top_I.branch[6].block[11].um_I.iw[8] ;
 wire \top_I.branch[6].block[11].um_I.iw[9] ;
 wire \top_I.branch[6].block[11].um_I.k_zero ;
 wire \top_I.branch[6].block[11].um_I.pg_vdd ;
 wire \top_I.branch[6].block[12].um_I.ana[2] ;
 wire \top_I.branch[6].block[12].um_I.ana[3] ;
 wire \top_I.branch[6].block[12].um_I.ana[4] ;
 wire \top_I.branch[6].block[12].um_I.ana[5] ;
 wire \top_I.branch[6].block[12].um_I.ana[6] ;
 wire \top_I.branch[6].block[12].um_I.ana[7] ;
 wire \top_I.branch[6].block[12].um_I.clk ;
 wire \top_I.branch[6].block[12].um_I.ena ;
 wire \top_I.branch[6].block[12].um_I.iw[10] ;
 wire \top_I.branch[6].block[12].um_I.iw[11] ;
 wire \top_I.branch[6].block[12].um_I.iw[12] ;
 wire \top_I.branch[6].block[12].um_I.iw[13] ;
 wire \top_I.branch[6].block[12].um_I.iw[14] ;
 wire \top_I.branch[6].block[12].um_I.iw[15] ;
 wire \top_I.branch[6].block[12].um_I.iw[16] ;
 wire \top_I.branch[6].block[12].um_I.iw[17] ;
 wire \top_I.branch[6].block[12].um_I.iw[1] ;
 wire \top_I.branch[6].block[12].um_I.iw[2] ;
 wire \top_I.branch[6].block[12].um_I.iw[3] ;
 wire \top_I.branch[6].block[12].um_I.iw[4] ;
 wire \top_I.branch[6].block[12].um_I.iw[5] ;
 wire \top_I.branch[6].block[12].um_I.iw[6] ;
 wire \top_I.branch[6].block[12].um_I.iw[7] ;
 wire \top_I.branch[6].block[12].um_I.iw[8] ;
 wire \top_I.branch[6].block[12].um_I.iw[9] ;
 wire \top_I.branch[6].block[12].um_I.k_zero ;
 wire \top_I.branch[6].block[12].um_I.pg_vdd ;
 wire \top_I.branch[6].block[13].um_I.ana[2] ;
 wire \top_I.branch[6].block[13].um_I.ana[3] ;
 wire \top_I.branch[6].block[13].um_I.ana[4] ;
 wire \top_I.branch[6].block[13].um_I.ana[5] ;
 wire \top_I.branch[6].block[13].um_I.ana[6] ;
 wire \top_I.branch[6].block[13].um_I.ana[7] ;
 wire \top_I.branch[6].block[13].um_I.clk ;
 wire \top_I.branch[6].block[13].um_I.ena ;
 wire \top_I.branch[6].block[13].um_I.iw[10] ;
 wire \top_I.branch[6].block[13].um_I.iw[11] ;
 wire \top_I.branch[6].block[13].um_I.iw[12] ;
 wire \top_I.branch[6].block[13].um_I.iw[13] ;
 wire \top_I.branch[6].block[13].um_I.iw[14] ;
 wire \top_I.branch[6].block[13].um_I.iw[15] ;
 wire \top_I.branch[6].block[13].um_I.iw[16] ;
 wire \top_I.branch[6].block[13].um_I.iw[17] ;
 wire \top_I.branch[6].block[13].um_I.iw[1] ;
 wire \top_I.branch[6].block[13].um_I.iw[2] ;
 wire \top_I.branch[6].block[13].um_I.iw[3] ;
 wire \top_I.branch[6].block[13].um_I.iw[4] ;
 wire \top_I.branch[6].block[13].um_I.iw[5] ;
 wire \top_I.branch[6].block[13].um_I.iw[6] ;
 wire \top_I.branch[6].block[13].um_I.iw[7] ;
 wire \top_I.branch[6].block[13].um_I.iw[8] ;
 wire \top_I.branch[6].block[13].um_I.iw[9] ;
 wire \top_I.branch[6].block[13].um_I.k_zero ;
 wire \top_I.branch[6].block[13].um_I.pg_vdd ;
 wire \top_I.branch[6].block[14].um_I.ana[2] ;
 wire \top_I.branch[6].block[14].um_I.ana[3] ;
 wire \top_I.branch[6].block[14].um_I.ana[4] ;
 wire \top_I.branch[6].block[14].um_I.ana[5] ;
 wire \top_I.branch[6].block[14].um_I.ana[6] ;
 wire \top_I.branch[6].block[14].um_I.ana[7] ;
 wire \top_I.branch[6].block[14].um_I.clk ;
 wire \top_I.branch[6].block[14].um_I.ena ;
 wire \top_I.branch[6].block[14].um_I.iw[10] ;
 wire \top_I.branch[6].block[14].um_I.iw[11] ;
 wire \top_I.branch[6].block[14].um_I.iw[12] ;
 wire \top_I.branch[6].block[14].um_I.iw[13] ;
 wire \top_I.branch[6].block[14].um_I.iw[14] ;
 wire \top_I.branch[6].block[14].um_I.iw[15] ;
 wire \top_I.branch[6].block[14].um_I.iw[16] ;
 wire \top_I.branch[6].block[14].um_I.iw[17] ;
 wire \top_I.branch[6].block[14].um_I.iw[1] ;
 wire \top_I.branch[6].block[14].um_I.iw[2] ;
 wire \top_I.branch[6].block[14].um_I.iw[3] ;
 wire \top_I.branch[6].block[14].um_I.iw[4] ;
 wire \top_I.branch[6].block[14].um_I.iw[5] ;
 wire \top_I.branch[6].block[14].um_I.iw[6] ;
 wire \top_I.branch[6].block[14].um_I.iw[7] ;
 wire \top_I.branch[6].block[14].um_I.iw[8] ;
 wire \top_I.branch[6].block[14].um_I.iw[9] ;
 wire \top_I.branch[6].block[14].um_I.k_zero ;
 wire \top_I.branch[6].block[14].um_I.pg_vdd ;
 wire \top_I.branch[6].block[15].um_I.ana[2] ;
 wire \top_I.branch[6].block[15].um_I.ana[3] ;
 wire \top_I.branch[6].block[15].um_I.ana[4] ;
 wire \top_I.branch[6].block[15].um_I.ana[5] ;
 wire \top_I.branch[6].block[15].um_I.ana[6] ;
 wire \top_I.branch[6].block[15].um_I.ana[7] ;
 wire \top_I.branch[6].block[15].um_I.clk ;
 wire \top_I.branch[6].block[15].um_I.ena ;
 wire \top_I.branch[6].block[15].um_I.iw[10] ;
 wire \top_I.branch[6].block[15].um_I.iw[11] ;
 wire \top_I.branch[6].block[15].um_I.iw[12] ;
 wire \top_I.branch[6].block[15].um_I.iw[13] ;
 wire \top_I.branch[6].block[15].um_I.iw[14] ;
 wire \top_I.branch[6].block[15].um_I.iw[15] ;
 wire \top_I.branch[6].block[15].um_I.iw[16] ;
 wire \top_I.branch[6].block[15].um_I.iw[17] ;
 wire \top_I.branch[6].block[15].um_I.iw[1] ;
 wire \top_I.branch[6].block[15].um_I.iw[2] ;
 wire \top_I.branch[6].block[15].um_I.iw[3] ;
 wire \top_I.branch[6].block[15].um_I.iw[4] ;
 wire \top_I.branch[6].block[15].um_I.iw[5] ;
 wire \top_I.branch[6].block[15].um_I.iw[6] ;
 wire \top_I.branch[6].block[15].um_I.iw[7] ;
 wire \top_I.branch[6].block[15].um_I.iw[8] ;
 wire \top_I.branch[6].block[15].um_I.iw[9] ;
 wire \top_I.branch[6].block[15].um_I.k_zero ;
 wire \top_I.branch[6].block[15].um_I.pg_vdd ;
 wire \top_I.branch[6].block[1].um_I.ana[2] ;
 wire \top_I.branch[6].block[1].um_I.ana[3] ;
 wire \top_I.branch[6].block[1].um_I.ana[4] ;
 wire \top_I.branch[6].block[1].um_I.ana[5] ;
 wire \top_I.branch[6].block[1].um_I.ana[6] ;
 wire \top_I.branch[6].block[1].um_I.ana[7] ;
 wire \top_I.branch[6].block[1].um_I.clk ;
 wire \top_I.branch[6].block[1].um_I.ena ;
 wire \top_I.branch[6].block[1].um_I.iw[10] ;
 wire \top_I.branch[6].block[1].um_I.iw[11] ;
 wire \top_I.branch[6].block[1].um_I.iw[12] ;
 wire \top_I.branch[6].block[1].um_I.iw[13] ;
 wire \top_I.branch[6].block[1].um_I.iw[14] ;
 wire \top_I.branch[6].block[1].um_I.iw[15] ;
 wire \top_I.branch[6].block[1].um_I.iw[16] ;
 wire \top_I.branch[6].block[1].um_I.iw[17] ;
 wire \top_I.branch[6].block[1].um_I.iw[1] ;
 wire \top_I.branch[6].block[1].um_I.iw[2] ;
 wire \top_I.branch[6].block[1].um_I.iw[3] ;
 wire \top_I.branch[6].block[1].um_I.iw[4] ;
 wire \top_I.branch[6].block[1].um_I.iw[5] ;
 wire \top_I.branch[6].block[1].um_I.iw[6] ;
 wire \top_I.branch[6].block[1].um_I.iw[7] ;
 wire \top_I.branch[6].block[1].um_I.iw[8] ;
 wire \top_I.branch[6].block[1].um_I.iw[9] ;
 wire \top_I.branch[6].block[1].um_I.k_zero ;
 wire \top_I.branch[6].block[1].um_I.pg_vdd ;
 wire \top_I.branch[6].block[2].um_I.ana[2] ;
 wire \top_I.branch[6].block[2].um_I.ana[3] ;
 wire \top_I.branch[6].block[2].um_I.ana[4] ;
 wire \top_I.branch[6].block[2].um_I.ana[5] ;
 wire \top_I.branch[6].block[2].um_I.ana[6] ;
 wire \top_I.branch[6].block[2].um_I.ana[7] ;
 wire \top_I.branch[6].block[2].um_I.clk ;
 wire \top_I.branch[6].block[2].um_I.ena ;
 wire \top_I.branch[6].block[2].um_I.iw[10] ;
 wire \top_I.branch[6].block[2].um_I.iw[11] ;
 wire \top_I.branch[6].block[2].um_I.iw[12] ;
 wire \top_I.branch[6].block[2].um_I.iw[13] ;
 wire \top_I.branch[6].block[2].um_I.iw[14] ;
 wire \top_I.branch[6].block[2].um_I.iw[15] ;
 wire \top_I.branch[6].block[2].um_I.iw[16] ;
 wire \top_I.branch[6].block[2].um_I.iw[17] ;
 wire \top_I.branch[6].block[2].um_I.iw[1] ;
 wire \top_I.branch[6].block[2].um_I.iw[2] ;
 wire \top_I.branch[6].block[2].um_I.iw[3] ;
 wire \top_I.branch[6].block[2].um_I.iw[4] ;
 wire \top_I.branch[6].block[2].um_I.iw[5] ;
 wire \top_I.branch[6].block[2].um_I.iw[6] ;
 wire \top_I.branch[6].block[2].um_I.iw[7] ;
 wire \top_I.branch[6].block[2].um_I.iw[8] ;
 wire \top_I.branch[6].block[2].um_I.iw[9] ;
 wire \top_I.branch[6].block[2].um_I.k_zero ;
 wire \top_I.branch[6].block[2].um_I.pg_vdd ;
 wire \top_I.branch[6].block[3].um_I.ana[2] ;
 wire \top_I.branch[6].block[3].um_I.ana[3] ;
 wire \top_I.branch[6].block[3].um_I.ana[4] ;
 wire \top_I.branch[6].block[3].um_I.ana[5] ;
 wire \top_I.branch[6].block[3].um_I.ana[6] ;
 wire \top_I.branch[6].block[3].um_I.ana[7] ;
 wire \top_I.branch[6].block[3].um_I.clk ;
 wire \top_I.branch[6].block[3].um_I.ena ;
 wire \top_I.branch[6].block[3].um_I.iw[10] ;
 wire \top_I.branch[6].block[3].um_I.iw[11] ;
 wire \top_I.branch[6].block[3].um_I.iw[12] ;
 wire \top_I.branch[6].block[3].um_I.iw[13] ;
 wire \top_I.branch[6].block[3].um_I.iw[14] ;
 wire \top_I.branch[6].block[3].um_I.iw[15] ;
 wire \top_I.branch[6].block[3].um_I.iw[16] ;
 wire \top_I.branch[6].block[3].um_I.iw[17] ;
 wire \top_I.branch[6].block[3].um_I.iw[1] ;
 wire \top_I.branch[6].block[3].um_I.iw[2] ;
 wire \top_I.branch[6].block[3].um_I.iw[3] ;
 wire \top_I.branch[6].block[3].um_I.iw[4] ;
 wire \top_I.branch[6].block[3].um_I.iw[5] ;
 wire \top_I.branch[6].block[3].um_I.iw[6] ;
 wire \top_I.branch[6].block[3].um_I.iw[7] ;
 wire \top_I.branch[6].block[3].um_I.iw[8] ;
 wire \top_I.branch[6].block[3].um_I.iw[9] ;
 wire \top_I.branch[6].block[3].um_I.k_zero ;
 wire \top_I.branch[6].block[3].um_I.pg_vdd ;
 wire \top_I.branch[6].block[4].um_I.ana[2] ;
 wire \top_I.branch[6].block[4].um_I.ana[3] ;
 wire \top_I.branch[6].block[4].um_I.ana[4] ;
 wire \top_I.branch[6].block[4].um_I.ana[5] ;
 wire \top_I.branch[6].block[4].um_I.ana[6] ;
 wire \top_I.branch[6].block[4].um_I.ana[7] ;
 wire \top_I.branch[6].block[4].um_I.clk ;
 wire \top_I.branch[6].block[4].um_I.ena ;
 wire \top_I.branch[6].block[4].um_I.iw[10] ;
 wire \top_I.branch[6].block[4].um_I.iw[11] ;
 wire \top_I.branch[6].block[4].um_I.iw[12] ;
 wire \top_I.branch[6].block[4].um_I.iw[13] ;
 wire \top_I.branch[6].block[4].um_I.iw[14] ;
 wire \top_I.branch[6].block[4].um_I.iw[15] ;
 wire \top_I.branch[6].block[4].um_I.iw[16] ;
 wire \top_I.branch[6].block[4].um_I.iw[17] ;
 wire \top_I.branch[6].block[4].um_I.iw[1] ;
 wire \top_I.branch[6].block[4].um_I.iw[2] ;
 wire \top_I.branch[6].block[4].um_I.iw[3] ;
 wire \top_I.branch[6].block[4].um_I.iw[4] ;
 wire \top_I.branch[6].block[4].um_I.iw[5] ;
 wire \top_I.branch[6].block[4].um_I.iw[6] ;
 wire \top_I.branch[6].block[4].um_I.iw[7] ;
 wire \top_I.branch[6].block[4].um_I.iw[8] ;
 wire \top_I.branch[6].block[4].um_I.iw[9] ;
 wire \top_I.branch[6].block[4].um_I.k_zero ;
 wire \top_I.branch[6].block[4].um_I.pg_vdd ;
 wire \top_I.branch[6].block[5].um_I.ana[2] ;
 wire \top_I.branch[6].block[5].um_I.ana[3] ;
 wire \top_I.branch[6].block[5].um_I.ana[4] ;
 wire \top_I.branch[6].block[5].um_I.ana[5] ;
 wire \top_I.branch[6].block[5].um_I.ana[6] ;
 wire \top_I.branch[6].block[5].um_I.ana[7] ;
 wire \top_I.branch[6].block[5].um_I.clk ;
 wire \top_I.branch[6].block[5].um_I.ena ;
 wire \top_I.branch[6].block[5].um_I.iw[10] ;
 wire \top_I.branch[6].block[5].um_I.iw[11] ;
 wire \top_I.branch[6].block[5].um_I.iw[12] ;
 wire \top_I.branch[6].block[5].um_I.iw[13] ;
 wire \top_I.branch[6].block[5].um_I.iw[14] ;
 wire \top_I.branch[6].block[5].um_I.iw[15] ;
 wire \top_I.branch[6].block[5].um_I.iw[16] ;
 wire \top_I.branch[6].block[5].um_I.iw[17] ;
 wire \top_I.branch[6].block[5].um_I.iw[1] ;
 wire \top_I.branch[6].block[5].um_I.iw[2] ;
 wire \top_I.branch[6].block[5].um_I.iw[3] ;
 wire \top_I.branch[6].block[5].um_I.iw[4] ;
 wire \top_I.branch[6].block[5].um_I.iw[5] ;
 wire \top_I.branch[6].block[5].um_I.iw[6] ;
 wire \top_I.branch[6].block[5].um_I.iw[7] ;
 wire \top_I.branch[6].block[5].um_I.iw[8] ;
 wire \top_I.branch[6].block[5].um_I.iw[9] ;
 wire \top_I.branch[6].block[5].um_I.k_zero ;
 wire \top_I.branch[6].block[5].um_I.pg_vdd ;
 wire \top_I.branch[6].block[6].um_I.ana[2] ;
 wire \top_I.branch[6].block[6].um_I.ana[3] ;
 wire \top_I.branch[6].block[6].um_I.ana[4] ;
 wire \top_I.branch[6].block[6].um_I.ana[5] ;
 wire \top_I.branch[6].block[6].um_I.ana[6] ;
 wire \top_I.branch[6].block[6].um_I.ana[7] ;
 wire \top_I.branch[6].block[6].um_I.clk ;
 wire \top_I.branch[6].block[6].um_I.ena ;
 wire \top_I.branch[6].block[6].um_I.iw[10] ;
 wire \top_I.branch[6].block[6].um_I.iw[11] ;
 wire \top_I.branch[6].block[6].um_I.iw[12] ;
 wire \top_I.branch[6].block[6].um_I.iw[13] ;
 wire \top_I.branch[6].block[6].um_I.iw[14] ;
 wire \top_I.branch[6].block[6].um_I.iw[15] ;
 wire \top_I.branch[6].block[6].um_I.iw[16] ;
 wire \top_I.branch[6].block[6].um_I.iw[17] ;
 wire \top_I.branch[6].block[6].um_I.iw[1] ;
 wire \top_I.branch[6].block[6].um_I.iw[2] ;
 wire \top_I.branch[6].block[6].um_I.iw[3] ;
 wire \top_I.branch[6].block[6].um_I.iw[4] ;
 wire \top_I.branch[6].block[6].um_I.iw[5] ;
 wire \top_I.branch[6].block[6].um_I.iw[6] ;
 wire \top_I.branch[6].block[6].um_I.iw[7] ;
 wire \top_I.branch[6].block[6].um_I.iw[8] ;
 wire \top_I.branch[6].block[6].um_I.iw[9] ;
 wire \top_I.branch[6].block[6].um_I.k_zero ;
 wire \top_I.branch[6].block[6].um_I.pg_vdd ;
 wire \top_I.branch[6].block[7].um_I.ana[2] ;
 wire \top_I.branch[6].block[7].um_I.ana[3] ;
 wire \top_I.branch[6].block[7].um_I.ana[4] ;
 wire \top_I.branch[6].block[7].um_I.ana[5] ;
 wire \top_I.branch[6].block[7].um_I.ana[6] ;
 wire \top_I.branch[6].block[7].um_I.ana[7] ;
 wire \top_I.branch[6].block[7].um_I.clk ;
 wire \top_I.branch[6].block[7].um_I.ena ;
 wire \top_I.branch[6].block[7].um_I.iw[10] ;
 wire \top_I.branch[6].block[7].um_I.iw[11] ;
 wire \top_I.branch[6].block[7].um_I.iw[12] ;
 wire \top_I.branch[6].block[7].um_I.iw[13] ;
 wire \top_I.branch[6].block[7].um_I.iw[14] ;
 wire \top_I.branch[6].block[7].um_I.iw[15] ;
 wire \top_I.branch[6].block[7].um_I.iw[16] ;
 wire \top_I.branch[6].block[7].um_I.iw[17] ;
 wire \top_I.branch[6].block[7].um_I.iw[1] ;
 wire \top_I.branch[6].block[7].um_I.iw[2] ;
 wire \top_I.branch[6].block[7].um_I.iw[3] ;
 wire \top_I.branch[6].block[7].um_I.iw[4] ;
 wire \top_I.branch[6].block[7].um_I.iw[5] ;
 wire \top_I.branch[6].block[7].um_I.iw[6] ;
 wire \top_I.branch[6].block[7].um_I.iw[7] ;
 wire \top_I.branch[6].block[7].um_I.iw[8] ;
 wire \top_I.branch[6].block[7].um_I.iw[9] ;
 wire \top_I.branch[6].block[7].um_I.k_zero ;
 wire \top_I.branch[6].block[7].um_I.pg_vdd ;
 wire \top_I.branch[6].block[8].um_I.ana[2] ;
 wire \top_I.branch[6].block[8].um_I.ana[3] ;
 wire \top_I.branch[6].block[8].um_I.ana[4] ;
 wire \top_I.branch[6].block[8].um_I.ana[5] ;
 wire \top_I.branch[6].block[8].um_I.ana[6] ;
 wire \top_I.branch[6].block[8].um_I.ana[7] ;
 wire \top_I.branch[6].block[8].um_I.clk ;
 wire \top_I.branch[6].block[8].um_I.ena ;
 wire \top_I.branch[6].block[8].um_I.iw[10] ;
 wire \top_I.branch[6].block[8].um_I.iw[11] ;
 wire \top_I.branch[6].block[8].um_I.iw[12] ;
 wire \top_I.branch[6].block[8].um_I.iw[13] ;
 wire \top_I.branch[6].block[8].um_I.iw[14] ;
 wire \top_I.branch[6].block[8].um_I.iw[15] ;
 wire \top_I.branch[6].block[8].um_I.iw[16] ;
 wire \top_I.branch[6].block[8].um_I.iw[17] ;
 wire \top_I.branch[6].block[8].um_I.iw[1] ;
 wire \top_I.branch[6].block[8].um_I.iw[2] ;
 wire \top_I.branch[6].block[8].um_I.iw[3] ;
 wire \top_I.branch[6].block[8].um_I.iw[4] ;
 wire \top_I.branch[6].block[8].um_I.iw[5] ;
 wire \top_I.branch[6].block[8].um_I.iw[6] ;
 wire \top_I.branch[6].block[8].um_I.iw[7] ;
 wire \top_I.branch[6].block[8].um_I.iw[8] ;
 wire \top_I.branch[6].block[8].um_I.iw[9] ;
 wire \top_I.branch[6].block[8].um_I.k_zero ;
 wire \top_I.branch[6].block[8].um_I.pg_vdd ;
 wire \top_I.branch[6].block[9].um_I.ana[2] ;
 wire \top_I.branch[6].block[9].um_I.ana[3] ;
 wire \top_I.branch[6].block[9].um_I.ana[4] ;
 wire \top_I.branch[6].block[9].um_I.ana[5] ;
 wire \top_I.branch[6].block[9].um_I.ana[6] ;
 wire \top_I.branch[6].block[9].um_I.ana[7] ;
 wire \top_I.branch[6].block[9].um_I.clk ;
 wire \top_I.branch[6].block[9].um_I.ena ;
 wire \top_I.branch[6].block[9].um_I.iw[10] ;
 wire \top_I.branch[6].block[9].um_I.iw[11] ;
 wire \top_I.branch[6].block[9].um_I.iw[12] ;
 wire \top_I.branch[6].block[9].um_I.iw[13] ;
 wire \top_I.branch[6].block[9].um_I.iw[14] ;
 wire \top_I.branch[6].block[9].um_I.iw[15] ;
 wire \top_I.branch[6].block[9].um_I.iw[16] ;
 wire \top_I.branch[6].block[9].um_I.iw[17] ;
 wire \top_I.branch[6].block[9].um_I.iw[1] ;
 wire \top_I.branch[6].block[9].um_I.iw[2] ;
 wire \top_I.branch[6].block[9].um_I.iw[3] ;
 wire \top_I.branch[6].block[9].um_I.iw[4] ;
 wire \top_I.branch[6].block[9].um_I.iw[5] ;
 wire \top_I.branch[6].block[9].um_I.iw[6] ;
 wire \top_I.branch[6].block[9].um_I.iw[7] ;
 wire \top_I.branch[6].block[9].um_I.iw[8] ;
 wire \top_I.branch[6].block[9].um_I.iw[9] ;
 wire \top_I.branch[6].block[9].um_I.k_zero ;
 wire \top_I.branch[6].block[9].um_I.pg_vdd ;
 wire \top_I.branch[6].l_addr[0] ;
 wire \top_I.branch[6].l_addr[2] ;
 wire \top_I.branch[7].block[0].um_I.ana[2] ;
 wire \top_I.branch[7].block[0].um_I.ana[3] ;
 wire \top_I.branch[7].block[0].um_I.ana[4] ;
 wire \top_I.branch[7].block[0].um_I.ana[5] ;
 wire \top_I.branch[7].block[0].um_I.ana[6] ;
 wire \top_I.branch[7].block[0].um_I.ana[7] ;
 wire \top_I.branch[7].block[0].um_I.clk ;
 wire \top_I.branch[7].block[0].um_I.ena ;
 wire \top_I.branch[7].block[0].um_I.iw[10] ;
 wire \top_I.branch[7].block[0].um_I.iw[11] ;
 wire \top_I.branch[7].block[0].um_I.iw[12] ;
 wire \top_I.branch[7].block[0].um_I.iw[13] ;
 wire \top_I.branch[7].block[0].um_I.iw[14] ;
 wire \top_I.branch[7].block[0].um_I.iw[15] ;
 wire \top_I.branch[7].block[0].um_I.iw[16] ;
 wire \top_I.branch[7].block[0].um_I.iw[17] ;
 wire \top_I.branch[7].block[0].um_I.iw[1] ;
 wire \top_I.branch[7].block[0].um_I.iw[2] ;
 wire \top_I.branch[7].block[0].um_I.iw[3] ;
 wire \top_I.branch[7].block[0].um_I.iw[4] ;
 wire \top_I.branch[7].block[0].um_I.iw[5] ;
 wire \top_I.branch[7].block[0].um_I.iw[6] ;
 wire \top_I.branch[7].block[0].um_I.iw[7] ;
 wire \top_I.branch[7].block[0].um_I.iw[8] ;
 wire \top_I.branch[7].block[0].um_I.iw[9] ;
 wire \top_I.branch[7].block[0].um_I.k_zero ;
 wire \top_I.branch[7].block[0].um_I.pg_vdd ;
 wire \top_I.branch[7].block[10].um_I.ana[2] ;
 wire \top_I.branch[7].block[10].um_I.ana[3] ;
 wire \top_I.branch[7].block[10].um_I.ana[4] ;
 wire \top_I.branch[7].block[10].um_I.ana[5] ;
 wire \top_I.branch[7].block[10].um_I.ana[6] ;
 wire \top_I.branch[7].block[10].um_I.ana[7] ;
 wire \top_I.branch[7].block[10].um_I.clk ;
 wire \top_I.branch[7].block[10].um_I.ena ;
 wire \top_I.branch[7].block[10].um_I.iw[10] ;
 wire \top_I.branch[7].block[10].um_I.iw[11] ;
 wire \top_I.branch[7].block[10].um_I.iw[12] ;
 wire \top_I.branch[7].block[10].um_I.iw[13] ;
 wire \top_I.branch[7].block[10].um_I.iw[14] ;
 wire \top_I.branch[7].block[10].um_I.iw[15] ;
 wire \top_I.branch[7].block[10].um_I.iw[16] ;
 wire \top_I.branch[7].block[10].um_I.iw[17] ;
 wire \top_I.branch[7].block[10].um_I.iw[1] ;
 wire \top_I.branch[7].block[10].um_I.iw[2] ;
 wire \top_I.branch[7].block[10].um_I.iw[3] ;
 wire \top_I.branch[7].block[10].um_I.iw[4] ;
 wire \top_I.branch[7].block[10].um_I.iw[5] ;
 wire \top_I.branch[7].block[10].um_I.iw[6] ;
 wire \top_I.branch[7].block[10].um_I.iw[7] ;
 wire \top_I.branch[7].block[10].um_I.iw[8] ;
 wire \top_I.branch[7].block[10].um_I.iw[9] ;
 wire \top_I.branch[7].block[10].um_I.k_zero ;
 wire \top_I.branch[7].block[10].um_I.pg_vdd ;
 wire \top_I.branch[7].block[11].um_I.ana[2] ;
 wire \top_I.branch[7].block[11].um_I.ana[3] ;
 wire \top_I.branch[7].block[11].um_I.ana[4] ;
 wire \top_I.branch[7].block[11].um_I.ana[5] ;
 wire \top_I.branch[7].block[11].um_I.ana[6] ;
 wire \top_I.branch[7].block[11].um_I.ana[7] ;
 wire \top_I.branch[7].block[11].um_I.clk ;
 wire \top_I.branch[7].block[11].um_I.ena ;
 wire \top_I.branch[7].block[11].um_I.iw[10] ;
 wire \top_I.branch[7].block[11].um_I.iw[11] ;
 wire \top_I.branch[7].block[11].um_I.iw[12] ;
 wire \top_I.branch[7].block[11].um_I.iw[13] ;
 wire \top_I.branch[7].block[11].um_I.iw[14] ;
 wire \top_I.branch[7].block[11].um_I.iw[15] ;
 wire \top_I.branch[7].block[11].um_I.iw[16] ;
 wire \top_I.branch[7].block[11].um_I.iw[17] ;
 wire \top_I.branch[7].block[11].um_I.iw[1] ;
 wire \top_I.branch[7].block[11].um_I.iw[2] ;
 wire \top_I.branch[7].block[11].um_I.iw[3] ;
 wire \top_I.branch[7].block[11].um_I.iw[4] ;
 wire \top_I.branch[7].block[11].um_I.iw[5] ;
 wire \top_I.branch[7].block[11].um_I.iw[6] ;
 wire \top_I.branch[7].block[11].um_I.iw[7] ;
 wire \top_I.branch[7].block[11].um_I.iw[8] ;
 wire \top_I.branch[7].block[11].um_I.iw[9] ;
 wire \top_I.branch[7].block[11].um_I.k_zero ;
 wire \top_I.branch[7].block[11].um_I.pg_vdd ;
 wire \top_I.branch[7].block[12].um_I.ana[2] ;
 wire \top_I.branch[7].block[12].um_I.ana[3] ;
 wire \top_I.branch[7].block[12].um_I.ana[4] ;
 wire \top_I.branch[7].block[12].um_I.ana[5] ;
 wire \top_I.branch[7].block[12].um_I.ana[6] ;
 wire \top_I.branch[7].block[12].um_I.ana[7] ;
 wire \top_I.branch[7].block[12].um_I.clk ;
 wire \top_I.branch[7].block[12].um_I.ena ;
 wire \top_I.branch[7].block[12].um_I.iw[10] ;
 wire \top_I.branch[7].block[12].um_I.iw[11] ;
 wire \top_I.branch[7].block[12].um_I.iw[12] ;
 wire \top_I.branch[7].block[12].um_I.iw[13] ;
 wire \top_I.branch[7].block[12].um_I.iw[14] ;
 wire \top_I.branch[7].block[12].um_I.iw[15] ;
 wire \top_I.branch[7].block[12].um_I.iw[16] ;
 wire \top_I.branch[7].block[12].um_I.iw[17] ;
 wire \top_I.branch[7].block[12].um_I.iw[1] ;
 wire \top_I.branch[7].block[12].um_I.iw[2] ;
 wire \top_I.branch[7].block[12].um_I.iw[3] ;
 wire \top_I.branch[7].block[12].um_I.iw[4] ;
 wire \top_I.branch[7].block[12].um_I.iw[5] ;
 wire \top_I.branch[7].block[12].um_I.iw[6] ;
 wire \top_I.branch[7].block[12].um_I.iw[7] ;
 wire \top_I.branch[7].block[12].um_I.iw[8] ;
 wire \top_I.branch[7].block[12].um_I.iw[9] ;
 wire \top_I.branch[7].block[12].um_I.k_zero ;
 wire \top_I.branch[7].block[12].um_I.pg_vdd ;
 wire \top_I.branch[7].block[13].um_I.ana[2] ;
 wire \top_I.branch[7].block[13].um_I.ana[3] ;
 wire \top_I.branch[7].block[13].um_I.ana[4] ;
 wire \top_I.branch[7].block[13].um_I.ana[5] ;
 wire \top_I.branch[7].block[13].um_I.ana[6] ;
 wire \top_I.branch[7].block[13].um_I.ana[7] ;
 wire \top_I.branch[7].block[13].um_I.clk ;
 wire \top_I.branch[7].block[13].um_I.ena ;
 wire \top_I.branch[7].block[13].um_I.iw[10] ;
 wire \top_I.branch[7].block[13].um_I.iw[11] ;
 wire \top_I.branch[7].block[13].um_I.iw[12] ;
 wire \top_I.branch[7].block[13].um_I.iw[13] ;
 wire \top_I.branch[7].block[13].um_I.iw[14] ;
 wire \top_I.branch[7].block[13].um_I.iw[15] ;
 wire \top_I.branch[7].block[13].um_I.iw[16] ;
 wire \top_I.branch[7].block[13].um_I.iw[17] ;
 wire \top_I.branch[7].block[13].um_I.iw[1] ;
 wire \top_I.branch[7].block[13].um_I.iw[2] ;
 wire \top_I.branch[7].block[13].um_I.iw[3] ;
 wire \top_I.branch[7].block[13].um_I.iw[4] ;
 wire \top_I.branch[7].block[13].um_I.iw[5] ;
 wire \top_I.branch[7].block[13].um_I.iw[6] ;
 wire \top_I.branch[7].block[13].um_I.iw[7] ;
 wire \top_I.branch[7].block[13].um_I.iw[8] ;
 wire \top_I.branch[7].block[13].um_I.iw[9] ;
 wire \top_I.branch[7].block[13].um_I.k_zero ;
 wire \top_I.branch[7].block[13].um_I.pg_vdd ;
 wire \top_I.branch[7].block[14].um_I.ana[2] ;
 wire \top_I.branch[7].block[14].um_I.ana[3] ;
 wire \top_I.branch[7].block[14].um_I.ana[4] ;
 wire \top_I.branch[7].block[14].um_I.ana[5] ;
 wire \top_I.branch[7].block[14].um_I.ana[6] ;
 wire \top_I.branch[7].block[14].um_I.ana[7] ;
 wire \top_I.branch[7].block[14].um_I.clk ;
 wire \top_I.branch[7].block[14].um_I.ena ;
 wire \top_I.branch[7].block[14].um_I.iw[10] ;
 wire \top_I.branch[7].block[14].um_I.iw[11] ;
 wire \top_I.branch[7].block[14].um_I.iw[12] ;
 wire \top_I.branch[7].block[14].um_I.iw[13] ;
 wire \top_I.branch[7].block[14].um_I.iw[14] ;
 wire \top_I.branch[7].block[14].um_I.iw[15] ;
 wire \top_I.branch[7].block[14].um_I.iw[16] ;
 wire \top_I.branch[7].block[14].um_I.iw[17] ;
 wire \top_I.branch[7].block[14].um_I.iw[1] ;
 wire \top_I.branch[7].block[14].um_I.iw[2] ;
 wire \top_I.branch[7].block[14].um_I.iw[3] ;
 wire \top_I.branch[7].block[14].um_I.iw[4] ;
 wire \top_I.branch[7].block[14].um_I.iw[5] ;
 wire \top_I.branch[7].block[14].um_I.iw[6] ;
 wire \top_I.branch[7].block[14].um_I.iw[7] ;
 wire \top_I.branch[7].block[14].um_I.iw[8] ;
 wire \top_I.branch[7].block[14].um_I.iw[9] ;
 wire \top_I.branch[7].block[14].um_I.k_zero ;
 wire \top_I.branch[7].block[14].um_I.pg_vdd ;
 wire \top_I.branch[7].block[15].um_I.ana[2] ;
 wire \top_I.branch[7].block[15].um_I.ana[3] ;
 wire \top_I.branch[7].block[15].um_I.ana[4] ;
 wire \top_I.branch[7].block[15].um_I.ana[5] ;
 wire \top_I.branch[7].block[15].um_I.ana[6] ;
 wire \top_I.branch[7].block[15].um_I.ana[7] ;
 wire \top_I.branch[7].block[15].um_I.clk ;
 wire \top_I.branch[7].block[15].um_I.ena ;
 wire \top_I.branch[7].block[15].um_I.iw[10] ;
 wire \top_I.branch[7].block[15].um_I.iw[11] ;
 wire \top_I.branch[7].block[15].um_I.iw[12] ;
 wire \top_I.branch[7].block[15].um_I.iw[13] ;
 wire \top_I.branch[7].block[15].um_I.iw[14] ;
 wire \top_I.branch[7].block[15].um_I.iw[15] ;
 wire \top_I.branch[7].block[15].um_I.iw[16] ;
 wire \top_I.branch[7].block[15].um_I.iw[17] ;
 wire \top_I.branch[7].block[15].um_I.iw[1] ;
 wire \top_I.branch[7].block[15].um_I.iw[2] ;
 wire \top_I.branch[7].block[15].um_I.iw[3] ;
 wire \top_I.branch[7].block[15].um_I.iw[4] ;
 wire \top_I.branch[7].block[15].um_I.iw[5] ;
 wire \top_I.branch[7].block[15].um_I.iw[6] ;
 wire \top_I.branch[7].block[15].um_I.iw[7] ;
 wire \top_I.branch[7].block[15].um_I.iw[8] ;
 wire \top_I.branch[7].block[15].um_I.iw[9] ;
 wire \top_I.branch[7].block[15].um_I.k_zero ;
 wire \top_I.branch[7].block[15].um_I.pg_vdd ;
 wire \top_I.branch[7].block[1].um_I.ana[2] ;
 wire \top_I.branch[7].block[1].um_I.ana[3] ;
 wire \top_I.branch[7].block[1].um_I.ana[4] ;
 wire \top_I.branch[7].block[1].um_I.ana[5] ;
 wire \top_I.branch[7].block[1].um_I.ana[6] ;
 wire \top_I.branch[7].block[1].um_I.ana[7] ;
 wire \top_I.branch[7].block[1].um_I.clk ;
 wire \top_I.branch[7].block[1].um_I.ena ;
 wire \top_I.branch[7].block[1].um_I.iw[10] ;
 wire \top_I.branch[7].block[1].um_I.iw[11] ;
 wire \top_I.branch[7].block[1].um_I.iw[12] ;
 wire \top_I.branch[7].block[1].um_I.iw[13] ;
 wire \top_I.branch[7].block[1].um_I.iw[14] ;
 wire \top_I.branch[7].block[1].um_I.iw[15] ;
 wire \top_I.branch[7].block[1].um_I.iw[16] ;
 wire \top_I.branch[7].block[1].um_I.iw[17] ;
 wire \top_I.branch[7].block[1].um_I.iw[1] ;
 wire \top_I.branch[7].block[1].um_I.iw[2] ;
 wire \top_I.branch[7].block[1].um_I.iw[3] ;
 wire \top_I.branch[7].block[1].um_I.iw[4] ;
 wire \top_I.branch[7].block[1].um_I.iw[5] ;
 wire \top_I.branch[7].block[1].um_I.iw[6] ;
 wire \top_I.branch[7].block[1].um_I.iw[7] ;
 wire \top_I.branch[7].block[1].um_I.iw[8] ;
 wire \top_I.branch[7].block[1].um_I.iw[9] ;
 wire \top_I.branch[7].block[1].um_I.k_zero ;
 wire \top_I.branch[7].block[1].um_I.pg_vdd ;
 wire \top_I.branch[7].block[2].um_I.ana[2] ;
 wire \top_I.branch[7].block[2].um_I.ana[3] ;
 wire \top_I.branch[7].block[2].um_I.ana[4] ;
 wire \top_I.branch[7].block[2].um_I.ana[5] ;
 wire \top_I.branch[7].block[2].um_I.ana[6] ;
 wire \top_I.branch[7].block[2].um_I.ana[7] ;
 wire \top_I.branch[7].block[2].um_I.clk ;
 wire \top_I.branch[7].block[2].um_I.ena ;
 wire \top_I.branch[7].block[2].um_I.iw[10] ;
 wire \top_I.branch[7].block[2].um_I.iw[11] ;
 wire \top_I.branch[7].block[2].um_I.iw[12] ;
 wire \top_I.branch[7].block[2].um_I.iw[13] ;
 wire \top_I.branch[7].block[2].um_I.iw[14] ;
 wire \top_I.branch[7].block[2].um_I.iw[15] ;
 wire \top_I.branch[7].block[2].um_I.iw[16] ;
 wire \top_I.branch[7].block[2].um_I.iw[17] ;
 wire \top_I.branch[7].block[2].um_I.iw[1] ;
 wire \top_I.branch[7].block[2].um_I.iw[2] ;
 wire \top_I.branch[7].block[2].um_I.iw[3] ;
 wire \top_I.branch[7].block[2].um_I.iw[4] ;
 wire \top_I.branch[7].block[2].um_I.iw[5] ;
 wire \top_I.branch[7].block[2].um_I.iw[6] ;
 wire \top_I.branch[7].block[2].um_I.iw[7] ;
 wire \top_I.branch[7].block[2].um_I.iw[8] ;
 wire \top_I.branch[7].block[2].um_I.iw[9] ;
 wire \top_I.branch[7].block[2].um_I.k_zero ;
 wire \top_I.branch[7].block[2].um_I.pg_vdd ;
 wire \top_I.branch[7].block[3].um_I.ana[2] ;
 wire \top_I.branch[7].block[3].um_I.ana[3] ;
 wire \top_I.branch[7].block[3].um_I.ana[4] ;
 wire \top_I.branch[7].block[3].um_I.ana[5] ;
 wire \top_I.branch[7].block[3].um_I.ana[6] ;
 wire \top_I.branch[7].block[3].um_I.ana[7] ;
 wire \top_I.branch[7].block[3].um_I.clk ;
 wire \top_I.branch[7].block[3].um_I.ena ;
 wire \top_I.branch[7].block[3].um_I.iw[10] ;
 wire \top_I.branch[7].block[3].um_I.iw[11] ;
 wire \top_I.branch[7].block[3].um_I.iw[12] ;
 wire \top_I.branch[7].block[3].um_I.iw[13] ;
 wire \top_I.branch[7].block[3].um_I.iw[14] ;
 wire \top_I.branch[7].block[3].um_I.iw[15] ;
 wire \top_I.branch[7].block[3].um_I.iw[16] ;
 wire \top_I.branch[7].block[3].um_I.iw[17] ;
 wire \top_I.branch[7].block[3].um_I.iw[1] ;
 wire \top_I.branch[7].block[3].um_I.iw[2] ;
 wire \top_I.branch[7].block[3].um_I.iw[3] ;
 wire \top_I.branch[7].block[3].um_I.iw[4] ;
 wire \top_I.branch[7].block[3].um_I.iw[5] ;
 wire \top_I.branch[7].block[3].um_I.iw[6] ;
 wire \top_I.branch[7].block[3].um_I.iw[7] ;
 wire \top_I.branch[7].block[3].um_I.iw[8] ;
 wire \top_I.branch[7].block[3].um_I.iw[9] ;
 wire \top_I.branch[7].block[3].um_I.k_zero ;
 wire \top_I.branch[7].block[3].um_I.pg_vdd ;
 wire \top_I.branch[7].block[4].um_I.ana[2] ;
 wire \top_I.branch[7].block[4].um_I.ana[3] ;
 wire \top_I.branch[7].block[4].um_I.ana[4] ;
 wire \top_I.branch[7].block[4].um_I.ana[5] ;
 wire \top_I.branch[7].block[4].um_I.ana[6] ;
 wire \top_I.branch[7].block[4].um_I.ana[7] ;
 wire \top_I.branch[7].block[4].um_I.clk ;
 wire \top_I.branch[7].block[4].um_I.ena ;
 wire \top_I.branch[7].block[4].um_I.iw[10] ;
 wire \top_I.branch[7].block[4].um_I.iw[11] ;
 wire \top_I.branch[7].block[4].um_I.iw[12] ;
 wire \top_I.branch[7].block[4].um_I.iw[13] ;
 wire \top_I.branch[7].block[4].um_I.iw[14] ;
 wire \top_I.branch[7].block[4].um_I.iw[15] ;
 wire \top_I.branch[7].block[4].um_I.iw[16] ;
 wire \top_I.branch[7].block[4].um_I.iw[17] ;
 wire \top_I.branch[7].block[4].um_I.iw[1] ;
 wire \top_I.branch[7].block[4].um_I.iw[2] ;
 wire \top_I.branch[7].block[4].um_I.iw[3] ;
 wire \top_I.branch[7].block[4].um_I.iw[4] ;
 wire \top_I.branch[7].block[4].um_I.iw[5] ;
 wire \top_I.branch[7].block[4].um_I.iw[6] ;
 wire \top_I.branch[7].block[4].um_I.iw[7] ;
 wire \top_I.branch[7].block[4].um_I.iw[8] ;
 wire \top_I.branch[7].block[4].um_I.iw[9] ;
 wire \top_I.branch[7].block[4].um_I.k_zero ;
 wire \top_I.branch[7].block[4].um_I.pg_vdd ;
 wire \top_I.branch[7].block[5].um_I.ana[2] ;
 wire \top_I.branch[7].block[5].um_I.ana[3] ;
 wire \top_I.branch[7].block[5].um_I.ana[4] ;
 wire \top_I.branch[7].block[5].um_I.ana[5] ;
 wire \top_I.branch[7].block[5].um_I.ana[6] ;
 wire \top_I.branch[7].block[5].um_I.ana[7] ;
 wire \top_I.branch[7].block[5].um_I.clk ;
 wire \top_I.branch[7].block[5].um_I.ena ;
 wire \top_I.branch[7].block[5].um_I.iw[10] ;
 wire \top_I.branch[7].block[5].um_I.iw[11] ;
 wire \top_I.branch[7].block[5].um_I.iw[12] ;
 wire \top_I.branch[7].block[5].um_I.iw[13] ;
 wire \top_I.branch[7].block[5].um_I.iw[14] ;
 wire \top_I.branch[7].block[5].um_I.iw[15] ;
 wire \top_I.branch[7].block[5].um_I.iw[16] ;
 wire \top_I.branch[7].block[5].um_I.iw[17] ;
 wire \top_I.branch[7].block[5].um_I.iw[1] ;
 wire \top_I.branch[7].block[5].um_I.iw[2] ;
 wire \top_I.branch[7].block[5].um_I.iw[3] ;
 wire \top_I.branch[7].block[5].um_I.iw[4] ;
 wire \top_I.branch[7].block[5].um_I.iw[5] ;
 wire \top_I.branch[7].block[5].um_I.iw[6] ;
 wire \top_I.branch[7].block[5].um_I.iw[7] ;
 wire \top_I.branch[7].block[5].um_I.iw[8] ;
 wire \top_I.branch[7].block[5].um_I.iw[9] ;
 wire \top_I.branch[7].block[5].um_I.k_zero ;
 wire \top_I.branch[7].block[5].um_I.pg_vdd ;
 wire \top_I.branch[7].block[6].um_I.ana[2] ;
 wire \top_I.branch[7].block[6].um_I.ana[3] ;
 wire \top_I.branch[7].block[6].um_I.ana[4] ;
 wire \top_I.branch[7].block[6].um_I.ana[5] ;
 wire \top_I.branch[7].block[6].um_I.ana[6] ;
 wire \top_I.branch[7].block[6].um_I.ana[7] ;
 wire \top_I.branch[7].block[6].um_I.clk ;
 wire \top_I.branch[7].block[6].um_I.ena ;
 wire \top_I.branch[7].block[6].um_I.iw[10] ;
 wire \top_I.branch[7].block[6].um_I.iw[11] ;
 wire \top_I.branch[7].block[6].um_I.iw[12] ;
 wire \top_I.branch[7].block[6].um_I.iw[13] ;
 wire \top_I.branch[7].block[6].um_I.iw[14] ;
 wire \top_I.branch[7].block[6].um_I.iw[15] ;
 wire \top_I.branch[7].block[6].um_I.iw[16] ;
 wire \top_I.branch[7].block[6].um_I.iw[17] ;
 wire \top_I.branch[7].block[6].um_I.iw[1] ;
 wire \top_I.branch[7].block[6].um_I.iw[2] ;
 wire \top_I.branch[7].block[6].um_I.iw[3] ;
 wire \top_I.branch[7].block[6].um_I.iw[4] ;
 wire \top_I.branch[7].block[6].um_I.iw[5] ;
 wire \top_I.branch[7].block[6].um_I.iw[6] ;
 wire \top_I.branch[7].block[6].um_I.iw[7] ;
 wire \top_I.branch[7].block[6].um_I.iw[8] ;
 wire \top_I.branch[7].block[6].um_I.iw[9] ;
 wire \top_I.branch[7].block[6].um_I.k_zero ;
 wire \top_I.branch[7].block[6].um_I.pg_vdd ;
 wire \top_I.branch[7].block[7].um_I.ana[2] ;
 wire \top_I.branch[7].block[7].um_I.ana[3] ;
 wire \top_I.branch[7].block[7].um_I.ana[4] ;
 wire \top_I.branch[7].block[7].um_I.ana[5] ;
 wire \top_I.branch[7].block[7].um_I.ana[6] ;
 wire \top_I.branch[7].block[7].um_I.ana[7] ;
 wire \top_I.branch[7].block[7].um_I.clk ;
 wire \top_I.branch[7].block[7].um_I.ena ;
 wire \top_I.branch[7].block[7].um_I.iw[10] ;
 wire \top_I.branch[7].block[7].um_I.iw[11] ;
 wire \top_I.branch[7].block[7].um_I.iw[12] ;
 wire \top_I.branch[7].block[7].um_I.iw[13] ;
 wire \top_I.branch[7].block[7].um_I.iw[14] ;
 wire \top_I.branch[7].block[7].um_I.iw[15] ;
 wire \top_I.branch[7].block[7].um_I.iw[16] ;
 wire \top_I.branch[7].block[7].um_I.iw[17] ;
 wire \top_I.branch[7].block[7].um_I.iw[1] ;
 wire \top_I.branch[7].block[7].um_I.iw[2] ;
 wire \top_I.branch[7].block[7].um_I.iw[3] ;
 wire \top_I.branch[7].block[7].um_I.iw[4] ;
 wire \top_I.branch[7].block[7].um_I.iw[5] ;
 wire \top_I.branch[7].block[7].um_I.iw[6] ;
 wire \top_I.branch[7].block[7].um_I.iw[7] ;
 wire \top_I.branch[7].block[7].um_I.iw[8] ;
 wire \top_I.branch[7].block[7].um_I.iw[9] ;
 wire \top_I.branch[7].block[7].um_I.k_zero ;
 wire \top_I.branch[7].block[7].um_I.pg_vdd ;
 wire \top_I.branch[7].block[8].um_I.ana[2] ;
 wire \top_I.branch[7].block[8].um_I.ana[3] ;
 wire \top_I.branch[7].block[8].um_I.ana[4] ;
 wire \top_I.branch[7].block[8].um_I.ana[5] ;
 wire \top_I.branch[7].block[8].um_I.ana[6] ;
 wire \top_I.branch[7].block[8].um_I.ana[7] ;
 wire \top_I.branch[7].block[8].um_I.clk ;
 wire \top_I.branch[7].block[8].um_I.ena ;
 wire \top_I.branch[7].block[8].um_I.iw[10] ;
 wire \top_I.branch[7].block[8].um_I.iw[11] ;
 wire \top_I.branch[7].block[8].um_I.iw[12] ;
 wire \top_I.branch[7].block[8].um_I.iw[13] ;
 wire \top_I.branch[7].block[8].um_I.iw[14] ;
 wire \top_I.branch[7].block[8].um_I.iw[15] ;
 wire \top_I.branch[7].block[8].um_I.iw[16] ;
 wire \top_I.branch[7].block[8].um_I.iw[17] ;
 wire \top_I.branch[7].block[8].um_I.iw[1] ;
 wire \top_I.branch[7].block[8].um_I.iw[2] ;
 wire \top_I.branch[7].block[8].um_I.iw[3] ;
 wire \top_I.branch[7].block[8].um_I.iw[4] ;
 wire \top_I.branch[7].block[8].um_I.iw[5] ;
 wire \top_I.branch[7].block[8].um_I.iw[6] ;
 wire \top_I.branch[7].block[8].um_I.iw[7] ;
 wire \top_I.branch[7].block[8].um_I.iw[8] ;
 wire \top_I.branch[7].block[8].um_I.iw[9] ;
 wire \top_I.branch[7].block[8].um_I.k_zero ;
 wire \top_I.branch[7].block[8].um_I.pg_vdd ;
 wire \top_I.branch[7].block[9].um_I.ana[2] ;
 wire \top_I.branch[7].block[9].um_I.ana[3] ;
 wire \top_I.branch[7].block[9].um_I.ana[4] ;
 wire \top_I.branch[7].block[9].um_I.ana[5] ;
 wire \top_I.branch[7].block[9].um_I.ana[6] ;
 wire \top_I.branch[7].block[9].um_I.ana[7] ;
 wire \top_I.branch[7].block[9].um_I.clk ;
 wire \top_I.branch[7].block[9].um_I.ena ;
 wire \top_I.branch[7].block[9].um_I.iw[10] ;
 wire \top_I.branch[7].block[9].um_I.iw[11] ;
 wire \top_I.branch[7].block[9].um_I.iw[12] ;
 wire \top_I.branch[7].block[9].um_I.iw[13] ;
 wire \top_I.branch[7].block[9].um_I.iw[14] ;
 wire \top_I.branch[7].block[9].um_I.iw[15] ;
 wire \top_I.branch[7].block[9].um_I.iw[16] ;
 wire \top_I.branch[7].block[9].um_I.iw[17] ;
 wire \top_I.branch[7].block[9].um_I.iw[1] ;
 wire \top_I.branch[7].block[9].um_I.iw[2] ;
 wire \top_I.branch[7].block[9].um_I.iw[3] ;
 wire \top_I.branch[7].block[9].um_I.iw[4] ;
 wire \top_I.branch[7].block[9].um_I.iw[5] ;
 wire \top_I.branch[7].block[9].um_I.iw[6] ;
 wire \top_I.branch[7].block[9].um_I.iw[7] ;
 wire \top_I.branch[7].block[9].um_I.iw[8] ;
 wire \top_I.branch[7].block[9].um_I.iw[9] ;
 wire \top_I.branch[7].block[9].um_I.k_zero ;
 wire \top_I.branch[7].block[9].um_I.pg_vdd ;
 wire \top_I.branch[7].l_addr[0] ;
 wire \top_I.branch[7].l_addr[2] ;
 wire \top_I.branch[8].block[0].um_I.ana[2] ;
 wire \top_I.branch[8].block[0].um_I.ana[3] ;
 wire \top_I.branch[8].block[0].um_I.ana[4] ;
 wire \top_I.branch[8].block[0].um_I.ana[5] ;
 wire \top_I.branch[8].block[0].um_I.ana[6] ;
 wire \top_I.branch[8].block[0].um_I.ana[7] ;
 wire \top_I.branch[8].block[0].um_I.clk ;
 wire \top_I.branch[8].block[0].um_I.ena ;
 wire \top_I.branch[8].block[0].um_I.iw[10] ;
 wire \top_I.branch[8].block[0].um_I.iw[11] ;
 wire \top_I.branch[8].block[0].um_I.iw[12] ;
 wire \top_I.branch[8].block[0].um_I.iw[13] ;
 wire \top_I.branch[8].block[0].um_I.iw[14] ;
 wire \top_I.branch[8].block[0].um_I.iw[15] ;
 wire \top_I.branch[8].block[0].um_I.iw[16] ;
 wire \top_I.branch[8].block[0].um_I.iw[17] ;
 wire \top_I.branch[8].block[0].um_I.iw[1] ;
 wire \top_I.branch[8].block[0].um_I.iw[2] ;
 wire \top_I.branch[8].block[0].um_I.iw[3] ;
 wire \top_I.branch[8].block[0].um_I.iw[4] ;
 wire \top_I.branch[8].block[0].um_I.iw[5] ;
 wire \top_I.branch[8].block[0].um_I.iw[6] ;
 wire \top_I.branch[8].block[0].um_I.iw[7] ;
 wire \top_I.branch[8].block[0].um_I.iw[8] ;
 wire \top_I.branch[8].block[0].um_I.iw[9] ;
 wire \top_I.branch[8].block[0].um_I.k_zero ;
 wire \top_I.branch[8].block[0].um_I.pg_vdd ;
 wire \top_I.branch[8].block[10].um_I.ana[2] ;
 wire \top_I.branch[8].block[10].um_I.ana[3] ;
 wire \top_I.branch[8].block[10].um_I.ana[4] ;
 wire \top_I.branch[8].block[10].um_I.ana[5] ;
 wire \top_I.branch[8].block[10].um_I.ana[6] ;
 wire \top_I.branch[8].block[10].um_I.ana[7] ;
 wire \top_I.branch[8].block[10].um_I.clk ;
 wire \top_I.branch[8].block[10].um_I.ena ;
 wire \top_I.branch[8].block[10].um_I.iw[10] ;
 wire \top_I.branch[8].block[10].um_I.iw[11] ;
 wire \top_I.branch[8].block[10].um_I.iw[12] ;
 wire \top_I.branch[8].block[10].um_I.iw[13] ;
 wire \top_I.branch[8].block[10].um_I.iw[14] ;
 wire \top_I.branch[8].block[10].um_I.iw[15] ;
 wire \top_I.branch[8].block[10].um_I.iw[16] ;
 wire \top_I.branch[8].block[10].um_I.iw[17] ;
 wire \top_I.branch[8].block[10].um_I.iw[1] ;
 wire \top_I.branch[8].block[10].um_I.iw[2] ;
 wire \top_I.branch[8].block[10].um_I.iw[3] ;
 wire \top_I.branch[8].block[10].um_I.iw[4] ;
 wire \top_I.branch[8].block[10].um_I.iw[5] ;
 wire \top_I.branch[8].block[10].um_I.iw[6] ;
 wire \top_I.branch[8].block[10].um_I.iw[7] ;
 wire \top_I.branch[8].block[10].um_I.iw[8] ;
 wire \top_I.branch[8].block[10].um_I.iw[9] ;
 wire \top_I.branch[8].block[10].um_I.k_zero ;
 wire \top_I.branch[8].block[10].um_I.pg_vdd ;
 wire \top_I.branch[8].block[11].um_I.ana[2] ;
 wire \top_I.branch[8].block[11].um_I.ana[3] ;
 wire \top_I.branch[8].block[11].um_I.ana[4] ;
 wire \top_I.branch[8].block[11].um_I.ana[5] ;
 wire \top_I.branch[8].block[11].um_I.ana[6] ;
 wire \top_I.branch[8].block[11].um_I.ana[7] ;
 wire \top_I.branch[8].block[11].um_I.clk ;
 wire \top_I.branch[8].block[11].um_I.ena ;
 wire \top_I.branch[8].block[11].um_I.iw[10] ;
 wire \top_I.branch[8].block[11].um_I.iw[11] ;
 wire \top_I.branch[8].block[11].um_I.iw[12] ;
 wire \top_I.branch[8].block[11].um_I.iw[13] ;
 wire \top_I.branch[8].block[11].um_I.iw[14] ;
 wire \top_I.branch[8].block[11].um_I.iw[15] ;
 wire \top_I.branch[8].block[11].um_I.iw[16] ;
 wire \top_I.branch[8].block[11].um_I.iw[17] ;
 wire \top_I.branch[8].block[11].um_I.iw[1] ;
 wire \top_I.branch[8].block[11].um_I.iw[2] ;
 wire \top_I.branch[8].block[11].um_I.iw[3] ;
 wire \top_I.branch[8].block[11].um_I.iw[4] ;
 wire \top_I.branch[8].block[11].um_I.iw[5] ;
 wire \top_I.branch[8].block[11].um_I.iw[6] ;
 wire \top_I.branch[8].block[11].um_I.iw[7] ;
 wire \top_I.branch[8].block[11].um_I.iw[8] ;
 wire \top_I.branch[8].block[11].um_I.iw[9] ;
 wire \top_I.branch[8].block[11].um_I.k_zero ;
 wire \top_I.branch[8].block[11].um_I.pg_vdd ;
 wire \top_I.branch[8].block[12].um_I.ana[2] ;
 wire \top_I.branch[8].block[12].um_I.ana[3] ;
 wire \top_I.branch[8].block[12].um_I.ana[4] ;
 wire \top_I.branch[8].block[12].um_I.ana[5] ;
 wire \top_I.branch[8].block[12].um_I.ana[6] ;
 wire \top_I.branch[8].block[12].um_I.ana[7] ;
 wire \top_I.branch[8].block[12].um_I.clk ;
 wire \top_I.branch[8].block[12].um_I.ena ;
 wire \top_I.branch[8].block[12].um_I.iw[10] ;
 wire \top_I.branch[8].block[12].um_I.iw[11] ;
 wire \top_I.branch[8].block[12].um_I.iw[12] ;
 wire \top_I.branch[8].block[12].um_I.iw[13] ;
 wire \top_I.branch[8].block[12].um_I.iw[14] ;
 wire \top_I.branch[8].block[12].um_I.iw[15] ;
 wire \top_I.branch[8].block[12].um_I.iw[16] ;
 wire \top_I.branch[8].block[12].um_I.iw[17] ;
 wire \top_I.branch[8].block[12].um_I.iw[1] ;
 wire \top_I.branch[8].block[12].um_I.iw[2] ;
 wire \top_I.branch[8].block[12].um_I.iw[3] ;
 wire \top_I.branch[8].block[12].um_I.iw[4] ;
 wire \top_I.branch[8].block[12].um_I.iw[5] ;
 wire \top_I.branch[8].block[12].um_I.iw[6] ;
 wire \top_I.branch[8].block[12].um_I.iw[7] ;
 wire \top_I.branch[8].block[12].um_I.iw[8] ;
 wire \top_I.branch[8].block[12].um_I.iw[9] ;
 wire \top_I.branch[8].block[12].um_I.k_zero ;
 wire \top_I.branch[8].block[12].um_I.pg_vdd ;
 wire \top_I.branch[8].block[13].um_I.ana[2] ;
 wire \top_I.branch[8].block[13].um_I.ana[3] ;
 wire \top_I.branch[8].block[13].um_I.ana[4] ;
 wire \top_I.branch[8].block[13].um_I.ana[5] ;
 wire \top_I.branch[8].block[13].um_I.ana[6] ;
 wire \top_I.branch[8].block[13].um_I.ana[7] ;
 wire \top_I.branch[8].block[13].um_I.clk ;
 wire \top_I.branch[8].block[13].um_I.ena ;
 wire \top_I.branch[8].block[13].um_I.iw[10] ;
 wire \top_I.branch[8].block[13].um_I.iw[11] ;
 wire \top_I.branch[8].block[13].um_I.iw[12] ;
 wire \top_I.branch[8].block[13].um_I.iw[13] ;
 wire \top_I.branch[8].block[13].um_I.iw[14] ;
 wire \top_I.branch[8].block[13].um_I.iw[15] ;
 wire \top_I.branch[8].block[13].um_I.iw[16] ;
 wire \top_I.branch[8].block[13].um_I.iw[17] ;
 wire \top_I.branch[8].block[13].um_I.iw[1] ;
 wire \top_I.branch[8].block[13].um_I.iw[2] ;
 wire \top_I.branch[8].block[13].um_I.iw[3] ;
 wire \top_I.branch[8].block[13].um_I.iw[4] ;
 wire \top_I.branch[8].block[13].um_I.iw[5] ;
 wire \top_I.branch[8].block[13].um_I.iw[6] ;
 wire \top_I.branch[8].block[13].um_I.iw[7] ;
 wire \top_I.branch[8].block[13].um_I.iw[8] ;
 wire \top_I.branch[8].block[13].um_I.iw[9] ;
 wire \top_I.branch[8].block[13].um_I.k_zero ;
 wire \top_I.branch[8].block[13].um_I.pg_vdd ;
 wire \top_I.branch[8].block[14].um_I.ana[2] ;
 wire \top_I.branch[8].block[14].um_I.ana[3] ;
 wire \top_I.branch[8].block[14].um_I.ana[4] ;
 wire \top_I.branch[8].block[14].um_I.ana[5] ;
 wire \top_I.branch[8].block[14].um_I.ana[6] ;
 wire \top_I.branch[8].block[14].um_I.ana[7] ;
 wire \top_I.branch[8].block[14].um_I.clk ;
 wire \top_I.branch[8].block[14].um_I.ena ;
 wire \top_I.branch[8].block[14].um_I.iw[10] ;
 wire \top_I.branch[8].block[14].um_I.iw[11] ;
 wire \top_I.branch[8].block[14].um_I.iw[12] ;
 wire \top_I.branch[8].block[14].um_I.iw[13] ;
 wire \top_I.branch[8].block[14].um_I.iw[14] ;
 wire \top_I.branch[8].block[14].um_I.iw[15] ;
 wire \top_I.branch[8].block[14].um_I.iw[16] ;
 wire \top_I.branch[8].block[14].um_I.iw[17] ;
 wire \top_I.branch[8].block[14].um_I.iw[1] ;
 wire \top_I.branch[8].block[14].um_I.iw[2] ;
 wire \top_I.branch[8].block[14].um_I.iw[3] ;
 wire \top_I.branch[8].block[14].um_I.iw[4] ;
 wire \top_I.branch[8].block[14].um_I.iw[5] ;
 wire \top_I.branch[8].block[14].um_I.iw[6] ;
 wire \top_I.branch[8].block[14].um_I.iw[7] ;
 wire \top_I.branch[8].block[14].um_I.iw[8] ;
 wire \top_I.branch[8].block[14].um_I.iw[9] ;
 wire \top_I.branch[8].block[14].um_I.k_zero ;
 wire \top_I.branch[8].block[14].um_I.pg_vdd ;
 wire \top_I.branch[8].block[15].um_I.ana[2] ;
 wire \top_I.branch[8].block[15].um_I.ana[3] ;
 wire \top_I.branch[8].block[15].um_I.ana[4] ;
 wire \top_I.branch[8].block[15].um_I.ana[5] ;
 wire \top_I.branch[8].block[15].um_I.ana[6] ;
 wire \top_I.branch[8].block[15].um_I.ana[7] ;
 wire \top_I.branch[8].block[15].um_I.clk ;
 wire \top_I.branch[8].block[15].um_I.ena ;
 wire \top_I.branch[8].block[15].um_I.iw[10] ;
 wire \top_I.branch[8].block[15].um_I.iw[11] ;
 wire \top_I.branch[8].block[15].um_I.iw[12] ;
 wire \top_I.branch[8].block[15].um_I.iw[13] ;
 wire \top_I.branch[8].block[15].um_I.iw[14] ;
 wire \top_I.branch[8].block[15].um_I.iw[15] ;
 wire \top_I.branch[8].block[15].um_I.iw[16] ;
 wire \top_I.branch[8].block[15].um_I.iw[17] ;
 wire \top_I.branch[8].block[15].um_I.iw[1] ;
 wire \top_I.branch[8].block[15].um_I.iw[2] ;
 wire \top_I.branch[8].block[15].um_I.iw[3] ;
 wire \top_I.branch[8].block[15].um_I.iw[4] ;
 wire \top_I.branch[8].block[15].um_I.iw[5] ;
 wire \top_I.branch[8].block[15].um_I.iw[6] ;
 wire \top_I.branch[8].block[15].um_I.iw[7] ;
 wire \top_I.branch[8].block[15].um_I.iw[8] ;
 wire \top_I.branch[8].block[15].um_I.iw[9] ;
 wire \top_I.branch[8].block[15].um_I.k_zero ;
 wire \top_I.branch[8].block[15].um_I.pg_vdd ;
 wire \top_I.branch[8].block[1].um_I.ana[2] ;
 wire \top_I.branch[8].block[1].um_I.ana[3] ;
 wire \top_I.branch[8].block[1].um_I.ana[4] ;
 wire \top_I.branch[8].block[1].um_I.ana[5] ;
 wire \top_I.branch[8].block[1].um_I.ana[6] ;
 wire \top_I.branch[8].block[1].um_I.ana[7] ;
 wire \top_I.branch[8].block[1].um_I.clk ;
 wire \top_I.branch[8].block[1].um_I.ena ;
 wire \top_I.branch[8].block[1].um_I.iw[10] ;
 wire \top_I.branch[8].block[1].um_I.iw[11] ;
 wire \top_I.branch[8].block[1].um_I.iw[12] ;
 wire \top_I.branch[8].block[1].um_I.iw[13] ;
 wire \top_I.branch[8].block[1].um_I.iw[14] ;
 wire \top_I.branch[8].block[1].um_I.iw[15] ;
 wire \top_I.branch[8].block[1].um_I.iw[16] ;
 wire \top_I.branch[8].block[1].um_I.iw[17] ;
 wire \top_I.branch[8].block[1].um_I.iw[1] ;
 wire \top_I.branch[8].block[1].um_I.iw[2] ;
 wire \top_I.branch[8].block[1].um_I.iw[3] ;
 wire \top_I.branch[8].block[1].um_I.iw[4] ;
 wire \top_I.branch[8].block[1].um_I.iw[5] ;
 wire \top_I.branch[8].block[1].um_I.iw[6] ;
 wire \top_I.branch[8].block[1].um_I.iw[7] ;
 wire \top_I.branch[8].block[1].um_I.iw[8] ;
 wire \top_I.branch[8].block[1].um_I.iw[9] ;
 wire \top_I.branch[8].block[1].um_I.k_zero ;
 wire \top_I.branch[8].block[1].um_I.pg_vdd ;
 wire \top_I.branch[8].block[2].um_I.ana[2] ;
 wire \top_I.branch[8].block[2].um_I.ana[3] ;
 wire \top_I.branch[8].block[2].um_I.ana[4] ;
 wire \top_I.branch[8].block[2].um_I.ana[5] ;
 wire \top_I.branch[8].block[2].um_I.ana[6] ;
 wire \top_I.branch[8].block[2].um_I.ana[7] ;
 wire \top_I.branch[8].block[2].um_I.clk ;
 wire \top_I.branch[8].block[2].um_I.ena ;
 wire \top_I.branch[8].block[2].um_I.iw[10] ;
 wire \top_I.branch[8].block[2].um_I.iw[11] ;
 wire \top_I.branch[8].block[2].um_I.iw[12] ;
 wire \top_I.branch[8].block[2].um_I.iw[13] ;
 wire \top_I.branch[8].block[2].um_I.iw[14] ;
 wire \top_I.branch[8].block[2].um_I.iw[15] ;
 wire \top_I.branch[8].block[2].um_I.iw[16] ;
 wire \top_I.branch[8].block[2].um_I.iw[17] ;
 wire \top_I.branch[8].block[2].um_I.iw[1] ;
 wire \top_I.branch[8].block[2].um_I.iw[2] ;
 wire \top_I.branch[8].block[2].um_I.iw[3] ;
 wire \top_I.branch[8].block[2].um_I.iw[4] ;
 wire \top_I.branch[8].block[2].um_I.iw[5] ;
 wire \top_I.branch[8].block[2].um_I.iw[6] ;
 wire \top_I.branch[8].block[2].um_I.iw[7] ;
 wire \top_I.branch[8].block[2].um_I.iw[8] ;
 wire \top_I.branch[8].block[2].um_I.iw[9] ;
 wire \top_I.branch[8].block[2].um_I.k_zero ;
 wire \top_I.branch[8].block[2].um_I.pg_vdd ;
 wire \top_I.branch[8].block[3].um_I.ana[2] ;
 wire \top_I.branch[8].block[3].um_I.ana[3] ;
 wire \top_I.branch[8].block[3].um_I.ana[4] ;
 wire \top_I.branch[8].block[3].um_I.ana[5] ;
 wire \top_I.branch[8].block[3].um_I.ana[6] ;
 wire \top_I.branch[8].block[3].um_I.ana[7] ;
 wire \top_I.branch[8].block[3].um_I.clk ;
 wire \top_I.branch[8].block[3].um_I.ena ;
 wire \top_I.branch[8].block[3].um_I.iw[10] ;
 wire \top_I.branch[8].block[3].um_I.iw[11] ;
 wire \top_I.branch[8].block[3].um_I.iw[12] ;
 wire \top_I.branch[8].block[3].um_I.iw[13] ;
 wire \top_I.branch[8].block[3].um_I.iw[14] ;
 wire \top_I.branch[8].block[3].um_I.iw[15] ;
 wire \top_I.branch[8].block[3].um_I.iw[16] ;
 wire \top_I.branch[8].block[3].um_I.iw[17] ;
 wire \top_I.branch[8].block[3].um_I.iw[1] ;
 wire \top_I.branch[8].block[3].um_I.iw[2] ;
 wire \top_I.branch[8].block[3].um_I.iw[3] ;
 wire \top_I.branch[8].block[3].um_I.iw[4] ;
 wire \top_I.branch[8].block[3].um_I.iw[5] ;
 wire \top_I.branch[8].block[3].um_I.iw[6] ;
 wire \top_I.branch[8].block[3].um_I.iw[7] ;
 wire \top_I.branch[8].block[3].um_I.iw[8] ;
 wire \top_I.branch[8].block[3].um_I.iw[9] ;
 wire \top_I.branch[8].block[3].um_I.k_zero ;
 wire \top_I.branch[8].block[3].um_I.pg_vdd ;
 wire \top_I.branch[8].block[4].um_I.ana[2] ;
 wire \top_I.branch[8].block[4].um_I.ana[3] ;
 wire \top_I.branch[8].block[4].um_I.ana[4] ;
 wire \top_I.branch[8].block[4].um_I.ana[5] ;
 wire \top_I.branch[8].block[4].um_I.ana[6] ;
 wire \top_I.branch[8].block[4].um_I.ana[7] ;
 wire \top_I.branch[8].block[4].um_I.clk ;
 wire \top_I.branch[8].block[4].um_I.ena ;
 wire \top_I.branch[8].block[4].um_I.iw[10] ;
 wire \top_I.branch[8].block[4].um_I.iw[11] ;
 wire \top_I.branch[8].block[4].um_I.iw[12] ;
 wire \top_I.branch[8].block[4].um_I.iw[13] ;
 wire \top_I.branch[8].block[4].um_I.iw[14] ;
 wire \top_I.branch[8].block[4].um_I.iw[15] ;
 wire \top_I.branch[8].block[4].um_I.iw[16] ;
 wire \top_I.branch[8].block[4].um_I.iw[17] ;
 wire \top_I.branch[8].block[4].um_I.iw[1] ;
 wire \top_I.branch[8].block[4].um_I.iw[2] ;
 wire \top_I.branch[8].block[4].um_I.iw[3] ;
 wire \top_I.branch[8].block[4].um_I.iw[4] ;
 wire \top_I.branch[8].block[4].um_I.iw[5] ;
 wire \top_I.branch[8].block[4].um_I.iw[6] ;
 wire \top_I.branch[8].block[4].um_I.iw[7] ;
 wire \top_I.branch[8].block[4].um_I.iw[8] ;
 wire \top_I.branch[8].block[4].um_I.iw[9] ;
 wire \top_I.branch[8].block[4].um_I.k_zero ;
 wire \top_I.branch[8].block[4].um_I.pg_vdd ;
 wire \top_I.branch[8].block[5].um_I.ana[2] ;
 wire \top_I.branch[8].block[5].um_I.ana[3] ;
 wire \top_I.branch[8].block[5].um_I.ana[4] ;
 wire \top_I.branch[8].block[5].um_I.ana[5] ;
 wire \top_I.branch[8].block[5].um_I.ana[6] ;
 wire \top_I.branch[8].block[5].um_I.ana[7] ;
 wire \top_I.branch[8].block[5].um_I.clk ;
 wire \top_I.branch[8].block[5].um_I.ena ;
 wire \top_I.branch[8].block[5].um_I.iw[10] ;
 wire \top_I.branch[8].block[5].um_I.iw[11] ;
 wire \top_I.branch[8].block[5].um_I.iw[12] ;
 wire \top_I.branch[8].block[5].um_I.iw[13] ;
 wire \top_I.branch[8].block[5].um_I.iw[14] ;
 wire \top_I.branch[8].block[5].um_I.iw[15] ;
 wire \top_I.branch[8].block[5].um_I.iw[16] ;
 wire \top_I.branch[8].block[5].um_I.iw[17] ;
 wire \top_I.branch[8].block[5].um_I.iw[1] ;
 wire \top_I.branch[8].block[5].um_I.iw[2] ;
 wire \top_I.branch[8].block[5].um_I.iw[3] ;
 wire \top_I.branch[8].block[5].um_I.iw[4] ;
 wire \top_I.branch[8].block[5].um_I.iw[5] ;
 wire \top_I.branch[8].block[5].um_I.iw[6] ;
 wire \top_I.branch[8].block[5].um_I.iw[7] ;
 wire \top_I.branch[8].block[5].um_I.iw[8] ;
 wire \top_I.branch[8].block[5].um_I.iw[9] ;
 wire \top_I.branch[8].block[5].um_I.k_zero ;
 wire \top_I.branch[8].block[5].um_I.pg_vdd ;
 wire \top_I.branch[8].block[6].um_I.ana[2] ;
 wire \top_I.branch[8].block[6].um_I.ana[3] ;
 wire \top_I.branch[8].block[6].um_I.ana[4] ;
 wire \top_I.branch[8].block[6].um_I.ana[5] ;
 wire \top_I.branch[8].block[6].um_I.ana[6] ;
 wire \top_I.branch[8].block[6].um_I.ana[7] ;
 wire \top_I.branch[8].block[6].um_I.clk ;
 wire \top_I.branch[8].block[6].um_I.ena ;
 wire \top_I.branch[8].block[6].um_I.iw[10] ;
 wire \top_I.branch[8].block[6].um_I.iw[11] ;
 wire \top_I.branch[8].block[6].um_I.iw[12] ;
 wire \top_I.branch[8].block[6].um_I.iw[13] ;
 wire \top_I.branch[8].block[6].um_I.iw[14] ;
 wire \top_I.branch[8].block[6].um_I.iw[15] ;
 wire \top_I.branch[8].block[6].um_I.iw[16] ;
 wire \top_I.branch[8].block[6].um_I.iw[17] ;
 wire \top_I.branch[8].block[6].um_I.iw[1] ;
 wire \top_I.branch[8].block[6].um_I.iw[2] ;
 wire \top_I.branch[8].block[6].um_I.iw[3] ;
 wire \top_I.branch[8].block[6].um_I.iw[4] ;
 wire \top_I.branch[8].block[6].um_I.iw[5] ;
 wire \top_I.branch[8].block[6].um_I.iw[6] ;
 wire \top_I.branch[8].block[6].um_I.iw[7] ;
 wire \top_I.branch[8].block[6].um_I.iw[8] ;
 wire \top_I.branch[8].block[6].um_I.iw[9] ;
 wire \top_I.branch[8].block[6].um_I.k_zero ;
 wire \top_I.branch[8].block[6].um_I.pg_vdd ;
 wire \top_I.branch[8].block[7].um_I.ana[2] ;
 wire \top_I.branch[8].block[7].um_I.ana[3] ;
 wire \top_I.branch[8].block[7].um_I.ana[4] ;
 wire \top_I.branch[8].block[7].um_I.ana[5] ;
 wire \top_I.branch[8].block[7].um_I.ana[6] ;
 wire \top_I.branch[8].block[7].um_I.ana[7] ;
 wire \top_I.branch[8].block[7].um_I.clk ;
 wire \top_I.branch[8].block[7].um_I.ena ;
 wire \top_I.branch[8].block[7].um_I.iw[10] ;
 wire \top_I.branch[8].block[7].um_I.iw[11] ;
 wire \top_I.branch[8].block[7].um_I.iw[12] ;
 wire \top_I.branch[8].block[7].um_I.iw[13] ;
 wire \top_I.branch[8].block[7].um_I.iw[14] ;
 wire \top_I.branch[8].block[7].um_I.iw[15] ;
 wire \top_I.branch[8].block[7].um_I.iw[16] ;
 wire \top_I.branch[8].block[7].um_I.iw[17] ;
 wire \top_I.branch[8].block[7].um_I.iw[1] ;
 wire \top_I.branch[8].block[7].um_I.iw[2] ;
 wire \top_I.branch[8].block[7].um_I.iw[3] ;
 wire \top_I.branch[8].block[7].um_I.iw[4] ;
 wire \top_I.branch[8].block[7].um_I.iw[5] ;
 wire \top_I.branch[8].block[7].um_I.iw[6] ;
 wire \top_I.branch[8].block[7].um_I.iw[7] ;
 wire \top_I.branch[8].block[7].um_I.iw[8] ;
 wire \top_I.branch[8].block[7].um_I.iw[9] ;
 wire \top_I.branch[8].block[7].um_I.k_zero ;
 wire \top_I.branch[8].block[7].um_I.pg_vdd ;
 wire \top_I.branch[8].block[8].um_I.ana[2] ;
 wire \top_I.branch[8].block[8].um_I.ana[3] ;
 wire \top_I.branch[8].block[8].um_I.ana[4] ;
 wire \top_I.branch[8].block[8].um_I.ana[5] ;
 wire \top_I.branch[8].block[8].um_I.ana[6] ;
 wire \top_I.branch[8].block[8].um_I.ana[7] ;
 wire \top_I.branch[8].block[8].um_I.clk ;
 wire \top_I.branch[8].block[8].um_I.ena ;
 wire \top_I.branch[8].block[8].um_I.iw[10] ;
 wire \top_I.branch[8].block[8].um_I.iw[11] ;
 wire \top_I.branch[8].block[8].um_I.iw[12] ;
 wire \top_I.branch[8].block[8].um_I.iw[13] ;
 wire \top_I.branch[8].block[8].um_I.iw[14] ;
 wire \top_I.branch[8].block[8].um_I.iw[15] ;
 wire \top_I.branch[8].block[8].um_I.iw[16] ;
 wire \top_I.branch[8].block[8].um_I.iw[17] ;
 wire \top_I.branch[8].block[8].um_I.iw[1] ;
 wire \top_I.branch[8].block[8].um_I.iw[2] ;
 wire \top_I.branch[8].block[8].um_I.iw[3] ;
 wire \top_I.branch[8].block[8].um_I.iw[4] ;
 wire \top_I.branch[8].block[8].um_I.iw[5] ;
 wire \top_I.branch[8].block[8].um_I.iw[6] ;
 wire \top_I.branch[8].block[8].um_I.iw[7] ;
 wire \top_I.branch[8].block[8].um_I.iw[8] ;
 wire \top_I.branch[8].block[8].um_I.iw[9] ;
 wire \top_I.branch[8].block[8].um_I.k_zero ;
 wire \top_I.branch[8].block[8].um_I.pg_vdd ;
 wire \top_I.branch[8].block[9].um_I.ana[2] ;
 wire \top_I.branch[8].block[9].um_I.ana[3] ;
 wire \top_I.branch[8].block[9].um_I.ana[4] ;
 wire \top_I.branch[8].block[9].um_I.ana[5] ;
 wire \top_I.branch[8].block[9].um_I.ana[6] ;
 wire \top_I.branch[8].block[9].um_I.ana[7] ;
 wire \top_I.branch[8].block[9].um_I.clk ;
 wire \top_I.branch[8].block[9].um_I.ena ;
 wire \top_I.branch[8].block[9].um_I.iw[10] ;
 wire \top_I.branch[8].block[9].um_I.iw[11] ;
 wire \top_I.branch[8].block[9].um_I.iw[12] ;
 wire \top_I.branch[8].block[9].um_I.iw[13] ;
 wire \top_I.branch[8].block[9].um_I.iw[14] ;
 wire \top_I.branch[8].block[9].um_I.iw[15] ;
 wire \top_I.branch[8].block[9].um_I.iw[16] ;
 wire \top_I.branch[8].block[9].um_I.iw[17] ;
 wire \top_I.branch[8].block[9].um_I.iw[1] ;
 wire \top_I.branch[8].block[9].um_I.iw[2] ;
 wire \top_I.branch[8].block[9].um_I.iw[3] ;
 wire \top_I.branch[8].block[9].um_I.iw[4] ;
 wire \top_I.branch[8].block[9].um_I.iw[5] ;
 wire \top_I.branch[8].block[9].um_I.iw[6] ;
 wire \top_I.branch[8].block[9].um_I.iw[7] ;
 wire \top_I.branch[8].block[9].um_I.iw[8] ;
 wire \top_I.branch[8].block[9].um_I.iw[9] ;
 wire \top_I.branch[8].block[9].um_I.k_zero ;
 wire \top_I.branch[8].block[9].um_I.pg_vdd ;
 wire \top_I.branch[8].l_addr[0] ;
 wire \top_I.branch[8].l_addr[2] ;
 wire \top_I.branch[9].block[0].um_I.ana[2] ;
 wire \top_I.branch[9].block[0].um_I.ana[3] ;
 wire \top_I.branch[9].block[0].um_I.ana[4] ;
 wire \top_I.branch[9].block[0].um_I.ana[5] ;
 wire \top_I.branch[9].block[0].um_I.ana[6] ;
 wire \top_I.branch[9].block[0].um_I.ana[7] ;
 wire \top_I.branch[9].block[0].um_I.clk ;
 wire \top_I.branch[9].block[0].um_I.ena ;
 wire \top_I.branch[9].block[0].um_I.iw[10] ;
 wire \top_I.branch[9].block[0].um_I.iw[11] ;
 wire \top_I.branch[9].block[0].um_I.iw[12] ;
 wire \top_I.branch[9].block[0].um_I.iw[13] ;
 wire \top_I.branch[9].block[0].um_I.iw[14] ;
 wire \top_I.branch[9].block[0].um_I.iw[15] ;
 wire \top_I.branch[9].block[0].um_I.iw[16] ;
 wire \top_I.branch[9].block[0].um_I.iw[17] ;
 wire \top_I.branch[9].block[0].um_I.iw[1] ;
 wire \top_I.branch[9].block[0].um_I.iw[2] ;
 wire \top_I.branch[9].block[0].um_I.iw[3] ;
 wire \top_I.branch[9].block[0].um_I.iw[4] ;
 wire \top_I.branch[9].block[0].um_I.iw[5] ;
 wire \top_I.branch[9].block[0].um_I.iw[6] ;
 wire \top_I.branch[9].block[0].um_I.iw[7] ;
 wire \top_I.branch[9].block[0].um_I.iw[8] ;
 wire \top_I.branch[9].block[0].um_I.iw[9] ;
 wire \top_I.branch[9].block[0].um_I.k_zero ;
 wire \top_I.branch[9].block[0].um_I.pg_vdd ;
 wire \top_I.branch[9].block[10].um_I.ana[2] ;
 wire \top_I.branch[9].block[10].um_I.ana[3] ;
 wire \top_I.branch[9].block[10].um_I.ana[4] ;
 wire \top_I.branch[9].block[10].um_I.ana[5] ;
 wire \top_I.branch[9].block[10].um_I.ana[6] ;
 wire \top_I.branch[9].block[10].um_I.ana[7] ;
 wire \top_I.branch[9].block[10].um_I.clk ;
 wire \top_I.branch[9].block[10].um_I.ena ;
 wire \top_I.branch[9].block[10].um_I.iw[10] ;
 wire \top_I.branch[9].block[10].um_I.iw[11] ;
 wire \top_I.branch[9].block[10].um_I.iw[12] ;
 wire \top_I.branch[9].block[10].um_I.iw[13] ;
 wire \top_I.branch[9].block[10].um_I.iw[14] ;
 wire \top_I.branch[9].block[10].um_I.iw[15] ;
 wire \top_I.branch[9].block[10].um_I.iw[16] ;
 wire \top_I.branch[9].block[10].um_I.iw[17] ;
 wire \top_I.branch[9].block[10].um_I.iw[1] ;
 wire \top_I.branch[9].block[10].um_I.iw[2] ;
 wire \top_I.branch[9].block[10].um_I.iw[3] ;
 wire \top_I.branch[9].block[10].um_I.iw[4] ;
 wire \top_I.branch[9].block[10].um_I.iw[5] ;
 wire \top_I.branch[9].block[10].um_I.iw[6] ;
 wire \top_I.branch[9].block[10].um_I.iw[7] ;
 wire \top_I.branch[9].block[10].um_I.iw[8] ;
 wire \top_I.branch[9].block[10].um_I.iw[9] ;
 wire \top_I.branch[9].block[10].um_I.k_zero ;
 wire \top_I.branch[9].block[10].um_I.pg_vdd ;
 wire \top_I.branch[9].block[11].um_I.ana[2] ;
 wire \top_I.branch[9].block[11].um_I.ana[3] ;
 wire \top_I.branch[9].block[11].um_I.ana[4] ;
 wire \top_I.branch[9].block[11].um_I.ana[5] ;
 wire \top_I.branch[9].block[11].um_I.ana[6] ;
 wire \top_I.branch[9].block[11].um_I.ana[7] ;
 wire \top_I.branch[9].block[11].um_I.clk ;
 wire \top_I.branch[9].block[11].um_I.ena ;
 wire \top_I.branch[9].block[11].um_I.iw[10] ;
 wire \top_I.branch[9].block[11].um_I.iw[11] ;
 wire \top_I.branch[9].block[11].um_I.iw[12] ;
 wire \top_I.branch[9].block[11].um_I.iw[13] ;
 wire \top_I.branch[9].block[11].um_I.iw[14] ;
 wire \top_I.branch[9].block[11].um_I.iw[15] ;
 wire \top_I.branch[9].block[11].um_I.iw[16] ;
 wire \top_I.branch[9].block[11].um_I.iw[17] ;
 wire \top_I.branch[9].block[11].um_I.iw[1] ;
 wire \top_I.branch[9].block[11].um_I.iw[2] ;
 wire \top_I.branch[9].block[11].um_I.iw[3] ;
 wire \top_I.branch[9].block[11].um_I.iw[4] ;
 wire \top_I.branch[9].block[11].um_I.iw[5] ;
 wire \top_I.branch[9].block[11].um_I.iw[6] ;
 wire \top_I.branch[9].block[11].um_I.iw[7] ;
 wire \top_I.branch[9].block[11].um_I.iw[8] ;
 wire \top_I.branch[9].block[11].um_I.iw[9] ;
 wire \top_I.branch[9].block[11].um_I.k_zero ;
 wire \top_I.branch[9].block[11].um_I.pg_vdd ;
 wire \top_I.branch[9].block[12].um_I.ana[2] ;
 wire \top_I.branch[9].block[12].um_I.ana[3] ;
 wire \top_I.branch[9].block[12].um_I.ana[4] ;
 wire \top_I.branch[9].block[12].um_I.ana[5] ;
 wire \top_I.branch[9].block[12].um_I.ana[6] ;
 wire \top_I.branch[9].block[12].um_I.ana[7] ;
 wire \top_I.branch[9].block[12].um_I.clk ;
 wire \top_I.branch[9].block[12].um_I.ena ;
 wire \top_I.branch[9].block[12].um_I.iw[10] ;
 wire \top_I.branch[9].block[12].um_I.iw[11] ;
 wire \top_I.branch[9].block[12].um_I.iw[12] ;
 wire \top_I.branch[9].block[12].um_I.iw[13] ;
 wire \top_I.branch[9].block[12].um_I.iw[14] ;
 wire \top_I.branch[9].block[12].um_I.iw[15] ;
 wire \top_I.branch[9].block[12].um_I.iw[16] ;
 wire \top_I.branch[9].block[12].um_I.iw[17] ;
 wire \top_I.branch[9].block[12].um_I.iw[1] ;
 wire \top_I.branch[9].block[12].um_I.iw[2] ;
 wire \top_I.branch[9].block[12].um_I.iw[3] ;
 wire \top_I.branch[9].block[12].um_I.iw[4] ;
 wire \top_I.branch[9].block[12].um_I.iw[5] ;
 wire \top_I.branch[9].block[12].um_I.iw[6] ;
 wire \top_I.branch[9].block[12].um_I.iw[7] ;
 wire \top_I.branch[9].block[12].um_I.iw[8] ;
 wire \top_I.branch[9].block[12].um_I.iw[9] ;
 wire \top_I.branch[9].block[12].um_I.k_zero ;
 wire \top_I.branch[9].block[12].um_I.pg_vdd ;
 wire \top_I.branch[9].block[13].um_I.ana[2] ;
 wire \top_I.branch[9].block[13].um_I.ana[3] ;
 wire \top_I.branch[9].block[13].um_I.ana[4] ;
 wire \top_I.branch[9].block[13].um_I.ana[5] ;
 wire \top_I.branch[9].block[13].um_I.ana[6] ;
 wire \top_I.branch[9].block[13].um_I.ana[7] ;
 wire \top_I.branch[9].block[13].um_I.clk ;
 wire \top_I.branch[9].block[13].um_I.ena ;
 wire \top_I.branch[9].block[13].um_I.iw[10] ;
 wire \top_I.branch[9].block[13].um_I.iw[11] ;
 wire \top_I.branch[9].block[13].um_I.iw[12] ;
 wire \top_I.branch[9].block[13].um_I.iw[13] ;
 wire \top_I.branch[9].block[13].um_I.iw[14] ;
 wire \top_I.branch[9].block[13].um_I.iw[15] ;
 wire \top_I.branch[9].block[13].um_I.iw[16] ;
 wire \top_I.branch[9].block[13].um_I.iw[17] ;
 wire \top_I.branch[9].block[13].um_I.iw[1] ;
 wire \top_I.branch[9].block[13].um_I.iw[2] ;
 wire \top_I.branch[9].block[13].um_I.iw[3] ;
 wire \top_I.branch[9].block[13].um_I.iw[4] ;
 wire \top_I.branch[9].block[13].um_I.iw[5] ;
 wire \top_I.branch[9].block[13].um_I.iw[6] ;
 wire \top_I.branch[9].block[13].um_I.iw[7] ;
 wire \top_I.branch[9].block[13].um_I.iw[8] ;
 wire \top_I.branch[9].block[13].um_I.iw[9] ;
 wire \top_I.branch[9].block[13].um_I.k_zero ;
 wire \top_I.branch[9].block[13].um_I.pg_vdd ;
 wire \top_I.branch[9].block[14].um_I.ana[2] ;
 wire \top_I.branch[9].block[14].um_I.ana[3] ;
 wire \top_I.branch[9].block[14].um_I.ana[4] ;
 wire \top_I.branch[9].block[14].um_I.ana[5] ;
 wire \top_I.branch[9].block[14].um_I.ana[6] ;
 wire \top_I.branch[9].block[14].um_I.ana[7] ;
 wire \top_I.branch[9].block[14].um_I.clk ;
 wire \top_I.branch[9].block[14].um_I.ena ;
 wire \top_I.branch[9].block[14].um_I.iw[10] ;
 wire \top_I.branch[9].block[14].um_I.iw[11] ;
 wire \top_I.branch[9].block[14].um_I.iw[12] ;
 wire \top_I.branch[9].block[14].um_I.iw[13] ;
 wire \top_I.branch[9].block[14].um_I.iw[14] ;
 wire \top_I.branch[9].block[14].um_I.iw[15] ;
 wire \top_I.branch[9].block[14].um_I.iw[16] ;
 wire \top_I.branch[9].block[14].um_I.iw[17] ;
 wire \top_I.branch[9].block[14].um_I.iw[1] ;
 wire \top_I.branch[9].block[14].um_I.iw[2] ;
 wire \top_I.branch[9].block[14].um_I.iw[3] ;
 wire \top_I.branch[9].block[14].um_I.iw[4] ;
 wire \top_I.branch[9].block[14].um_I.iw[5] ;
 wire \top_I.branch[9].block[14].um_I.iw[6] ;
 wire \top_I.branch[9].block[14].um_I.iw[7] ;
 wire \top_I.branch[9].block[14].um_I.iw[8] ;
 wire \top_I.branch[9].block[14].um_I.iw[9] ;
 wire \top_I.branch[9].block[14].um_I.k_zero ;
 wire \top_I.branch[9].block[14].um_I.pg_vdd ;
 wire \top_I.branch[9].block[15].um_I.ana[2] ;
 wire \top_I.branch[9].block[15].um_I.ana[3] ;
 wire \top_I.branch[9].block[15].um_I.ana[4] ;
 wire \top_I.branch[9].block[15].um_I.ana[5] ;
 wire \top_I.branch[9].block[15].um_I.ana[6] ;
 wire \top_I.branch[9].block[15].um_I.ana[7] ;
 wire \top_I.branch[9].block[15].um_I.clk ;
 wire \top_I.branch[9].block[15].um_I.ena ;
 wire \top_I.branch[9].block[15].um_I.iw[10] ;
 wire \top_I.branch[9].block[15].um_I.iw[11] ;
 wire \top_I.branch[9].block[15].um_I.iw[12] ;
 wire \top_I.branch[9].block[15].um_I.iw[13] ;
 wire \top_I.branch[9].block[15].um_I.iw[14] ;
 wire \top_I.branch[9].block[15].um_I.iw[15] ;
 wire \top_I.branch[9].block[15].um_I.iw[16] ;
 wire \top_I.branch[9].block[15].um_I.iw[17] ;
 wire \top_I.branch[9].block[15].um_I.iw[1] ;
 wire \top_I.branch[9].block[15].um_I.iw[2] ;
 wire \top_I.branch[9].block[15].um_I.iw[3] ;
 wire \top_I.branch[9].block[15].um_I.iw[4] ;
 wire \top_I.branch[9].block[15].um_I.iw[5] ;
 wire \top_I.branch[9].block[15].um_I.iw[6] ;
 wire \top_I.branch[9].block[15].um_I.iw[7] ;
 wire \top_I.branch[9].block[15].um_I.iw[8] ;
 wire \top_I.branch[9].block[15].um_I.iw[9] ;
 wire \top_I.branch[9].block[15].um_I.k_zero ;
 wire \top_I.branch[9].block[15].um_I.pg_vdd ;
 wire \top_I.branch[9].block[1].um_I.ana[2] ;
 wire \top_I.branch[9].block[1].um_I.ana[3] ;
 wire \top_I.branch[9].block[1].um_I.ana[4] ;
 wire \top_I.branch[9].block[1].um_I.ana[5] ;
 wire \top_I.branch[9].block[1].um_I.ana[6] ;
 wire \top_I.branch[9].block[1].um_I.ana[7] ;
 wire \top_I.branch[9].block[1].um_I.clk ;
 wire \top_I.branch[9].block[1].um_I.ena ;
 wire \top_I.branch[9].block[1].um_I.iw[10] ;
 wire \top_I.branch[9].block[1].um_I.iw[11] ;
 wire \top_I.branch[9].block[1].um_I.iw[12] ;
 wire \top_I.branch[9].block[1].um_I.iw[13] ;
 wire \top_I.branch[9].block[1].um_I.iw[14] ;
 wire \top_I.branch[9].block[1].um_I.iw[15] ;
 wire \top_I.branch[9].block[1].um_I.iw[16] ;
 wire \top_I.branch[9].block[1].um_I.iw[17] ;
 wire \top_I.branch[9].block[1].um_I.iw[1] ;
 wire \top_I.branch[9].block[1].um_I.iw[2] ;
 wire \top_I.branch[9].block[1].um_I.iw[3] ;
 wire \top_I.branch[9].block[1].um_I.iw[4] ;
 wire \top_I.branch[9].block[1].um_I.iw[5] ;
 wire \top_I.branch[9].block[1].um_I.iw[6] ;
 wire \top_I.branch[9].block[1].um_I.iw[7] ;
 wire \top_I.branch[9].block[1].um_I.iw[8] ;
 wire \top_I.branch[9].block[1].um_I.iw[9] ;
 wire \top_I.branch[9].block[1].um_I.k_zero ;
 wire \top_I.branch[9].block[1].um_I.pg_vdd ;
 wire \top_I.branch[9].block[2].um_I.ana[2] ;
 wire \top_I.branch[9].block[2].um_I.ana[3] ;
 wire \top_I.branch[9].block[2].um_I.ana[4] ;
 wire \top_I.branch[9].block[2].um_I.ana[5] ;
 wire \top_I.branch[9].block[2].um_I.ana[6] ;
 wire \top_I.branch[9].block[2].um_I.ana[7] ;
 wire \top_I.branch[9].block[2].um_I.clk ;
 wire \top_I.branch[9].block[2].um_I.ena ;
 wire \top_I.branch[9].block[2].um_I.iw[10] ;
 wire \top_I.branch[9].block[2].um_I.iw[11] ;
 wire \top_I.branch[9].block[2].um_I.iw[12] ;
 wire \top_I.branch[9].block[2].um_I.iw[13] ;
 wire \top_I.branch[9].block[2].um_I.iw[14] ;
 wire \top_I.branch[9].block[2].um_I.iw[15] ;
 wire \top_I.branch[9].block[2].um_I.iw[16] ;
 wire \top_I.branch[9].block[2].um_I.iw[17] ;
 wire \top_I.branch[9].block[2].um_I.iw[1] ;
 wire \top_I.branch[9].block[2].um_I.iw[2] ;
 wire \top_I.branch[9].block[2].um_I.iw[3] ;
 wire \top_I.branch[9].block[2].um_I.iw[4] ;
 wire \top_I.branch[9].block[2].um_I.iw[5] ;
 wire \top_I.branch[9].block[2].um_I.iw[6] ;
 wire \top_I.branch[9].block[2].um_I.iw[7] ;
 wire \top_I.branch[9].block[2].um_I.iw[8] ;
 wire \top_I.branch[9].block[2].um_I.iw[9] ;
 wire \top_I.branch[9].block[2].um_I.k_zero ;
 wire \top_I.branch[9].block[2].um_I.pg_vdd ;
 wire \top_I.branch[9].block[3].um_I.ana[2] ;
 wire \top_I.branch[9].block[3].um_I.ana[3] ;
 wire \top_I.branch[9].block[3].um_I.ana[4] ;
 wire \top_I.branch[9].block[3].um_I.ana[5] ;
 wire \top_I.branch[9].block[3].um_I.ana[6] ;
 wire \top_I.branch[9].block[3].um_I.ana[7] ;
 wire \top_I.branch[9].block[3].um_I.clk ;
 wire \top_I.branch[9].block[3].um_I.ena ;
 wire \top_I.branch[9].block[3].um_I.iw[10] ;
 wire \top_I.branch[9].block[3].um_I.iw[11] ;
 wire \top_I.branch[9].block[3].um_I.iw[12] ;
 wire \top_I.branch[9].block[3].um_I.iw[13] ;
 wire \top_I.branch[9].block[3].um_I.iw[14] ;
 wire \top_I.branch[9].block[3].um_I.iw[15] ;
 wire \top_I.branch[9].block[3].um_I.iw[16] ;
 wire \top_I.branch[9].block[3].um_I.iw[17] ;
 wire \top_I.branch[9].block[3].um_I.iw[1] ;
 wire \top_I.branch[9].block[3].um_I.iw[2] ;
 wire \top_I.branch[9].block[3].um_I.iw[3] ;
 wire \top_I.branch[9].block[3].um_I.iw[4] ;
 wire \top_I.branch[9].block[3].um_I.iw[5] ;
 wire \top_I.branch[9].block[3].um_I.iw[6] ;
 wire \top_I.branch[9].block[3].um_I.iw[7] ;
 wire \top_I.branch[9].block[3].um_I.iw[8] ;
 wire \top_I.branch[9].block[3].um_I.iw[9] ;
 wire \top_I.branch[9].block[3].um_I.k_zero ;
 wire \top_I.branch[9].block[3].um_I.pg_vdd ;
 wire \top_I.branch[9].block[4].um_I.ana[2] ;
 wire \top_I.branch[9].block[4].um_I.ana[3] ;
 wire \top_I.branch[9].block[4].um_I.ana[4] ;
 wire \top_I.branch[9].block[4].um_I.ana[5] ;
 wire \top_I.branch[9].block[4].um_I.ana[6] ;
 wire \top_I.branch[9].block[4].um_I.ana[7] ;
 wire \top_I.branch[9].block[4].um_I.clk ;
 wire \top_I.branch[9].block[4].um_I.ena ;
 wire \top_I.branch[9].block[4].um_I.iw[10] ;
 wire \top_I.branch[9].block[4].um_I.iw[11] ;
 wire \top_I.branch[9].block[4].um_I.iw[12] ;
 wire \top_I.branch[9].block[4].um_I.iw[13] ;
 wire \top_I.branch[9].block[4].um_I.iw[14] ;
 wire \top_I.branch[9].block[4].um_I.iw[15] ;
 wire \top_I.branch[9].block[4].um_I.iw[16] ;
 wire \top_I.branch[9].block[4].um_I.iw[17] ;
 wire \top_I.branch[9].block[4].um_I.iw[1] ;
 wire \top_I.branch[9].block[4].um_I.iw[2] ;
 wire \top_I.branch[9].block[4].um_I.iw[3] ;
 wire \top_I.branch[9].block[4].um_I.iw[4] ;
 wire \top_I.branch[9].block[4].um_I.iw[5] ;
 wire \top_I.branch[9].block[4].um_I.iw[6] ;
 wire \top_I.branch[9].block[4].um_I.iw[7] ;
 wire \top_I.branch[9].block[4].um_I.iw[8] ;
 wire \top_I.branch[9].block[4].um_I.iw[9] ;
 wire \top_I.branch[9].block[4].um_I.k_zero ;
 wire \top_I.branch[9].block[4].um_I.pg_vdd ;
 wire \top_I.branch[9].block[5].um_I.ana[2] ;
 wire \top_I.branch[9].block[5].um_I.ana[3] ;
 wire \top_I.branch[9].block[5].um_I.ana[4] ;
 wire \top_I.branch[9].block[5].um_I.ana[5] ;
 wire \top_I.branch[9].block[5].um_I.ana[6] ;
 wire \top_I.branch[9].block[5].um_I.ana[7] ;
 wire \top_I.branch[9].block[5].um_I.clk ;
 wire \top_I.branch[9].block[5].um_I.ena ;
 wire \top_I.branch[9].block[5].um_I.iw[10] ;
 wire \top_I.branch[9].block[5].um_I.iw[11] ;
 wire \top_I.branch[9].block[5].um_I.iw[12] ;
 wire \top_I.branch[9].block[5].um_I.iw[13] ;
 wire \top_I.branch[9].block[5].um_I.iw[14] ;
 wire \top_I.branch[9].block[5].um_I.iw[15] ;
 wire \top_I.branch[9].block[5].um_I.iw[16] ;
 wire \top_I.branch[9].block[5].um_I.iw[17] ;
 wire \top_I.branch[9].block[5].um_I.iw[1] ;
 wire \top_I.branch[9].block[5].um_I.iw[2] ;
 wire \top_I.branch[9].block[5].um_I.iw[3] ;
 wire \top_I.branch[9].block[5].um_I.iw[4] ;
 wire \top_I.branch[9].block[5].um_I.iw[5] ;
 wire \top_I.branch[9].block[5].um_I.iw[6] ;
 wire \top_I.branch[9].block[5].um_I.iw[7] ;
 wire \top_I.branch[9].block[5].um_I.iw[8] ;
 wire \top_I.branch[9].block[5].um_I.iw[9] ;
 wire \top_I.branch[9].block[5].um_I.k_zero ;
 wire \top_I.branch[9].block[5].um_I.pg_vdd ;
 wire \top_I.branch[9].block[6].um_I.ana[2] ;
 wire \top_I.branch[9].block[6].um_I.ana[3] ;
 wire \top_I.branch[9].block[6].um_I.ana[4] ;
 wire \top_I.branch[9].block[6].um_I.ana[5] ;
 wire \top_I.branch[9].block[6].um_I.ana[6] ;
 wire \top_I.branch[9].block[6].um_I.ana[7] ;
 wire \top_I.branch[9].block[6].um_I.clk ;
 wire \top_I.branch[9].block[6].um_I.ena ;
 wire \top_I.branch[9].block[6].um_I.iw[10] ;
 wire \top_I.branch[9].block[6].um_I.iw[11] ;
 wire \top_I.branch[9].block[6].um_I.iw[12] ;
 wire \top_I.branch[9].block[6].um_I.iw[13] ;
 wire \top_I.branch[9].block[6].um_I.iw[14] ;
 wire \top_I.branch[9].block[6].um_I.iw[15] ;
 wire \top_I.branch[9].block[6].um_I.iw[16] ;
 wire \top_I.branch[9].block[6].um_I.iw[17] ;
 wire \top_I.branch[9].block[6].um_I.iw[1] ;
 wire \top_I.branch[9].block[6].um_I.iw[2] ;
 wire \top_I.branch[9].block[6].um_I.iw[3] ;
 wire \top_I.branch[9].block[6].um_I.iw[4] ;
 wire \top_I.branch[9].block[6].um_I.iw[5] ;
 wire \top_I.branch[9].block[6].um_I.iw[6] ;
 wire \top_I.branch[9].block[6].um_I.iw[7] ;
 wire \top_I.branch[9].block[6].um_I.iw[8] ;
 wire \top_I.branch[9].block[6].um_I.iw[9] ;
 wire \top_I.branch[9].block[6].um_I.k_zero ;
 wire \top_I.branch[9].block[6].um_I.pg_vdd ;
 wire \top_I.branch[9].block[7].um_I.ana[2] ;
 wire \top_I.branch[9].block[7].um_I.ana[3] ;
 wire \top_I.branch[9].block[7].um_I.ana[4] ;
 wire \top_I.branch[9].block[7].um_I.ana[5] ;
 wire \top_I.branch[9].block[7].um_I.ana[6] ;
 wire \top_I.branch[9].block[7].um_I.ana[7] ;
 wire \top_I.branch[9].block[7].um_I.clk ;
 wire \top_I.branch[9].block[7].um_I.ena ;
 wire \top_I.branch[9].block[7].um_I.iw[10] ;
 wire \top_I.branch[9].block[7].um_I.iw[11] ;
 wire \top_I.branch[9].block[7].um_I.iw[12] ;
 wire \top_I.branch[9].block[7].um_I.iw[13] ;
 wire \top_I.branch[9].block[7].um_I.iw[14] ;
 wire \top_I.branch[9].block[7].um_I.iw[15] ;
 wire \top_I.branch[9].block[7].um_I.iw[16] ;
 wire \top_I.branch[9].block[7].um_I.iw[17] ;
 wire \top_I.branch[9].block[7].um_I.iw[1] ;
 wire \top_I.branch[9].block[7].um_I.iw[2] ;
 wire \top_I.branch[9].block[7].um_I.iw[3] ;
 wire \top_I.branch[9].block[7].um_I.iw[4] ;
 wire \top_I.branch[9].block[7].um_I.iw[5] ;
 wire \top_I.branch[9].block[7].um_I.iw[6] ;
 wire \top_I.branch[9].block[7].um_I.iw[7] ;
 wire \top_I.branch[9].block[7].um_I.iw[8] ;
 wire \top_I.branch[9].block[7].um_I.iw[9] ;
 wire \top_I.branch[9].block[7].um_I.k_zero ;
 wire \top_I.branch[9].block[7].um_I.pg_vdd ;
 wire \top_I.branch[9].block[8].um_I.ana[2] ;
 wire \top_I.branch[9].block[8].um_I.ana[3] ;
 wire \top_I.branch[9].block[8].um_I.ana[4] ;
 wire \top_I.branch[9].block[8].um_I.ana[5] ;
 wire \top_I.branch[9].block[8].um_I.ana[6] ;
 wire \top_I.branch[9].block[8].um_I.ana[7] ;
 wire \top_I.branch[9].block[8].um_I.clk ;
 wire \top_I.branch[9].block[8].um_I.ena ;
 wire \top_I.branch[9].block[8].um_I.iw[10] ;
 wire \top_I.branch[9].block[8].um_I.iw[11] ;
 wire \top_I.branch[9].block[8].um_I.iw[12] ;
 wire \top_I.branch[9].block[8].um_I.iw[13] ;
 wire \top_I.branch[9].block[8].um_I.iw[14] ;
 wire \top_I.branch[9].block[8].um_I.iw[15] ;
 wire \top_I.branch[9].block[8].um_I.iw[16] ;
 wire \top_I.branch[9].block[8].um_I.iw[17] ;
 wire \top_I.branch[9].block[8].um_I.iw[1] ;
 wire \top_I.branch[9].block[8].um_I.iw[2] ;
 wire \top_I.branch[9].block[8].um_I.iw[3] ;
 wire \top_I.branch[9].block[8].um_I.iw[4] ;
 wire \top_I.branch[9].block[8].um_I.iw[5] ;
 wire \top_I.branch[9].block[8].um_I.iw[6] ;
 wire \top_I.branch[9].block[8].um_I.iw[7] ;
 wire \top_I.branch[9].block[8].um_I.iw[8] ;
 wire \top_I.branch[9].block[8].um_I.iw[9] ;
 wire \top_I.branch[9].block[8].um_I.k_zero ;
 wire \top_I.branch[9].block[8].um_I.pg_vdd ;
 wire \top_I.branch[9].block[9].um_I.ana[2] ;
 wire \top_I.branch[9].block[9].um_I.ana[3] ;
 wire \top_I.branch[9].block[9].um_I.ana[4] ;
 wire \top_I.branch[9].block[9].um_I.ana[5] ;
 wire \top_I.branch[9].block[9].um_I.ana[6] ;
 wire \top_I.branch[9].block[9].um_I.ana[7] ;
 wire \top_I.branch[9].block[9].um_I.clk ;
 wire \top_I.branch[9].block[9].um_I.ena ;
 wire \top_I.branch[9].block[9].um_I.iw[10] ;
 wire \top_I.branch[9].block[9].um_I.iw[11] ;
 wire \top_I.branch[9].block[9].um_I.iw[12] ;
 wire \top_I.branch[9].block[9].um_I.iw[13] ;
 wire \top_I.branch[9].block[9].um_I.iw[14] ;
 wire \top_I.branch[9].block[9].um_I.iw[15] ;
 wire \top_I.branch[9].block[9].um_I.iw[16] ;
 wire \top_I.branch[9].block[9].um_I.iw[17] ;
 wire \top_I.branch[9].block[9].um_I.iw[1] ;
 wire \top_I.branch[9].block[9].um_I.iw[2] ;
 wire \top_I.branch[9].block[9].um_I.iw[3] ;
 wire \top_I.branch[9].block[9].um_I.iw[4] ;
 wire \top_I.branch[9].block[9].um_I.iw[5] ;
 wire \top_I.branch[9].block[9].um_I.iw[6] ;
 wire \top_I.branch[9].block[9].um_I.iw[7] ;
 wire \top_I.branch[9].block[9].um_I.iw[8] ;
 wire \top_I.branch[9].block[9].um_I.iw[9] ;
 wire \top_I.branch[9].block[9].um_I.k_zero ;
 wire \top_I.branch[9].block[9].um_I.pg_vdd ;
 wire \top_I.branch[9].l_addr[0] ;
 wire \top_I.branch[9].l_addr[2] ;
 wire \top_I.io_ana[0] ;
 wire \top_I.io_ana[1] ;
 wire \top_I.io_ana[2] ;
 wire \top_I.io_ana[36] ;
 wire \top_I.io_ana[37] ;
 wire \top_I.io_ana[3] ;
 wire \top_I.io_ana[4] ;
 wire \top_I.io_ana[5] ;
 wire \top_I.io_ana[6] ;
 wire \top_I.io_oeb[0] ;

 tt_um_chip_rom \top_I.branch[0].block[0].um_I.block_0_0.tt_um_I  (.clk(\top_I.branch[0].block[0].um_I.clk ),
    .ena(\top_I.branch[0].block[0].um_I.ena ),
    .rst_n(\top_I.branch[0].block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].block[0].um_I.iw[9] ,
    \top_I.branch[0].block[0].um_I.iw[8] ,
    \top_I.branch[0].block[0].um_I.iw[7] ,
    \top_I.branch[0].block[0].um_I.iw[6] ,
    \top_I.branch[0].block[0].um_I.iw[5] ,
    \top_I.branch[0].block[0].um_I.iw[4] ,
    \top_I.branch[0].block[0].um_I.iw[3] ,
    \top_I.branch[0].block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].block[0].um_I.iw[17] ,
    \top_I.branch[0].block[0].um_I.iw[16] ,
    \top_I.branch[0].block[0].um_I.iw[15] ,
    \top_I.branch[0].block[0].um_I.iw[14] ,
    \top_I.branch[0].block[0].um_I.iw[13] ,
    \top_I.branch[0].block[0].um_I.iw[12] ,
    \top_I.branch[0].block[0].um_I.iw[11] ,
    \top_I.branch[0].block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].block[0].um_I.ow[23] ,
    \top_I.branch[0].block[0].um_I.ow[22] ,
    \top_I.branch[0].block[0].um_I.ow[21] ,
    \top_I.branch[0].block[0].um_I.ow[20] ,
    \top_I.branch[0].block[0].um_I.ow[19] ,
    \top_I.branch[0].block[0].um_I.ow[18] ,
    \top_I.branch[0].block[0].um_I.ow[17] ,
    \top_I.branch[0].block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].block[0].um_I.ow[15] ,
    \top_I.branch[0].block[0].um_I.ow[14] ,
    \top_I.branch[0].block[0].um_I.ow[13] ,
    \top_I.branch[0].block[0].um_I.ow[12] ,
    \top_I.branch[0].block[0].um_I.ow[11] ,
    \top_I.branch[0].block[0].um_I.ow[10] ,
    \top_I.branch[0].block[0].um_I.ow[9] ,
    \top_I.branch[0].block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].block[0].um_I.ow[7] ,
    \top_I.branch[0].block[0].um_I.ow[6] ,
    \top_I.branch[0].block[0].um_I.ow[5] ,
    \top_I.branch[0].block[0].um_I.ow[4] ,
    \top_I.branch[0].block[0].um_I.ow[3] ,
    \top_I.branch[0].block[0].um_I.ow[2] ,
    \top_I.branch[0].block[0].um_I.ow[1] ,
    \top_I.branch[0].block[0].um_I.ow[0] }));
 tt_um_factory_test \top_I.branch[0].block[1].um_I.block_0_1.tt_um_I  (.clk(\top_I.branch[0].block[1].um_I.clk ),
    .ena(\top_I.branch[0].block[1].um_I.ena ),
    .rst_n(\top_I.branch[0].block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].block[1].um_I.iw[9] ,
    \top_I.branch[0].block[1].um_I.iw[8] ,
    \top_I.branch[0].block[1].um_I.iw[7] ,
    \top_I.branch[0].block[1].um_I.iw[6] ,
    \top_I.branch[0].block[1].um_I.iw[5] ,
    \top_I.branch[0].block[1].um_I.iw[4] ,
    \top_I.branch[0].block[1].um_I.iw[3] ,
    \top_I.branch[0].block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].block[1].um_I.iw[17] ,
    \top_I.branch[0].block[1].um_I.iw[16] ,
    \top_I.branch[0].block[1].um_I.iw[15] ,
    \top_I.branch[0].block[1].um_I.iw[14] ,
    \top_I.branch[0].block[1].um_I.iw[13] ,
    \top_I.branch[0].block[1].um_I.iw[12] ,
    \top_I.branch[0].block[1].um_I.iw[11] ,
    \top_I.branch[0].block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].block[1].um_I.ow[23] ,
    \top_I.branch[0].block[1].um_I.ow[22] ,
    \top_I.branch[0].block[1].um_I.ow[21] ,
    \top_I.branch[0].block[1].um_I.ow[20] ,
    \top_I.branch[0].block[1].um_I.ow[19] ,
    \top_I.branch[0].block[1].um_I.ow[18] ,
    \top_I.branch[0].block[1].um_I.ow[17] ,
    \top_I.branch[0].block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].block[1].um_I.ow[15] ,
    \top_I.branch[0].block[1].um_I.ow[14] ,
    \top_I.branch[0].block[1].um_I.ow[13] ,
    \top_I.branch[0].block[1].um_I.ow[12] ,
    \top_I.branch[0].block[1].um_I.ow[11] ,
    \top_I.branch[0].block[1].um_I.ow[10] ,
    \top_I.branch[0].block[1].um_I.ow[9] ,
    \top_I.branch[0].block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].block[1].um_I.ow[7] ,
    \top_I.branch[0].block[1].um_I.ow[6] ,
    \top_I.branch[0].block[1].um_I.ow[5] ,
    \top_I.branch[0].block[1].um_I.ow[4] ,
    \top_I.branch[0].block[1].um_I.ow[3] ,
    \top_I.branch[0].block[1].um_I.ow[2] ,
    \top_I.branch[0].block[1].um_I.ow[1] ,
    \top_I.branch[0].block[1].um_I.ow[0] }));
 tt_mux \top_I.branch[0].mux_I  (.k_one(\top_I.branch[0].l_k_one ),
    .k_zero(\top_I.branch[0].l_addr[0] ),
    .addr({\top_I.branch[0].l_addr[0] ,
    \top_I.branch[0].l_addr[0] ,
    \top_I.branch[0].l_addr[0] ,
    \top_I.branch[0].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[0].block[15].um_I.ena ,
    \top_I.branch[0].block[14].um_I.ena ,
    \top_I.branch[0].block[13].um_I.ena ,
    \top_I.branch[0].block[12].um_I.ena ,
    \top_I.branch[0].block[11].um_I.ena ,
    \top_I.branch[0].block[10].um_I.ena ,
    \top_I.branch[0].block[9].um_I.ena ,
    \top_I.branch[0].block[8].um_I.ena ,
    \top_I.branch[0].block[7].um_I.ena ,
    \top_I.branch[0].block[6].um_I.ena ,
    \top_I.branch[0].block[5].um_I.ena ,
    \top_I.branch[0].block[4].um_I.ena ,
    \top_I.branch[0].block[3].um_I.ena ,
    \top_I.branch[0].block[2].um_I.ena ,
    \top_I.branch[0].block[1].um_I.ena ,
    \top_I.branch[0].block[0].um_I.ena }),
    .um_iw({\top_I.branch[0].block[15].um_I.iw[17] ,
    \top_I.branch[0].block[15].um_I.iw[16] ,
    \top_I.branch[0].block[15].um_I.iw[15] ,
    \top_I.branch[0].block[15].um_I.iw[14] ,
    \top_I.branch[0].block[15].um_I.iw[13] ,
    \top_I.branch[0].block[15].um_I.iw[12] ,
    \top_I.branch[0].block[15].um_I.iw[11] ,
    \top_I.branch[0].block[15].um_I.iw[10] ,
    \top_I.branch[0].block[15].um_I.iw[9] ,
    \top_I.branch[0].block[15].um_I.iw[8] ,
    \top_I.branch[0].block[15].um_I.iw[7] ,
    \top_I.branch[0].block[15].um_I.iw[6] ,
    \top_I.branch[0].block[15].um_I.iw[5] ,
    \top_I.branch[0].block[15].um_I.iw[4] ,
    \top_I.branch[0].block[15].um_I.iw[3] ,
    \top_I.branch[0].block[15].um_I.iw[2] ,
    \top_I.branch[0].block[15].um_I.iw[1] ,
    \top_I.branch[0].block[15].um_I.clk ,
    \top_I.branch[0].block[14].um_I.iw[17] ,
    \top_I.branch[0].block[14].um_I.iw[16] ,
    \top_I.branch[0].block[14].um_I.iw[15] ,
    \top_I.branch[0].block[14].um_I.iw[14] ,
    \top_I.branch[0].block[14].um_I.iw[13] ,
    \top_I.branch[0].block[14].um_I.iw[12] ,
    \top_I.branch[0].block[14].um_I.iw[11] ,
    \top_I.branch[0].block[14].um_I.iw[10] ,
    \top_I.branch[0].block[14].um_I.iw[9] ,
    \top_I.branch[0].block[14].um_I.iw[8] ,
    \top_I.branch[0].block[14].um_I.iw[7] ,
    \top_I.branch[0].block[14].um_I.iw[6] ,
    \top_I.branch[0].block[14].um_I.iw[5] ,
    \top_I.branch[0].block[14].um_I.iw[4] ,
    \top_I.branch[0].block[14].um_I.iw[3] ,
    \top_I.branch[0].block[14].um_I.iw[2] ,
    \top_I.branch[0].block[14].um_I.iw[1] ,
    \top_I.branch[0].block[14].um_I.clk ,
    \top_I.branch[0].block[13].um_I.iw[17] ,
    \top_I.branch[0].block[13].um_I.iw[16] ,
    \top_I.branch[0].block[13].um_I.iw[15] ,
    \top_I.branch[0].block[13].um_I.iw[14] ,
    \top_I.branch[0].block[13].um_I.iw[13] ,
    \top_I.branch[0].block[13].um_I.iw[12] ,
    \top_I.branch[0].block[13].um_I.iw[11] ,
    \top_I.branch[0].block[13].um_I.iw[10] ,
    \top_I.branch[0].block[13].um_I.iw[9] ,
    \top_I.branch[0].block[13].um_I.iw[8] ,
    \top_I.branch[0].block[13].um_I.iw[7] ,
    \top_I.branch[0].block[13].um_I.iw[6] ,
    \top_I.branch[0].block[13].um_I.iw[5] ,
    \top_I.branch[0].block[13].um_I.iw[4] ,
    \top_I.branch[0].block[13].um_I.iw[3] ,
    \top_I.branch[0].block[13].um_I.iw[2] ,
    \top_I.branch[0].block[13].um_I.iw[1] ,
    \top_I.branch[0].block[13].um_I.clk ,
    \top_I.branch[0].block[12].um_I.iw[17] ,
    \top_I.branch[0].block[12].um_I.iw[16] ,
    \top_I.branch[0].block[12].um_I.iw[15] ,
    \top_I.branch[0].block[12].um_I.iw[14] ,
    \top_I.branch[0].block[12].um_I.iw[13] ,
    \top_I.branch[0].block[12].um_I.iw[12] ,
    \top_I.branch[0].block[12].um_I.iw[11] ,
    \top_I.branch[0].block[12].um_I.iw[10] ,
    \top_I.branch[0].block[12].um_I.iw[9] ,
    \top_I.branch[0].block[12].um_I.iw[8] ,
    \top_I.branch[0].block[12].um_I.iw[7] ,
    \top_I.branch[0].block[12].um_I.iw[6] ,
    \top_I.branch[0].block[12].um_I.iw[5] ,
    \top_I.branch[0].block[12].um_I.iw[4] ,
    \top_I.branch[0].block[12].um_I.iw[3] ,
    \top_I.branch[0].block[12].um_I.iw[2] ,
    \top_I.branch[0].block[12].um_I.iw[1] ,
    \top_I.branch[0].block[12].um_I.clk ,
    \top_I.branch[0].block[11].um_I.iw[17] ,
    \top_I.branch[0].block[11].um_I.iw[16] ,
    \top_I.branch[0].block[11].um_I.iw[15] ,
    \top_I.branch[0].block[11].um_I.iw[14] ,
    \top_I.branch[0].block[11].um_I.iw[13] ,
    \top_I.branch[0].block[11].um_I.iw[12] ,
    \top_I.branch[0].block[11].um_I.iw[11] ,
    \top_I.branch[0].block[11].um_I.iw[10] ,
    \top_I.branch[0].block[11].um_I.iw[9] ,
    \top_I.branch[0].block[11].um_I.iw[8] ,
    \top_I.branch[0].block[11].um_I.iw[7] ,
    \top_I.branch[0].block[11].um_I.iw[6] ,
    \top_I.branch[0].block[11].um_I.iw[5] ,
    \top_I.branch[0].block[11].um_I.iw[4] ,
    \top_I.branch[0].block[11].um_I.iw[3] ,
    \top_I.branch[0].block[11].um_I.iw[2] ,
    \top_I.branch[0].block[11].um_I.iw[1] ,
    \top_I.branch[0].block[11].um_I.clk ,
    \top_I.branch[0].block[10].um_I.iw[17] ,
    \top_I.branch[0].block[10].um_I.iw[16] ,
    \top_I.branch[0].block[10].um_I.iw[15] ,
    \top_I.branch[0].block[10].um_I.iw[14] ,
    \top_I.branch[0].block[10].um_I.iw[13] ,
    \top_I.branch[0].block[10].um_I.iw[12] ,
    \top_I.branch[0].block[10].um_I.iw[11] ,
    \top_I.branch[0].block[10].um_I.iw[10] ,
    \top_I.branch[0].block[10].um_I.iw[9] ,
    \top_I.branch[0].block[10].um_I.iw[8] ,
    \top_I.branch[0].block[10].um_I.iw[7] ,
    \top_I.branch[0].block[10].um_I.iw[6] ,
    \top_I.branch[0].block[10].um_I.iw[5] ,
    \top_I.branch[0].block[10].um_I.iw[4] ,
    \top_I.branch[0].block[10].um_I.iw[3] ,
    \top_I.branch[0].block[10].um_I.iw[2] ,
    \top_I.branch[0].block[10].um_I.iw[1] ,
    \top_I.branch[0].block[10].um_I.clk ,
    \top_I.branch[0].block[9].um_I.iw[17] ,
    \top_I.branch[0].block[9].um_I.iw[16] ,
    \top_I.branch[0].block[9].um_I.iw[15] ,
    \top_I.branch[0].block[9].um_I.iw[14] ,
    \top_I.branch[0].block[9].um_I.iw[13] ,
    \top_I.branch[0].block[9].um_I.iw[12] ,
    \top_I.branch[0].block[9].um_I.iw[11] ,
    \top_I.branch[0].block[9].um_I.iw[10] ,
    \top_I.branch[0].block[9].um_I.iw[9] ,
    \top_I.branch[0].block[9].um_I.iw[8] ,
    \top_I.branch[0].block[9].um_I.iw[7] ,
    \top_I.branch[0].block[9].um_I.iw[6] ,
    \top_I.branch[0].block[9].um_I.iw[5] ,
    \top_I.branch[0].block[9].um_I.iw[4] ,
    \top_I.branch[0].block[9].um_I.iw[3] ,
    \top_I.branch[0].block[9].um_I.iw[2] ,
    \top_I.branch[0].block[9].um_I.iw[1] ,
    \top_I.branch[0].block[9].um_I.clk ,
    \top_I.branch[0].block[8].um_I.iw[17] ,
    \top_I.branch[0].block[8].um_I.iw[16] ,
    \top_I.branch[0].block[8].um_I.iw[15] ,
    \top_I.branch[0].block[8].um_I.iw[14] ,
    \top_I.branch[0].block[8].um_I.iw[13] ,
    \top_I.branch[0].block[8].um_I.iw[12] ,
    \top_I.branch[0].block[8].um_I.iw[11] ,
    \top_I.branch[0].block[8].um_I.iw[10] ,
    \top_I.branch[0].block[8].um_I.iw[9] ,
    \top_I.branch[0].block[8].um_I.iw[8] ,
    \top_I.branch[0].block[8].um_I.iw[7] ,
    \top_I.branch[0].block[8].um_I.iw[6] ,
    \top_I.branch[0].block[8].um_I.iw[5] ,
    \top_I.branch[0].block[8].um_I.iw[4] ,
    \top_I.branch[0].block[8].um_I.iw[3] ,
    \top_I.branch[0].block[8].um_I.iw[2] ,
    \top_I.branch[0].block[8].um_I.iw[1] ,
    \top_I.branch[0].block[8].um_I.clk ,
    \top_I.branch[0].block[7].um_I.iw[17] ,
    \top_I.branch[0].block[7].um_I.iw[16] ,
    \top_I.branch[0].block[7].um_I.iw[15] ,
    \top_I.branch[0].block[7].um_I.iw[14] ,
    \top_I.branch[0].block[7].um_I.iw[13] ,
    \top_I.branch[0].block[7].um_I.iw[12] ,
    \top_I.branch[0].block[7].um_I.iw[11] ,
    \top_I.branch[0].block[7].um_I.iw[10] ,
    \top_I.branch[0].block[7].um_I.iw[9] ,
    \top_I.branch[0].block[7].um_I.iw[8] ,
    \top_I.branch[0].block[7].um_I.iw[7] ,
    \top_I.branch[0].block[7].um_I.iw[6] ,
    \top_I.branch[0].block[7].um_I.iw[5] ,
    \top_I.branch[0].block[7].um_I.iw[4] ,
    \top_I.branch[0].block[7].um_I.iw[3] ,
    \top_I.branch[0].block[7].um_I.iw[2] ,
    \top_I.branch[0].block[7].um_I.iw[1] ,
    \top_I.branch[0].block[7].um_I.clk ,
    \top_I.branch[0].block[6].um_I.iw[17] ,
    \top_I.branch[0].block[6].um_I.iw[16] ,
    \top_I.branch[0].block[6].um_I.iw[15] ,
    \top_I.branch[0].block[6].um_I.iw[14] ,
    \top_I.branch[0].block[6].um_I.iw[13] ,
    \top_I.branch[0].block[6].um_I.iw[12] ,
    \top_I.branch[0].block[6].um_I.iw[11] ,
    \top_I.branch[0].block[6].um_I.iw[10] ,
    \top_I.branch[0].block[6].um_I.iw[9] ,
    \top_I.branch[0].block[6].um_I.iw[8] ,
    \top_I.branch[0].block[6].um_I.iw[7] ,
    \top_I.branch[0].block[6].um_I.iw[6] ,
    \top_I.branch[0].block[6].um_I.iw[5] ,
    \top_I.branch[0].block[6].um_I.iw[4] ,
    \top_I.branch[0].block[6].um_I.iw[3] ,
    \top_I.branch[0].block[6].um_I.iw[2] ,
    \top_I.branch[0].block[6].um_I.iw[1] ,
    \top_I.branch[0].block[6].um_I.clk ,
    \top_I.branch[0].block[5].um_I.iw[17] ,
    \top_I.branch[0].block[5].um_I.iw[16] ,
    \top_I.branch[0].block[5].um_I.iw[15] ,
    \top_I.branch[0].block[5].um_I.iw[14] ,
    \top_I.branch[0].block[5].um_I.iw[13] ,
    \top_I.branch[0].block[5].um_I.iw[12] ,
    \top_I.branch[0].block[5].um_I.iw[11] ,
    \top_I.branch[0].block[5].um_I.iw[10] ,
    \top_I.branch[0].block[5].um_I.iw[9] ,
    \top_I.branch[0].block[5].um_I.iw[8] ,
    \top_I.branch[0].block[5].um_I.iw[7] ,
    \top_I.branch[0].block[5].um_I.iw[6] ,
    \top_I.branch[0].block[5].um_I.iw[5] ,
    \top_I.branch[0].block[5].um_I.iw[4] ,
    \top_I.branch[0].block[5].um_I.iw[3] ,
    \top_I.branch[0].block[5].um_I.iw[2] ,
    \top_I.branch[0].block[5].um_I.iw[1] ,
    \top_I.branch[0].block[5].um_I.clk ,
    \top_I.branch[0].block[4].um_I.iw[17] ,
    \top_I.branch[0].block[4].um_I.iw[16] ,
    \top_I.branch[0].block[4].um_I.iw[15] ,
    \top_I.branch[0].block[4].um_I.iw[14] ,
    \top_I.branch[0].block[4].um_I.iw[13] ,
    \top_I.branch[0].block[4].um_I.iw[12] ,
    \top_I.branch[0].block[4].um_I.iw[11] ,
    \top_I.branch[0].block[4].um_I.iw[10] ,
    \top_I.branch[0].block[4].um_I.iw[9] ,
    \top_I.branch[0].block[4].um_I.iw[8] ,
    \top_I.branch[0].block[4].um_I.iw[7] ,
    \top_I.branch[0].block[4].um_I.iw[6] ,
    \top_I.branch[0].block[4].um_I.iw[5] ,
    \top_I.branch[0].block[4].um_I.iw[4] ,
    \top_I.branch[0].block[4].um_I.iw[3] ,
    \top_I.branch[0].block[4].um_I.iw[2] ,
    \top_I.branch[0].block[4].um_I.iw[1] ,
    \top_I.branch[0].block[4].um_I.clk ,
    \top_I.branch[0].block[3].um_I.iw[17] ,
    \top_I.branch[0].block[3].um_I.iw[16] ,
    \top_I.branch[0].block[3].um_I.iw[15] ,
    \top_I.branch[0].block[3].um_I.iw[14] ,
    \top_I.branch[0].block[3].um_I.iw[13] ,
    \top_I.branch[0].block[3].um_I.iw[12] ,
    \top_I.branch[0].block[3].um_I.iw[11] ,
    \top_I.branch[0].block[3].um_I.iw[10] ,
    \top_I.branch[0].block[3].um_I.iw[9] ,
    \top_I.branch[0].block[3].um_I.iw[8] ,
    \top_I.branch[0].block[3].um_I.iw[7] ,
    \top_I.branch[0].block[3].um_I.iw[6] ,
    \top_I.branch[0].block[3].um_I.iw[5] ,
    \top_I.branch[0].block[3].um_I.iw[4] ,
    \top_I.branch[0].block[3].um_I.iw[3] ,
    \top_I.branch[0].block[3].um_I.iw[2] ,
    \top_I.branch[0].block[3].um_I.iw[1] ,
    \top_I.branch[0].block[3].um_I.clk ,
    \top_I.branch[0].block[2].um_I.iw[17] ,
    \top_I.branch[0].block[2].um_I.iw[16] ,
    \top_I.branch[0].block[2].um_I.iw[15] ,
    \top_I.branch[0].block[2].um_I.iw[14] ,
    \top_I.branch[0].block[2].um_I.iw[13] ,
    \top_I.branch[0].block[2].um_I.iw[12] ,
    \top_I.branch[0].block[2].um_I.iw[11] ,
    \top_I.branch[0].block[2].um_I.iw[10] ,
    \top_I.branch[0].block[2].um_I.iw[9] ,
    \top_I.branch[0].block[2].um_I.iw[8] ,
    \top_I.branch[0].block[2].um_I.iw[7] ,
    \top_I.branch[0].block[2].um_I.iw[6] ,
    \top_I.branch[0].block[2].um_I.iw[5] ,
    \top_I.branch[0].block[2].um_I.iw[4] ,
    \top_I.branch[0].block[2].um_I.iw[3] ,
    \top_I.branch[0].block[2].um_I.iw[2] ,
    \top_I.branch[0].block[2].um_I.iw[1] ,
    \top_I.branch[0].block[2].um_I.clk ,
    \top_I.branch[0].block[1].um_I.iw[17] ,
    \top_I.branch[0].block[1].um_I.iw[16] ,
    \top_I.branch[0].block[1].um_I.iw[15] ,
    \top_I.branch[0].block[1].um_I.iw[14] ,
    \top_I.branch[0].block[1].um_I.iw[13] ,
    \top_I.branch[0].block[1].um_I.iw[12] ,
    \top_I.branch[0].block[1].um_I.iw[11] ,
    \top_I.branch[0].block[1].um_I.iw[10] ,
    \top_I.branch[0].block[1].um_I.iw[9] ,
    \top_I.branch[0].block[1].um_I.iw[8] ,
    \top_I.branch[0].block[1].um_I.iw[7] ,
    \top_I.branch[0].block[1].um_I.iw[6] ,
    \top_I.branch[0].block[1].um_I.iw[5] ,
    \top_I.branch[0].block[1].um_I.iw[4] ,
    \top_I.branch[0].block[1].um_I.iw[3] ,
    \top_I.branch[0].block[1].um_I.iw[2] ,
    \top_I.branch[0].block[1].um_I.iw[1] ,
    \top_I.branch[0].block[1].um_I.clk ,
    \top_I.branch[0].block[0].um_I.iw[17] ,
    \top_I.branch[0].block[0].um_I.iw[16] ,
    \top_I.branch[0].block[0].um_I.iw[15] ,
    \top_I.branch[0].block[0].um_I.iw[14] ,
    \top_I.branch[0].block[0].um_I.iw[13] ,
    \top_I.branch[0].block[0].um_I.iw[12] ,
    \top_I.branch[0].block[0].um_I.iw[11] ,
    \top_I.branch[0].block[0].um_I.iw[10] ,
    \top_I.branch[0].block[0].um_I.iw[9] ,
    \top_I.branch[0].block[0].um_I.iw[8] ,
    \top_I.branch[0].block[0].um_I.iw[7] ,
    \top_I.branch[0].block[0].um_I.iw[6] ,
    \top_I.branch[0].block[0].um_I.iw[5] ,
    \top_I.branch[0].block[0].um_I.iw[4] ,
    \top_I.branch[0].block[0].um_I.iw[3] ,
    \top_I.branch[0].block[0].um_I.iw[2] ,
    \top_I.branch[0].block[0].um_I.iw[1] ,
    \top_I.branch[0].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[1].um_I.k_zero ,
    \top_I.branch[0].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[1].um_I.ow[23] ,
    \top_I.branch[0].block[1].um_I.ow[22] ,
    \top_I.branch[0].block[1].um_I.ow[21] ,
    \top_I.branch[0].block[1].um_I.ow[20] ,
    \top_I.branch[0].block[1].um_I.ow[19] ,
    \top_I.branch[0].block[1].um_I.ow[18] ,
    \top_I.branch[0].block[1].um_I.ow[17] ,
    \top_I.branch[0].block[1].um_I.ow[16] ,
    \top_I.branch[0].block[1].um_I.ow[15] ,
    \top_I.branch[0].block[1].um_I.ow[14] ,
    \top_I.branch[0].block[1].um_I.ow[13] ,
    \top_I.branch[0].block[1].um_I.ow[12] ,
    \top_I.branch[0].block[1].um_I.ow[11] ,
    \top_I.branch[0].block[1].um_I.ow[10] ,
    \top_I.branch[0].block[1].um_I.ow[9] ,
    \top_I.branch[0].block[1].um_I.ow[8] ,
    \top_I.branch[0].block[1].um_I.ow[7] ,
    \top_I.branch[0].block[1].um_I.ow[6] ,
    \top_I.branch[0].block[1].um_I.ow[5] ,
    \top_I.branch[0].block[1].um_I.ow[4] ,
    \top_I.branch[0].block[1].um_I.ow[3] ,
    \top_I.branch[0].block[1].um_I.ow[2] ,
    \top_I.branch[0].block[1].um_I.ow[1] ,
    \top_I.branch[0].block[1].um_I.ow[0] ,
    \top_I.branch[0].block[0].um_I.ow[23] ,
    \top_I.branch[0].block[0].um_I.ow[22] ,
    \top_I.branch[0].block[0].um_I.ow[21] ,
    \top_I.branch[0].block[0].um_I.ow[20] ,
    \top_I.branch[0].block[0].um_I.ow[19] ,
    \top_I.branch[0].block[0].um_I.ow[18] ,
    \top_I.branch[0].block[0].um_I.ow[17] ,
    \top_I.branch[0].block[0].um_I.ow[16] ,
    \top_I.branch[0].block[0].um_I.ow[15] ,
    \top_I.branch[0].block[0].um_I.ow[14] ,
    \top_I.branch[0].block[0].um_I.ow[13] ,
    \top_I.branch[0].block[0].um_I.ow[12] ,
    \top_I.branch[0].block[0].um_I.ow[11] ,
    \top_I.branch[0].block[0].um_I.ow[10] ,
    \top_I.branch[0].block[0].um_I.ow[9] ,
    \top_I.branch[0].block[0].um_I.ow[8] ,
    \top_I.branch[0].block[0].um_I.ow[7] ,
    \top_I.branch[0].block[0].um_I.ow[6] ,
    \top_I.branch[0].block[0].um_I.ow[5] ,
    \top_I.branch[0].block[0].um_I.ow[4] ,
    \top_I.branch[0].block[0].um_I.ow[3] ,
    \top_I.branch[0].block[0].um_I.ow[2] ,
    \top_I.branch[0].block[0].um_I.ow[1] ,
    \top_I.branch[0].block[0].um_I.ow[0] }),
    .um_pg_vdd({\top_I.branch[0].block[15].um_I.pg_vdd ,
    \top_I.branch[0].block[14].um_I.pg_vdd ,
    \top_I.branch[0].block[13].um_I.pg_vdd ,
    \top_I.branch[0].block[12].um_I.pg_vdd ,
    \top_I.branch[0].block[11].um_I.pg_vdd ,
    \top_I.branch[0].block[10].um_I.pg_vdd ,
    \top_I.branch[0].block[9].um_I.pg_vdd ,
    \top_I.branch[0].block[8].um_I.pg_vdd ,
    \top_I.branch[0].block[7].um_I.pg_vdd ,
    \top_I.branch[0].block[6].um_I.pg_vdd ,
    \top_I.branch[0].block[5].um_I.pg_vdd ,
    \top_I.branch[0].block[4].um_I.pg_vdd ,
    \top_I.branch[0].block[3].um_I.pg_vdd ,
    \top_I.branch[0].block[2].um_I.pg_vdd ,
    \top_I.branch[0].block[1].um_I.pg_vdd ,
    \top_I.branch[0].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[10].mux_I  (.k_one(\top_I.branch[10].l_addr[0] ),
    .k_zero(\top_I.branch[10].l_addr[1] ),
    .addr({\top_I.branch[10].l_addr[1] ,
    \top_I.branch[10].l_addr[0] ,
    \top_I.branch[10].l_addr[1] ,
    \top_I.branch[10].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[10].block[15].um_I.ena ,
    \top_I.branch[10].block[14].um_I.ena ,
    \top_I.branch[10].block[13].um_I.ena ,
    \top_I.branch[10].block[12].um_I.ena ,
    \top_I.branch[10].block[11].um_I.ena ,
    \top_I.branch[10].block[10].um_I.ena ,
    \top_I.branch[10].block[9].um_I.ena ,
    \top_I.branch[10].block[8].um_I.ena ,
    \top_I.branch[10].block[7].um_I.ena ,
    \top_I.branch[10].block[6].um_I.ena ,
    \top_I.branch[10].block[5].um_I.ena ,
    \top_I.branch[10].block[4].um_I.ena ,
    \top_I.branch[10].block[3].um_I.ena ,
    \top_I.branch[10].block[2].um_I.ena ,
    \top_I.branch[10].block[1].um_I.ena ,
    \top_I.branch[10].block[0].um_I.ena }),
    .um_iw({\top_I.branch[10].block[15].um_I.iw[17] ,
    \top_I.branch[10].block[15].um_I.iw[16] ,
    \top_I.branch[10].block[15].um_I.iw[15] ,
    \top_I.branch[10].block[15].um_I.iw[14] ,
    \top_I.branch[10].block[15].um_I.iw[13] ,
    \top_I.branch[10].block[15].um_I.iw[12] ,
    \top_I.branch[10].block[15].um_I.iw[11] ,
    \top_I.branch[10].block[15].um_I.iw[10] ,
    \top_I.branch[10].block[15].um_I.iw[9] ,
    \top_I.branch[10].block[15].um_I.iw[8] ,
    \top_I.branch[10].block[15].um_I.iw[7] ,
    \top_I.branch[10].block[15].um_I.iw[6] ,
    \top_I.branch[10].block[15].um_I.iw[5] ,
    \top_I.branch[10].block[15].um_I.iw[4] ,
    \top_I.branch[10].block[15].um_I.iw[3] ,
    \top_I.branch[10].block[15].um_I.iw[2] ,
    \top_I.branch[10].block[15].um_I.iw[1] ,
    \top_I.branch[10].block[15].um_I.clk ,
    \top_I.branch[10].block[14].um_I.iw[17] ,
    \top_I.branch[10].block[14].um_I.iw[16] ,
    \top_I.branch[10].block[14].um_I.iw[15] ,
    \top_I.branch[10].block[14].um_I.iw[14] ,
    \top_I.branch[10].block[14].um_I.iw[13] ,
    \top_I.branch[10].block[14].um_I.iw[12] ,
    \top_I.branch[10].block[14].um_I.iw[11] ,
    \top_I.branch[10].block[14].um_I.iw[10] ,
    \top_I.branch[10].block[14].um_I.iw[9] ,
    \top_I.branch[10].block[14].um_I.iw[8] ,
    \top_I.branch[10].block[14].um_I.iw[7] ,
    \top_I.branch[10].block[14].um_I.iw[6] ,
    \top_I.branch[10].block[14].um_I.iw[5] ,
    \top_I.branch[10].block[14].um_I.iw[4] ,
    \top_I.branch[10].block[14].um_I.iw[3] ,
    \top_I.branch[10].block[14].um_I.iw[2] ,
    \top_I.branch[10].block[14].um_I.iw[1] ,
    \top_I.branch[10].block[14].um_I.clk ,
    \top_I.branch[10].block[13].um_I.iw[17] ,
    \top_I.branch[10].block[13].um_I.iw[16] ,
    \top_I.branch[10].block[13].um_I.iw[15] ,
    \top_I.branch[10].block[13].um_I.iw[14] ,
    \top_I.branch[10].block[13].um_I.iw[13] ,
    \top_I.branch[10].block[13].um_I.iw[12] ,
    \top_I.branch[10].block[13].um_I.iw[11] ,
    \top_I.branch[10].block[13].um_I.iw[10] ,
    \top_I.branch[10].block[13].um_I.iw[9] ,
    \top_I.branch[10].block[13].um_I.iw[8] ,
    \top_I.branch[10].block[13].um_I.iw[7] ,
    \top_I.branch[10].block[13].um_I.iw[6] ,
    \top_I.branch[10].block[13].um_I.iw[5] ,
    \top_I.branch[10].block[13].um_I.iw[4] ,
    \top_I.branch[10].block[13].um_I.iw[3] ,
    \top_I.branch[10].block[13].um_I.iw[2] ,
    \top_I.branch[10].block[13].um_I.iw[1] ,
    \top_I.branch[10].block[13].um_I.clk ,
    \top_I.branch[10].block[12].um_I.iw[17] ,
    \top_I.branch[10].block[12].um_I.iw[16] ,
    \top_I.branch[10].block[12].um_I.iw[15] ,
    \top_I.branch[10].block[12].um_I.iw[14] ,
    \top_I.branch[10].block[12].um_I.iw[13] ,
    \top_I.branch[10].block[12].um_I.iw[12] ,
    \top_I.branch[10].block[12].um_I.iw[11] ,
    \top_I.branch[10].block[12].um_I.iw[10] ,
    \top_I.branch[10].block[12].um_I.iw[9] ,
    \top_I.branch[10].block[12].um_I.iw[8] ,
    \top_I.branch[10].block[12].um_I.iw[7] ,
    \top_I.branch[10].block[12].um_I.iw[6] ,
    \top_I.branch[10].block[12].um_I.iw[5] ,
    \top_I.branch[10].block[12].um_I.iw[4] ,
    \top_I.branch[10].block[12].um_I.iw[3] ,
    \top_I.branch[10].block[12].um_I.iw[2] ,
    \top_I.branch[10].block[12].um_I.iw[1] ,
    \top_I.branch[10].block[12].um_I.clk ,
    \top_I.branch[10].block[11].um_I.iw[17] ,
    \top_I.branch[10].block[11].um_I.iw[16] ,
    \top_I.branch[10].block[11].um_I.iw[15] ,
    \top_I.branch[10].block[11].um_I.iw[14] ,
    \top_I.branch[10].block[11].um_I.iw[13] ,
    \top_I.branch[10].block[11].um_I.iw[12] ,
    \top_I.branch[10].block[11].um_I.iw[11] ,
    \top_I.branch[10].block[11].um_I.iw[10] ,
    \top_I.branch[10].block[11].um_I.iw[9] ,
    \top_I.branch[10].block[11].um_I.iw[8] ,
    \top_I.branch[10].block[11].um_I.iw[7] ,
    \top_I.branch[10].block[11].um_I.iw[6] ,
    \top_I.branch[10].block[11].um_I.iw[5] ,
    \top_I.branch[10].block[11].um_I.iw[4] ,
    \top_I.branch[10].block[11].um_I.iw[3] ,
    \top_I.branch[10].block[11].um_I.iw[2] ,
    \top_I.branch[10].block[11].um_I.iw[1] ,
    \top_I.branch[10].block[11].um_I.clk ,
    \top_I.branch[10].block[10].um_I.iw[17] ,
    \top_I.branch[10].block[10].um_I.iw[16] ,
    \top_I.branch[10].block[10].um_I.iw[15] ,
    \top_I.branch[10].block[10].um_I.iw[14] ,
    \top_I.branch[10].block[10].um_I.iw[13] ,
    \top_I.branch[10].block[10].um_I.iw[12] ,
    \top_I.branch[10].block[10].um_I.iw[11] ,
    \top_I.branch[10].block[10].um_I.iw[10] ,
    \top_I.branch[10].block[10].um_I.iw[9] ,
    \top_I.branch[10].block[10].um_I.iw[8] ,
    \top_I.branch[10].block[10].um_I.iw[7] ,
    \top_I.branch[10].block[10].um_I.iw[6] ,
    \top_I.branch[10].block[10].um_I.iw[5] ,
    \top_I.branch[10].block[10].um_I.iw[4] ,
    \top_I.branch[10].block[10].um_I.iw[3] ,
    \top_I.branch[10].block[10].um_I.iw[2] ,
    \top_I.branch[10].block[10].um_I.iw[1] ,
    \top_I.branch[10].block[10].um_I.clk ,
    \top_I.branch[10].block[9].um_I.iw[17] ,
    \top_I.branch[10].block[9].um_I.iw[16] ,
    \top_I.branch[10].block[9].um_I.iw[15] ,
    \top_I.branch[10].block[9].um_I.iw[14] ,
    \top_I.branch[10].block[9].um_I.iw[13] ,
    \top_I.branch[10].block[9].um_I.iw[12] ,
    \top_I.branch[10].block[9].um_I.iw[11] ,
    \top_I.branch[10].block[9].um_I.iw[10] ,
    \top_I.branch[10].block[9].um_I.iw[9] ,
    \top_I.branch[10].block[9].um_I.iw[8] ,
    \top_I.branch[10].block[9].um_I.iw[7] ,
    \top_I.branch[10].block[9].um_I.iw[6] ,
    \top_I.branch[10].block[9].um_I.iw[5] ,
    \top_I.branch[10].block[9].um_I.iw[4] ,
    \top_I.branch[10].block[9].um_I.iw[3] ,
    \top_I.branch[10].block[9].um_I.iw[2] ,
    \top_I.branch[10].block[9].um_I.iw[1] ,
    \top_I.branch[10].block[9].um_I.clk ,
    \top_I.branch[10].block[8].um_I.iw[17] ,
    \top_I.branch[10].block[8].um_I.iw[16] ,
    \top_I.branch[10].block[8].um_I.iw[15] ,
    \top_I.branch[10].block[8].um_I.iw[14] ,
    \top_I.branch[10].block[8].um_I.iw[13] ,
    \top_I.branch[10].block[8].um_I.iw[12] ,
    \top_I.branch[10].block[8].um_I.iw[11] ,
    \top_I.branch[10].block[8].um_I.iw[10] ,
    \top_I.branch[10].block[8].um_I.iw[9] ,
    \top_I.branch[10].block[8].um_I.iw[8] ,
    \top_I.branch[10].block[8].um_I.iw[7] ,
    \top_I.branch[10].block[8].um_I.iw[6] ,
    \top_I.branch[10].block[8].um_I.iw[5] ,
    \top_I.branch[10].block[8].um_I.iw[4] ,
    \top_I.branch[10].block[8].um_I.iw[3] ,
    \top_I.branch[10].block[8].um_I.iw[2] ,
    \top_I.branch[10].block[8].um_I.iw[1] ,
    \top_I.branch[10].block[8].um_I.clk ,
    \top_I.branch[10].block[7].um_I.iw[17] ,
    \top_I.branch[10].block[7].um_I.iw[16] ,
    \top_I.branch[10].block[7].um_I.iw[15] ,
    \top_I.branch[10].block[7].um_I.iw[14] ,
    \top_I.branch[10].block[7].um_I.iw[13] ,
    \top_I.branch[10].block[7].um_I.iw[12] ,
    \top_I.branch[10].block[7].um_I.iw[11] ,
    \top_I.branch[10].block[7].um_I.iw[10] ,
    \top_I.branch[10].block[7].um_I.iw[9] ,
    \top_I.branch[10].block[7].um_I.iw[8] ,
    \top_I.branch[10].block[7].um_I.iw[7] ,
    \top_I.branch[10].block[7].um_I.iw[6] ,
    \top_I.branch[10].block[7].um_I.iw[5] ,
    \top_I.branch[10].block[7].um_I.iw[4] ,
    \top_I.branch[10].block[7].um_I.iw[3] ,
    \top_I.branch[10].block[7].um_I.iw[2] ,
    \top_I.branch[10].block[7].um_I.iw[1] ,
    \top_I.branch[10].block[7].um_I.clk ,
    \top_I.branch[10].block[6].um_I.iw[17] ,
    \top_I.branch[10].block[6].um_I.iw[16] ,
    \top_I.branch[10].block[6].um_I.iw[15] ,
    \top_I.branch[10].block[6].um_I.iw[14] ,
    \top_I.branch[10].block[6].um_I.iw[13] ,
    \top_I.branch[10].block[6].um_I.iw[12] ,
    \top_I.branch[10].block[6].um_I.iw[11] ,
    \top_I.branch[10].block[6].um_I.iw[10] ,
    \top_I.branch[10].block[6].um_I.iw[9] ,
    \top_I.branch[10].block[6].um_I.iw[8] ,
    \top_I.branch[10].block[6].um_I.iw[7] ,
    \top_I.branch[10].block[6].um_I.iw[6] ,
    \top_I.branch[10].block[6].um_I.iw[5] ,
    \top_I.branch[10].block[6].um_I.iw[4] ,
    \top_I.branch[10].block[6].um_I.iw[3] ,
    \top_I.branch[10].block[6].um_I.iw[2] ,
    \top_I.branch[10].block[6].um_I.iw[1] ,
    \top_I.branch[10].block[6].um_I.clk ,
    \top_I.branch[10].block[5].um_I.iw[17] ,
    \top_I.branch[10].block[5].um_I.iw[16] ,
    \top_I.branch[10].block[5].um_I.iw[15] ,
    \top_I.branch[10].block[5].um_I.iw[14] ,
    \top_I.branch[10].block[5].um_I.iw[13] ,
    \top_I.branch[10].block[5].um_I.iw[12] ,
    \top_I.branch[10].block[5].um_I.iw[11] ,
    \top_I.branch[10].block[5].um_I.iw[10] ,
    \top_I.branch[10].block[5].um_I.iw[9] ,
    \top_I.branch[10].block[5].um_I.iw[8] ,
    \top_I.branch[10].block[5].um_I.iw[7] ,
    \top_I.branch[10].block[5].um_I.iw[6] ,
    \top_I.branch[10].block[5].um_I.iw[5] ,
    \top_I.branch[10].block[5].um_I.iw[4] ,
    \top_I.branch[10].block[5].um_I.iw[3] ,
    \top_I.branch[10].block[5].um_I.iw[2] ,
    \top_I.branch[10].block[5].um_I.iw[1] ,
    \top_I.branch[10].block[5].um_I.clk ,
    \top_I.branch[10].block[4].um_I.iw[17] ,
    \top_I.branch[10].block[4].um_I.iw[16] ,
    \top_I.branch[10].block[4].um_I.iw[15] ,
    \top_I.branch[10].block[4].um_I.iw[14] ,
    \top_I.branch[10].block[4].um_I.iw[13] ,
    \top_I.branch[10].block[4].um_I.iw[12] ,
    \top_I.branch[10].block[4].um_I.iw[11] ,
    \top_I.branch[10].block[4].um_I.iw[10] ,
    \top_I.branch[10].block[4].um_I.iw[9] ,
    \top_I.branch[10].block[4].um_I.iw[8] ,
    \top_I.branch[10].block[4].um_I.iw[7] ,
    \top_I.branch[10].block[4].um_I.iw[6] ,
    \top_I.branch[10].block[4].um_I.iw[5] ,
    \top_I.branch[10].block[4].um_I.iw[4] ,
    \top_I.branch[10].block[4].um_I.iw[3] ,
    \top_I.branch[10].block[4].um_I.iw[2] ,
    \top_I.branch[10].block[4].um_I.iw[1] ,
    \top_I.branch[10].block[4].um_I.clk ,
    \top_I.branch[10].block[3].um_I.iw[17] ,
    \top_I.branch[10].block[3].um_I.iw[16] ,
    \top_I.branch[10].block[3].um_I.iw[15] ,
    \top_I.branch[10].block[3].um_I.iw[14] ,
    \top_I.branch[10].block[3].um_I.iw[13] ,
    \top_I.branch[10].block[3].um_I.iw[12] ,
    \top_I.branch[10].block[3].um_I.iw[11] ,
    \top_I.branch[10].block[3].um_I.iw[10] ,
    \top_I.branch[10].block[3].um_I.iw[9] ,
    \top_I.branch[10].block[3].um_I.iw[8] ,
    \top_I.branch[10].block[3].um_I.iw[7] ,
    \top_I.branch[10].block[3].um_I.iw[6] ,
    \top_I.branch[10].block[3].um_I.iw[5] ,
    \top_I.branch[10].block[3].um_I.iw[4] ,
    \top_I.branch[10].block[3].um_I.iw[3] ,
    \top_I.branch[10].block[3].um_I.iw[2] ,
    \top_I.branch[10].block[3].um_I.iw[1] ,
    \top_I.branch[10].block[3].um_I.clk ,
    \top_I.branch[10].block[2].um_I.iw[17] ,
    \top_I.branch[10].block[2].um_I.iw[16] ,
    \top_I.branch[10].block[2].um_I.iw[15] ,
    \top_I.branch[10].block[2].um_I.iw[14] ,
    \top_I.branch[10].block[2].um_I.iw[13] ,
    \top_I.branch[10].block[2].um_I.iw[12] ,
    \top_I.branch[10].block[2].um_I.iw[11] ,
    \top_I.branch[10].block[2].um_I.iw[10] ,
    \top_I.branch[10].block[2].um_I.iw[9] ,
    \top_I.branch[10].block[2].um_I.iw[8] ,
    \top_I.branch[10].block[2].um_I.iw[7] ,
    \top_I.branch[10].block[2].um_I.iw[6] ,
    \top_I.branch[10].block[2].um_I.iw[5] ,
    \top_I.branch[10].block[2].um_I.iw[4] ,
    \top_I.branch[10].block[2].um_I.iw[3] ,
    \top_I.branch[10].block[2].um_I.iw[2] ,
    \top_I.branch[10].block[2].um_I.iw[1] ,
    \top_I.branch[10].block[2].um_I.clk ,
    \top_I.branch[10].block[1].um_I.iw[17] ,
    \top_I.branch[10].block[1].um_I.iw[16] ,
    \top_I.branch[10].block[1].um_I.iw[15] ,
    \top_I.branch[10].block[1].um_I.iw[14] ,
    \top_I.branch[10].block[1].um_I.iw[13] ,
    \top_I.branch[10].block[1].um_I.iw[12] ,
    \top_I.branch[10].block[1].um_I.iw[11] ,
    \top_I.branch[10].block[1].um_I.iw[10] ,
    \top_I.branch[10].block[1].um_I.iw[9] ,
    \top_I.branch[10].block[1].um_I.iw[8] ,
    \top_I.branch[10].block[1].um_I.iw[7] ,
    \top_I.branch[10].block[1].um_I.iw[6] ,
    \top_I.branch[10].block[1].um_I.iw[5] ,
    \top_I.branch[10].block[1].um_I.iw[4] ,
    \top_I.branch[10].block[1].um_I.iw[3] ,
    \top_I.branch[10].block[1].um_I.iw[2] ,
    \top_I.branch[10].block[1].um_I.iw[1] ,
    \top_I.branch[10].block[1].um_I.clk ,
    \top_I.branch[10].block[0].um_I.iw[17] ,
    \top_I.branch[10].block[0].um_I.iw[16] ,
    \top_I.branch[10].block[0].um_I.iw[15] ,
    \top_I.branch[10].block[0].um_I.iw[14] ,
    \top_I.branch[10].block[0].um_I.iw[13] ,
    \top_I.branch[10].block[0].um_I.iw[12] ,
    \top_I.branch[10].block[0].um_I.iw[11] ,
    \top_I.branch[10].block[0].um_I.iw[10] ,
    \top_I.branch[10].block[0].um_I.iw[9] ,
    \top_I.branch[10].block[0].um_I.iw[8] ,
    \top_I.branch[10].block[0].um_I.iw[7] ,
    \top_I.branch[10].block[0].um_I.iw[6] ,
    \top_I.branch[10].block[0].um_I.iw[5] ,
    \top_I.branch[10].block[0].um_I.iw[4] ,
    \top_I.branch[10].block[0].um_I.iw[3] ,
    \top_I.branch[10].block[0].um_I.iw[2] ,
    \top_I.branch[10].block[0].um_I.iw[1] ,
    \top_I.branch[10].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[10].block[15].um_I.pg_vdd ,
    \top_I.branch[10].block[14].um_I.pg_vdd ,
    \top_I.branch[10].block[13].um_I.pg_vdd ,
    \top_I.branch[10].block[12].um_I.pg_vdd ,
    \top_I.branch[10].block[11].um_I.pg_vdd ,
    \top_I.branch[10].block[10].um_I.pg_vdd ,
    \top_I.branch[10].block[9].um_I.pg_vdd ,
    \top_I.branch[10].block[8].um_I.pg_vdd ,
    \top_I.branch[10].block[7].um_I.pg_vdd ,
    \top_I.branch[10].block[6].um_I.pg_vdd ,
    \top_I.branch[10].block[5].um_I.pg_vdd ,
    \top_I.branch[10].block[4].um_I.pg_vdd ,
    \top_I.branch[10].block[3].um_I.pg_vdd ,
    \top_I.branch[10].block[2].um_I.pg_vdd ,
    \top_I.branch[10].block[1].um_I.pg_vdd ,
    \top_I.branch[10].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[11].mux_I  (.k_one(\top_I.branch[11].l_addr[0] ),
    .k_zero(\top_I.branch[11].l_addr[1] ),
    .addr({\top_I.branch[11].l_addr[1] ,
    \top_I.branch[11].l_addr[0] ,
    \top_I.branch[11].l_addr[1] ,
    \top_I.branch[11].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[11].block[15].um_I.ena ,
    \top_I.branch[11].block[14].um_I.ena ,
    \top_I.branch[11].block[13].um_I.ena ,
    \top_I.branch[11].block[12].um_I.ena ,
    \top_I.branch[11].block[11].um_I.ena ,
    \top_I.branch[11].block[10].um_I.ena ,
    \top_I.branch[11].block[9].um_I.ena ,
    \top_I.branch[11].block[8].um_I.ena ,
    \top_I.branch[11].block[7].um_I.ena ,
    \top_I.branch[11].block[6].um_I.ena ,
    \top_I.branch[11].block[5].um_I.ena ,
    \top_I.branch[11].block[4].um_I.ena ,
    \top_I.branch[11].block[3].um_I.ena ,
    \top_I.branch[11].block[2].um_I.ena ,
    \top_I.branch[11].block[1].um_I.ena ,
    \top_I.branch[11].block[0].um_I.ena }),
    .um_iw({\top_I.branch[11].block[15].um_I.iw[17] ,
    \top_I.branch[11].block[15].um_I.iw[16] ,
    \top_I.branch[11].block[15].um_I.iw[15] ,
    \top_I.branch[11].block[15].um_I.iw[14] ,
    \top_I.branch[11].block[15].um_I.iw[13] ,
    \top_I.branch[11].block[15].um_I.iw[12] ,
    \top_I.branch[11].block[15].um_I.iw[11] ,
    \top_I.branch[11].block[15].um_I.iw[10] ,
    \top_I.branch[11].block[15].um_I.iw[9] ,
    \top_I.branch[11].block[15].um_I.iw[8] ,
    \top_I.branch[11].block[15].um_I.iw[7] ,
    \top_I.branch[11].block[15].um_I.iw[6] ,
    \top_I.branch[11].block[15].um_I.iw[5] ,
    \top_I.branch[11].block[15].um_I.iw[4] ,
    \top_I.branch[11].block[15].um_I.iw[3] ,
    \top_I.branch[11].block[15].um_I.iw[2] ,
    \top_I.branch[11].block[15].um_I.iw[1] ,
    \top_I.branch[11].block[15].um_I.clk ,
    \top_I.branch[11].block[14].um_I.iw[17] ,
    \top_I.branch[11].block[14].um_I.iw[16] ,
    \top_I.branch[11].block[14].um_I.iw[15] ,
    \top_I.branch[11].block[14].um_I.iw[14] ,
    \top_I.branch[11].block[14].um_I.iw[13] ,
    \top_I.branch[11].block[14].um_I.iw[12] ,
    \top_I.branch[11].block[14].um_I.iw[11] ,
    \top_I.branch[11].block[14].um_I.iw[10] ,
    \top_I.branch[11].block[14].um_I.iw[9] ,
    \top_I.branch[11].block[14].um_I.iw[8] ,
    \top_I.branch[11].block[14].um_I.iw[7] ,
    \top_I.branch[11].block[14].um_I.iw[6] ,
    \top_I.branch[11].block[14].um_I.iw[5] ,
    \top_I.branch[11].block[14].um_I.iw[4] ,
    \top_I.branch[11].block[14].um_I.iw[3] ,
    \top_I.branch[11].block[14].um_I.iw[2] ,
    \top_I.branch[11].block[14].um_I.iw[1] ,
    \top_I.branch[11].block[14].um_I.clk ,
    \top_I.branch[11].block[13].um_I.iw[17] ,
    \top_I.branch[11].block[13].um_I.iw[16] ,
    \top_I.branch[11].block[13].um_I.iw[15] ,
    \top_I.branch[11].block[13].um_I.iw[14] ,
    \top_I.branch[11].block[13].um_I.iw[13] ,
    \top_I.branch[11].block[13].um_I.iw[12] ,
    \top_I.branch[11].block[13].um_I.iw[11] ,
    \top_I.branch[11].block[13].um_I.iw[10] ,
    \top_I.branch[11].block[13].um_I.iw[9] ,
    \top_I.branch[11].block[13].um_I.iw[8] ,
    \top_I.branch[11].block[13].um_I.iw[7] ,
    \top_I.branch[11].block[13].um_I.iw[6] ,
    \top_I.branch[11].block[13].um_I.iw[5] ,
    \top_I.branch[11].block[13].um_I.iw[4] ,
    \top_I.branch[11].block[13].um_I.iw[3] ,
    \top_I.branch[11].block[13].um_I.iw[2] ,
    \top_I.branch[11].block[13].um_I.iw[1] ,
    \top_I.branch[11].block[13].um_I.clk ,
    \top_I.branch[11].block[12].um_I.iw[17] ,
    \top_I.branch[11].block[12].um_I.iw[16] ,
    \top_I.branch[11].block[12].um_I.iw[15] ,
    \top_I.branch[11].block[12].um_I.iw[14] ,
    \top_I.branch[11].block[12].um_I.iw[13] ,
    \top_I.branch[11].block[12].um_I.iw[12] ,
    \top_I.branch[11].block[12].um_I.iw[11] ,
    \top_I.branch[11].block[12].um_I.iw[10] ,
    \top_I.branch[11].block[12].um_I.iw[9] ,
    \top_I.branch[11].block[12].um_I.iw[8] ,
    \top_I.branch[11].block[12].um_I.iw[7] ,
    \top_I.branch[11].block[12].um_I.iw[6] ,
    \top_I.branch[11].block[12].um_I.iw[5] ,
    \top_I.branch[11].block[12].um_I.iw[4] ,
    \top_I.branch[11].block[12].um_I.iw[3] ,
    \top_I.branch[11].block[12].um_I.iw[2] ,
    \top_I.branch[11].block[12].um_I.iw[1] ,
    \top_I.branch[11].block[12].um_I.clk ,
    \top_I.branch[11].block[11].um_I.iw[17] ,
    \top_I.branch[11].block[11].um_I.iw[16] ,
    \top_I.branch[11].block[11].um_I.iw[15] ,
    \top_I.branch[11].block[11].um_I.iw[14] ,
    \top_I.branch[11].block[11].um_I.iw[13] ,
    \top_I.branch[11].block[11].um_I.iw[12] ,
    \top_I.branch[11].block[11].um_I.iw[11] ,
    \top_I.branch[11].block[11].um_I.iw[10] ,
    \top_I.branch[11].block[11].um_I.iw[9] ,
    \top_I.branch[11].block[11].um_I.iw[8] ,
    \top_I.branch[11].block[11].um_I.iw[7] ,
    \top_I.branch[11].block[11].um_I.iw[6] ,
    \top_I.branch[11].block[11].um_I.iw[5] ,
    \top_I.branch[11].block[11].um_I.iw[4] ,
    \top_I.branch[11].block[11].um_I.iw[3] ,
    \top_I.branch[11].block[11].um_I.iw[2] ,
    \top_I.branch[11].block[11].um_I.iw[1] ,
    \top_I.branch[11].block[11].um_I.clk ,
    \top_I.branch[11].block[10].um_I.iw[17] ,
    \top_I.branch[11].block[10].um_I.iw[16] ,
    \top_I.branch[11].block[10].um_I.iw[15] ,
    \top_I.branch[11].block[10].um_I.iw[14] ,
    \top_I.branch[11].block[10].um_I.iw[13] ,
    \top_I.branch[11].block[10].um_I.iw[12] ,
    \top_I.branch[11].block[10].um_I.iw[11] ,
    \top_I.branch[11].block[10].um_I.iw[10] ,
    \top_I.branch[11].block[10].um_I.iw[9] ,
    \top_I.branch[11].block[10].um_I.iw[8] ,
    \top_I.branch[11].block[10].um_I.iw[7] ,
    \top_I.branch[11].block[10].um_I.iw[6] ,
    \top_I.branch[11].block[10].um_I.iw[5] ,
    \top_I.branch[11].block[10].um_I.iw[4] ,
    \top_I.branch[11].block[10].um_I.iw[3] ,
    \top_I.branch[11].block[10].um_I.iw[2] ,
    \top_I.branch[11].block[10].um_I.iw[1] ,
    \top_I.branch[11].block[10].um_I.clk ,
    \top_I.branch[11].block[9].um_I.iw[17] ,
    \top_I.branch[11].block[9].um_I.iw[16] ,
    \top_I.branch[11].block[9].um_I.iw[15] ,
    \top_I.branch[11].block[9].um_I.iw[14] ,
    \top_I.branch[11].block[9].um_I.iw[13] ,
    \top_I.branch[11].block[9].um_I.iw[12] ,
    \top_I.branch[11].block[9].um_I.iw[11] ,
    \top_I.branch[11].block[9].um_I.iw[10] ,
    \top_I.branch[11].block[9].um_I.iw[9] ,
    \top_I.branch[11].block[9].um_I.iw[8] ,
    \top_I.branch[11].block[9].um_I.iw[7] ,
    \top_I.branch[11].block[9].um_I.iw[6] ,
    \top_I.branch[11].block[9].um_I.iw[5] ,
    \top_I.branch[11].block[9].um_I.iw[4] ,
    \top_I.branch[11].block[9].um_I.iw[3] ,
    \top_I.branch[11].block[9].um_I.iw[2] ,
    \top_I.branch[11].block[9].um_I.iw[1] ,
    \top_I.branch[11].block[9].um_I.clk ,
    \top_I.branch[11].block[8].um_I.iw[17] ,
    \top_I.branch[11].block[8].um_I.iw[16] ,
    \top_I.branch[11].block[8].um_I.iw[15] ,
    \top_I.branch[11].block[8].um_I.iw[14] ,
    \top_I.branch[11].block[8].um_I.iw[13] ,
    \top_I.branch[11].block[8].um_I.iw[12] ,
    \top_I.branch[11].block[8].um_I.iw[11] ,
    \top_I.branch[11].block[8].um_I.iw[10] ,
    \top_I.branch[11].block[8].um_I.iw[9] ,
    \top_I.branch[11].block[8].um_I.iw[8] ,
    \top_I.branch[11].block[8].um_I.iw[7] ,
    \top_I.branch[11].block[8].um_I.iw[6] ,
    \top_I.branch[11].block[8].um_I.iw[5] ,
    \top_I.branch[11].block[8].um_I.iw[4] ,
    \top_I.branch[11].block[8].um_I.iw[3] ,
    \top_I.branch[11].block[8].um_I.iw[2] ,
    \top_I.branch[11].block[8].um_I.iw[1] ,
    \top_I.branch[11].block[8].um_I.clk ,
    \top_I.branch[11].block[7].um_I.iw[17] ,
    \top_I.branch[11].block[7].um_I.iw[16] ,
    \top_I.branch[11].block[7].um_I.iw[15] ,
    \top_I.branch[11].block[7].um_I.iw[14] ,
    \top_I.branch[11].block[7].um_I.iw[13] ,
    \top_I.branch[11].block[7].um_I.iw[12] ,
    \top_I.branch[11].block[7].um_I.iw[11] ,
    \top_I.branch[11].block[7].um_I.iw[10] ,
    \top_I.branch[11].block[7].um_I.iw[9] ,
    \top_I.branch[11].block[7].um_I.iw[8] ,
    \top_I.branch[11].block[7].um_I.iw[7] ,
    \top_I.branch[11].block[7].um_I.iw[6] ,
    \top_I.branch[11].block[7].um_I.iw[5] ,
    \top_I.branch[11].block[7].um_I.iw[4] ,
    \top_I.branch[11].block[7].um_I.iw[3] ,
    \top_I.branch[11].block[7].um_I.iw[2] ,
    \top_I.branch[11].block[7].um_I.iw[1] ,
    \top_I.branch[11].block[7].um_I.clk ,
    \top_I.branch[11].block[6].um_I.iw[17] ,
    \top_I.branch[11].block[6].um_I.iw[16] ,
    \top_I.branch[11].block[6].um_I.iw[15] ,
    \top_I.branch[11].block[6].um_I.iw[14] ,
    \top_I.branch[11].block[6].um_I.iw[13] ,
    \top_I.branch[11].block[6].um_I.iw[12] ,
    \top_I.branch[11].block[6].um_I.iw[11] ,
    \top_I.branch[11].block[6].um_I.iw[10] ,
    \top_I.branch[11].block[6].um_I.iw[9] ,
    \top_I.branch[11].block[6].um_I.iw[8] ,
    \top_I.branch[11].block[6].um_I.iw[7] ,
    \top_I.branch[11].block[6].um_I.iw[6] ,
    \top_I.branch[11].block[6].um_I.iw[5] ,
    \top_I.branch[11].block[6].um_I.iw[4] ,
    \top_I.branch[11].block[6].um_I.iw[3] ,
    \top_I.branch[11].block[6].um_I.iw[2] ,
    \top_I.branch[11].block[6].um_I.iw[1] ,
    \top_I.branch[11].block[6].um_I.clk ,
    \top_I.branch[11].block[5].um_I.iw[17] ,
    \top_I.branch[11].block[5].um_I.iw[16] ,
    \top_I.branch[11].block[5].um_I.iw[15] ,
    \top_I.branch[11].block[5].um_I.iw[14] ,
    \top_I.branch[11].block[5].um_I.iw[13] ,
    \top_I.branch[11].block[5].um_I.iw[12] ,
    \top_I.branch[11].block[5].um_I.iw[11] ,
    \top_I.branch[11].block[5].um_I.iw[10] ,
    \top_I.branch[11].block[5].um_I.iw[9] ,
    \top_I.branch[11].block[5].um_I.iw[8] ,
    \top_I.branch[11].block[5].um_I.iw[7] ,
    \top_I.branch[11].block[5].um_I.iw[6] ,
    \top_I.branch[11].block[5].um_I.iw[5] ,
    \top_I.branch[11].block[5].um_I.iw[4] ,
    \top_I.branch[11].block[5].um_I.iw[3] ,
    \top_I.branch[11].block[5].um_I.iw[2] ,
    \top_I.branch[11].block[5].um_I.iw[1] ,
    \top_I.branch[11].block[5].um_I.clk ,
    \top_I.branch[11].block[4].um_I.iw[17] ,
    \top_I.branch[11].block[4].um_I.iw[16] ,
    \top_I.branch[11].block[4].um_I.iw[15] ,
    \top_I.branch[11].block[4].um_I.iw[14] ,
    \top_I.branch[11].block[4].um_I.iw[13] ,
    \top_I.branch[11].block[4].um_I.iw[12] ,
    \top_I.branch[11].block[4].um_I.iw[11] ,
    \top_I.branch[11].block[4].um_I.iw[10] ,
    \top_I.branch[11].block[4].um_I.iw[9] ,
    \top_I.branch[11].block[4].um_I.iw[8] ,
    \top_I.branch[11].block[4].um_I.iw[7] ,
    \top_I.branch[11].block[4].um_I.iw[6] ,
    \top_I.branch[11].block[4].um_I.iw[5] ,
    \top_I.branch[11].block[4].um_I.iw[4] ,
    \top_I.branch[11].block[4].um_I.iw[3] ,
    \top_I.branch[11].block[4].um_I.iw[2] ,
    \top_I.branch[11].block[4].um_I.iw[1] ,
    \top_I.branch[11].block[4].um_I.clk ,
    \top_I.branch[11].block[3].um_I.iw[17] ,
    \top_I.branch[11].block[3].um_I.iw[16] ,
    \top_I.branch[11].block[3].um_I.iw[15] ,
    \top_I.branch[11].block[3].um_I.iw[14] ,
    \top_I.branch[11].block[3].um_I.iw[13] ,
    \top_I.branch[11].block[3].um_I.iw[12] ,
    \top_I.branch[11].block[3].um_I.iw[11] ,
    \top_I.branch[11].block[3].um_I.iw[10] ,
    \top_I.branch[11].block[3].um_I.iw[9] ,
    \top_I.branch[11].block[3].um_I.iw[8] ,
    \top_I.branch[11].block[3].um_I.iw[7] ,
    \top_I.branch[11].block[3].um_I.iw[6] ,
    \top_I.branch[11].block[3].um_I.iw[5] ,
    \top_I.branch[11].block[3].um_I.iw[4] ,
    \top_I.branch[11].block[3].um_I.iw[3] ,
    \top_I.branch[11].block[3].um_I.iw[2] ,
    \top_I.branch[11].block[3].um_I.iw[1] ,
    \top_I.branch[11].block[3].um_I.clk ,
    \top_I.branch[11].block[2].um_I.iw[17] ,
    \top_I.branch[11].block[2].um_I.iw[16] ,
    \top_I.branch[11].block[2].um_I.iw[15] ,
    \top_I.branch[11].block[2].um_I.iw[14] ,
    \top_I.branch[11].block[2].um_I.iw[13] ,
    \top_I.branch[11].block[2].um_I.iw[12] ,
    \top_I.branch[11].block[2].um_I.iw[11] ,
    \top_I.branch[11].block[2].um_I.iw[10] ,
    \top_I.branch[11].block[2].um_I.iw[9] ,
    \top_I.branch[11].block[2].um_I.iw[8] ,
    \top_I.branch[11].block[2].um_I.iw[7] ,
    \top_I.branch[11].block[2].um_I.iw[6] ,
    \top_I.branch[11].block[2].um_I.iw[5] ,
    \top_I.branch[11].block[2].um_I.iw[4] ,
    \top_I.branch[11].block[2].um_I.iw[3] ,
    \top_I.branch[11].block[2].um_I.iw[2] ,
    \top_I.branch[11].block[2].um_I.iw[1] ,
    \top_I.branch[11].block[2].um_I.clk ,
    \top_I.branch[11].block[1].um_I.iw[17] ,
    \top_I.branch[11].block[1].um_I.iw[16] ,
    \top_I.branch[11].block[1].um_I.iw[15] ,
    \top_I.branch[11].block[1].um_I.iw[14] ,
    \top_I.branch[11].block[1].um_I.iw[13] ,
    \top_I.branch[11].block[1].um_I.iw[12] ,
    \top_I.branch[11].block[1].um_I.iw[11] ,
    \top_I.branch[11].block[1].um_I.iw[10] ,
    \top_I.branch[11].block[1].um_I.iw[9] ,
    \top_I.branch[11].block[1].um_I.iw[8] ,
    \top_I.branch[11].block[1].um_I.iw[7] ,
    \top_I.branch[11].block[1].um_I.iw[6] ,
    \top_I.branch[11].block[1].um_I.iw[5] ,
    \top_I.branch[11].block[1].um_I.iw[4] ,
    \top_I.branch[11].block[1].um_I.iw[3] ,
    \top_I.branch[11].block[1].um_I.iw[2] ,
    \top_I.branch[11].block[1].um_I.iw[1] ,
    \top_I.branch[11].block[1].um_I.clk ,
    \top_I.branch[11].block[0].um_I.iw[17] ,
    \top_I.branch[11].block[0].um_I.iw[16] ,
    \top_I.branch[11].block[0].um_I.iw[15] ,
    \top_I.branch[11].block[0].um_I.iw[14] ,
    \top_I.branch[11].block[0].um_I.iw[13] ,
    \top_I.branch[11].block[0].um_I.iw[12] ,
    \top_I.branch[11].block[0].um_I.iw[11] ,
    \top_I.branch[11].block[0].um_I.iw[10] ,
    \top_I.branch[11].block[0].um_I.iw[9] ,
    \top_I.branch[11].block[0].um_I.iw[8] ,
    \top_I.branch[11].block[0].um_I.iw[7] ,
    \top_I.branch[11].block[0].um_I.iw[6] ,
    \top_I.branch[11].block[0].um_I.iw[5] ,
    \top_I.branch[11].block[0].um_I.iw[4] ,
    \top_I.branch[11].block[0].um_I.iw[3] ,
    \top_I.branch[11].block[0].um_I.iw[2] ,
    \top_I.branch[11].block[0].um_I.iw[1] ,
    \top_I.branch[11].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[11].block[15].um_I.pg_vdd ,
    \top_I.branch[11].block[14].um_I.pg_vdd ,
    \top_I.branch[11].block[13].um_I.pg_vdd ,
    \top_I.branch[11].block[12].um_I.pg_vdd ,
    \top_I.branch[11].block[11].um_I.pg_vdd ,
    \top_I.branch[11].block[10].um_I.pg_vdd ,
    \top_I.branch[11].block[9].um_I.pg_vdd ,
    \top_I.branch[11].block[8].um_I.pg_vdd ,
    \top_I.branch[11].block[7].um_I.pg_vdd ,
    \top_I.branch[11].block[6].um_I.pg_vdd ,
    \top_I.branch[11].block[5].um_I.pg_vdd ,
    \top_I.branch[11].block[4].um_I.pg_vdd ,
    \top_I.branch[11].block[3].um_I.pg_vdd ,
    \top_I.branch[11].block[2].um_I.pg_vdd ,
    \top_I.branch[11].block[1].um_I.pg_vdd ,
    \top_I.branch[11].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[12].mux_I  (.k_one(\top_I.branch[12].l_addr[1] ),
    .k_zero(\top_I.branch[12].l_addr[0] ),
    .addr({\top_I.branch[12].l_addr[0] ,
    \top_I.branch[12].l_addr[1] ,
    \top_I.branch[12].l_addr[1] ,
    \top_I.branch[12].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[12].block[15].um_I.ena ,
    \top_I.branch[12].block[14].um_I.ena ,
    \top_I.branch[12].block[13].um_I.ena ,
    \top_I.branch[12].block[12].um_I.ena ,
    \top_I.branch[12].block[11].um_I.ena ,
    \top_I.branch[12].block[10].um_I.ena ,
    \top_I.branch[12].block[9].um_I.ena ,
    \top_I.branch[12].block[8].um_I.ena ,
    \top_I.branch[12].block[7].um_I.ena ,
    \top_I.branch[12].block[6].um_I.ena ,
    \top_I.branch[12].block[5].um_I.ena ,
    \top_I.branch[12].block[4].um_I.ena ,
    \top_I.branch[12].block[3].um_I.ena ,
    \top_I.branch[12].block[2].um_I.ena ,
    \top_I.branch[12].block[1].um_I.ena ,
    \top_I.branch[12].block[0].um_I.ena }),
    .um_iw({\top_I.branch[12].block[15].um_I.iw[17] ,
    \top_I.branch[12].block[15].um_I.iw[16] ,
    \top_I.branch[12].block[15].um_I.iw[15] ,
    \top_I.branch[12].block[15].um_I.iw[14] ,
    \top_I.branch[12].block[15].um_I.iw[13] ,
    \top_I.branch[12].block[15].um_I.iw[12] ,
    \top_I.branch[12].block[15].um_I.iw[11] ,
    \top_I.branch[12].block[15].um_I.iw[10] ,
    \top_I.branch[12].block[15].um_I.iw[9] ,
    \top_I.branch[12].block[15].um_I.iw[8] ,
    \top_I.branch[12].block[15].um_I.iw[7] ,
    \top_I.branch[12].block[15].um_I.iw[6] ,
    \top_I.branch[12].block[15].um_I.iw[5] ,
    \top_I.branch[12].block[15].um_I.iw[4] ,
    \top_I.branch[12].block[15].um_I.iw[3] ,
    \top_I.branch[12].block[15].um_I.iw[2] ,
    \top_I.branch[12].block[15].um_I.iw[1] ,
    \top_I.branch[12].block[15].um_I.clk ,
    \top_I.branch[12].block[14].um_I.iw[17] ,
    \top_I.branch[12].block[14].um_I.iw[16] ,
    \top_I.branch[12].block[14].um_I.iw[15] ,
    \top_I.branch[12].block[14].um_I.iw[14] ,
    \top_I.branch[12].block[14].um_I.iw[13] ,
    \top_I.branch[12].block[14].um_I.iw[12] ,
    \top_I.branch[12].block[14].um_I.iw[11] ,
    \top_I.branch[12].block[14].um_I.iw[10] ,
    \top_I.branch[12].block[14].um_I.iw[9] ,
    \top_I.branch[12].block[14].um_I.iw[8] ,
    \top_I.branch[12].block[14].um_I.iw[7] ,
    \top_I.branch[12].block[14].um_I.iw[6] ,
    \top_I.branch[12].block[14].um_I.iw[5] ,
    \top_I.branch[12].block[14].um_I.iw[4] ,
    \top_I.branch[12].block[14].um_I.iw[3] ,
    \top_I.branch[12].block[14].um_I.iw[2] ,
    \top_I.branch[12].block[14].um_I.iw[1] ,
    \top_I.branch[12].block[14].um_I.clk ,
    \top_I.branch[12].block[13].um_I.iw[17] ,
    \top_I.branch[12].block[13].um_I.iw[16] ,
    \top_I.branch[12].block[13].um_I.iw[15] ,
    \top_I.branch[12].block[13].um_I.iw[14] ,
    \top_I.branch[12].block[13].um_I.iw[13] ,
    \top_I.branch[12].block[13].um_I.iw[12] ,
    \top_I.branch[12].block[13].um_I.iw[11] ,
    \top_I.branch[12].block[13].um_I.iw[10] ,
    \top_I.branch[12].block[13].um_I.iw[9] ,
    \top_I.branch[12].block[13].um_I.iw[8] ,
    \top_I.branch[12].block[13].um_I.iw[7] ,
    \top_I.branch[12].block[13].um_I.iw[6] ,
    \top_I.branch[12].block[13].um_I.iw[5] ,
    \top_I.branch[12].block[13].um_I.iw[4] ,
    \top_I.branch[12].block[13].um_I.iw[3] ,
    \top_I.branch[12].block[13].um_I.iw[2] ,
    \top_I.branch[12].block[13].um_I.iw[1] ,
    \top_I.branch[12].block[13].um_I.clk ,
    \top_I.branch[12].block[12].um_I.iw[17] ,
    \top_I.branch[12].block[12].um_I.iw[16] ,
    \top_I.branch[12].block[12].um_I.iw[15] ,
    \top_I.branch[12].block[12].um_I.iw[14] ,
    \top_I.branch[12].block[12].um_I.iw[13] ,
    \top_I.branch[12].block[12].um_I.iw[12] ,
    \top_I.branch[12].block[12].um_I.iw[11] ,
    \top_I.branch[12].block[12].um_I.iw[10] ,
    \top_I.branch[12].block[12].um_I.iw[9] ,
    \top_I.branch[12].block[12].um_I.iw[8] ,
    \top_I.branch[12].block[12].um_I.iw[7] ,
    \top_I.branch[12].block[12].um_I.iw[6] ,
    \top_I.branch[12].block[12].um_I.iw[5] ,
    \top_I.branch[12].block[12].um_I.iw[4] ,
    \top_I.branch[12].block[12].um_I.iw[3] ,
    \top_I.branch[12].block[12].um_I.iw[2] ,
    \top_I.branch[12].block[12].um_I.iw[1] ,
    \top_I.branch[12].block[12].um_I.clk ,
    \top_I.branch[12].block[11].um_I.iw[17] ,
    \top_I.branch[12].block[11].um_I.iw[16] ,
    \top_I.branch[12].block[11].um_I.iw[15] ,
    \top_I.branch[12].block[11].um_I.iw[14] ,
    \top_I.branch[12].block[11].um_I.iw[13] ,
    \top_I.branch[12].block[11].um_I.iw[12] ,
    \top_I.branch[12].block[11].um_I.iw[11] ,
    \top_I.branch[12].block[11].um_I.iw[10] ,
    \top_I.branch[12].block[11].um_I.iw[9] ,
    \top_I.branch[12].block[11].um_I.iw[8] ,
    \top_I.branch[12].block[11].um_I.iw[7] ,
    \top_I.branch[12].block[11].um_I.iw[6] ,
    \top_I.branch[12].block[11].um_I.iw[5] ,
    \top_I.branch[12].block[11].um_I.iw[4] ,
    \top_I.branch[12].block[11].um_I.iw[3] ,
    \top_I.branch[12].block[11].um_I.iw[2] ,
    \top_I.branch[12].block[11].um_I.iw[1] ,
    \top_I.branch[12].block[11].um_I.clk ,
    \top_I.branch[12].block[10].um_I.iw[17] ,
    \top_I.branch[12].block[10].um_I.iw[16] ,
    \top_I.branch[12].block[10].um_I.iw[15] ,
    \top_I.branch[12].block[10].um_I.iw[14] ,
    \top_I.branch[12].block[10].um_I.iw[13] ,
    \top_I.branch[12].block[10].um_I.iw[12] ,
    \top_I.branch[12].block[10].um_I.iw[11] ,
    \top_I.branch[12].block[10].um_I.iw[10] ,
    \top_I.branch[12].block[10].um_I.iw[9] ,
    \top_I.branch[12].block[10].um_I.iw[8] ,
    \top_I.branch[12].block[10].um_I.iw[7] ,
    \top_I.branch[12].block[10].um_I.iw[6] ,
    \top_I.branch[12].block[10].um_I.iw[5] ,
    \top_I.branch[12].block[10].um_I.iw[4] ,
    \top_I.branch[12].block[10].um_I.iw[3] ,
    \top_I.branch[12].block[10].um_I.iw[2] ,
    \top_I.branch[12].block[10].um_I.iw[1] ,
    \top_I.branch[12].block[10].um_I.clk ,
    \top_I.branch[12].block[9].um_I.iw[17] ,
    \top_I.branch[12].block[9].um_I.iw[16] ,
    \top_I.branch[12].block[9].um_I.iw[15] ,
    \top_I.branch[12].block[9].um_I.iw[14] ,
    \top_I.branch[12].block[9].um_I.iw[13] ,
    \top_I.branch[12].block[9].um_I.iw[12] ,
    \top_I.branch[12].block[9].um_I.iw[11] ,
    \top_I.branch[12].block[9].um_I.iw[10] ,
    \top_I.branch[12].block[9].um_I.iw[9] ,
    \top_I.branch[12].block[9].um_I.iw[8] ,
    \top_I.branch[12].block[9].um_I.iw[7] ,
    \top_I.branch[12].block[9].um_I.iw[6] ,
    \top_I.branch[12].block[9].um_I.iw[5] ,
    \top_I.branch[12].block[9].um_I.iw[4] ,
    \top_I.branch[12].block[9].um_I.iw[3] ,
    \top_I.branch[12].block[9].um_I.iw[2] ,
    \top_I.branch[12].block[9].um_I.iw[1] ,
    \top_I.branch[12].block[9].um_I.clk ,
    \top_I.branch[12].block[8].um_I.iw[17] ,
    \top_I.branch[12].block[8].um_I.iw[16] ,
    \top_I.branch[12].block[8].um_I.iw[15] ,
    \top_I.branch[12].block[8].um_I.iw[14] ,
    \top_I.branch[12].block[8].um_I.iw[13] ,
    \top_I.branch[12].block[8].um_I.iw[12] ,
    \top_I.branch[12].block[8].um_I.iw[11] ,
    \top_I.branch[12].block[8].um_I.iw[10] ,
    \top_I.branch[12].block[8].um_I.iw[9] ,
    \top_I.branch[12].block[8].um_I.iw[8] ,
    \top_I.branch[12].block[8].um_I.iw[7] ,
    \top_I.branch[12].block[8].um_I.iw[6] ,
    \top_I.branch[12].block[8].um_I.iw[5] ,
    \top_I.branch[12].block[8].um_I.iw[4] ,
    \top_I.branch[12].block[8].um_I.iw[3] ,
    \top_I.branch[12].block[8].um_I.iw[2] ,
    \top_I.branch[12].block[8].um_I.iw[1] ,
    \top_I.branch[12].block[8].um_I.clk ,
    \top_I.branch[12].block[7].um_I.iw[17] ,
    \top_I.branch[12].block[7].um_I.iw[16] ,
    \top_I.branch[12].block[7].um_I.iw[15] ,
    \top_I.branch[12].block[7].um_I.iw[14] ,
    \top_I.branch[12].block[7].um_I.iw[13] ,
    \top_I.branch[12].block[7].um_I.iw[12] ,
    \top_I.branch[12].block[7].um_I.iw[11] ,
    \top_I.branch[12].block[7].um_I.iw[10] ,
    \top_I.branch[12].block[7].um_I.iw[9] ,
    \top_I.branch[12].block[7].um_I.iw[8] ,
    \top_I.branch[12].block[7].um_I.iw[7] ,
    \top_I.branch[12].block[7].um_I.iw[6] ,
    \top_I.branch[12].block[7].um_I.iw[5] ,
    \top_I.branch[12].block[7].um_I.iw[4] ,
    \top_I.branch[12].block[7].um_I.iw[3] ,
    \top_I.branch[12].block[7].um_I.iw[2] ,
    \top_I.branch[12].block[7].um_I.iw[1] ,
    \top_I.branch[12].block[7].um_I.clk ,
    \top_I.branch[12].block[6].um_I.iw[17] ,
    \top_I.branch[12].block[6].um_I.iw[16] ,
    \top_I.branch[12].block[6].um_I.iw[15] ,
    \top_I.branch[12].block[6].um_I.iw[14] ,
    \top_I.branch[12].block[6].um_I.iw[13] ,
    \top_I.branch[12].block[6].um_I.iw[12] ,
    \top_I.branch[12].block[6].um_I.iw[11] ,
    \top_I.branch[12].block[6].um_I.iw[10] ,
    \top_I.branch[12].block[6].um_I.iw[9] ,
    \top_I.branch[12].block[6].um_I.iw[8] ,
    \top_I.branch[12].block[6].um_I.iw[7] ,
    \top_I.branch[12].block[6].um_I.iw[6] ,
    \top_I.branch[12].block[6].um_I.iw[5] ,
    \top_I.branch[12].block[6].um_I.iw[4] ,
    \top_I.branch[12].block[6].um_I.iw[3] ,
    \top_I.branch[12].block[6].um_I.iw[2] ,
    \top_I.branch[12].block[6].um_I.iw[1] ,
    \top_I.branch[12].block[6].um_I.clk ,
    \top_I.branch[12].block[5].um_I.iw[17] ,
    \top_I.branch[12].block[5].um_I.iw[16] ,
    \top_I.branch[12].block[5].um_I.iw[15] ,
    \top_I.branch[12].block[5].um_I.iw[14] ,
    \top_I.branch[12].block[5].um_I.iw[13] ,
    \top_I.branch[12].block[5].um_I.iw[12] ,
    \top_I.branch[12].block[5].um_I.iw[11] ,
    \top_I.branch[12].block[5].um_I.iw[10] ,
    \top_I.branch[12].block[5].um_I.iw[9] ,
    \top_I.branch[12].block[5].um_I.iw[8] ,
    \top_I.branch[12].block[5].um_I.iw[7] ,
    \top_I.branch[12].block[5].um_I.iw[6] ,
    \top_I.branch[12].block[5].um_I.iw[5] ,
    \top_I.branch[12].block[5].um_I.iw[4] ,
    \top_I.branch[12].block[5].um_I.iw[3] ,
    \top_I.branch[12].block[5].um_I.iw[2] ,
    \top_I.branch[12].block[5].um_I.iw[1] ,
    \top_I.branch[12].block[5].um_I.clk ,
    \top_I.branch[12].block[4].um_I.iw[17] ,
    \top_I.branch[12].block[4].um_I.iw[16] ,
    \top_I.branch[12].block[4].um_I.iw[15] ,
    \top_I.branch[12].block[4].um_I.iw[14] ,
    \top_I.branch[12].block[4].um_I.iw[13] ,
    \top_I.branch[12].block[4].um_I.iw[12] ,
    \top_I.branch[12].block[4].um_I.iw[11] ,
    \top_I.branch[12].block[4].um_I.iw[10] ,
    \top_I.branch[12].block[4].um_I.iw[9] ,
    \top_I.branch[12].block[4].um_I.iw[8] ,
    \top_I.branch[12].block[4].um_I.iw[7] ,
    \top_I.branch[12].block[4].um_I.iw[6] ,
    \top_I.branch[12].block[4].um_I.iw[5] ,
    \top_I.branch[12].block[4].um_I.iw[4] ,
    \top_I.branch[12].block[4].um_I.iw[3] ,
    \top_I.branch[12].block[4].um_I.iw[2] ,
    \top_I.branch[12].block[4].um_I.iw[1] ,
    \top_I.branch[12].block[4].um_I.clk ,
    \top_I.branch[12].block[3].um_I.iw[17] ,
    \top_I.branch[12].block[3].um_I.iw[16] ,
    \top_I.branch[12].block[3].um_I.iw[15] ,
    \top_I.branch[12].block[3].um_I.iw[14] ,
    \top_I.branch[12].block[3].um_I.iw[13] ,
    \top_I.branch[12].block[3].um_I.iw[12] ,
    \top_I.branch[12].block[3].um_I.iw[11] ,
    \top_I.branch[12].block[3].um_I.iw[10] ,
    \top_I.branch[12].block[3].um_I.iw[9] ,
    \top_I.branch[12].block[3].um_I.iw[8] ,
    \top_I.branch[12].block[3].um_I.iw[7] ,
    \top_I.branch[12].block[3].um_I.iw[6] ,
    \top_I.branch[12].block[3].um_I.iw[5] ,
    \top_I.branch[12].block[3].um_I.iw[4] ,
    \top_I.branch[12].block[3].um_I.iw[3] ,
    \top_I.branch[12].block[3].um_I.iw[2] ,
    \top_I.branch[12].block[3].um_I.iw[1] ,
    \top_I.branch[12].block[3].um_I.clk ,
    \top_I.branch[12].block[2].um_I.iw[17] ,
    \top_I.branch[12].block[2].um_I.iw[16] ,
    \top_I.branch[12].block[2].um_I.iw[15] ,
    \top_I.branch[12].block[2].um_I.iw[14] ,
    \top_I.branch[12].block[2].um_I.iw[13] ,
    \top_I.branch[12].block[2].um_I.iw[12] ,
    \top_I.branch[12].block[2].um_I.iw[11] ,
    \top_I.branch[12].block[2].um_I.iw[10] ,
    \top_I.branch[12].block[2].um_I.iw[9] ,
    \top_I.branch[12].block[2].um_I.iw[8] ,
    \top_I.branch[12].block[2].um_I.iw[7] ,
    \top_I.branch[12].block[2].um_I.iw[6] ,
    \top_I.branch[12].block[2].um_I.iw[5] ,
    \top_I.branch[12].block[2].um_I.iw[4] ,
    \top_I.branch[12].block[2].um_I.iw[3] ,
    \top_I.branch[12].block[2].um_I.iw[2] ,
    \top_I.branch[12].block[2].um_I.iw[1] ,
    \top_I.branch[12].block[2].um_I.clk ,
    \top_I.branch[12].block[1].um_I.iw[17] ,
    \top_I.branch[12].block[1].um_I.iw[16] ,
    \top_I.branch[12].block[1].um_I.iw[15] ,
    \top_I.branch[12].block[1].um_I.iw[14] ,
    \top_I.branch[12].block[1].um_I.iw[13] ,
    \top_I.branch[12].block[1].um_I.iw[12] ,
    \top_I.branch[12].block[1].um_I.iw[11] ,
    \top_I.branch[12].block[1].um_I.iw[10] ,
    \top_I.branch[12].block[1].um_I.iw[9] ,
    \top_I.branch[12].block[1].um_I.iw[8] ,
    \top_I.branch[12].block[1].um_I.iw[7] ,
    \top_I.branch[12].block[1].um_I.iw[6] ,
    \top_I.branch[12].block[1].um_I.iw[5] ,
    \top_I.branch[12].block[1].um_I.iw[4] ,
    \top_I.branch[12].block[1].um_I.iw[3] ,
    \top_I.branch[12].block[1].um_I.iw[2] ,
    \top_I.branch[12].block[1].um_I.iw[1] ,
    \top_I.branch[12].block[1].um_I.clk ,
    \top_I.branch[12].block[0].um_I.iw[17] ,
    \top_I.branch[12].block[0].um_I.iw[16] ,
    \top_I.branch[12].block[0].um_I.iw[15] ,
    \top_I.branch[12].block[0].um_I.iw[14] ,
    \top_I.branch[12].block[0].um_I.iw[13] ,
    \top_I.branch[12].block[0].um_I.iw[12] ,
    \top_I.branch[12].block[0].um_I.iw[11] ,
    \top_I.branch[12].block[0].um_I.iw[10] ,
    \top_I.branch[12].block[0].um_I.iw[9] ,
    \top_I.branch[12].block[0].um_I.iw[8] ,
    \top_I.branch[12].block[0].um_I.iw[7] ,
    \top_I.branch[12].block[0].um_I.iw[6] ,
    \top_I.branch[12].block[0].um_I.iw[5] ,
    \top_I.branch[12].block[0].um_I.iw[4] ,
    \top_I.branch[12].block[0].um_I.iw[3] ,
    \top_I.branch[12].block[0].um_I.iw[2] ,
    \top_I.branch[12].block[0].um_I.iw[1] ,
    \top_I.branch[12].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[12].block[15].um_I.pg_vdd ,
    \top_I.branch[12].block[14].um_I.pg_vdd ,
    \top_I.branch[12].block[13].um_I.pg_vdd ,
    \top_I.branch[12].block[12].um_I.pg_vdd ,
    \top_I.branch[12].block[11].um_I.pg_vdd ,
    \top_I.branch[12].block[10].um_I.pg_vdd ,
    \top_I.branch[12].block[9].um_I.pg_vdd ,
    \top_I.branch[12].block[8].um_I.pg_vdd ,
    \top_I.branch[12].block[7].um_I.pg_vdd ,
    \top_I.branch[12].block[6].um_I.pg_vdd ,
    \top_I.branch[12].block[5].um_I.pg_vdd ,
    \top_I.branch[12].block[4].um_I.pg_vdd ,
    \top_I.branch[12].block[3].um_I.pg_vdd ,
    \top_I.branch[12].block[2].um_I.pg_vdd ,
    \top_I.branch[12].block[1].um_I.pg_vdd ,
    \top_I.branch[12].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[13].mux_I  (.k_one(\top_I.branch[13].l_addr[1] ),
    .k_zero(\top_I.branch[13].l_addr[0] ),
    .addr({\top_I.branch[13].l_addr[0] ,
    \top_I.branch[13].l_addr[1] ,
    \top_I.branch[13].l_addr[1] ,
    \top_I.branch[13].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[13].block[15].um_I.ena ,
    \top_I.branch[13].block[14].um_I.ena ,
    \top_I.branch[13].block[13].um_I.ena ,
    \top_I.branch[13].block[12].um_I.ena ,
    \top_I.branch[13].block[11].um_I.ena ,
    \top_I.branch[13].block[10].um_I.ena ,
    \top_I.branch[13].block[9].um_I.ena ,
    \top_I.branch[13].block[8].um_I.ena ,
    \top_I.branch[13].block[7].um_I.ena ,
    \top_I.branch[13].block[6].um_I.ena ,
    \top_I.branch[13].block[5].um_I.ena ,
    \top_I.branch[13].block[4].um_I.ena ,
    \top_I.branch[13].block[3].um_I.ena ,
    \top_I.branch[13].block[2].um_I.ena ,
    \top_I.branch[13].block[1].um_I.ena ,
    \top_I.branch[13].block[0].um_I.ena }),
    .um_iw({\top_I.branch[13].block[15].um_I.iw[17] ,
    \top_I.branch[13].block[15].um_I.iw[16] ,
    \top_I.branch[13].block[15].um_I.iw[15] ,
    \top_I.branch[13].block[15].um_I.iw[14] ,
    \top_I.branch[13].block[15].um_I.iw[13] ,
    \top_I.branch[13].block[15].um_I.iw[12] ,
    \top_I.branch[13].block[15].um_I.iw[11] ,
    \top_I.branch[13].block[15].um_I.iw[10] ,
    \top_I.branch[13].block[15].um_I.iw[9] ,
    \top_I.branch[13].block[15].um_I.iw[8] ,
    \top_I.branch[13].block[15].um_I.iw[7] ,
    \top_I.branch[13].block[15].um_I.iw[6] ,
    \top_I.branch[13].block[15].um_I.iw[5] ,
    \top_I.branch[13].block[15].um_I.iw[4] ,
    \top_I.branch[13].block[15].um_I.iw[3] ,
    \top_I.branch[13].block[15].um_I.iw[2] ,
    \top_I.branch[13].block[15].um_I.iw[1] ,
    \top_I.branch[13].block[15].um_I.clk ,
    \top_I.branch[13].block[14].um_I.iw[17] ,
    \top_I.branch[13].block[14].um_I.iw[16] ,
    \top_I.branch[13].block[14].um_I.iw[15] ,
    \top_I.branch[13].block[14].um_I.iw[14] ,
    \top_I.branch[13].block[14].um_I.iw[13] ,
    \top_I.branch[13].block[14].um_I.iw[12] ,
    \top_I.branch[13].block[14].um_I.iw[11] ,
    \top_I.branch[13].block[14].um_I.iw[10] ,
    \top_I.branch[13].block[14].um_I.iw[9] ,
    \top_I.branch[13].block[14].um_I.iw[8] ,
    \top_I.branch[13].block[14].um_I.iw[7] ,
    \top_I.branch[13].block[14].um_I.iw[6] ,
    \top_I.branch[13].block[14].um_I.iw[5] ,
    \top_I.branch[13].block[14].um_I.iw[4] ,
    \top_I.branch[13].block[14].um_I.iw[3] ,
    \top_I.branch[13].block[14].um_I.iw[2] ,
    \top_I.branch[13].block[14].um_I.iw[1] ,
    \top_I.branch[13].block[14].um_I.clk ,
    \top_I.branch[13].block[13].um_I.iw[17] ,
    \top_I.branch[13].block[13].um_I.iw[16] ,
    \top_I.branch[13].block[13].um_I.iw[15] ,
    \top_I.branch[13].block[13].um_I.iw[14] ,
    \top_I.branch[13].block[13].um_I.iw[13] ,
    \top_I.branch[13].block[13].um_I.iw[12] ,
    \top_I.branch[13].block[13].um_I.iw[11] ,
    \top_I.branch[13].block[13].um_I.iw[10] ,
    \top_I.branch[13].block[13].um_I.iw[9] ,
    \top_I.branch[13].block[13].um_I.iw[8] ,
    \top_I.branch[13].block[13].um_I.iw[7] ,
    \top_I.branch[13].block[13].um_I.iw[6] ,
    \top_I.branch[13].block[13].um_I.iw[5] ,
    \top_I.branch[13].block[13].um_I.iw[4] ,
    \top_I.branch[13].block[13].um_I.iw[3] ,
    \top_I.branch[13].block[13].um_I.iw[2] ,
    \top_I.branch[13].block[13].um_I.iw[1] ,
    \top_I.branch[13].block[13].um_I.clk ,
    \top_I.branch[13].block[12].um_I.iw[17] ,
    \top_I.branch[13].block[12].um_I.iw[16] ,
    \top_I.branch[13].block[12].um_I.iw[15] ,
    \top_I.branch[13].block[12].um_I.iw[14] ,
    \top_I.branch[13].block[12].um_I.iw[13] ,
    \top_I.branch[13].block[12].um_I.iw[12] ,
    \top_I.branch[13].block[12].um_I.iw[11] ,
    \top_I.branch[13].block[12].um_I.iw[10] ,
    \top_I.branch[13].block[12].um_I.iw[9] ,
    \top_I.branch[13].block[12].um_I.iw[8] ,
    \top_I.branch[13].block[12].um_I.iw[7] ,
    \top_I.branch[13].block[12].um_I.iw[6] ,
    \top_I.branch[13].block[12].um_I.iw[5] ,
    \top_I.branch[13].block[12].um_I.iw[4] ,
    \top_I.branch[13].block[12].um_I.iw[3] ,
    \top_I.branch[13].block[12].um_I.iw[2] ,
    \top_I.branch[13].block[12].um_I.iw[1] ,
    \top_I.branch[13].block[12].um_I.clk ,
    \top_I.branch[13].block[11].um_I.iw[17] ,
    \top_I.branch[13].block[11].um_I.iw[16] ,
    \top_I.branch[13].block[11].um_I.iw[15] ,
    \top_I.branch[13].block[11].um_I.iw[14] ,
    \top_I.branch[13].block[11].um_I.iw[13] ,
    \top_I.branch[13].block[11].um_I.iw[12] ,
    \top_I.branch[13].block[11].um_I.iw[11] ,
    \top_I.branch[13].block[11].um_I.iw[10] ,
    \top_I.branch[13].block[11].um_I.iw[9] ,
    \top_I.branch[13].block[11].um_I.iw[8] ,
    \top_I.branch[13].block[11].um_I.iw[7] ,
    \top_I.branch[13].block[11].um_I.iw[6] ,
    \top_I.branch[13].block[11].um_I.iw[5] ,
    \top_I.branch[13].block[11].um_I.iw[4] ,
    \top_I.branch[13].block[11].um_I.iw[3] ,
    \top_I.branch[13].block[11].um_I.iw[2] ,
    \top_I.branch[13].block[11].um_I.iw[1] ,
    \top_I.branch[13].block[11].um_I.clk ,
    \top_I.branch[13].block[10].um_I.iw[17] ,
    \top_I.branch[13].block[10].um_I.iw[16] ,
    \top_I.branch[13].block[10].um_I.iw[15] ,
    \top_I.branch[13].block[10].um_I.iw[14] ,
    \top_I.branch[13].block[10].um_I.iw[13] ,
    \top_I.branch[13].block[10].um_I.iw[12] ,
    \top_I.branch[13].block[10].um_I.iw[11] ,
    \top_I.branch[13].block[10].um_I.iw[10] ,
    \top_I.branch[13].block[10].um_I.iw[9] ,
    \top_I.branch[13].block[10].um_I.iw[8] ,
    \top_I.branch[13].block[10].um_I.iw[7] ,
    \top_I.branch[13].block[10].um_I.iw[6] ,
    \top_I.branch[13].block[10].um_I.iw[5] ,
    \top_I.branch[13].block[10].um_I.iw[4] ,
    \top_I.branch[13].block[10].um_I.iw[3] ,
    \top_I.branch[13].block[10].um_I.iw[2] ,
    \top_I.branch[13].block[10].um_I.iw[1] ,
    \top_I.branch[13].block[10].um_I.clk ,
    \top_I.branch[13].block[9].um_I.iw[17] ,
    \top_I.branch[13].block[9].um_I.iw[16] ,
    \top_I.branch[13].block[9].um_I.iw[15] ,
    \top_I.branch[13].block[9].um_I.iw[14] ,
    \top_I.branch[13].block[9].um_I.iw[13] ,
    \top_I.branch[13].block[9].um_I.iw[12] ,
    \top_I.branch[13].block[9].um_I.iw[11] ,
    \top_I.branch[13].block[9].um_I.iw[10] ,
    \top_I.branch[13].block[9].um_I.iw[9] ,
    \top_I.branch[13].block[9].um_I.iw[8] ,
    \top_I.branch[13].block[9].um_I.iw[7] ,
    \top_I.branch[13].block[9].um_I.iw[6] ,
    \top_I.branch[13].block[9].um_I.iw[5] ,
    \top_I.branch[13].block[9].um_I.iw[4] ,
    \top_I.branch[13].block[9].um_I.iw[3] ,
    \top_I.branch[13].block[9].um_I.iw[2] ,
    \top_I.branch[13].block[9].um_I.iw[1] ,
    \top_I.branch[13].block[9].um_I.clk ,
    \top_I.branch[13].block[8].um_I.iw[17] ,
    \top_I.branch[13].block[8].um_I.iw[16] ,
    \top_I.branch[13].block[8].um_I.iw[15] ,
    \top_I.branch[13].block[8].um_I.iw[14] ,
    \top_I.branch[13].block[8].um_I.iw[13] ,
    \top_I.branch[13].block[8].um_I.iw[12] ,
    \top_I.branch[13].block[8].um_I.iw[11] ,
    \top_I.branch[13].block[8].um_I.iw[10] ,
    \top_I.branch[13].block[8].um_I.iw[9] ,
    \top_I.branch[13].block[8].um_I.iw[8] ,
    \top_I.branch[13].block[8].um_I.iw[7] ,
    \top_I.branch[13].block[8].um_I.iw[6] ,
    \top_I.branch[13].block[8].um_I.iw[5] ,
    \top_I.branch[13].block[8].um_I.iw[4] ,
    \top_I.branch[13].block[8].um_I.iw[3] ,
    \top_I.branch[13].block[8].um_I.iw[2] ,
    \top_I.branch[13].block[8].um_I.iw[1] ,
    \top_I.branch[13].block[8].um_I.clk ,
    \top_I.branch[13].block[7].um_I.iw[17] ,
    \top_I.branch[13].block[7].um_I.iw[16] ,
    \top_I.branch[13].block[7].um_I.iw[15] ,
    \top_I.branch[13].block[7].um_I.iw[14] ,
    \top_I.branch[13].block[7].um_I.iw[13] ,
    \top_I.branch[13].block[7].um_I.iw[12] ,
    \top_I.branch[13].block[7].um_I.iw[11] ,
    \top_I.branch[13].block[7].um_I.iw[10] ,
    \top_I.branch[13].block[7].um_I.iw[9] ,
    \top_I.branch[13].block[7].um_I.iw[8] ,
    \top_I.branch[13].block[7].um_I.iw[7] ,
    \top_I.branch[13].block[7].um_I.iw[6] ,
    \top_I.branch[13].block[7].um_I.iw[5] ,
    \top_I.branch[13].block[7].um_I.iw[4] ,
    \top_I.branch[13].block[7].um_I.iw[3] ,
    \top_I.branch[13].block[7].um_I.iw[2] ,
    \top_I.branch[13].block[7].um_I.iw[1] ,
    \top_I.branch[13].block[7].um_I.clk ,
    \top_I.branch[13].block[6].um_I.iw[17] ,
    \top_I.branch[13].block[6].um_I.iw[16] ,
    \top_I.branch[13].block[6].um_I.iw[15] ,
    \top_I.branch[13].block[6].um_I.iw[14] ,
    \top_I.branch[13].block[6].um_I.iw[13] ,
    \top_I.branch[13].block[6].um_I.iw[12] ,
    \top_I.branch[13].block[6].um_I.iw[11] ,
    \top_I.branch[13].block[6].um_I.iw[10] ,
    \top_I.branch[13].block[6].um_I.iw[9] ,
    \top_I.branch[13].block[6].um_I.iw[8] ,
    \top_I.branch[13].block[6].um_I.iw[7] ,
    \top_I.branch[13].block[6].um_I.iw[6] ,
    \top_I.branch[13].block[6].um_I.iw[5] ,
    \top_I.branch[13].block[6].um_I.iw[4] ,
    \top_I.branch[13].block[6].um_I.iw[3] ,
    \top_I.branch[13].block[6].um_I.iw[2] ,
    \top_I.branch[13].block[6].um_I.iw[1] ,
    \top_I.branch[13].block[6].um_I.clk ,
    \top_I.branch[13].block[5].um_I.iw[17] ,
    \top_I.branch[13].block[5].um_I.iw[16] ,
    \top_I.branch[13].block[5].um_I.iw[15] ,
    \top_I.branch[13].block[5].um_I.iw[14] ,
    \top_I.branch[13].block[5].um_I.iw[13] ,
    \top_I.branch[13].block[5].um_I.iw[12] ,
    \top_I.branch[13].block[5].um_I.iw[11] ,
    \top_I.branch[13].block[5].um_I.iw[10] ,
    \top_I.branch[13].block[5].um_I.iw[9] ,
    \top_I.branch[13].block[5].um_I.iw[8] ,
    \top_I.branch[13].block[5].um_I.iw[7] ,
    \top_I.branch[13].block[5].um_I.iw[6] ,
    \top_I.branch[13].block[5].um_I.iw[5] ,
    \top_I.branch[13].block[5].um_I.iw[4] ,
    \top_I.branch[13].block[5].um_I.iw[3] ,
    \top_I.branch[13].block[5].um_I.iw[2] ,
    \top_I.branch[13].block[5].um_I.iw[1] ,
    \top_I.branch[13].block[5].um_I.clk ,
    \top_I.branch[13].block[4].um_I.iw[17] ,
    \top_I.branch[13].block[4].um_I.iw[16] ,
    \top_I.branch[13].block[4].um_I.iw[15] ,
    \top_I.branch[13].block[4].um_I.iw[14] ,
    \top_I.branch[13].block[4].um_I.iw[13] ,
    \top_I.branch[13].block[4].um_I.iw[12] ,
    \top_I.branch[13].block[4].um_I.iw[11] ,
    \top_I.branch[13].block[4].um_I.iw[10] ,
    \top_I.branch[13].block[4].um_I.iw[9] ,
    \top_I.branch[13].block[4].um_I.iw[8] ,
    \top_I.branch[13].block[4].um_I.iw[7] ,
    \top_I.branch[13].block[4].um_I.iw[6] ,
    \top_I.branch[13].block[4].um_I.iw[5] ,
    \top_I.branch[13].block[4].um_I.iw[4] ,
    \top_I.branch[13].block[4].um_I.iw[3] ,
    \top_I.branch[13].block[4].um_I.iw[2] ,
    \top_I.branch[13].block[4].um_I.iw[1] ,
    \top_I.branch[13].block[4].um_I.clk ,
    \top_I.branch[13].block[3].um_I.iw[17] ,
    \top_I.branch[13].block[3].um_I.iw[16] ,
    \top_I.branch[13].block[3].um_I.iw[15] ,
    \top_I.branch[13].block[3].um_I.iw[14] ,
    \top_I.branch[13].block[3].um_I.iw[13] ,
    \top_I.branch[13].block[3].um_I.iw[12] ,
    \top_I.branch[13].block[3].um_I.iw[11] ,
    \top_I.branch[13].block[3].um_I.iw[10] ,
    \top_I.branch[13].block[3].um_I.iw[9] ,
    \top_I.branch[13].block[3].um_I.iw[8] ,
    \top_I.branch[13].block[3].um_I.iw[7] ,
    \top_I.branch[13].block[3].um_I.iw[6] ,
    \top_I.branch[13].block[3].um_I.iw[5] ,
    \top_I.branch[13].block[3].um_I.iw[4] ,
    \top_I.branch[13].block[3].um_I.iw[3] ,
    \top_I.branch[13].block[3].um_I.iw[2] ,
    \top_I.branch[13].block[3].um_I.iw[1] ,
    \top_I.branch[13].block[3].um_I.clk ,
    \top_I.branch[13].block[2].um_I.iw[17] ,
    \top_I.branch[13].block[2].um_I.iw[16] ,
    \top_I.branch[13].block[2].um_I.iw[15] ,
    \top_I.branch[13].block[2].um_I.iw[14] ,
    \top_I.branch[13].block[2].um_I.iw[13] ,
    \top_I.branch[13].block[2].um_I.iw[12] ,
    \top_I.branch[13].block[2].um_I.iw[11] ,
    \top_I.branch[13].block[2].um_I.iw[10] ,
    \top_I.branch[13].block[2].um_I.iw[9] ,
    \top_I.branch[13].block[2].um_I.iw[8] ,
    \top_I.branch[13].block[2].um_I.iw[7] ,
    \top_I.branch[13].block[2].um_I.iw[6] ,
    \top_I.branch[13].block[2].um_I.iw[5] ,
    \top_I.branch[13].block[2].um_I.iw[4] ,
    \top_I.branch[13].block[2].um_I.iw[3] ,
    \top_I.branch[13].block[2].um_I.iw[2] ,
    \top_I.branch[13].block[2].um_I.iw[1] ,
    \top_I.branch[13].block[2].um_I.clk ,
    \top_I.branch[13].block[1].um_I.iw[17] ,
    \top_I.branch[13].block[1].um_I.iw[16] ,
    \top_I.branch[13].block[1].um_I.iw[15] ,
    \top_I.branch[13].block[1].um_I.iw[14] ,
    \top_I.branch[13].block[1].um_I.iw[13] ,
    \top_I.branch[13].block[1].um_I.iw[12] ,
    \top_I.branch[13].block[1].um_I.iw[11] ,
    \top_I.branch[13].block[1].um_I.iw[10] ,
    \top_I.branch[13].block[1].um_I.iw[9] ,
    \top_I.branch[13].block[1].um_I.iw[8] ,
    \top_I.branch[13].block[1].um_I.iw[7] ,
    \top_I.branch[13].block[1].um_I.iw[6] ,
    \top_I.branch[13].block[1].um_I.iw[5] ,
    \top_I.branch[13].block[1].um_I.iw[4] ,
    \top_I.branch[13].block[1].um_I.iw[3] ,
    \top_I.branch[13].block[1].um_I.iw[2] ,
    \top_I.branch[13].block[1].um_I.iw[1] ,
    \top_I.branch[13].block[1].um_I.clk ,
    \top_I.branch[13].block[0].um_I.iw[17] ,
    \top_I.branch[13].block[0].um_I.iw[16] ,
    \top_I.branch[13].block[0].um_I.iw[15] ,
    \top_I.branch[13].block[0].um_I.iw[14] ,
    \top_I.branch[13].block[0].um_I.iw[13] ,
    \top_I.branch[13].block[0].um_I.iw[12] ,
    \top_I.branch[13].block[0].um_I.iw[11] ,
    \top_I.branch[13].block[0].um_I.iw[10] ,
    \top_I.branch[13].block[0].um_I.iw[9] ,
    \top_I.branch[13].block[0].um_I.iw[8] ,
    \top_I.branch[13].block[0].um_I.iw[7] ,
    \top_I.branch[13].block[0].um_I.iw[6] ,
    \top_I.branch[13].block[0].um_I.iw[5] ,
    \top_I.branch[13].block[0].um_I.iw[4] ,
    \top_I.branch[13].block[0].um_I.iw[3] ,
    \top_I.branch[13].block[0].um_I.iw[2] ,
    \top_I.branch[13].block[0].um_I.iw[1] ,
    \top_I.branch[13].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[13].block[15].um_I.pg_vdd ,
    \top_I.branch[13].block[14].um_I.pg_vdd ,
    \top_I.branch[13].block[13].um_I.pg_vdd ,
    \top_I.branch[13].block[12].um_I.pg_vdd ,
    \top_I.branch[13].block[11].um_I.pg_vdd ,
    \top_I.branch[13].block[10].um_I.pg_vdd ,
    \top_I.branch[13].block[9].um_I.pg_vdd ,
    \top_I.branch[13].block[8].um_I.pg_vdd ,
    \top_I.branch[13].block[7].um_I.pg_vdd ,
    \top_I.branch[13].block[6].um_I.pg_vdd ,
    \top_I.branch[13].block[5].um_I.pg_vdd ,
    \top_I.branch[13].block[4].um_I.pg_vdd ,
    \top_I.branch[13].block[3].um_I.pg_vdd ,
    \top_I.branch[13].block[2].um_I.pg_vdd ,
    \top_I.branch[13].block[1].um_I.pg_vdd ,
    \top_I.branch[13].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[14].mux_I  (.k_one(\top_I.branch[14].l_addr[0] ),
    .k_zero(\top_I.branch[14].l_addr[3] ),
    .addr({\top_I.branch[14].l_addr[3] ,
    \top_I.branch[14].l_addr[0] ,
    \top_I.branch[14].l_addr[0] ,
    \top_I.branch[14].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[14].block[15].um_I.ena ,
    \top_I.branch[14].block[14].um_I.ena ,
    \top_I.branch[14].block[13].um_I.ena ,
    \top_I.branch[14].block[12].um_I.ena ,
    \top_I.branch[14].block[11].um_I.ena ,
    \top_I.branch[14].block[10].um_I.ena ,
    \top_I.branch[14].block[9].um_I.ena ,
    \top_I.branch[14].block[8].um_I.ena ,
    \top_I.branch[14].block[7].um_I.ena ,
    \top_I.branch[14].block[6].um_I.ena ,
    \top_I.branch[14].block[5].um_I.ena ,
    \top_I.branch[14].block[4].um_I.ena ,
    \top_I.branch[14].block[3].um_I.ena ,
    \top_I.branch[14].block[2].um_I.ena ,
    \top_I.branch[14].block[1].um_I.ena ,
    \top_I.branch[14].block[0].um_I.ena }),
    .um_iw({\top_I.branch[14].block[15].um_I.iw[17] ,
    \top_I.branch[14].block[15].um_I.iw[16] ,
    \top_I.branch[14].block[15].um_I.iw[15] ,
    \top_I.branch[14].block[15].um_I.iw[14] ,
    \top_I.branch[14].block[15].um_I.iw[13] ,
    \top_I.branch[14].block[15].um_I.iw[12] ,
    \top_I.branch[14].block[15].um_I.iw[11] ,
    \top_I.branch[14].block[15].um_I.iw[10] ,
    \top_I.branch[14].block[15].um_I.iw[9] ,
    \top_I.branch[14].block[15].um_I.iw[8] ,
    \top_I.branch[14].block[15].um_I.iw[7] ,
    \top_I.branch[14].block[15].um_I.iw[6] ,
    \top_I.branch[14].block[15].um_I.iw[5] ,
    \top_I.branch[14].block[15].um_I.iw[4] ,
    \top_I.branch[14].block[15].um_I.iw[3] ,
    \top_I.branch[14].block[15].um_I.iw[2] ,
    \top_I.branch[14].block[15].um_I.iw[1] ,
    \top_I.branch[14].block[15].um_I.clk ,
    \top_I.branch[14].block[14].um_I.iw[17] ,
    \top_I.branch[14].block[14].um_I.iw[16] ,
    \top_I.branch[14].block[14].um_I.iw[15] ,
    \top_I.branch[14].block[14].um_I.iw[14] ,
    \top_I.branch[14].block[14].um_I.iw[13] ,
    \top_I.branch[14].block[14].um_I.iw[12] ,
    \top_I.branch[14].block[14].um_I.iw[11] ,
    \top_I.branch[14].block[14].um_I.iw[10] ,
    \top_I.branch[14].block[14].um_I.iw[9] ,
    \top_I.branch[14].block[14].um_I.iw[8] ,
    \top_I.branch[14].block[14].um_I.iw[7] ,
    \top_I.branch[14].block[14].um_I.iw[6] ,
    \top_I.branch[14].block[14].um_I.iw[5] ,
    \top_I.branch[14].block[14].um_I.iw[4] ,
    \top_I.branch[14].block[14].um_I.iw[3] ,
    \top_I.branch[14].block[14].um_I.iw[2] ,
    \top_I.branch[14].block[14].um_I.iw[1] ,
    \top_I.branch[14].block[14].um_I.clk ,
    \top_I.branch[14].block[13].um_I.iw[17] ,
    \top_I.branch[14].block[13].um_I.iw[16] ,
    \top_I.branch[14].block[13].um_I.iw[15] ,
    \top_I.branch[14].block[13].um_I.iw[14] ,
    \top_I.branch[14].block[13].um_I.iw[13] ,
    \top_I.branch[14].block[13].um_I.iw[12] ,
    \top_I.branch[14].block[13].um_I.iw[11] ,
    \top_I.branch[14].block[13].um_I.iw[10] ,
    \top_I.branch[14].block[13].um_I.iw[9] ,
    \top_I.branch[14].block[13].um_I.iw[8] ,
    \top_I.branch[14].block[13].um_I.iw[7] ,
    \top_I.branch[14].block[13].um_I.iw[6] ,
    \top_I.branch[14].block[13].um_I.iw[5] ,
    \top_I.branch[14].block[13].um_I.iw[4] ,
    \top_I.branch[14].block[13].um_I.iw[3] ,
    \top_I.branch[14].block[13].um_I.iw[2] ,
    \top_I.branch[14].block[13].um_I.iw[1] ,
    \top_I.branch[14].block[13].um_I.clk ,
    \top_I.branch[14].block[12].um_I.iw[17] ,
    \top_I.branch[14].block[12].um_I.iw[16] ,
    \top_I.branch[14].block[12].um_I.iw[15] ,
    \top_I.branch[14].block[12].um_I.iw[14] ,
    \top_I.branch[14].block[12].um_I.iw[13] ,
    \top_I.branch[14].block[12].um_I.iw[12] ,
    \top_I.branch[14].block[12].um_I.iw[11] ,
    \top_I.branch[14].block[12].um_I.iw[10] ,
    \top_I.branch[14].block[12].um_I.iw[9] ,
    \top_I.branch[14].block[12].um_I.iw[8] ,
    \top_I.branch[14].block[12].um_I.iw[7] ,
    \top_I.branch[14].block[12].um_I.iw[6] ,
    \top_I.branch[14].block[12].um_I.iw[5] ,
    \top_I.branch[14].block[12].um_I.iw[4] ,
    \top_I.branch[14].block[12].um_I.iw[3] ,
    \top_I.branch[14].block[12].um_I.iw[2] ,
    \top_I.branch[14].block[12].um_I.iw[1] ,
    \top_I.branch[14].block[12].um_I.clk ,
    \top_I.branch[14].block[11].um_I.iw[17] ,
    \top_I.branch[14].block[11].um_I.iw[16] ,
    \top_I.branch[14].block[11].um_I.iw[15] ,
    \top_I.branch[14].block[11].um_I.iw[14] ,
    \top_I.branch[14].block[11].um_I.iw[13] ,
    \top_I.branch[14].block[11].um_I.iw[12] ,
    \top_I.branch[14].block[11].um_I.iw[11] ,
    \top_I.branch[14].block[11].um_I.iw[10] ,
    \top_I.branch[14].block[11].um_I.iw[9] ,
    \top_I.branch[14].block[11].um_I.iw[8] ,
    \top_I.branch[14].block[11].um_I.iw[7] ,
    \top_I.branch[14].block[11].um_I.iw[6] ,
    \top_I.branch[14].block[11].um_I.iw[5] ,
    \top_I.branch[14].block[11].um_I.iw[4] ,
    \top_I.branch[14].block[11].um_I.iw[3] ,
    \top_I.branch[14].block[11].um_I.iw[2] ,
    \top_I.branch[14].block[11].um_I.iw[1] ,
    \top_I.branch[14].block[11].um_I.clk ,
    \top_I.branch[14].block[10].um_I.iw[17] ,
    \top_I.branch[14].block[10].um_I.iw[16] ,
    \top_I.branch[14].block[10].um_I.iw[15] ,
    \top_I.branch[14].block[10].um_I.iw[14] ,
    \top_I.branch[14].block[10].um_I.iw[13] ,
    \top_I.branch[14].block[10].um_I.iw[12] ,
    \top_I.branch[14].block[10].um_I.iw[11] ,
    \top_I.branch[14].block[10].um_I.iw[10] ,
    \top_I.branch[14].block[10].um_I.iw[9] ,
    \top_I.branch[14].block[10].um_I.iw[8] ,
    \top_I.branch[14].block[10].um_I.iw[7] ,
    \top_I.branch[14].block[10].um_I.iw[6] ,
    \top_I.branch[14].block[10].um_I.iw[5] ,
    \top_I.branch[14].block[10].um_I.iw[4] ,
    \top_I.branch[14].block[10].um_I.iw[3] ,
    \top_I.branch[14].block[10].um_I.iw[2] ,
    \top_I.branch[14].block[10].um_I.iw[1] ,
    \top_I.branch[14].block[10].um_I.clk ,
    \top_I.branch[14].block[9].um_I.iw[17] ,
    \top_I.branch[14].block[9].um_I.iw[16] ,
    \top_I.branch[14].block[9].um_I.iw[15] ,
    \top_I.branch[14].block[9].um_I.iw[14] ,
    \top_I.branch[14].block[9].um_I.iw[13] ,
    \top_I.branch[14].block[9].um_I.iw[12] ,
    \top_I.branch[14].block[9].um_I.iw[11] ,
    \top_I.branch[14].block[9].um_I.iw[10] ,
    \top_I.branch[14].block[9].um_I.iw[9] ,
    \top_I.branch[14].block[9].um_I.iw[8] ,
    \top_I.branch[14].block[9].um_I.iw[7] ,
    \top_I.branch[14].block[9].um_I.iw[6] ,
    \top_I.branch[14].block[9].um_I.iw[5] ,
    \top_I.branch[14].block[9].um_I.iw[4] ,
    \top_I.branch[14].block[9].um_I.iw[3] ,
    \top_I.branch[14].block[9].um_I.iw[2] ,
    \top_I.branch[14].block[9].um_I.iw[1] ,
    \top_I.branch[14].block[9].um_I.clk ,
    \top_I.branch[14].block[8].um_I.iw[17] ,
    \top_I.branch[14].block[8].um_I.iw[16] ,
    \top_I.branch[14].block[8].um_I.iw[15] ,
    \top_I.branch[14].block[8].um_I.iw[14] ,
    \top_I.branch[14].block[8].um_I.iw[13] ,
    \top_I.branch[14].block[8].um_I.iw[12] ,
    \top_I.branch[14].block[8].um_I.iw[11] ,
    \top_I.branch[14].block[8].um_I.iw[10] ,
    \top_I.branch[14].block[8].um_I.iw[9] ,
    \top_I.branch[14].block[8].um_I.iw[8] ,
    \top_I.branch[14].block[8].um_I.iw[7] ,
    \top_I.branch[14].block[8].um_I.iw[6] ,
    \top_I.branch[14].block[8].um_I.iw[5] ,
    \top_I.branch[14].block[8].um_I.iw[4] ,
    \top_I.branch[14].block[8].um_I.iw[3] ,
    \top_I.branch[14].block[8].um_I.iw[2] ,
    \top_I.branch[14].block[8].um_I.iw[1] ,
    \top_I.branch[14].block[8].um_I.clk ,
    \top_I.branch[14].block[7].um_I.iw[17] ,
    \top_I.branch[14].block[7].um_I.iw[16] ,
    \top_I.branch[14].block[7].um_I.iw[15] ,
    \top_I.branch[14].block[7].um_I.iw[14] ,
    \top_I.branch[14].block[7].um_I.iw[13] ,
    \top_I.branch[14].block[7].um_I.iw[12] ,
    \top_I.branch[14].block[7].um_I.iw[11] ,
    \top_I.branch[14].block[7].um_I.iw[10] ,
    \top_I.branch[14].block[7].um_I.iw[9] ,
    \top_I.branch[14].block[7].um_I.iw[8] ,
    \top_I.branch[14].block[7].um_I.iw[7] ,
    \top_I.branch[14].block[7].um_I.iw[6] ,
    \top_I.branch[14].block[7].um_I.iw[5] ,
    \top_I.branch[14].block[7].um_I.iw[4] ,
    \top_I.branch[14].block[7].um_I.iw[3] ,
    \top_I.branch[14].block[7].um_I.iw[2] ,
    \top_I.branch[14].block[7].um_I.iw[1] ,
    \top_I.branch[14].block[7].um_I.clk ,
    \top_I.branch[14].block[6].um_I.iw[17] ,
    \top_I.branch[14].block[6].um_I.iw[16] ,
    \top_I.branch[14].block[6].um_I.iw[15] ,
    \top_I.branch[14].block[6].um_I.iw[14] ,
    \top_I.branch[14].block[6].um_I.iw[13] ,
    \top_I.branch[14].block[6].um_I.iw[12] ,
    \top_I.branch[14].block[6].um_I.iw[11] ,
    \top_I.branch[14].block[6].um_I.iw[10] ,
    \top_I.branch[14].block[6].um_I.iw[9] ,
    \top_I.branch[14].block[6].um_I.iw[8] ,
    \top_I.branch[14].block[6].um_I.iw[7] ,
    \top_I.branch[14].block[6].um_I.iw[6] ,
    \top_I.branch[14].block[6].um_I.iw[5] ,
    \top_I.branch[14].block[6].um_I.iw[4] ,
    \top_I.branch[14].block[6].um_I.iw[3] ,
    \top_I.branch[14].block[6].um_I.iw[2] ,
    \top_I.branch[14].block[6].um_I.iw[1] ,
    \top_I.branch[14].block[6].um_I.clk ,
    \top_I.branch[14].block[5].um_I.iw[17] ,
    \top_I.branch[14].block[5].um_I.iw[16] ,
    \top_I.branch[14].block[5].um_I.iw[15] ,
    \top_I.branch[14].block[5].um_I.iw[14] ,
    \top_I.branch[14].block[5].um_I.iw[13] ,
    \top_I.branch[14].block[5].um_I.iw[12] ,
    \top_I.branch[14].block[5].um_I.iw[11] ,
    \top_I.branch[14].block[5].um_I.iw[10] ,
    \top_I.branch[14].block[5].um_I.iw[9] ,
    \top_I.branch[14].block[5].um_I.iw[8] ,
    \top_I.branch[14].block[5].um_I.iw[7] ,
    \top_I.branch[14].block[5].um_I.iw[6] ,
    \top_I.branch[14].block[5].um_I.iw[5] ,
    \top_I.branch[14].block[5].um_I.iw[4] ,
    \top_I.branch[14].block[5].um_I.iw[3] ,
    \top_I.branch[14].block[5].um_I.iw[2] ,
    \top_I.branch[14].block[5].um_I.iw[1] ,
    \top_I.branch[14].block[5].um_I.clk ,
    \top_I.branch[14].block[4].um_I.iw[17] ,
    \top_I.branch[14].block[4].um_I.iw[16] ,
    \top_I.branch[14].block[4].um_I.iw[15] ,
    \top_I.branch[14].block[4].um_I.iw[14] ,
    \top_I.branch[14].block[4].um_I.iw[13] ,
    \top_I.branch[14].block[4].um_I.iw[12] ,
    \top_I.branch[14].block[4].um_I.iw[11] ,
    \top_I.branch[14].block[4].um_I.iw[10] ,
    \top_I.branch[14].block[4].um_I.iw[9] ,
    \top_I.branch[14].block[4].um_I.iw[8] ,
    \top_I.branch[14].block[4].um_I.iw[7] ,
    \top_I.branch[14].block[4].um_I.iw[6] ,
    \top_I.branch[14].block[4].um_I.iw[5] ,
    \top_I.branch[14].block[4].um_I.iw[4] ,
    \top_I.branch[14].block[4].um_I.iw[3] ,
    \top_I.branch[14].block[4].um_I.iw[2] ,
    \top_I.branch[14].block[4].um_I.iw[1] ,
    \top_I.branch[14].block[4].um_I.clk ,
    \top_I.branch[14].block[3].um_I.iw[17] ,
    \top_I.branch[14].block[3].um_I.iw[16] ,
    \top_I.branch[14].block[3].um_I.iw[15] ,
    \top_I.branch[14].block[3].um_I.iw[14] ,
    \top_I.branch[14].block[3].um_I.iw[13] ,
    \top_I.branch[14].block[3].um_I.iw[12] ,
    \top_I.branch[14].block[3].um_I.iw[11] ,
    \top_I.branch[14].block[3].um_I.iw[10] ,
    \top_I.branch[14].block[3].um_I.iw[9] ,
    \top_I.branch[14].block[3].um_I.iw[8] ,
    \top_I.branch[14].block[3].um_I.iw[7] ,
    \top_I.branch[14].block[3].um_I.iw[6] ,
    \top_I.branch[14].block[3].um_I.iw[5] ,
    \top_I.branch[14].block[3].um_I.iw[4] ,
    \top_I.branch[14].block[3].um_I.iw[3] ,
    \top_I.branch[14].block[3].um_I.iw[2] ,
    \top_I.branch[14].block[3].um_I.iw[1] ,
    \top_I.branch[14].block[3].um_I.clk ,
    \top_I.branch[14].block[2].um_I.iw[17] ,
    \top_I.branch[14].block[2].um_I.iw[16] ,
    \top_I.branch[14].block[2].um_I.iw[15] ,
    \top_I.branch[14].block[2].um_I.iw[14] ,
    \top_I.branch[14].block[2].um_I.iw[13] ,
    \top_I.branch[14].block[2].um_I.iw[12] ,
    \top_I.branch[14].block[2].um_I.iw[11] ,
    \top_I.branch[14].block[2].um_I.iw[10] ,
    \top_I.branch[14].block[2].um_I.iw[9] ,
    \top_I.branch[14].block[2].um_I.iw[8] ,
    \top_I.branch[14].block[2].um_I.iw[7] ,
    \top_I.branch[14].block[2].um_I.iw[6] ,
    \top_I.branch[14].block[2].um_I.iw[5] ,
    \top_I.branch[14].block[2].um_I.iw[4] ,
    \top_I.branch[14].block[2].um_I.iw[3] ,
    \top_I.branch[14].block[2].um_I.iw[2] ,
    \top_I.branch[14].block[2].um_I.iw[1] ,
    \top_I.branch[14].block[2].um_I.clk ,
    \top_I.branch[14].block[1].um_I.iw[17] ,
    \top_I.branch[14].block[1].um_I.iw[16] ,
    \top_I.branch[14].block[1].um_I.iw[15] ,
    \top_I.branch[14].block[1].um_I.iw[14] ,
    \top_I.branch[14].block[1].um_I.iw[13] ,
    \top_I.branch[14].block[1].um_I.iw[12] ,
    \top_I.branch[14].block[1].um_I.iw[11] ,
    \top_I.branch[14].block[1].um_I.iw[10] ,
    \top_I.branch[14].block[1].um_I.iw[9] ,
    \top_I.branch[14].block[1].um_I.iw[8] ,
    \top_I.branch[14].block[1].um_I.iw[7] ,
    \top_I.branch[14].block[1].um_I.iw[6] ,
    \top_I.branch[14].block[1].um_I.iw[5] ,
    \top_I.branch[14].block[1].um_I.iw[4] ,
    \top_I.branch[14].block[1].um_I.iw[3] ,
    \top_I.branch[14].block[1].um_I.iw[2] ,
    \top_I.branch[14].block[1].um_I.iw[1] ,
    \top_I.branch[14].block[1].um_I.clk ,
    \top_I.branch[14].block[0].um_I.iw[17] ,
    \top_I.branch[14].block[0].um_I.iw[16] ,
    \top_I.branch[14].block[0].um_I.iw[15] ,
    \top_I.branch[14].block[0].um_I.iw[14] ,
    \top_I.branch[14].block[0].um_I.iw[13] ,
    \top_I.branch[14].block[0].um_I.iw[12] ,
    \top_I.branch[14].block[0].um_I.iw[11] ,
    \top_I.branch[14].block[0].um_I.iw[10] ,
    \top_I.branch[14].block[0].um_I.iw[9] ,
    \top_I.branch[14].block[0].um_I.iw[8] ,
    \top_I.branch[14].block[0].um_I.iw[7] ,
    \top_I.branch[14].block[0].um_I.iw[6] ,
    \top_I.branch[14].block[0].um_I.iw[5] ,
    \top_I.branch[14].block[0].um_I.iw[4] ,
    \top_I.branch[14].block[0].um_I.iw[3] ,
    \top_I.branch[14].block[0].um_I.iw[2] ,
    \top_I.branch[14].block[0].um_I.iw[1] ,
    \top_I.branch[14].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[14].block[15].um_I.pg_vdd ,
    \top_I.branch[14].block[14].um_I.pg_vdd ,
    \top_I.branch[14].block[13].um_I.pg_vdd ,
    \top_I.branch[14].block[12].um_I.pg_vdd ,
    \top_I.branch[14].block[11].um_I.pg_vdd ,
    \top_I.branch[14].block[10].um_I.pg_vdd ,
    \top_I.branch[14].block[9].um_I.pg_vdd ,
    \top_I.branch[14].block[8].um_I.pg_vdd ,
    \top_I.branch[14].block[7].um_I.pg_vdd ,
    \top_I.branch[14].block[6].um_I.pg_vdd ,
    \top_I.branch[14].block[5].um_I.pg_vdd ,
    \top_I.branch[14].block[4].um_I.pg_vdd ,
    \top_I.branch[14].block[3].um_I.pg_vdd ,
    \top_I.branch[14].block[2].um_I.pg_vdd ,
    \top_I.branch[14].block[1].um_I.pg_vdd ,
    \top_I.branch[14].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[15].mux_I  (.k_one(\top_I.branch[15].l_addr[0] ),
    .k_zero(\top_I.branch[15].l_addr[3] ),
    .addr({\top_I.branch[15].l_addr[3] ,
    \top_I.branch[15].l_addr[0] ,
    \top_I.branch[15].l_addr[0] ,
    \top_I.branch[15].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[15].block[15].um_I.ena ,
    \top_I.branch[15].block[14].um_I.ena ,
    \top_I.branch[15].block[13].um_I.ena ,
    \top_I.branch[15].block[12].um_I.ena ,
    \top_I.branch[15].block[11].um_I.ena ,
    \top_I.branch[15].block[10].um_I.ena ,
    \top_I.branch[15].block[9].um_I.ena ,
    \top_I.branch[15].block[8].um_I.ena ,
    \top_I.branch[15].block[7].um_I.ena ,
    \top_I.branch[15].block[6].um_I.ena ,
    \top_I.branch[15].block[5].um_I.ena ,
    \top_I.branch[15].block[4].um_I.ena ,
    \top_I.branch[15].block[3].um_I.ena ,
    \top_I.branch[15].block[2].um_I.ena ,
    \top_I.branch[15].block[1].um_I.ena ,
    \top_I.branch[15].block[0].um_I.ena }),
    .um_iw({\top_I.branch[15].block[15].um_I.iw[17] ,
    \top_I.branch[15].block[15].um_I.iw[16] ,
    \top_I.branch[15].block[15].um_I.iw[15] ,
    \top_I.branch[15].block[15].um_I.iw[14] ,
    \top_I.branch[15].block[15].um_I.iw[13] ,
    \top_I.branch[15].block[15].um_I.iw[12] ,
    \top_I.branch[15].block[15].um_I.iw[11] ,
    \top_I.branch[15].block[15].um_I.iw[10] ,
    \top_I.branch[15].block[15].um_I.iw[9] ,
    \top_I.branch[15].block[15].um_I.iw[8] ,
    \top_I.branch[15].block[15].um_I.iw[7] ,
    \top_I.branch[15].block[15].um_I.iw[6] ,
    \top_I.branch[15].block[15].um_I.iw[5] ,
    \top_I.branch[15].block[15].um_I.iw[4] ,
    \top_I.branch[15].block[15].um_I.iw[3] ,
    \top_I.branch[15].block[15].um_I.iw[2] ,
    \top_I.branch[15].block[15].um_I.iw[1] ,
    \top_I.branch[15].block[15].um_I.clk ,
    \top_I.branch[15].block[14].um_I.iw[17] ,
    \top_I.branch[15].block[14].um_I.iw[16] ,
    \top_I.branch[15].block[14].um_I.iw[15] ,
    \top_I.branch[15].block[14].um_I.iw[14] ,
    \top_I.branch[15].block[14].um_I.iw[13] ,
    \top_I.branch[15].block[14].um_I.iw[12] ,
    \top_I.branch[15].block[14].um_I.iw[11] ,
    \top_I.branch[15].block[14].um_I.iw[10] ,
    \top_I.branch[15].block[14].um_I.iw[9] ,
    \top_I.branch[15].block[14].um_I.iw[8] ,
    \top_I.branch[15].block[14].um_I.iw[7] ,
    \top_I.branch[15].block[14].um_I.iw[6] ,
    \top_I.branch[15].block[14].um_I.iw[5] ,
    \top_I.branch[15].block[14].um_I.iw[4] ,
    \top_I.branch[15].block[14].um_I.iw[3] ,
    \top_I.branch[15].block[14].um_I.iw[2] ,
    \top_I.branch[15].block[14].um_I.iw[1] ,
    \top_I.branch[15].block[14].um_I.clk ,
    \top_I.branch[15].block[13].um_I.iw[17] ,
    \top_I.branch[15].block[13].um_I.iw[16] ,
    \top_I.branch[15].block[13].um_I.iw[15] ,
    \top_I.branch[15].block[13].um_I.iw[14] ,
    \top_I.branch[15].block[13].um_I.iw[13] ,
    \top_I.branch[15].block[13].um_I.iw[12] ,
    \top_I.branch[15].block[13].um_I.iw[11] ,
    \top_I.branch[15].block[13].um_I.iw[10] ,
    \top_I.branch[15].block[13].um_I.iw[9] ,
    \top_I.branch[15].block[13].um_I.iw[8] ,
    \top_I.branch[15].block[13].um_I.iw[7] ,
    \top_I.branch[15].block[13].um_I.iw[6] ,
    \top_I.branch[15].block[13].um_I.iw[5] ,
    \top_I.branch[15].block[13].um_I.iw[4] ,
    \top_I.branch[15].block[13].um_I.iw[3] ,
    \top_I.branch[15].block[13].um_I.iw[2] ,
    \top_I.branch[15].block[13].um_I.iw[1] ,
    \top_I.branch[15].block[13].um_I.clk ,
    \top_I.branch[15].block[12].um_I.iw[17] ,
    \top_I.branch[15].block[12].um_I.iw[16] ,
    \top_I.branch[15].block[12].um_I.iw[15] ,
    \top_I.branch[15].block[12].um_I.iw[14] ,
    \top_I.branch[15].block[12].um_I.iw[13] ,
    \top_I.branch[15].block[12].um_I.iw[12] ,
    \top_I.branch[15].block[12].um_I.iw[11] ,
    \top_I.branch[15].block[12].um_I.iw[10] ,
    \top_I.branch[15].block[12].um_I.iw[9] ,
    \top_I.branch[15].block[12].um_I.iw[8] ,
    \top_I.branch[15].block[12].um_I.iw[7] ,
    \top_I.branch[15].block[12].um_I.iw[6] ,
    \top_I.branch[15].block[12].um_I.iw[5] ,
    \top_I.branch[15].block[12].um_I.iw[4] ,
    \top_I.branch[15].block[12].um_I.iw[3] ,
    \top_I.branch[15].block[12].um_I.iw[2] ,
    \top_I.branch[15].block[12].um_I.iw[1] ,
    \top_I.branch[15].block[12].um_I.clk ,
    \top_I.branch[15].block[11].um_I.iw[17] ,
    \top_I.branch[15].block[11].um_I.iw[16] ,
    \top_I.branch[15].block[11].um_I.iw[15] ,
    \top_I.branch[15].block[11].um_I.iw[14] ,
    \top_I.branch[15].block[11].um_I.iw[13] ,
    \top_I.branch[15].block[11].um_I.iw[12] ,
    \top_I.branch[15].block[11].um_I.iw[11] ,
    \top_I.branch[15].block[11].um_I.iw[10] ,
    \top_I.branch[15].block[11].um_I.iw[9] ,
    \top_I.branch[15].block[11].um_I.iw[8] ,
    \top_I.branch[15].block[11].um_I.iw[7] ,
    \top_I.branch[15].block[11].um_I.iw[6] ,
    \top_I.branch[15].block[11].um_I.iw[5] ,
    \top_I.branch[15].block[11].um_I.iw[4] ,
    \top_I.branch[15].block[11].um_I.iw[3] ,
    \top_I.branch[15].block[11].um_I.iw[2] ,
    \top_I.branch[15].block[11].um_I.iw[1] ,
    \top_I.branch[15].block[11].um_I.clk ,
    \top_I.branch[15].block[10].um_I.iw[17] ,
    \top_I.branch[15].block[10].um_I.iw[16] ,
    \top_I.branch[15].block[10].um_I.iw[15] ,
    \top_I.branch[15].block[10].um_I.iw[14] ,
    \top_I.branch[15].block[10].um_I.iw[13] ,
    \top_I.branch[15].block[10].um_I.iw[12] ,
    \top_I.branch[15].block[10].um_I.iw[11] ,
    \top_I.branch[15].block[10].um_I.iw[10] ,
    \top_I.branch[15].block[10].um_I.iw[9] ,
    \top_I.branch[15].block[10].um_I.iw[8] ,
    \top_I.branch[15].block[10].um_I.iw[7] ,
    \top_I.branch[15].block[10].um_I.iw[6] ,
    \top_I.branch[15].block[10].um_I.iw[5] ,
    \top_I.branch[15].block[10].um_I.iw[4] ,
    \top_I.branch[15].block[10].um_I.iw[3] ,
    \top_I.branch[15].block[10].um_I.iw[2] ,
    \top_I.branch[15].block[10].um_I.iw[1] ,
    \top_I.branch[15].block[10].um_I.clk ,
    \top_I.branch[15].block[9].um_I.iw[17] ,
    \top_I.branch[15].block[9].um_I.iw[16] ,
    \top_I.branch[15].block[9].um_I.iw[15] ,
    \top_I.branch[15].block[9].um_I.iw[14] ,
    \top_I.branch[15].block[9].um_I.iw[13] ,
    \top_I.branch[15].block[9].um_I.iw[12] ,
    \top_I.branch[15].block[9].um_I.iw[11] ,
    \top_I.branch[15].block[9].um_I.iw[10] ,
    \top_I.branch[15].block[9].um_I.iw[9] ,
    \top_I.branch[15].block[9].um_I.iw[8] ,
    \top_I.branch[15].block[9].um_I.iw[7] ,
    \top_I.branch[15].block[9].um_I.iw[6] ,
    \top_I.branch[15].block[9].um_I.iw[5] ,
    \top_I.branch[15].block[9].um_I.iw[4] ,
    \top_I.branch[15].block[9].um_I.iw[3] ,
    \top_I.branch[15].block[9].um_I.iw[2] ,
    \top_I.branch[15].block[9].um_I.iw[1] ,
    \top_I.branch[15].block[9].um_I.clk ,
    \top_I.branch[15].block[8].um_I.iw[17] ,
    \top_I.branch[15].block[8].um_I.iw[16] ,
    \top_I.branch[15].block[8].um_I.iw[15] ,
    \top_I.branch[15].block[8].um_I.iw[14] ,
    \top_I.branch[15].block[8].um_I.iw[13] ,
    \top_I.branch[15].block[8].um_I.iw[12] ,
    \top_I.branch[15].block[8].um_I.iw[11] ,
    \top_I.branch[15].block[8].um_I.iw[10] ,
    \top_I.branch[15].block[8].um_I.iw[9] ,
    \top_I.branch[15].block[8].um_I.iw[8] ,
    \top_I.branch[15].block[8].um_I.iw[7] ,
    \top_I.branch[15].block[8].um_I.iw[6] ,
    \top_I.branch[15].block[8].um_I.iw[5] ,
    \top_I.branch[15].block[8].um_I.iw[4] ,
    \top_I.branch[15].block[8].um_I.iw[3] ,
    \top_I.branch[15].block[8].um_I.iw[2] ,
    \top_I.branch[15].block[8].um_I.iw[1] ,
    \top_I.branch[15].block[8].um_I.clk ,
    \top_I.branch[15].block[7].um_I.iw[17] ,
    \top_I.branch[15].block[7].um_I.iw[16] ,
    \top_I.branch[15].block[7].um_I.iw[15] ,
    \top_I.branch[15].block[7].um_I.iw[14] ,
    \top_I.branch[15].block[7].um_I.iw[13] ,
    \top_I.branch[15].block[7].um_I.iw[12] ,
    \top_I.branch[15].block[7].um_I.iw[11] ,
    \top_I.branch[15].block[7].um_I.iw[10] ,
    \top_I.branch[15].block[7].um_I.iw[9] ,
    \top_I.branch[15].block[7].um_I.iw[8] ,
    \top_I.branch[15].block[7].um_I.iw[7] ,
    \top_I.branch[15].block[7].um_I.iw[6] ,
    \top_I.branch[15].block[7].um_I.iw[5] ,
    \top_I.branch[15].block[7].um_I.iw[4] ,
    \top_I.branch[15].block[7].um_I.iw[3] ,
    \top_I.branch[15].block[7].um_I.iw[2] ,
    \top_I.branch[15].block[7].um_I.iw[1] ,
    \top_I.branch[15].block[7].um_I.clk ,
    \top_I.branch[15].block[6].um_I.iw[17] ,
    \top_I.branch[15].block[6].um_I.iw[16] ,
    \top_I.branch[15].block[6].um_I.iw[15] ,
    \top_I.branch[15].block[6].um_I.iw[14] ,
    \top_I.branch[15].block[6].um_I.iw[13] ,
    \top_I.branch[15].block[6].um_I.iw[12] ,
    \top_I.branch[15].block[6].um_I.iw[11] ,
    \top_I.branch[15].block[6].um_I.iw[10] ,
    \top_I.branch[15].block[6].um_I.iw[9] ,
    \top_I.branch[15].block[6].um_I.iw[8] ,
    \top_I.branch[15].block[6].um_I.iw[7] ,
    \top_I.branch[15].block[6].um_I.iw[6] ,
    \top_I.branch[15].block[6].um_I.iw[5] ,
    \top_I.branch[15].block[6].um_I.iw[4] ,
    \top_I.branch[15].block[6].um_I.iw[3] ,
    \top_I.branch[15].block[6].um_I.iw[2] ,
    \top_I.branch[15].block[6].um_I.iw[1] ,
    \top_I.branch[15].block[6].um_I.clk ,
    \top_I.branch[15].block[5].um_I.iw[17] ,
    \top_I.branch[15].block[5].um_I.iw[16] ,
    \top_I.branch[15].block[5].um_I.iw[15] ,
    \top_I.branch[15].block[5].um_I.iw[14] ,
    \top_I.branch[15].block[5].um_I.iw[13] ,
    \top_I.branch[15].block[5].um_I.iw[12] ,
    \top_I.branch[15].block[5].um_I.iw[11] ,
    \top_I.branch[15].block[5].um_I.iw[10] ,
    \top_I.branch[15].block[5].um_I.iw[9] ,
    \top_I.branch[15].block[5].um_I.iw[8] ,
    \top_I.branch[15].block[5].um_I.iw[7] ,
    \top_I.branch[15].block[5].um_I.iw[6] ,
    \top_I.branch[15].block[5].um_I.iw[5] ,
    \top_I.branch[15].block[5].um_I.iw[4] ,
    \top_I.branch[15].block[5].um_I.iw[3] ,
    \top_I.branch[15].block[5].um_I.iw[2] ,
    \top_I.branch[15].block[5].um_I.iw[1] ,
    \top_I.branch[15].block[5].um_I.clk ,
    \top_I.branch[15].block[4].um_I.iw[17] ,
    \top_I.branch[15].block[4].um_I.iw[16] ,
    \top_I.branch[15].block[4].um_I.iw[15] ,
    \top_I.branch[15].block[4].um_I.iw[14] ,
    \top_I.branch[15].block[4].um_I.iw[13] ,
    \top_I.branch[15].block[4].um_I.iw[12] ,
    \top_I.branch[15].block[4].um_I.iw[11] ,
    \top_I.branch[15].block[4].um_I.iw[10] ,
    \top_I.branch[15].block[4].um_I.iw[9] ,
    \top_I.branch[15].block[4].um_I.iw[8] ,
    \top_I.branch[15].block[4].um_I.iw[7] ,
    \top_I.branch[15].block[4].um_I.iw[6] ,
    \top_I.branch[15].block[4].um_I.iw[5] ,
    \top_I.branch[15].block[4].um_I.iw[4] ,
    \top_I.branch[15].block[4].um_I.iw[3] ,
    \top_I.branch[15].block[4].um_I.iw[2] ,
    \top_I.branch[15].block[4].um_I.iw[1] ,
    \top_I.branch[15].block[4].um_I.clk ,
    \top_I.branch[15].block[3].um_I.iw[17] ,
    \top_I.branch[15].block[3].um_I.iw[16] ,
    \top_I.branch[15].block[3].um_I.iw[15] ,
    \top_I.branch[15].block[3].um_I.iw[14] ,
    \top_I.branch[15].block[3].um_I.iw[13] ,
    \top_I.branch[15].block[3].um_I.iw[12] ,
    \top_I.branch[15].block[3].um_I.iw[11] ,
    \top_I.branch[15].block[3].um_I.iw[10] ,
    \top_I.branch[15].block[3].um_I.iw[9] ,
    \top_I.branch[15].block[3].um_I.iw[8] ,
    \top_I.branch[15].block[3].um_I.iw[7] ,
    \top_I.branch[15].block[3].um_I.iw[6] ,
    \top_I.branch[15].block[3].um_I.iw[5] ,
    \top_I.branch[15].block[3].um_I.iw[4] ,
    \top_I.branch[15].block[3].um_I.iw[3] ,
    \top_I.branch[15].block[3].um_I.iw[2] ,
    \top_I.branch[15].block[3].um_I.iw[1] ,
    \top_I.branch[15].block[3].um_I.clk ,
    \top_I.branch[15].block[2].um_I.iw[17] ,
    \top_I.branch[15].block[2].um_I.iw[16] ,
    \top_I.branch[15].block[2].um_I.iw[15] ,
    \top_I.branch[15].block[2].um_I.iw[14] ,
    \top_I.branch[15].block[2].um_I.iw[13] ,
    \top_I.branch[15].block[2].um_I.iw[12] ,
    \top_I.branch[15].block[2].um_I.iw[11] ,
    \top_I.branch[15].block[2].um_I.iw[10] ,
    \top_I.branch[15].block[2].um_I.iw[9] ,
    \top_I.branch[15].block[2].um_I.iw[8] ,
    \top_I.branch[15].block[2].um_I.iw[7] ,
    \top_I.branch[15].block[2].um_I.iw[6] ,
    \top_I.branch[15].block[2].um_I.iw[5] ,
    \top_I.branch[15].block[2].um_I.iw[4] ,
    \top_I.branch[15].block[2].um_I.iw[3] ,
    \top_I.branch[15].block[2].um_I.iw[2] ,
    \top_I.branch[15].block[2].um_I.iw[1] ,
    \top_I.branch[15].block[2].um_I.clk ,
    \top_I.branch[15].block[1].um_I.iw[17] ,
    \top_I.branch[15].block[1].um_I.iw[16] ,
    \top_I.branch[15].block[1].um_I.iw[15] ,
    \top_I.branch[15].block[1].um_I.iw[14] ,
    \top_I.branch[15].block[1].um_I.iw[13] ,
    \top_I.branch[15].block[1].um_I.iw[12] ,
    \top_I.branch[15].block[1].um_I.iw[11] ,
    \top_I.branch[15].block[1].um_I.iw[10] ,
    \top_I.branch[15].block[1].um_I.iw[9] ,
    \top_I.branch[15].block[1].um_I.iw[8] ,
    \top_I.branch[15].block[1].um_I.iw[7] ,
    \top_I.branch[15].block[1].um_I.iw[6] ,
    \top_I.branch[15].block[1].um_I.iw[5] ,
    \top_I.branch[15].block[1].um_I.iw[4] ,
    \top_I.branch[15].block[1].um_I.iw[3] ,
    \top_I.branch[15].block[1].um_I.iw[2] ,
    \top_I.branch[15].block[1].um_I.iw[1] ,
    \top_I.branch[15].block[1].um_I.clk ,
    \top_I.branch[15].block[0].um_I.iw[17] ,
    \top_I.branch[15].block[0].um_I.iw[16] ,
    \top_I.branch[15].block[0].um_I.iw[15] ,
    \top_I.branch[15].block[0].um_I.iw[14] ,
    \top_I.branch[15].block[0].um_I.iw[13] ,
    \top_I.branch[15].block[0].um_I.iw[12] ,
    \top_I.branch[15].block[0].um_I.iw[11] ,
    \top_I.branch[15].block[0].um_I.iw[10] ,
    \top_I.branch[15].block[0].um_I.iw[9] ,
    \top_I.branch[15].block[0].um_I.iw[8] ,
    \top_I.branch[15].block[0].um_I.iw[7] ,
    \top_I.branch[15].block[0].um_I.iw[6] ,
    \top_I.branch[15].block[0].um_I.iw[5] ,
    \top_I.branch[15].block[0].um_I.iw[4] ,
    \top_I.branch[15].block[0].um_I.iw[3] ,
    \top_I.branch[15].block[0].um_I.iw[2] ,
    \top_I.branch[15].block[0].um_I.iw[1] ,
    \top_I.branch[15].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[15].block[15].um_I.pg_vdd ,
    \top_I.branch[15].block[14].um_I.pg_vdd ,
    \top_I.branch[15].block[13].um_I.pg_vdd ,
    \top_I.branch[15].block[12].um_I.pg_vdd ,
    \top_I.branch[15].block[11].um_I.pg_vdd ,
    \top_I.branch[15].block[10].um_I.pg_vdd ,
    \top_I.branch[15].block[9].um_I.pg_vdd ,
    \top_I.branch[15].block[8].um_I.pg_vdd ,
    \top_I.branch[15].block[7].um_I.pg_vdd ,
    \top_I.branch[15].block[6].um_I.pg_vdd ,
    \top_I.branch[15].block[5].um_I.pg_vdd ,
    \top_I.branch[15].block[4].um_I.pg_vdd ,
    \top_I.branch[15].block[3].um_I.pg_vdd ,
    \top_I.branch[15].block[2].um_I.pg_vdd ,
    \top_I.branch[15].block[1].um_I.pg_vdd ,
    \top_I.branch[15].block[0].um_I.pg_vdd }));
 tt_um_factory_test \top_I.branch[16].block[4].um_I.block_16_4.tt_um_I  (.clk(\top_I.branch[16].block[4].um_I.clk ),
    .ena(\top_I.branch[16].block[4].um_I.ena ),
    .rst_n(\top_I.branch[16].block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[16].block[4].um_I.iw[9] ,
    \top_I.branch[16].block[4].um_I.iw[8] ,
    \top_I.branch[16].block[4].um_I.iw[7] ,
    \top_I.branch[16].block[4].um_I.iw[6] ,
    \top_I.branch[16].block[4].um_I.iw[5] ,
    \top_I.branch[16].block[4].um_I.iw[4] ,
    \top_I.branch[16].block[4].um_I.iw[3] ,
    \top_I.branch[16].block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[16].block[4].um_I.iw[17] ,
    \top_I.branch[16].block[4].um_I.iw[16] ,
    \top_I.branch[16].block[4].um_I.iw[15] ,
    \top_I.branch[16].block[4].um_I.iw[14] ,
    \top_I.branch[16].block[4].um_I.iw[13] ,
    \top_I.branch[16].block[4].um_I.iw[12] ,
    \top_I.branch[16].block[4].um_I.iw[11] ,
    \top_I.branch[16].block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[16].block[4].um_I.ow[23] ,
    \top_I.branch[16].block[4].um_I.ow[22] ,
    \top_I.branch[16].block[4].um_I.ow[21] ,
    \top_I.branch[16].block[4].um_I.ow[20] ,
    \top_I.branch[16].block[4].um_I.ow[19] ,
    \top_I.branch[16].block[4].um_I.ow[18] ,
    \top_I.branch[16].block[4].um_I.ow[17] ,
    \top_I.branch[16].block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[16].block[4].um_I.ow[15] ,
    \top_I.branch[16].block[4].um_I.ow[14] ,
    \top_I.branch[16].block[4].um_I.ow[13] ,
    \top_I.branch[16].block[4].um_I.ow[12] ,
    \top_I.branch[16].block[4].um_I.ow[11] ,
    \top_I.branch[16].block[4].um_I.ow[10] ,
    \top_I.branch[16].block[4].um_I.ow[9] ,
    \top_I.branch[16].block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[16].block[4].um_I.ow[7] ,
    \top_I.branch[16].block[4].um_I.ow[6] ,
    \top_I.branch[16].block[4].um_I.ow[5] ,
    \top_I.branch[16].block[4].um_I.ow[4] ,
    \top_I.branch[16].block[4].um_I.ow[3] ,
    \top_I.branch[16].block[4].um_I.ow[2] ,
    \top_I.branch[16].block[4].um_I.ow[1] ,
    \top_I.branch[16].block[4].um_I.ow[0] }));
 tt_mux \top_I.branch[16].mux_I  (.k_one(\top_I.branch[16].l_addr[3] ),
    .k_zero(\top_I.branch[16].l_addr[0] ),
    .addr({\top_I.branch[16].l_addr[3] ,
    \top_I.branch[16].l_addr[0] ,
    \top_I.branch[16].l_addr[0] ,
    \top_I.branch[16].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[16].block[15].um_I.ena ,
    \top_I.branch[16].block[14].um_I.ena ,
    \top_I.branch[16].block[13].um_I.ena ,
    \top_I.branch[16].block[12].um_I.ena ,
    \top_I.branch[16].block[11].um_I.ena ,
    \top_I.branch[16].block[10].um_I.ena ,
    \top_I.branch[16].block[9].um_I.ena ,
    \top_I.branch[16].block[8].um_I.ena ,
    \top_I.branch[16].block[7].um_I.ena ,
    \top_I.branch[16].block[6].um_I.ena ,
    \top_I.branch[16].block[5].um_I.ena ,
    \top_I.branch[16].block[4].um_I.ena ,
    \top_I.branch[16].block[3].um_I.ena ,
    \top_I.branch[16].block[2].um_I.ena ,
    \top_I.branch[16].block[1].um_I.ena ,
    \top_I.branch[16].block[0].um_I.ena }),
    .um_iw({\top_I.branch[16].block[15].um_I.iw[17] ,
    \top_I.branch[16].block[15].um_I.iw[16] ,
    \top_I.branch[16].block[15].um_I.iw[15] ,
    \top_I.branch[16].block[15].um_I.iw[14] ,
    \top_I.branch[16].block[15].um_I.iw[13] ,
    \top_I.branch[16].block[15].um_I.iw[12] ,
    \top_I.branch[16].block[15].um_I.iw[11] ,
    \top_I.branch[16].block[15].um_I.iw[10] ,
    \top_I.branch[16].block[15].um_I.iw[9] ,
    \top_I.branch[16].block[15].um_I.iw[8] ,
    \top_I.branch[16].block[15].um_I.iw[7] ,
    \top_I.branch[16].block[15].um_I.iw[6] ,
    \top_I.branch[16].block[15].um_I.iw[5] ,
    \top_I.branch[16].block[15].um_I.iw[4] ,
    \top_I.branch[16].block[15].um_I.iw[3] ,
    \top_I.branch[16].block[15].um_I.iw[2] ,
    \top_I.branch[16].block[15].um_I.iw[1] ,
    \top_I.branch[16].block[15].um_I.clk ,
    \top_I.branch[16].block[14].um_I.iw[17] ,
    \top_I.branch[16].block[14].um_I.iw[16] ,
    \top_I.branch[16].block[14].um_I.iw[15] ,
    \top_I.branch[16].block[14].um_I.iw[14] ,
    \top_I.branch[16].block[14].um_I.iw[13] ,
    \top_I.branch[16].block[14].um_I.iw[12] ,
    \top_I.branch[16].block[14].um_I.iw[11] ,
    \top_I.branch[16].block[14].um_I.iw[10] ,
    \top_I.branch[16].block[14].um_I.iw[9] ,
    \top_I.branch[16].block[14].um_I.iw[8] ,
    \top_I.branch[16].block[14].um_I.iw[7] ,
    \top_I.branch[16].block[14].um_I.iw[6] ,
    \top_I.branch[16].block[14].um_I.iw[5] ,
    \top_I.branch[16].block[14].um_I.iw[4] ,
    \top_I.branch[16].block[14].um_I.iw[3] ,
    \top_I.branch[16].block[14].um_I.iw[2] ,
    \top_I.branch[16].block[14].um_I.iw[1] ,
    \top_I.branch[16].block[14].um_I.clk ,
    \top_I.branch[16].block[13].um_I.iw[17] ,
    \top_I.branch[16].block[13].um_I.iw[16] ,
    \top_I.branch[16].block[13].um_I.iw[15] ,
    \top_I.branch[16].block[13].um_I.iw[14] ,
    \top_I.branch[16].block[13].um_I.iw[13] ,
    \top_I.branch[16].block[13].um_I.iw[12] ,
    \top_I.branch[16].block[13].um_I.iw[11] ,
    \top_I.branch[16].block[13].um_I.iw[10] ,
    \top_I.branch[16].block[13].um_I.iw[9] ,
    \top_I.branch[16].block[13].um_I.iw[8] ,
    \top_I.branch[16].block[13].um_I.iw[7] ,
    \top_I.branch[16].block[13].um_I.iw[6] ,
    \top_I.branch[16].block[13].um_I.iw[5] ,
    \top_I.branch[16].block[13].um_I.iw[4] ,
    \top_I.branch[16].block[13].um_I.iw[3] ,
    \top_I.branch[16].block[13].um_I.iw[2] ,
    \top_I.branch[16].block[13].um_I.iw[1] ,
    \top_I.branch[16].block[13].um_I.clk ,
    \top_I.branch[16].block[12].um_I.iw[17] ,
    \top_I.branch[16].block[12].um_I.iw[16] ,
    \top_I.branch[16].block[12].um_I.iw[15] ,
    \top_I.branch[16].block[12].um_I.iw[14] ,
    \top_I.branch[16].block[12].um_I.iw[13] ,
    \top_I.branch[16].block[12].um_I.iw[12] ,
    \top_I.branch[16].block[12].um_I.iw[11] ,
    \top_I.branch[16].block[12].um_I.iw[10] ,
    \top_I.branch[16].block[12].um_I.iw[9] ,
    \top_I.branch[16].block[12].um_I.iw[8] ,
    \top_I.branch[16].block[12].um_I.iw[7] ,
    \top_I.branch[16].block[12].um_I.iw[6] ,
    \top_I.branch[16].block[12].um_I.iw[5] ,
    \top_I.branch[16].block[12].um_I.iw[4] ,
    \top_I.branch[16].block[12].um_I.iw[3] ,
    \top_I.branch[16].block[12].um_I.iw[2] ,
    \top_I.branch[16].block[12].um_I.iw[1] ,
    \top_I.branch[16].block[12].um_I.clk ,
    \top_I.branch[16].block[11].um_I.iw[17] ,
    \top_I.branch[16].block[11].um_I.iw[16] ,
    \top_I.branch[16].block[11].um_I.iw[15] ,
    \top_I.branch[16].block[11].um_I.iw[14] ,
    \top_I.branch[16].block[11].um_I.iw[13] ,
    \top_I.branch[16].block[11].um_I.iw[12] ,
    \top_I.branch[16].block[11].um_I.iw[11] ,
    \top_I.branch[16].block[11].um_I.iw[10] ,
    \top_I.branch[16].block[11].um_I.iw[9] ,
    \top_I.branch[16].block[11].um_I.iw[8] ,
    \top_I.branch[16].block[11].um_I.iw[7] ,
    \top_I.branch[16].block[11].um_I.iw[6] ,
    \top_I.branch[16].block[11].um_I.iw[5] ,
    \top_I.branch[16].block[11].um_I.iw[4] ,
    \top_I.branch[16].block[11].um_I.iw[3] ,
    \top_I.branch[16].block[11].um_I.iw[2] ,
    \top_I.branch[16].block[11].um_I.iw[1] ,
    \top_I.branch[16].block[11].um_I.clk ,
    \top_I.branch[16].block[10].um_I.iw[17] ,
    \top_I.branch[16].block[10].um_I.iw[16] ,
    \top_I.branch[16].block[10].um_I.iw[15] ,
    \top_I.branch[16].block[10].um_I.iw[14] ,
    \top_I.branch[16].block[10].um_I.iw[13] ,
    \top_I.branch[16].block[10].um_I.iw[12] ,
    \top_I.branch[16].block[10].um_I.iw[11] ,
    \top_I.branch[16].block[10].um_I.iw[10] ,
    \top_I.branch[16].block[10].um_I.iw[9] ,
    \top_I.branch[16].block[10].um_I.iw[8] ,
    \top_I.branch[16].block[10].um_I.iw[7] ,
    \top_I.branch[16].block[10].um_I.iw[6] ,
    \top_I.branch[16].block[10].um_I.iw[5] ,
    \top_I.branch[16].block[10].um_I.iw[4] ,
    \top_I.branch[16].block[10].um_I.iw[3] ,
    \top_I.branch[16].block[10].um_I.iw[2] ,
    \top_I.branch[16].block[10].um_I.iw[1] ,
    \top_I.branch[16].block[10].um_I.clk ,
    \top_I.branch[16].block[9].um_I.iw[17] ,
    \top_I.branch[16].block[9].um_I.iw[16] ,
    \top_I.branch[16].block[9].um_I.iw[15] ,
    \top_I.branch[16].block[9].um_I.iw[14] ,
    \top_I.branch[16].block[9].um_I.iw[13] ,
    \top_I.branch[16].block[9].um_I.iw[12] ,
    \top_I.branch[16].block[9].um_I.iw[11] ,
    \top_I.branch[16].block[9].um_I.iw[10] ,
    \top_I.branch[16].block[9].um_I.iw[9] ,
    \top_I.branch[16].block[9].um_I.iw[8] ,
    \top_I.branch[16].block[9].um_I.iw[7] ,
    \top_I.branch[16].block[9].um_I.iw[6] ,
    \top_I.branch[16].block[9].um_I.iw[5] ,
    \top_I.branch[16].block[9].um_I.iw[4] ,
    \top_I.branch[16].block[9].um_I.iw[3] ,
    \top_I.branch[16].block[9].um_I.iw[2] ,
    \top_I.branch[16].block[9].um_I.iw[1] ,
    \top_I.branch[16].block[9].um_I.clk ,
    \top_I.branch[16].block[8].um_I.iw[17] ,
    \top_I.branch[16].block[8].um_I.iw[16] ,
    \top_I.branch[16].block[8].um_I.iw[15] ,
    \top_I.branch[16].block[8].um_I.iw[14] ,
    \top_I.branch[16].block[8].um_I.iw[13] ,
    \top_I.branch[16].block[8].um_I.iw[12] ,
    \top_I.branch[16].block[8].um_I.iw[11] ,
    \top_I.branch[16].block[8].um_I.iw[10] ,
    \top_I.branch[16].block[8].um_I.iw[9] ,
    \top_I.branch[16].block[8].um_I.iw[8] ,
    \top_I.branch[16].block[8].um_I.iw[7] ,
    \top_I.branch[16].block[8].um_I.iw[6] ,
    \top_I.branch[16].block[8].um_I.iw[5] ,
    \top_I.branch[16].block[8].um_I.iw[4] ,
    \top_I.branch[16].block[8].um_I.iw[3] ,
    \top_I.branch[16].block[8].um_I.iw[2] ,
    \top_I.branch[16].block[8].um_I.iw[1] ,
    \top_I.branch[16].block[8].um_I.clk ,
    \top_I.branch[16].block[7].um_I.iw[17] ,
    \top_I.branch[16].block[7].um_I.iw[16] ,
    \top_I.branch[16].block[7].um_I.iw[15] ,
    \top_I.branch[16].block[7].um_I.iw[14] ,
    \top_I.branch[16].block[7].um_I.iw[13] ,
    \top_I.branch[16].block[7].um_I.iw[12] ,
    \top_I.branch[16].block[7].um_I.iw[11] ,
    \top_I.branch[16].block[7].um_I.iw[10] ,
    \top_I.branch[16].block[7].um_I.iw[9] ,
    \top_I.branch[16].block[7].um_I.iw[8] ,
    \top_I.branch[16].block[7].um_I.iw[7] ,
    \top_I.branch[16].block[7].um_I.iw[6] ,
    \top_I.branch[16].block[7].um_I.iw[5] ,
    \top_I.branch[16].block[7].um_I.iw[4] ,
    \top_I.branch[16].block[7].um_I.iw[3] ,
    \top_I.branch[16].block[7].um_I.iw[2] ,
    \top_I.branch[16].block[7].um_I.iw[1] ,
    \top_I.branch[16].block[7].um_I.clk ,
    \top_I.branch[16].block[6].um_I.iw[17] ,
    \top_I.branch[16].block[6].um_I.iw[16] ,
    \top_I.branch[16].block[6].um_I.iw[15] ,
    \top_I.branch[16].block[6].um_I.iw[14] ,
    \top_I.branch[16].block[6].um_I.iw[13] ,
    \top_I.branch[16].block[6].um_I.iw[12] ,
    \top_I.branch[16].block[6].um_I.iw[11] ,
    \top_I.branch[16].block[6].um_I.iw[10] ,
    \top_I.branch[16].block[6].um_I.iw[9] ,
    \top_I.branch[16].block[6].um_I.iw[8] ,
    \top_I.branch[16].block[6].um_I.iw[7] ,
    \top_I.branch[16].block[6].um_I.iw[6] ,
    \top_I.branch[16].block[6].um_I.iw[5] ,
    \top_I.branch[16].block[6].um_I.iw[4] ,
    \top_I.branch[16].block[6].um_I.iw[3] ,
    \top_I.branch[16].block[6].um_I.iw[2] ,
    \top_I.branch[16].block[6].um_I.iw[1] ,
    \top_I.branch[16].block[6].um_I.clk ,
    \top_I.branch[16].block[5].um_I.iw[17] ,
    \top_I.branch[16].block[5].um_I.iw[16] ,
    \top_I.branch[16].block[5].um_I.iw[15] ,
    \top_I.branch[16].block[5].um_I.iw[14] ,
    \top_I.branch[16].block[5].um_I.iw[13] ,
    \top_I.branch[16].block[5].um_I.iw[12] ,
    \top_I.branch[16].block[5].um_I.iw[11] ,
    \top_I.branch[16].block[5].um_I.iw[10] ,
    \top_I.branch[16].block[5].um_I.iw[9] ,
    \top_I.branch[16].block[5].um_I.iw[8] ,
    \top_I.branch[16].block[5].um_I.iw[7] ,
    \top_I.branch[16].block[5].um_I.iw[6] ,
    \top_I.branch[16].block[5].um_I.iw[5] ,
    \top_I.branch[16].block[5].um_I.iw[4] ,
    \top_I.branch[16].block[5].um_I.iw[3] ,
    \top_I.branch[16].block[5].um_I.iw[2] ,
    \top_I.branch[16].block[5].um_I.iw[1] ,
    \top_I.branch[16].block[5].um_I.clk ,
    \top_I.branch[16].block[4].um_I.iw[17] ,
    \top_I.branch[16].block[4].um_I.iw[16] ,
    \top_I.branch[16].block[4].um_I.iw[15] ,
    \top_I.branch[16].block[4].um_I.iw[14] ,
    \top_I.branch[16].block[4].um_I.iw[13] ,
    \top_I.branch[16].block[4].um_I.iw[12] ,
    \top_I.branch[16].block[4].um_I.iw[11] ,
    \top_I.branch[16].block[4].um_I.iw[10] ,
    \top_I.branch[16].block[4].um_I.iw[9] ,
    \top_I.branch[16].block[4].um_I.iw[8] ,
    \top_I.branch[16].block[4].um_I.iw[7] ,
    \top_I.branch[16].block[4].um_I.iw[6] ,
    \top_I.branch[16].block[4].um_I.iw[5] ,
    \top_I.branch[16].block[4].um_I.iw[4] ,
    \top_I.branch[16].block[4].um_I.iw[3] ,
    \top_I.branch[16].block[4].um_I.iw[2] ,
    \top_I.branch[16].block[4].um_I.iw[1] ,
    \top_I.branch[16].block[4].um_I.clk ,
    \top_I.branch[16].block[3].um_I.iw[17] ,
    \top_I.branch[16].block[3].um_I.iw[16] ,
    \top_I.branch[16].block[3].um_I.iw[15] ,
    \top_I.branch[16].block[3].um_I.iw[14] ,
    \top_I.branch[16].block[3].um_I.iw[13] ,
    \top_I.branch[16].block[3].um_I.iw[12] ,
    \top_I.branch[16].block[3].um_I.iw[11] ,
    \top_I.branch[16].block[3].um_I.iw[10] ,
    \top_I.branch[16].block[3].um_I.iw[9] ,
    \top_I.branch[16].block[3].um_I.iw[8] ,
    \top_I.branch[16].block[3].um_I.iw[7] ,
    \top_I.branch[16].block[3].um_I.iw[6] ,
    \top_I.branch[16].block[3].um_I.iw[5] ,
    \top_I.branch[16].block[3].um_I.iw[4] ,
    \top_I.branch[16].block[3].um_I.iw[3] ,
    \top_I.branch[16].block[3].um_I.iw[2] ,
    \top_I.branch[16].block[3].um_I.iw[1] ,
    \top_I.branch[16].block[3].um_I.clk ,
    \top_I.branch[16].block[2].um_I.iw[17] ,
    \top_I.branch[16].block[2].um_I.iw[16] ,
    \top_I.branch[16].block[2].um_I.iw[15] ,
    \top_I.branch[16].block[2].um_I.iw[14] ,
    \top_I.branch[16].block[2].um_I.iw[13] ,
    \top_I.branch[16].block[2].um_I.iw[12] ,
    \top_I.branch[16].block[2].um_I.iw[11] ,
    \top_I.branch[16].block[2].um_I.iw[10] ,
    \top_I.branch[16].block[2].um_I.iw[9] ,
    \top_I.branch[16].block[2].um_I.iw[8] ,
    \top_I.branch[16].block[2].um_I.iw[7] ,
    \top_I.branch[16].block[2].um_I.iw[6] ,
    \top_I.branch[16].block[2].um_I.iw[5] ,
    \top_I.branch[16].block[2].um_I.iw[4] ,
    \top_I.branch[16].block[2].um_I.iw[3] ,
    \top_I.branch[16].block[2].um_I.iw[2] ,
    \top_I.branch[16].block[2].um_I.iw[1] ,
    \top_I.branch[16].block[2].um_I.clk ,
    \top_I.branch[16].block[1].um_I.iw[17] ,
    \top_I.branch[16].block[1].um_I.iw[16] ,
    \top_I.branch[16].block[1].um_I.iw[15] ,
    \top_I.branch[16].block[1].um_I.iw[14] ,
    \top_I.branch[16].block[1].um_I.iw[13] ,
    \top_I.branch[16].block[1].um_I.iw[12] ,
    \top_I.branch[16].block[1].um_I.iw[11] ,
    \top_I.branch[16].block[1].um_I.iw[10] ,
    \top_I.branch[16].block[1].um_I.iw[9] ,
    \top_I.branch[16].block[1].um_I.iw[8] ,
    \top_I.branch[16].block[1].um_I.iw[7] ,
    \top_I.branch[16].block[1].um_I.iw[6] ,
    \top_I.branch[16].block[1].um_I.iw[5] ,
    \top_I.branch[16].block[1].um_I.iw[4] ,
    \top_I.branch[16].block[1].um_I.iw[3] ,
    \top_I.branch[16].block[1].um_I.iw[2] ,
    \top_I.branch[16].block[1].um_I.iw[1] ,
    \top_I.branch[16].block[1].um_I.clk ,
    \top_I.branch[16].block[0].um_I.iw[17] ,
    \top_I.branch[16].block[0].um_I.iw[16] ,
    \top_I.branch[16].block[0].um_I.iw[15] ,
    \top_I.branch[16].block[0].um_I.iw[14] ,
    \top_I.branch[16].block[0].um_I.iw[13] ,
    \top_I.branch[16].block[0].um_I.iw[12] ,
    \top_I.branch[16].block[0].um_I.iw[11] ,
    \top_I.branch[16].block[0].um_I.iw[10] ,
    \top_I.branch[16].block[0].um_I.iw[9] ,
    \top_I.branch[16].block[0].um_I.iw[8] ,
    \top_I.branch[16].block[0].um_I.iw[7] ,
    \top_I.branch[16].block[0].um_I.iw[6] ,
    \top_I.branch[16].block[0].um_I.iw[5] ,
    \top_I.branch[16].block[0].um_I.iw[4] ,
    \top_I.branch[16].block[0].um_I.iw[3] ,
    \top_I.branch[16].block[0].um_I.iw[2] ,
    \top_I.branch[16].block[0].um_I.iw[1] ,
    \top_I.branch[16].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.ow[23] ,
    \top_I.branch[16].block[4].um_I.ow[22] ,
    \top_I.branch[16].block[4].um_I.ow[21] ,
    \top_I.branch[16].block[4].um_I.ow[20] ,
    \top_I.branch[16].block[4].um_I.ow[19] ,
    \top_I.branch[16].block[4].um_I.ow[18] ,
    \top_I.branch[16].block[4].um_I.ow[17] ,
    \top_I.branch[16].block[4].um_I.ow[16] ,
    \top_I.branch[16].block[4].um_I.ow[15] ,
    \top_I.branch[16].block[4].um_I.ow[14] ,
    \top_I.branch[16].block[4].um_I.ow[13] ,
    \top_I.branch[16].block[4].um_I.ow[12] ,
    \top_I.branch[16].block[4].um_I.ow[11] ,
    \top_I.branch[16].block[4].um_I.ow[10] ,
    \top_I.branch[16].block[4].um_I.ow[9] ,
    \top_I.branch[16].block[4].um_I.ow[8] ,
    \top_I.branch[16].block[4].um_I.ow[7] ,
    \top_I.branch[16].block[4].um_I.ow[6] ,
    \top_I.branch[16].block[4].um_I.ow[5] ,
    \top_I.branch[16].block[4].um_I.ow[4] ,
    \top_I.branch[16].block[4].um_I.ow[3] ,
    \top_I.branch[16].block[4].um_I.ow[2] ,
    \top_I.branch[16].block[4].um_I.ow[1] ,
    \top_I.branch[16].block[4].um_I.ow[0] ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[16].block[15].um_I.pg_vdd ,
    \top_I.branch[16].block[14].um_I.pg_vdd ,
    \top_I.branch[16].block[13].um_I.pg_vdd ,
    \top_I.branch[16].block[12].um_I.pg_vdd ,
    \top_I.branch[16].block[11].um_I.pg_vdd ,
    \top_I.branch[16].block[10].um_I.pg_vdd ,
    \top_I.branch[16].block[9].um_I.pg_vdd ,
    \top_I.branch[16].block[8].um_I.pg_vdd ,
    \top_I.branch[16].block[7].um_I.pg_vdd ,
    \top_I.branch[16].block[6].um_I.pg_vdd ,
    \top_I.branch[16].block[5].um_I.pg_vdd ,
    \top_I.branch[16].block[4].um_I.pg_vdd ,
    \top_I.branch[16].block[3].um_I.pg_vdd ,
    \top_I.branch[16].block[2].um_I.pg_vdd ,
    \top_I.branch[16].block[1].um_I.pg_vdd ,
    \top_I.branch[16].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[17].mux_I  (.k_one(\top_I.branch[17].l_addr[3] ),
    .k_zero(\top_I.branch[17].l_addr[0] ),
    .addr({\top_I.branch[17].l_addr[3] ,
    \top_I.branch[17].l_addr[0] ,
    \top_I.branch[17].l_addr[0] ,
    \top_I.branch[17].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[17].block[15].um_I.ena ,
    \top_I.branch[17].block[14].um_I.ena ,
    \top_I.branch[17].block[13].um_I.ena ,
    \top_I.branch[17].block[12].um_I.ena ,
    \top_I.branch[17].block[11].um_I.ena ,
    \top_I.branch[17].block[10].um_I.ena ,
    \top_I.branch[17].block[9].um_I.ena ,
    \top_I.branch[17].block[8].um_I.ena ,
    \top_I.branch[17].block[7].um_I.ena ,
    \top_I.branch[17].block[6].um_I.ena ,
    \top_I.branch[17].block[5].um_I.ena ,
    \top_I.branch[17].block[4].um_I.ena ,
    \top_I.branch[17].block[3].um_I.ena ,
    \top_I.branch[17].block[2].um_I.ena ,
    \top_I.branch[17].block[1].um_I.ena ,
    \top_I.branch[17].block[0].um_I.ena }),
    .um_iw({\top_I.branch[17].block[15].um_I.iw[17] ,
    \top_I.branch[17].block[15].um_I.iw[16] ,
    \top_I.branch[17].block[15].um_I.iw[15] ,
    \top_I.branch[17].block[15].um_I.iw[14] ,
    \top_I.branch[17].block[15].um_I.iw[13] ,
    \top_I.branch[17].block[15].um_I.iw[12] ,
    \top_I.branch[17].block[15].um_I.iw[11] ,
    \top_I.branch[17].block[15].um_I.iw[10] ,
    \top_I.branch[17].block[15].um_I.iw[9] ,
    \top_I.branch[17].block[15].um_I.iw[8] ,
    \top_I.branch[17].block[15].um_I.iw[7] ,
    \top_I.branch[17].block[15].um_I.iw[6] ,
    \top_I.branch[17].block[15].um_I.iw[5] ,
    \top_I.branch[17].block[15].um_I.iw[4] ,
    \top_I.branch[17].block[15].um_I.iw[3] ,
    \top_I.branch[17].block[15].um_I.iw[2] ,
    \top_I.branch[17].block[15].um_I.iw[1] ,
    \top_I.branch[17].block[15].um_I.clk ,
    \top_I.branch[17].block[14].um_I.iw[17] ,
    \top_I.branch[17].block[14].um_I.iw[16] ,
    \top_I.branch[17].block[14].um_I.iw[15] ,
    \top_I.branch[17].block[14].um_I.iw[14] ,
    \top_I.branch[17].block[14].um_I.iw[13] ,
    \top_I.branch[17].block[14].um_I.iw[12] ,
    \top_I.branch[17].block[14].um_I.iw[11] ,
    \top_I.branch[17].block[14].um_I.iw[10] ,
    \top_I.branch[17].block[14].um_I.iw[9] ,
    \top_I.branch[17].block[14].um_I.iw[8] ,
    \top_I.branch[17].block[14].um_I.iw[7] ,
    \top_I.branch[17].block[14].um_I.iw[6] ,
    \top_I.branch[17].block[14].um_I.iw[5] ,
    \top_I.branch[17].block[14].um_I.iw[4] ,
    \top_I.branch[17].block[14].um_I.iw[3] ,
    \top_I.branch[17].block[14].um_I.iw[2] ,
    \top_I.branch[17].block[14].um_I.iw[1] ,
    \top_I.branch[17].block[14].um_I.clk ,
    \top_I.branch[17].block[13].um_I.iw[17] ,
    \top_I.branch[17].block[13].um_I.iw[16] ,
    \top_I.branch[17].block[13].um_I.iw[15] ,
    \top_I.branch[17].block[13].um_I.iw[14] ,
    \top_I.branch[17].block[13].um_I.iw[13] ,
    \top_I.branch[17].block[13].um_I.iw[12] ,
    \top_I.branch[17].block[13].um_I.iw[11] ,
    \top_I.branch[17].block[13].um_I.iw[10] ,
    \top_I.branch[17].block[13].um_I.iw[9] ,
    \top_I.branch[17].block[13].um_I.iw[8] ,
    \top_I.branch[17].block[13].um_I.iw[7] ,
    \top_I.branch[17].block[13].um_I.iw[6] ,
    \top_I.branch[17].block[13].um_I.iw[5] ,
    \top_I.branch[17].block[13].um_I.iw[4] ,
    \top_I.branch[17].block[13].um_I.iw[3] ,
    \top_I.branch[17].block[13].um_I.iw[2] ,
    \top_I.branch[17].block[13].um_I.iw[1] ,
    \top_I.branch[17].block[13].um_I.clk ,
    \top_I.branch[17].block[12].um_I.iw[17] ,
    \top_I.branch[17].block[12].um_I.iw[16] ,
    \top_I.branch[17].block[12].um_I.iw[15] ,
    \top_I.branch[17].block[12].um_I.iw[14] ,
    \top_I.branch[17].block[12].um_I.iw[13] ,
    \top_I.branch[17].block[12].um_I.iw[12] ,
    \top_I.branch[17].block[12].um_I.iw[11] ,
    \top_I.branch[17].block[12].um_I.iw[10] ,
    \top_I.branch[17].block[12].um_I.iw[9] ,
    \top_I.branch[17].block[12].um_I.iw[8] ,
    \top_I.branch[17].block[12].um_I.iw[7] ,
    \top_I.branch[17].block[12].um_I.iw[6] ,
    \top_I.branch[17].block[12].um_I.iw[5] ,
    \top_I.branch[17].block[12].um_I.iw[4] ,
    \top_I.branch[17].block[12].um_I.iw[3] ,
    \top_I.branch[17].block[12].um_I.iw[2] ,
    \top_I.branch[17].block[12].um_I.iw[1] ,
    \top_I.branch[17].block[12].um_I.clk ,
    \top_I.branch[17].block[11].um_I.iw[17] ,
    \top_I.branch[17].block[11].um_I.iw[16] ,
    \top_I.branch[17].block[11].um_I.iw[15] ,
    \top_I.branch[17].block[11].um_I.iw[14] ,
    \top_I.branch[17].block[11].um_I.iw[13] ,
    \top_I.branch[17].block[11].um_I.iw[12] ,
    \top_I.branch[17].block[11].um_I.iw[11] ,
    \top_I.branch[17].block[11].um_I.iw[10] ,
    \top_I.branch[17].block[11].um_I.iw[9] ,
    \top_I.branch[17].block[11].um_I.iw[8] ,
    \top_I.branch[17].block[11].um_I.iw[7] ,
    \top_I.branch[17].block[11].um_I.iw[6] ,
    \top_I.branch[17].block[11].um_I.iw[5] ,
    \top_I.branch[17].block[11].um_I.iw[4] ,
    \top_I.branch[17].block[11].um_I.iw[3] ,
    \top_I.branch[17].block[11].um_I.iw[2] ,
    \top_I.branch[17].block[11].um_I.iw[1] ,
    \top_I.branch[17].block[11].um_I.clk ,
    \top_I.branch[17].block[10].um_I.iw[17] ,
    \top_I.branch[17].block[10].um_I.iw[16] ,
    \top_I.branch[17].block[10].um_I.iw[15] ,
    \top_I.branch[17].block[10].um_I.iw[14] ,
    \top_I.branch[17].block[10].um_I.iw[13] ,
    \top_I.branch[17].block[10].um_I.iw[12] ,
    \top_I.branch[17].block[10].um_I.iw[11] ,
    \top_I.branch[17].block[10].um_I.iw[10] ,
    \top_I.branch[17].block[10].um_I.iw[9] ,
    \top_I.branch[17].block[10].um_I.iw[8] ,
    \top_I.branch[17].block[10].um_I.iw[7] ,
    \top_I.branch[17].block[10].um_I.iw[6] ,
    \top_I.branch[17].block[10].um_I.iw[5] ,
    \top_I.branch[17].block[10].um_I.iw[4] ,
    \top_I.branch[17].block[10].um_I.iw[3] ,
    \top_I.branch[17].block[10].um_I.iw[2] ,
    \top_I.branch[17].block[10].um_I.iw[1] ,
    \top_I.branch[17].block[10].um_I.clk ,
    \top_I.branch[17].block[9].um_I.iw[17] ,
    \top_I.branch[17].block[9].um_I.iw[16] ,
    \top_I.branch[17].block[9].um_I.iw[15] ,
    \top_I.branch[17].block[9].um_I.iw[14] ,
    \top_I.branch[17].block[9].um_I.iw[13] ,
    \top_I.branch[17].block[9].um_I.iw[12] ,
    \top_I.branch[17].block[9].um_I.iw[11] ,
    \top_I.branch[17].block[9].um_I.iw[10] ,
    \top_I.branch[17].block[9].um_I.iw[9] ,
    \top_I.branch[17].block[9].um_I.iw[8] ,
    \top_I.branch[17].block[9].um_I.iw[7] ,
    \top_I.branch[17].block[9].um_I.iw[6] ,
    \top_I.branch[17].block[9].um_I.iw[5] ,
    \top_I.branch[17].block[9].um_I.iw[4] ,
    \top_I.branch[17].block[9].um_I.iw[3] ,
    \top_I.branch[17].block[9].um_I.iw[2] ,
    \top_I.branch[17].block[9].um_I.iw[1] ,
    \top_I.branch[17].block[9].um_I.clk ,
    \top_I.branch[17].block[8].um_I.iw[17] ,
    \top_I.branch[17].block[8].um_I.iw[16] ,
    \top_I.branch[17].block[8].um_I.iw[15] ,
    \top_I.branch[17].block[8].um_I.iw[14] ,
    \top_I.branch[17].block[8].um_I.iw[13] ,
    \top_I.branch[17].block[8].um_I.iw[12] ,
    \top_I.branch[17].block[8].um_I.iw[11] ,
    \top_I.branch[17].block[8].um_I.iw[10] ,
    \top_I.branch[17].block[8].um_I.iw[9] ,
    \top_I.branch[17].block[8].um_I.iw[8] ,
    \top_I.branch[17].block[8].um_I.iw[7] ,
    \top_I.branch[17].block[8].um_I.iw[6] ,
    \top_I.branch[17].block[8].um_I.iw[5] ,
    \top_I.branch[17].block[8].um_I.iw[4] ,
    \top_I.branch[17].block[8].um_I.iw[3] ,
    \top_I.branch[17].block[8].um_I.iw[2] ,
    \top_I.branch[17].block[8].um_I.iw[1] ,
    \top_I.branch[17].block[8].um_I.clk ,
    \top_I.branch[17].block[7].um_I.iw[17] ,
    \top_I.branch[17].block[7].um_I.iw[16] ,
    \top_I.branch[17].block[7].um_I.iw[15] ,
    \top_I.branch[17].block[7].um_I.iw[14] ,
    \top_I.branch[17].block[7].um_I.iw[13] ,
    \top_I.branch[17].block[7].um_I.iw[12] ,
    \top_I.branch[17].block[7].um_I.iw[11] ,
    \top_I.branch[17].block[7].um_I.iw[10] ,
    \top_I.branch[17].block[7].um_I.iw[9] ,
    \top_I.branch[17].block[7].um_I.iw[8] ,
    \top_I.branch[17].block[7].um_I.iw[7] ,
    \top_I.branch[17].block[7].um_I.iw[6] ,
    \top_I.branch[17].block[7].um_I.iw[5] ,
    \top_I.branch[17].block[7].um_I.iw[4] ,
    \top_I.branch[17].block[7].um_I.iw[3] ,
    \top_I.branch[17].block[7].um_I.iw[2] ,
    \top_I.branch[17].block[7].um_I.iw[1] ,
    \top_I.branch[17].block[7].um_I.clk ,
    \top_I.branch[17].block[6].um_I.iw[17] ,
    \top_I.branch[17].block[6].um_I.iw[16] ,
    \top_I.branch[17].block[6].um_I.iw[15] ,
    \top_I.branch[17].block[6].um_I.iw[14] ,
    \top_I.branch[17].block[6].um_I.iw[13] ,
    \top_I.branch[17].block[6].um_I.iw[12] ,
    \top_I.branch[17].block[6].um_I.iw[11] ,
    \top_I.branch[17].block[6].um_I.iw[10] ,
    \top_I.branch[17].block[6].um_I.iw[9] ,
    \top_I.branch[17].block[6].um_I.iw[8] ,
    \top_I.branch[17].block[6].um_I.iw[7] ,
    \top_I.branch[17].block[6].um_I.iw[6] ,
    \top_I.branch[17].block[6].um_I.iw[5] ,
    \top_I.branch[17].block[6].um_I.iw[4] ,
    \top_I.branch[17].block[6].um_I.iw[3] ,
    \top_I.branch[17].block[6].um_I.iw[2] ,
    \top_I.branch[17].block[6].um_I.iw[1] ,
    \top_I.branch[17].block[6].um_I.clk ,
    \top_I.branch[17].block[5].um_I.iw[17] ,
    \top_I.branch[17].block[5].um_I.iw[16] ,
    \top_I.branch[17].block[5].um_I.iw[15] ,
    \top_I.branch[17].block[5].um_I.iw[14] ,
    \top_I.branch[17].block[5].um_I.iw[13] ,
    \top_I.branch[17].block[5].um_I.iw[12] ,
    \top_I.branch[17].block[5].um_I.iw[11] ,
    \top_I.branch[17].block[5].um_I.iw[10] ,
    \top_I.branch[17].block[5].um_I.iw[9] ,
    \top_I.branch[17].block[5].um_I.iw[8] ,
    \top_I.branch[17].block[5].um_I.iw[7] ,
    \top_I.branch[17].block[5].um_I.iw[6] ,
    \top_I.branch[17].block[5].um_I.iw[5] ,
    \top_I.branch[17].block[5].um_I.iw[4] ,
    \top_I.branch[17].block[5].um_I.iw[3] ,
    \top_I.branch[17].block[5].um_I.iw[2] ,
    \top_I.branch[17].block[5].um_I.iw[1] ,
    \top_I.branch[17].block[5].um_I.clk ,
    \top_I.branch[17].block[4].um_I.iw[17] ,
    \top_I.branch[17].block[4].um_I.iw[16] ,
    \top_I.branch[17].block[4].um_I.iw[15] ,
    \top_I.branch[17].block[4].um_I.iw[14] ,
    \top_I.branch[17].block[4].um_I.iw[13] ,
    \top_I.branch[17].block[4].um_I.iw[12] ,
    \top_I.branch[17].block[4].um_I.iw[11] ,
    \top_I.branch[17].block[4].um_I.iw[10] ,
    \top_I.branch[17].block[4].um_I.iw[9] ,
    \top_I.branch[17].block[4].um_I.iw[8] ,
    \top_I.branch[17].block[4].um_I.iw[7] ,
    \top_I.branch[17].block[4].um_I.iw[6] ,
    \top_I.branch[17].block[4].um_I.iw[5] ,
    \top_I.branch[17].block[4].um_I.iw[4] ,
    \top_I.branch[17].block[4].um_I.iw[3] ,
    \top_I.branch[17].block[4].um_I.iw[2] ,
    \top_I.branch[17].block[4].um_I.iw[1] ,
    \top_I.branch[17].block[4].um_I.clk ,
    \top_I.branch[17].block[3].um_I.iw[17] ,
    \top_I.branch[17].block[3].um_I.iw[16] ,
    \top_I.branch[17].block[3].um_I.iw[15] ,
    \top_I.branch[17].block[3].um_I.iw[14] ,
    \top_I.branch[17].block[3].um_I.iw[13] ,
    \top_I.branch[17].block[3].um_I.iw[12] ,
    \top_I.branch[17].block[3].um_I.iw[11] ,
    \top_I.branch[17].block[3].um_I.iw[10] ,
    \top_I.branch[17].block[3].um_I.iw[9] ,
    \top_I.branch[17].block[3].um_I.iw[8] ,
    \top_I.branch[17].block[3].um_I.iw[7] ,
    \top_I.branch[17].block[3].um_I.iw[6] ,
    \top_I.branch[17].block[3].um_I.iw[5] ,
    \top_I.branch[17].block[3].um_I.iw[4] ,
    \top_I.branch[17].block[3].um_I.iw[3] ,
    \top_I.branch[17].block[3].um_I.iw[2] ,
    \top_I.branch[17].block[3].um_I.iw[1] ,
    \top_I.branch[17].block[3].um_I.clk ,
    \top_I.branch[17].block[2].um_I.iw[17] ,
    \top_I.branch[17].block[2].um_I.iw[16] ,
    \top_I.branch[17].block[2].um_I.iw[15] ,
    \top_I.branch[17].block[2].um_I.iw[14] ,
    \top_I.branch[17].block[2].um_I.iw[13] ,
    \top_I.branch[17].block[2].um_I.iw[12] ,
    \top_I.branch[17].block[2].um_I.iw[11] ,
    \top_I.branch[17].block[2].um_I.iw[10] ,
    \top_I.branch[17].block[2].um_I.iw[9] ,
    \top_I.branch[17].block[2].um_I.iw[8] ,
    \top_I.branch[17].block[2].um_I.iw[7] ,
    \top_I.branch[17].block[2].um_I.iw[6] ,
    \top_I.branch[17].block[2].um_I.iw[5] ,
    \top_I.branch[17].block[2].um_I.iw[4] ,
    \top_I.branch[17].block[2].um_I.iw[3] ,
    \top_I.branch[17].block[2].um_I.iw[2] ,
    \top_I.branch[17].block[2].um_I.iw[1] ,
    \top_I.branch[17].block[2].um_I.clk ,
    \top_I.branch[17].block[1].um_I.iw[17] ,
    \top_I.branch[17].block[1].um_I.iw[16] ,
    \top_I.branch[17].block[1].um_I.iw[15] ,
    \top_I.branch[17].block[1].um_I.iw[14] ,
    \top_I.branch[17].block[1].um_I.iw[13] ,
    \top_I.branch[17].block[1].um_I.iw[12] ,
    \top_I.branch[17].block[1].um_I.iw[11] ,
    \top_I.branch[17].block[1].um_I.iw[10] ,
    \top_I.branch[17].block[1].um_I.iw[9] ,
    \top_I.branch[17].block[1].um_I.iw[8] ,
    \top_I.branch[17].block[1].um_I.iw[7] ,
    \top_I.branch[17].block[1].um_I.iw[6] ,
    \top_I.branch[17].block[1].um_I.iw[5] ,
    \top_I.branch[17].block[1].um_I.iw[4] ,
    \top_I.branch[17].block[1].um_I.iw[3] ,
    \top_I.branch[17].block[1].um_I.iw[2] ,
    \top_I.branch[17].block[1].um_I.iw[1] ,
    \top_I.branch[17].block[1].um_I.clk ,
    \top_I.branch[17].block[0].um_I.iw[17] ,
    \top_I.branch[17].block[0].um_I.iw[16] ,
    \top_I.branch[17].block[0].um_I.iw[15] ,
    \top_I.branch[17].block[0].um_I.iw[14] ,
    \top_I.branch[17].block[0].um_I.iw[13] ,
    \top_I.branch[17].block[0].um_I.iw[12] ,
    \top_I.branch[17].block[0].um_I.iw[11] ,
    \top_I.branch[17].block[0].um_I.iw[10] ,
    \top_I.branch[17].block[0].um_I.iw[9] ,
    \top_I.branch[17].block[0].um_I.iw[8] ,
    \top_I.branch[17].block[0].um_I.iw[7] ,
    \top_I.branch[17].block[0].um_I.iw[6] ,
    \top_I.branch[17].block[0].um_I.iw[5] ,
    \top_I.branch[17].block[0].um_I.iw[4] ,
    \top_I.branch[17].block[0].um_I.iw[3] ,
    \top_I.branch[17].block[0].um_I.iw[2] ,
    \top_I.branch[17].block[0].um_I.iw[1] ,
    \top_I.branch[17].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[17].block[15].um_I.pg_vdd ,
    \top_I.branch[17].block[14].um_I.pg_vdd ,
    \top_I.branch[17].block[13].um_I.pg_vdd ,
    \top_I.branch[17].block[12].um_I.pg_vdd ,
    \top_I.branch[17].block[11].um_I.pg_vdd ,
    \top_I.branch[17].block[10].um_I.pg_vdd ,
    \top_I.branch[17].block[9].um_I.pg_vdd ,
    \top_I.branch[17].block[8].um_I.pg_vdd ,
    \top_I.branch[17].block[7].um_I.pg_vdd ,
    \top_I.branch[17].block[6].um_I.pg_vdd ,
    \top_I.branch[17].block[5].um_I.pg_vdd ,
    \top_I.branch[17].block[4].um_I.pg_vdd ,
    \top_I.branch[17].block[3].um_I.pg_vdd ,
    \top_I.branch[17].block[2].um_I.pg_vdd ,
    \top_I.branch[17].block[1].um_I.pg_vdd ,
    \top_I.branch[17].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[18].mux_I  (.k_one(\top_I.branch[18].l_addr[0] ),
    .k_zero(\top_I.branch[18].l_addr[1] ),
    .addr({\top_I.branch[18].l_addr[0] ,
    \top_I.branch[18].l_addr[1] ,
    \top_I.branch[18].l_addr[1] ,
    \top_I.branch[18].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[18].block[15].um_I.ena ,
    \top_I.branch[18].block[14].um_I.ena ,
    \top_I.branch[18].block[13].um_I.ena ,
    \top_I.branch[18].block[12].um_I.ena ,
    \top_I.branch[18].block[11].um_I.ena ,
    \top_I.branch[18].block[10].um_I.ena ,
    \top_I.branch[18].block[9].um_I.ena ,
    \top_I.branch[18].block[8].um_I.ena ,
    \top_I.branch[18].block[7].um_I.ena ,
    \top_I.branch[18].block[6].um_I.ena ,
    \top_I.branch[18].block[5].um_I.ena ,
    \top_I.branch[18].block[4].um_I.ena ,
    \top_I.branch[18].block[3].um_I.ena ,
    \top_I.branch[18].block[2].um_I.ena ,
    \top_I.branch[18].block[1].um_I.ena ,
    \top_I.branch[18].block[0].um_I.ena }),
    .um_iw({\top_I.branch[18].block[15].um_I.iw[17] ,
    \top_I.branch[18].block[15].um_I.iw[16] ,
    \top_I.branch[18].block[15].um_I.iw[15] ,
    \top_I.branch[18].block[15].um_I.iw[14] ,
    \top_I.branch[18].block[15].um_I.iw[13] ,
    \top_I.branch[18].block[15].um_I.iw[12] ,
    \top_I.branch[18].block[15].um_I.iw[11] ,
    \top_I.branch[18].block[15].um_I.iw[10] ,
    \top_I.branch[18].block[15].um_I.iw[9] ,
    \top_I.branch[18].block[15].um_I.iw[8] ,
    \top_I.branch[18].block[15].um_I.iw[7] ,
    \top_I.branch[18].block[15].um_I.iw[6] ,
    \top_I.branch[18].block[15].um_I.iw[5] ,
    \top_I.branch[18].block[15].um_I.iw[4] ,
    \top_I.branch[18].block[15].um_I.iw[3] ,
    \top_I.branch[18].block[15].um_I.iw[2] ,
    \top_I.branch[18].block[15].um_I.iw[1] ,
    \top_I.branch[18].block[15].um_I.clk ,
    \top_I.branch[18].block[14].um_I.iw[17] ,
    \top_I.branch[18].block[14].um_I.iw[16] ,
    \top_I.branch[18].block[14].um_I.iw[15] ,
    \top_I.branch[18].block[14].um_I.iw[14] ,
    \top_I.branch[18].block[14].um_I.iw[13] ,
    \top_I.branch[18].block[14].um_I.iw[12] ,
    \top_I.branch[18].block[14].um_I.iw[11] ,
    \top_I.branch[18].block[14].um_I.iw[10] ,
    \top_I.branch[18].block[14].um_I.iw[9] ,
    \top_I.branch[18].block[14].um_I.iw[8] ,
    \top_I.branch[18].block[14].um_I.iw[7] ,
    \top_I.branch[18].block[14].um_I.iw[6] ,
    \top_I.branch[18].block[14].um_I.iw[5] ,
    \top_I.branch[18].block[14].um_I.iw[4] ,
    \top_I.branch[18].block[14].um_I.iw[3] ,
    \top_I.branch[18].block[14].um_I.iw[2] ,
    \top_I.branch[18].block[14].um_I.iw[1] ,
    \top_I.branch[18].block[14].um_I.clk ,
    \top_I.branch[18].block[13].um_I.iw[17] ,
    \top_I.branch[18].block[13].um_I.iw[16] ,
    \top_I.branch[18].block[13].um_I.iw[15] ,
    \top_I.branch[18].block[13].um_I.iw[14] ,
    \top_I.branch[18].block[13].um_I.iw[13] ,
    \top_I.branch[18].block[13].um_I.iw[12] ,
    \top_I.branch[18].block[13].um_I.iw[11] ,
    \top_I.branch[18].block[13].um_I.iw[10] ,
    \top_I.branch[18].block[13].um_I.iw[9] ,
    \top_I.branch[18].block[13].um_I.iw[8] ,
    \top_I.branch[18].block[13].um_I.iw[7] ,
    \top_I.branch[18].block[13].um_I.iw[6] ,
    \top_I.branch[18].block[13].um_I.iw[5] ,
    \top_I.branch[18].block[13].um_I.iw[4] ,
    \top_I.branch[18].block[13].um_I.iw[3] ,
    \top_I.branch[18].block[13].um_I.iw[2] ,
    \top_I.branch[18].block[13].um_I.iw[1] ,
    \top_I.branch[18].block[13].um_I.clk ,
    \top_I.branch[18].block[12].um_I.iw[17] ,
    \top_I.branch[18].block[12].um_I.iw[16] ,
    \top_I.branch[18].block[12].um_I.iw[15] ,
    \top_I.branch[18].block[12].um_I.iw[14] ,
    \top_I.branch[18].block[12].um_I.iw[13] ,
    \top_I.branch[18].block[12].um_I.iw[12] ,
    \top_I.branch[18].block[12].um_I.iw[11] ,
    \top_I.branch[18].block[12].um_I.iw[10] ,
    \top_I.branch[18].block[12].um_I.iw[9] ,
    \top_I.branch[18].block[12].um_I.iw[8] ,
    \top_I.branch[18].block[12].um_I.iw[7] ,
    \top_I.branch[18].block[12].um_I.iw[6] ,
    \top_I.branch[18].block[12].um_I.iw[5] ,
    \top_I.branch[18].block[12].um_I.iw[4] ,
    \top_I.branch[18].block[12].um_I.iw[3] ,
    \top_I.branch[18].block[12].um_I.iw[2] ,
    \top_I.branch[18].block[12].um_I.iw[1] ,
    \top_I.branch[18].block[12].um_I.clk ,
    \top_I.branch[18].block[11].um_I.iw[17] ,
    \top_I.branch[18].block[11].um_I.iw[16] ,
    \top_I.branch[18].block[11].um_I.iw[15] ,
    \top_I.branch[18].block[11].um_I.iw[14] ,
    \top_I.branch[18].block[11].um_I.iw[13] ,
    \top_I.branch[18].block[11].um_I.iw[12] ,
    \top_I.branch[18].block[11].um_I.iw[11] ,
    \top_I.branch[18].block[11].um_I.iw[10] ,
    \top_I.branch[18].block[11].um_I.iw[9] ,
    \top_I.branch[18].block[11].um_I.iw[8] ,
    \top_I.branch[18].block[11].um_I.iw[7] ,
    \top_I.branch[18].block[11].um_I.iw[6] ,
    \top_I.branch[18].block[11].um_I.iw[5] ,
    \top_I.branch[18].block[11].um_I.iw[4] ,
    \top_I.branch[18].block[11].um_I.iw[3] ,
    \top_I.branch[18].block[11].um_I.iw[2] ,
    \top_I.branch[18].block[11].um_I.iw[1] ,
    \top_I.branch[18].block[11].um_I.clk ,
    \top_I.branch[18].block[10].um_I.iw[17] ,
    \top_I.branch[18].block[10].um_I.iw[16] ,
    \top_I.branch[18].block[10].um_I.iw[15] ,
    \top_I.branch[18].block[10].um_I.iw[14] ,
    \top_I.branch[18].block[10].um_I.iw[13] ,
    \top_I.branch[18].block[10].um_I.iw[12] ,
    \top_I.branch[18].block[10].um_I.iw[11] ,
    \top_I.branch[18].block[10].um_I.iw[10] ,
    \top_I.branch[18].block[10].um_I.iw[9] ,
    \top_I.branch[18].block[10].um_I.iw[8] ,
    \top_I.branch[18].block[10].um_I.iw[7] ,
    \top_I.branch[18].block[10].um_I.iw[6] ,
    \top_I.branch[18].block[10].um_I.iw[5] ,
    \top_I.branch[18].block[10].um_I.iw[4] ,
    \top_I.branch[18].block[10].um_I.iw[3] ,
    \top_I.branch[18].block[10].um_I.iw[2] ,
    \top_I.branch[18].block[10].um_I.iw[1] ,
    \top_I.branch[18].block[10].um_I.clk ,
    \top_I.branch[18].block[9].um_I.iw[17] ,
    \top_I.branch[18].block[9].um_I.iw[16] ,
    \top_I.branch[18].block[9].um_I.iw[15] ,
    \top_I.branch[18].block[9].um_I.iw[14] ,
    \top_I.branch[18].block[9].um_I.iw[13] ,
    \top_I.branch[18].block[9].um_I.iw[12] ,
    \top_I.branch[18].block[9].um_I.iw[11] ,
    \top_I.branch[18].block[9].um_I.iw[10] ,
    \top_I.branch[18].block[9].um_I.iw[9] ,
    \top_I.branch[18].block[9].um_I.iw[8] ,
    \top_I.branch[18].block[9].um_I.iw[7] ,
    \top_I.branch[18].block[9].um_I.iw[6] ,
    \top_I.branch[18].block[9].um_I.iw[5] ,
    \top_I.branch[18].block[9].um_I.iw[4] ,
    \top_I.branch[18].block[9].um_I.iw[3] ,
    \top_I.branch[18].block[9].um_I.iw[2] ,
    \top_I.branch[18].block[9].um_I.iw[1] ,
    \top_I.branch[18].block[9].um_I.clk ,
    \top_I.branch[18].block[8].um_I.iw[17] ,
    \top_I.branch[18].block[8].um_I.iw[16] ,
    \top_I.branch[18].block[8].um_I.iw[15] ,
    \top_I.branch[18].block[8].um_I.iw[14] ,
    \top_I.branch[18].block[8].um_I.iw[13] ,
    \top_I.branch[18].block[8].um_I.iw[12] ,
    \top_I.branch[18].block[8].um_I.iw[11] ,
    \top_I.branch[18].block[8].um_I.iw[10] ,
    \top_I.branch[18].block[8].um_I.iw[9] ,
    \top_I.branch[18].block[8].um_I.iw[8] ,
    \top_I.branch[18].block[8].um_I.iw[7] ,
    \top_I.branch[18].block[8].um_I.iw[6] ,
    \top_I.branch[18].block[8].um_I.iw[5] ,
    \top_I.branch[18].block[8].um_I.iw[4] ,
    \top_I.branch[18].block[8].um_I.iw[3] ,
    \top_I.branch[18].block[8].um_I.iw[2] ,
    \top_I.branch[18].block[8].um_I.iw[1] ,
    \top_I.branch[18].block[8].um_I.clk ,
    \top_I.branch[18].block[7].um_I.iw[17] ,
    \top_I.branch[18].block[7].um_I.iw[16] ,
    \top_I.branch[18].block[7].um_I.iw[15] ,
    \top_I.branch[18].block[7].um_I.iw[14] ,
    \top_I.branch[18].block[7].um_I.iw[13] ,
    \top_I.branch[18].block[7].um_I.iw[12] ,
    \top_I.branch[18].block[7].um_I.iw[11] ,
    \top_I.branch[18].block[7].um_I.iw[10] ,
    \top_I.branch[18].block[7].um_I.iw[9] ,
    \top_I.branch[18].block[7].um_I.iw[8] ,
    \top_I.branch[18].block[7].um_I.iw[7] ,
    \top_I.branch[18].block[7].um_I.iw[6] ,
    \top_I.branch[18].block[7].um_I.iw[5] ,
    \top_I.branch[18].block[7].um_I.iw[4] ,
    \top_I.branch[18].block[7].um_I.iw[3] ,
    \top_I.branch[18].block[7].um_I.iw[2] ,
    \top_I.branch[18].block[7].um_I.iw[1] ,
    \top_I.branch[18].block[7].um_I.clk ,
    \top_I.branch[18].block[6].um_I.iw[17] ,
    \top_I.branch[18].block[6].um_I.iw[16] ,
    \top_I.branch[18].block[6].um_I.iw[15] ,
    \top_I.branch[18].block[6].um_I.iw[14] ,
    \top_I.branch[18].block[6].um_I.iw[13] ,
    \top_I.branch[18].block[6].um_I.iw[12] ,
    \top_I.branch[18].block[6].um_I.iw[11] ,
    \top_I.branch[18].block[6].um_I.iw[10] ,
    \top_I.branch[18].block[6].um_I.iw[9] ,
    \top_I.branch[18].block[6].um_I.iw[8] ,
    \top_I.branch[18].block[6].um_I.iw[7] ,
    \top_I.branch[18].block[6].um_I.iw[6] ,
    \top_I.branch[18].block[6].um_I.iw[5] ,
    \top_I.branch[18].block[6].um_I.iw[4] ,
    \top_I.branch[18].block[6].um_I.iw[3] ,
    \top_I.branch[18].block[6].um_I.iw[2] ,
    \top_I.branch[18].block[6].um_I.iw[1] ,
    \top_I.branch[18].block[6].um_I.clk ,
    \top_I.branch[18].block[5].um_I.iw[17] ,
    \top_I.branch[18].block[5].um_I.iw[16] ,
    \top_I.branch[18].block[5].um_I.iw[15] ,
    \top_I.branch[18].block[5].um_I.iw[14] ,
    \top_I.branch[18].block[5].um_I.iw[13] ,
    \top_I.branch[18].block[5].um_I.iw[12] ,
    \top_I.branch[18].block[5].um_I.iw[11] ,
    \top_I.branch[18].block[5].um_I.iw[10] ,
    \top_I.branch[18].block[5].um_I.iw[9] ,
    \top_I.branch[18].block[5].um_I.iw[8] ,
    \top_I.branch[18].block[5].um_I.iw[7] ,
    \top_I.branch[18].block[5].um_I.iw[6] ,
    \top_I.branch[18].block[5].um_I.iw[5] ,
    \top_I.branch[18].block[5].um_I.iw[4] ,
    \top_I.branch[18].block[5].um_I.iw[3] ,
    \top_I.branch[18].block[5].um_I.iw[2] ,
    \top_I.branch[18].block[5].um_I.iw[1] ,
    \top_I.branch[18].block[5].um_I.clk ,
    \top_I.branch[18].block[4].um_I.iw[17] ,
    \top_I.branch[18].block[4].um_I.iw[16] ,
    \top_I.branch[18].block[4].um_I.iw[15] ,
    \top_I.branch[18].block[4].um_I.iw[14] ,
    \top_I.branch[18].block[4].um_I.iw[13] ,
    \top_I.branch[18].block[4].um_I.iw[12] ,
    \top_I.branch[18].block[4].um_I.iw[11] ,
    \top_I.branch[18].block[4].um_I.iw[10] ,
    \top_I.branch[18].block[4].um_I.iw[9] ,
    \top_I.branch[18].block[4].um_I.iw[8] ,
    \top_I.branch[18].block[4].um_I.iw[7] ,
    \top_I.branch[18].block[4].um_I.iw[6] ,
    \top_I.branch[18].block[4].um_I.iw[5] ,
    \top_I.branch[18].block[4].um_I.iw[4] ,
    \top_I.branch[18].block[4].um_I.iw[3] ,
    \top_I.branch[18].block[4].um_I.iw[2] ,
    \top_I.branch[18].block[4].um_I.iw[1] ,
    \top_I.branch[18].block[4].um_I.clk ,
    \top_I.branch[18].block[3].um_I.iw[17] ,
    \top_I.branch[18].block[3].um_I.iw[16] ,
    \top_I.branch[18].block[3].um_I.iw[15] ,
    \top_I.branch[18].block[3].um_I.iw[14] ,
    \top_I.branch[18].block[3].um_I.iw[13] ,
    \top_I.branch[18].block[3].um_I.iw[12] ,
    \top_I.branch[18].block[3].um_I.iw[11] ,
    \top_I.branch[18].block[3].um_I.iw[10] ,
    \top_I.branch[18].block[3].um_I.iw[9] ,
    \top_I.branch[18].block[3].um_I.iw[8] ,
    \top_I.branch[18].block[3].um_I.iw[7] ,
    \top_I.branch[18].block[3].um_I.iw[6] ,
    \top_I.branch[18].block[3].um_I.iw[5] ,
    \top_I.branch[18].block[3].um_I.iw[4] ,
    \top_I.branch[18].block[3].um_I.iw[3] ,
    \top_I.branch[18].block[3].um_I.iw[2] ,
    \top_I.branch[18].block[3].um_I.iw[1] ,
    \top_I.branch[18].block[3].um_I.clk ,
    \top_I.branch[18].block[2].um_I.iw[17] ,
    \top_I.branch[18].block[2].um_I.iw[16] ,
    \top_I.branch[18].block[2].um_I.iw[15] ,
    \top_I.branch[18].block[2].um_I.iw[14] ,
    \top_I.branch[18].block[2].um_I.iw[13] ,
    \top_I.branch[18].block[2].um_I.iw[12] ,
    \top_I.branch[18].block[2].um_I.iw[11] ,
    \top_I.branch[18].block[2].um_I.iw[10] ,
    \top_I.branch[18].block[2].um_I.iw[9] ,
    \top_I.branch[18].block[2].um_I.iw[8] ,
    \top_I.branch[18].block[2].um_I.iw[7] ,
    \top_I.branch[18].block[2].um_I.iw[6] ,
    \top_I.branch[18].block[2].um_I.iw[5] ,
    \top_I.branch[18].block[2].um_I.iw[4] ,
    \top_I.branch[18].block[2].um_I.iw[3] ,
    \top_I.branch[18].block[2].um_I.iw[2] ,
    \top_I.branch[18].block[2].um_I.iw[1] ,
    \top_I.branch[18].block[2].um_I.clk ,
    \top_I.branch[18].block[1].um_I.iw[17] ,
    \top_I.branch[18].block[1].um_I.iw[16] ,
    \top_I.branch[18].block[1].um_I.iw[15] ,
    \top_I.branch[18].block[1].um_I.iw[14] ,
    \top_I.branch[18].block[1].um_I.iw[13] ,
    \top_I.branch[18].block[1].um_I.iw[12] ,
    \top_I.branch[18].block[1].um_I.iw[11] ,
    \top_I.branch[18].block[1].um_I.iw[10] ,
    \top_I.branch[18].block[1].um_I.iw[9] ,
    \top_I.branch[18].block[1].um_I.iw[8] ,
    \top_I.branch[18].block[1].um_I.iw[7] ,
    \top_I.branch[18].block[1].um_I.iw[6] ,
    \top_I.branch[18].block[1].um_I.iw[5] ,
    \top_I.branch[18].block[1].um_I.iw[4] ,
    \top_I.branch[18].block[1].um_I.iw[3] ,
    \top_I.branch[18].block[1].um_I.iw[2] ,
    \top_I.branch[18].block[1].um_I.iw[1] ,
    \top_I.branch[18].block[1].um_I.clk ,
    \top_I.branch[18].block[0].um_I.iw[17] ,
    \top_I.branch[18].block[0].um_I.iw[16] ,
    \top_I.branch[18].block[0].um_I.iw[15] ,
    \top_I.branch[18].block[0].um_I.iw[14] ,
    \top_I.branch[18].block[0].um_I.iw[13] ,
    \top_I.branch[18].block[0].um_I.iw[12] ,
    \top_I.branch[18].block[0].um_I.iw[11] ,
    \top_I.branch[18].block[0].um_I.iw[10] ,
    \top_I.branch[18].block[0].um_I.iw[9] ,
    \top_I.branch[18].block[0].um_I.iw[8] ,
    \top_I.branch[18].block[0].um_I.iw[7] ,
    \top_I.branch[18].block[0].um_I.iw[6] ,
    \top_I.branch[18].block[0].um_I.iw[5] ,
    \top_I.branch[18].block[0].um_I.iw[4] ,
    \top_I.branch[18].block[0].um_I.iw[3] ,
    \top_I.branch[18].block[0].um_I.iw[2] ,
    \top_I.branch[18].block[0].um_I.iw[1] ,
    \top_I.branch[18].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[18].block[15].um_I.pg_vdd ,
    \top_I.branch[18].block[14].um_I.pg_vdd ,
    \top_I.branch[18].block[13].um_I.pg_vdd ,
    \top_I.branch[18].block[12].um_I.pg_vdd ,
    \top_I.branch[18].block[11].um_I.pg_vdd ,
    \top_I.branch[18].block[10].um_I.pg_vdd ,
    \top_I.branch[18].block[9].um_I.pg_vdd ,
    \top_I.branch[18].block[8].um_I.pg_vdd ,
    \top_I.branch[18].block[7].um_I.pg_vdd ,
    \top_I.branch[18].block[6].um_I.pg_vdd ,
    \top_I.branch[18].block[5].um_I.pg_vdd ,
    \top_I.branch[18].block[4].um_I.pg_vdd ,
    \top_I.branch[18].block[3].um_I.pg_vdd ,
    \top_I.branch[18].block[2].um_I.pg_vdd ,
    \top_I.branch[18].block[1].um_I.pg_vdd ,
    \top_I.branch[18].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[19].mux_I  (.k_one(\top_I.branch[19].l_addr[0] ),
    .k_zero(\top_I.branch[19].l_addr[1] ),
    .addr({\top_I.branch[19].l_addr[0] ,
    \top_I.branch[19].l_addr[1] ,
    \top_I.branch[19].l_addr[1] ,
    \top_I.branch[19].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[19].block[15].um_I.ena ,
    \top_I.branch[19].block[14].um_I.ena ,
    \top_I.branch[19].block[13].um_I.ena ,
    \top_I.branch[19].block[12].um_I.ena ,
    \top_I.branch[19].block[11].um_I.ena ,
    \top_I.branch[19].block[10].um_I.ena ,
    \top_I.branch[19].block[9].um_I.ena ,
    \top_I.branch[19].block[8].um_I.ena ,
    \top_I.branch[19].block[7].um_I.ena ,
    \top_I.branch[19].block[6].um_I.ena ,
    \top_I.branch[19].block[5].um_I.ena ,
    \top_I.branch[19].block[4].um_I.ena ,
    \top_I.branch[19].block[3].um_I.ena ,
    \top_I.branch[19].block[2].um_I.ena ,
    \top_I.branch[19].block[1].um_I.ena ,
    \top_I.branch[19].block[0].um_I.ena }),
    .um_iw({\top_I.branch[19].block[15].um_I.iw[17] ,
    \top_I.branch[19].block[15].um_I.iw[16] ,
    \top_I.branch[19].block[15].um_I.iw[15] ,
    \top_I.branch[19].block[15].um_I.iw[14] ,
    \top_I.branch[19].block[15].um_I.iw[13] ,
    \top_I.branch[19].block[15].um_I.iw[12] ,
    \top_I.branch[19].block[15].um_I.iw[11] ,
    \top_I.branch[19].block[15].um_I.iw[10] ,
    \top_I.branch[19].block[15].um_I.iw[9] ,
    \top_I.branch[19].block[15].um_I.iw[8] ,
    \top_I.branch[19].block[15].um_I.iw[7] ,
    \top_I.branch[19].block[15].um_I.iw[6] ,
    \top_I.branch[19].block[15].um_I.iw[5] ,
    \top_I.branch[19].block[15].um_I.iw[4] ,
    \top_I.branch[19].block[15].um_I.iw[3] ,
    \top_I.branch[19].block[15].um_I.iw[2] ,
    \top_I.branch[19].block[15].um_I.iw[1] ,
    \top_I.branch[19].block[15].um_I.clk ,
    \top_I.branch[19].block[14].um_I.iw[17] ,
    \top_I.branch[19].block[14].um_I.iw[16] ,
    \top_I.branch[19].block[14].um_I.iw[15] ,
    \top_I.branch[19].block[14].um_I.iw[14] ,
    \top_I.branch[19].block[14].um_I.iw[13] ,
    \top_I.branch[19].block[14].um_I.iw[12] ,
    \top_I.branch[19].block[14].um_I.iw[11] ,
    \top_I.branch[19].block[14].um_I.iw[10] ,
    \top_I.branch[19].block[14].um_I.iw[9] ,
    \top_I.branch[19].block[14].um_I.iw[8] ,
    \top_I.branch[19].block[14].um_I.iw[7] ,
    \top_I.branch[19].block[14].um_I.iw[6] ,
    \top_I.branch[19].block[14].um_I.iw[5] ,
    \top_I.branch[19].block[14].um_I.iw[4] ,
    \top_I.branch[19].block[14].um_I.iw[3] ,
    \top_I.branch[19].block[14].um_I.iw[2] ,
    \top_I.branch[19].block[14].um_I.iw[1] ,
    \top_I.branch[19].block[14].um_I.clk ,
    \top_I.branch[19].block[13].um_I.iw[17] ,
    \top_I.branch[19].block[13].um_I.iw[16] ,
    \top_I.branch[19].block[13].um_I.iw[15] ,
    \top_I.branch[19].block[13].um_I.iw[14] ,
    \top_I.branch[19].block[13].um_I.iw[13] ,
    \top_I.branch[19].block[13].um_I.iw[12] ,
    \top_I.branch[19].block[13].um_I.iw[11] ,
    \top_I.branch[19].block[13].um_I.iw[10] ,
    \top_I.branch[19].block[13].um_I.iw[9] ,
    \top_I.branch[19].block[13].um_I.iw[8] ,
    \top_I.branch[19].block[13].um_I.iw[7] ,
    \top_I.branch[19].block[13].um_I.iw[6] ,
    \top_I.branch[19].block[13].um_I.iw[5] ,
    \top_I.branch[19].block[13].um_I.iw[4] ,
    \top_I.branch[19].block[13].um_I.iw[3] ,
    \top_I.branch[19].block[13].um_I.iw[2] ,
    \top_I.branch[19].block[13].um_I.iw[1] ,
    \top_I.branch[19].block[13].um_I.clk ,
    \top_I.branch[19].block[12].um_I.iw[17] ,
    \top_I.branch[19].block[12].um_I.iw[16] ,
    \top_I.branch[19].block[12].um_I.iw[15] ,
    \top_I.branch[19].block[12].um_I.iw[14] ,
    \top_I.branch[19].block[12].um_I.iw[13] ,
    \top_I.branch[19].block[12].um_I.iw[12] ,
    \top_I.branch[19].block[12].um_I.iw[11] ,
    \top_I.branch[19].block[12].um_I.iw[10] ,
    \top_I.branch[19].block[12].um_I.iw[9] ,
    \top_I.branch[19].block[12].um_I.iw[8] ,
    \top_I.branch[19].block[12].um_I.iw[7] ,
    \top_I.branch[19].block[12].um_I.iw[6] ,
    \top_I.branch[19].block[12].um_I.iw[5] ,
    \top_I.branch[19].block[12].um_I.iw[4] ,
    \top_I.branch[19].block[12].um_I.iw[3] ,
    \top_I.branch[19].block[12].um_I.iw[2] ,
    \top_I.branch[19].block[12].um_I.iw[1] ,
    \top_I.branch[19].block[12].um_I.clk ,
    \top_I.branch[19].block[11].um_I.iw[17] ,
    \top_I.branch[19].block[11].um_I.iw[16] ,
    \top_I.branch[19].block[11].um_I.iw[15] ,
    \top_I.branch[19].block[11].um_I.iw[14] ,
    \top_I.branch[19].block[11].um_I.iw[13] ,
    \top_I.branch[19].block[11].um_I.iw[12] ,
    \top_I.branch[19].block[11].um_I.iw[11] ,
    \top_I.branch[19].block[11].um_I.iw[10] ,
    \top_I.branch[19].block[11].um_I.iw[9] ,
    \top_I.branch[19].block[11].um_I.iw[8] ,
    \top_I.branch[19].block[11].um_I.iw[7] ,
    \top_I.branch[19].block[11].um_I.iw[6] ,
    \top_I.branch[19].block[11].um_I.iw[5] ,
    \top_I.branch[19].block[11].um_I.iw[4] ,
    \top_I.branch[19].block[11].um_I.iw[3] ,
    \top_I.branch[19].block[11].um_I.iw[2] ,
    \top_I.branch[19].block[11].um_I.iw[1] ,
    \top_I.branch[19].block[11].um_I.clk ,
    \top_I.branch[19].block[10].um_I.iw[17] ,
    \top_I.branch[19].block[10].um_I.iw[16] ,
    \top_I.branch[19].block[10].um_I.iw[15] ,
    \top_I.branch[19].block[10].um_I.iw[14] ,
    \top_I.branch[19].block[10].um_I.iw[13] ,
    \top_I.branch[19].block[10].um_I.iw[12] ,
    \top_I.branch[19].block[10].um_I.iw[11] ,
    \top_I.branch[19].block[10].um_I.iw[10] ,
    \top_I.branch[19].block[10].um_I.iw[9] ,
    \top_I.branch[19].block[10].um_I.iw[8] ,
    \top_I.branch[19].block[10].um_I.iw[7] ,
    \top_I.branch[19].block[10].um_I.iw[6] ,
    \top_I.branch[19].block[10].um_I.iw[5] ,
    \top_I.branch[19].block[10].um_I.iw[4] ,
    \top_I.branch[19].block[10].um_I.iw[3] ,
    \top_I.branch[19].block[10].um_I.iw[2] ,
    \top_I.branch[19].block[10].um_I.iw[1] ,
    \top_I.branch[19].block[10].um_I.clk ,
    \top_I.branch[19].block[9].um_I.iw[17] ,
    \top_I.branch[19].block[9].um_I.iw[16] ,
    \top_I.branch[19].block[9].um_I.iw[15] ,
    \top_I.branch[19].block[9].um_I.iw[14] ,
    \top_I.branch[19].block[9].um_I.iw[13] ,
    \top_I.branch[19].block[9].um_I.iw[12] ,
    \top_I.branch[19].block[9].um_I.iw[11] ,
    \top_I.branch[19].block[9].um_I.iw[10] ,
    \top_I.branch[19].block[9].um_I.iw[9] ,
    \top_I.branch[19].block[9].um_I.iw[8] ,
    \top_I.branch[19].block[9].um_I.iw[7] ,
    \top_I.branch[19].block[9].um_I.iw[6] ,
    \top_I.branch[19].block[9].um_I.iw[5] ,
    \top_I.branch[19].block[9].um_I.iw[4] ,
    \top_I.branch[19].block[9].um_I.iw[3] ,
    \top_I.branch[19].block[9].um_I.iw[2] ,
    \top_I.branch[19].block[9].um_I.iw[1] ,
    \top_I.branch[19].block[9].um_I.clk ,
    \top_I.branch[19].block[8].um_I.iw[17] ,
    \top_I.branch[19].block[8].um_I.iw[16] ,
    \top_I.branch[19].block[8].um_I.iw[15] ,
    \top_I.branch[19].block[8].um_I.iw[14] ,
    \top_I.branch[19].block[8].um_I.iw[13] ,
    \top_I.branch[19].block[8].um_I.iw[12] ,
    \top_I.branch[19].block[8].um_I.iw[11] ,
    \top_I.branch[19].block[8].um_I.iw[10] ,
    \top_I.branch[19].block[8].um_I.iw[9] ,
    \top_I.branch[19].block[8].um_I.iw[8] ,
    \top_I.branch[19].block[8].um_I.iw[7] ,
    \top_I.branch[19].block[8].um_I.iw[6] ,
    \top_I.branch[19].block[8].um_I.iw[5] ,
    \top_I.branch[19].block[8].um_I.iw[4] ,
    \top_I.branch[19].block[8].um_I.iw[3] ,
    \top_I.branch[19].block[8].um_I.iw[2] ,
    \top_I.branch[19].block[8].um_I.iw[1] ,
    \top_I.branch[19].block[8].um_I.clk ,
    \top_I.branch[19].block[7].um_I.iw[17] ,
    \top_I.branch[19].block[7].um_I.iw[16] ,
    \top_I.branch[19].block[7].um_I.iw[15] ,
    \top_I.branch[19].block[7].um_I.iw[14] ,
    \top_I.branch[19].block[7].um_I.iw[13] ,
    \top_I.branch[19].block[7].um_I.iw[12] ,
    \top_I.branch[19].block[7].um_I.iw[11] ,
    \top_I.branch[19].block[7].um_I.iw[10] ,
    \top_I.branch[19].block[7].um_I.iw[9] ,
    \top_I.branch[19].block[7].um_I.iw[8] ,
    \top_I.branch[19].block[7].um_I.iw[7] ,
    \top_I.branch[19].block[7].um_I.iw[6] ,
    \top_I.branch[19].block[7].um_I.iw[5] ,
    \top_I.branch[19].block[7].um_I.iw[4] ,
    \top_I.branch[19].block[7].um_I.iw[3] ,
    \top_I.branch[19].block[7].um_I.iw[2] ,
    \top_I.branch[19].block[7].um_I.iw[1] ,
    \top_I.branch[19].block[7].um_I.clk ,
    \top_I.branch[19].block[6].um_I.iw[17] ,
    \top_I.branch[19].block[6].um_I.iw[16] ,
    \top_I.branch[19].block[6].um_I.iw[15] ,
    \top_I.branch[19].block[6].um_I.iw[14] ,
    \top_I.branch[19].block[6].um_I.iw[13] ,
    \top_I.branch[19].block[6].um_I.iw[12] ,
    \top_I.branch[19].block[6].um_I.iw[11] ,
    \top_I.branch[19].block[6].um_I.iw[10] ,
    \top_I.branch[19].block[6].um_I.iw[9] ,
    \top_I.branch[19].block[6].um_I.iw[8] ,
    \top_I.branch[19].block[6].um_I.iw[7] ,
    \top_I.branch[19].block[6].um_I.iw[6] ,
    \top_I.branch[19].block[6].um_I.iw[5] ,
    \top_I.branch[19].block[6].um_I.iw[4] ,
    \top_I.branch[19].block[6].um_I.iw[3] ,
    \top_I.branch[19].block[6].um_I.iw[2] ,
    \top_I.branch[19].block[6].um_I.iw[1] ,
    \top_I.branch[19].block[6].um_I.clk ,
    \top_I.branch[19].block[5].um_I.iw[17] ,
    \top_I.branch[19].block[5].um_I.iw[16] ,
    \top_I.branch[19].block[5].um_I.iw[15] ,
    \top_I.branch[19].block[5].um_I.iw[14] ,
    \top_I.branch[19].block[5].um_I.iw[13] ,
    \top_I.branch[19].block[5].um_I.iw[12] ,
    \top_I.branch[19].block[5].um_I.iw[11] ,
    \top_I.branch[19].block[5].um_I.iw[10] ,
    \top_I.branch[19].block[5].um_I.iw[9] ,
    \top_I.branch[19].block[5].um_I.iw[8] ,
    \top_I.branch[19].block[5].um_I.iw[7] ,
    \top_I.branch[19].block[5].um_I.iw[6] ,
    \top_I.branch[19].block[5].um_I.iw[5] ,
    \top_I.branch[19].block[5].um_I.iw[4] ,
    \top_I.branch[19].block[5].um_I.iw[3] ,
    \top_I.branch[19].block[5].um_I.iw[2] ,
    \top_I.branch[19].block[5].um_I.iw[1] ,
    \top_I.branch[19].block[5].um_I.clk ,
    \top_I.branch[19].block[4].um_I.iw[17] ,
    \top_I.branch[19].block[4].um_I.iw[16] ,
    \top_I.branch[19].block[4].um_I.iw[15] ,
    \top_I.branch[19].block[4].um_I.iw[14] ,
    \top_I.branch[19].block[4].um_I.iw[13] ,
    \top_I.branch[19].block[4].um_I.iw[12] ,
    \top_I.branch[19].block[4].um_I.iw[11] ,
    \top_I.branch[19].block[4].um_I.iw[10] ,
    \top_I.branch[19].block[4].um_I.iw[9] ,
    \top_I.branch[19].block[4].um_I.iw[8] ,
    \top_I.branch[19].block[4].um_I.iw[7] ,
    \top_I.branch[19].block[4].um_I.iw[6] ,
    \top_I.branch[19].block[4].um_I.iw[5] ,
    \top_I.branch[19].block[4].um_I.iw[4] ,
    \top_I.branch[19].block[4].um_I.iw[3] ,
    \top_I.branch[19].block[4].um_I.iw[2] ,
    \top_I.branch[19].block[4].um_I.iw[1] ,
    \top_I.branch[19].block[4].um_I.clk ,
    \top_I.branch[19].block[3].um_I.iw[17] ,
    \top_I.branch[19].block[3].um_I.iw[16] ,
    \top_I.branch[19].block[3].um_I.iw[15] ,
    \top_I.branch[19].block[3].um_I.iw[14] ,
    \top_I.branch[19].block[3].um_I.iw[13] ,
    \top_I.branch[19].block[3].um_I.iw[12] ,
    \top_I.branch[19].block[3].um_I.iw[11] ,
    \top_I.branch[19].block[3].um_I.iw[10] ,
    \top_I.branch[19].block[3].um_I.iw[9] ,
    \top_I.branch[19].block[3].um_I.iw[8] ,
    \top_I.branch[19].block[3].um_I.iw[7] ,
    \top_I.branch[19].block[3].um_I.iw[6] ,
    \top_I.branch[19].block[3].um_I.iw[5] ,
    \top_I.branch[19].block[3].um_I.iw[4] ,
    \top_I.branch[19].block[3].um_I.iw[3] ,
    \top_I.branch[19].block[3].um_I.iw[2] ,
    \top_I.branch[19].block[3].um_I.iw[1] ,
    \top_I.branch[19].block[3].um_I.clk ,
    \top_I.branch[19].block[2].um_I.iw[17] ,
    \top_I.branch[19].block[2].um_I.iw[16] ,
    \top_I.branch[19].block[2].um_I.iw[15] ,
    \top_I.branch[19].block[2].um_I.iw[14] ,
    \top_I.branch[19].block[2].um_I.iw[13] ,
    \top_I.branch[19].block[2].um_I.iw[12] ,
    \top_I.branch[19].block[2].um_I.iw[11] ,
    \top_I.branch[19].block[2].um_I.iw[10] ,
    \top_I.branch[19].block[2].um_I.iw[9] ,
    \top_I.branch[19].block[2].um_I.iw[8] ,
    \top_I.branch[19].block[2].um_I.iw[7] ,
    \top_I.branch[19].block[2].um_I.iw[6] ,
    \top_I.branch[19].block[2].um_I.iw[5] ,
    \top_I.branch[19].block[2].um_I.iw[4] ,
    \top_I.branch[19].block[2].um_I.iw[3] ,
    \top_I.branch[19].block[2].um_I.iw[2] ,
    \top_I.branch[19].block[2].um_I.iw[1] ,
    \top_I.branch[19].block[2].um_I.clk ,
    \top_I.branch[19].block[1].um_I.iw[17] ,
    \top_I.branch[19].block[1].um_I.iw[16] ,
    \top_I.branch[19].block[1].um_I.iw[15] ,
    \top_I.branch[19].block[1].um_I.iw[14] ,
    \top_I.branch[19].block[1].um_I.iw[13] ,
    \top_I.branch[19].block[1].um_I.iw[12] ,
    \top_I.branch[19].block[1].um_I.iw[11] ,
    \top_I.branch[19].block[1].um_I.iw[10] ,
    \top_I.branch[19].block[1].um_I.iw[9] ,
    \top_I.branch[19].block[1].um_I.iw[8] ,
    \top_I.branch[19].block[1].um_I.iw[7] ,
    \top_I.branch[19].block[1].um_I.iw[6] ,
    \top_I.branch[19].block[1].um_I.iw[5] ,
    \top_I.branch[19].block[1].um_I.iw[4] ,
    \top_I.branch[19].block[1].um_I.iw[3] ,
    \top_I.branch[19].block[1].um_I.iw[2] ,
    \top_I.branch[19].block[1].um_I.iw[1] ,
    \top_I.branch[19].block[1].um_I.clk ,
    \top_I.branch[19].block[0].um_I.iw[17] ,
    \top_I.branch[19].block[0].um_I.iw[16] ,
    \top_I.branch[19].block[0].um_I.iw[15] ,
    \top_I.branch[19].block[0].um_I.iw[14] ,
    \top_I.branch[19].block[0].um_I.iw[13] ,
    \top_I.branch[19].block[0].um_I.iw[12] ,
    \top_I.branch[19].block[0].um_I.iw[11] ,
    \top_I.branch[19].block[0].um_I.iw[10] ,
    \top_I.branch[19].block[0].um_I.iw[9] ,
    \top_I.branch[19].block[0].um_I.iw[8] ,
    \top_I.branch[19].block[0].um_I.iw[7] ,
    \top_I.branch[19].block[0].um_I.iw[6] ,
    \top_I.branch[19].block[0].um_I.iw[5] ,
    \top_I.branch[19].block[0].um_I.iw[4] ,
    \top_I.branch[19].block[0].um_I.iw[3] ,
    \top_I.branch[19].block[0].um_I.iw[2] ,
    \top_I.branch[19].block[0].um_I.iw[1] ,
    \top_I.branch[19].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[19].block[15].um_I.pg_vdd ,
    \top_I.branch[19].block[14].um_I.pg_vdd ,
    \top_I.branch[19].block[13].um_I.pg_vdd ,
    \top_I.branch[19].block[12].um_I.pg_vdd ,
    \top_I.branch[19].block[11].um_I.pg_vdd ,
    \top_I.branch[19].block[10].um_I.pg_vdd ,
    \top_I.branch[19].block[9].um_I.pg_vdd ,
    \top_I.branch[19].block[8].um_I.pg_vdd ,
    \top_I.branch[19].block[7].um_I.pg_vdd ,
    \top_I.branch[19].block[6].um_I.pg_vdd ,
    \top_I.branch[19].block[5].um_I.pg_vdd ,
    \top_I.branch[19].block[4].um_I.pg_vdd ,
    \top_I.branch[19].block[3].um_I.pg_vdd ,
    \top_I.branch[19].block[2].um_I.pg_vdd ,
    \top_I.branch[19].block[1].um_I.pg_vdd ,
    \top_I.branch[19].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[1].mux_I  (.k_one(\top_I.branch[1].l_k_one ),
    .k_zero(\top_I.branch[1].l_addr[0] ),
    .addr({\top_I.branch[1].l_addr[0] ,
    \top_I.branch[1].l_addr[0] ,
    \top_I.branch[1].l_addr[0] ,
    \top_I.branch[1].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[1].block[15].um_I.ena ,
    \top_I.branch[1].block[14].um_I.ena ,
    \top_I.branch[1].block[13].um_I.ena ,
    \top_I.branch[1].block[12].um_I.ena ,
    \top_I.branch[1].block[11].um_I.ena ,
    \top_I.branch[1].block[10].um_I.ena ,
    \top_I.branch[1].block[9].um_I.ena ,
    \top_I.branch[1].block[8].um_I.ena ,
    \top_I.branch[1].block[7].um_I.ena ,
    \top_I.branch[1].block[6].um_I.ena ,
    \top_I.branch[1].block[5].um_I.ena ,
    \top_I.branch[1].block[4].um_I.ena ,
    \top_I.branch[1].block[3].um_I.ena ,
    \top_I.branch[1].block[2].um_I.ena ,
    \top_I.branch[1].block[1].um_I.ena ,
    \top_I.branch[1].block[0].um_I.ena }),
    .um_iw({\top_I.branch[1].block[15].um_I.iw[17] ,
    \top_I.branch[1].block[15].um_I.iw[16] ,
    \top_I.branch[1].block[15].um_I.iw[15] ,
    \top_I.branch[1].block[15].um_I.iw[14] ,
    \top_I.branch[1].block[15].um_I.iw[13] ,
    \top_I.branch[1].block[15].um_I.iw[12] ,
    \top_I.branch[1].block[15].um_I.iw[11] ,
    \top_I.branch[1].block[15].um_I.iw[10] ,
    \top_I.branch[1].block[15].um_I.iw[9] ,
    \top_I.branch[1].block[15].um_I.iw[8] ,
    \top_I.branch[1].block[15].um_I.iw[7] ,
    \top_I.branch[1].block[15].um_I.iw[6] ,
    \top_I.branch[1].block[15].um_I.iw[5] ,
    \top_I.branch[1].block[15].um_I.iw[4] ,
    \top_I.branch[1].block[15].um_I.iw[3] ,
    \top_I.branch[1].block[15].um_I.iw[2] ,
    \top_I.branch[1].block[15].um_I.iw[1] ,
    \top_I.branch[1].block[15].um_I.clk ,
    \top_I.branch[1].block[14].um_I.iw[17] ,
    \top_I.branch[1].block[14].um_I.iw[16] ,
    \top_I.branch[1].block[14].um_I.iw[15] ,
    \top_I.branch[1].block[14].um_I.iw[14] ,
    \top_I.branch[1].block[14].um_I.iw[13] ,
    \top_I.branch[1].block[14].um_I.iw[12] ,
    \top_I.branch[1].block[14].um_I.iw[11] ,
    \top_I.branch[1].block[14].um_I.iw[10] ,
    \top_I.branch[1].block[14].um_I.iw[9] ,
    \top_I.branch[1].block[14].um_I.iw[8] ,
    \top_I.branch[1].block[14].um_I.iw[7] ,
    \top_I.branch[1].block[14].um_I.iw[6] ,
    \top_I.branch[1].block[14].um_I.iw[5] ,
    \top_I.branch[1].block[14].um_I.iw[4] ,
    \top_I.branch[1].block[14].um_I.iw[3] ,
    \top_I.branch[1].block[14].um_I.iw[2] ,
    \top_I.branch[1].block[14].um_I.iw[1] ,
    \top_I.branch[1].block[14].um_I.clk ,
    \top_I.branch[1].block[13].um_I.iw[17] ,
    \top_I.branch[1].block[13].um_I.iw[16] ,
    \top_I.branch[1].block[13].um_I.iw[15] ,
    \top_I.branch[1].block[13].um_I.iw[14] ,
    \top_I.branch[1].block[13].um_I.iw[13] ,
    \top_I.branch[1].block[13].um_I.iw[12] ,
    \top_I.branch[1].block[13].um_I.iw[11] ,
    \top_I.branch[1].block[13].um_I.iw[10] ,
    \top_I.branch[1].block[13].um_I.iw[9] ,
    \top_I.branch[1].block[13].um_I.iw[8] ,
    \top_I.branch[1].block[13].um_I.iw[7] ,
    \top_I.branch[1].block[13].um_I.iw[6] ,
    \top_I.branch[1].block[13].um_I.iw[5] ,
    \top_I.branch[1].block[13].um_I.iw[4] ,
    \top_I.branch[1].block[13].um_I.iw[3] ,
    \top_I.branch[1].block[13].um_I.iw[2] ,
    \top_I.branch[1].block[13].um_I.iw[1] ,
    \top_I.branch[1].block[13].um_I.clk ,
    \top_I.branch[1].block[12].um_I.iw[17] ,
    \top_I.branch[1].block[12].um_I.iw[16] ,
    \top_I.branch[1].block[12].um_I.iw[15] ,
    \top_I.branch[1].block[12].um_I.iw[14] ,
    \top_I.branch[1].block[12].um_I.iw[13] ,
    \top_I.branch[1].block[12].um_I.iw[12] ,
    \top_I.branch[1].block[12].um_I.iw[11] ,
    \top_I.branch[1].block[12].um_I.iw[10] ,
    \top_I.branch[1].block[12].um_I.iw[9] ,
    \top_I.branch[1].block[12].um_I.iw[8] ,
    \top_I.branch[1].block[12].um_I.iw[7] ,
    \top_I.branch[1].block[12].um_I.iw[6] ,
    \top_I.branch[1].block[12].um_I.iw[5] ,
    \top_I.branch[1].block[12].um_I.iw[4] ,
    \top_I.branch[1].block[12].um_I.iw[3] ,
    \top_I.branch[1].block[12].um_I.iw[2] ,
    \top_I.branch[1].block[12].um_I.iw[1] ,
    \top_I.branch[1].block[12].um_I.clk ,
    \top_I.branch[1].block[11].um_I.iw[17] ,
    \top_I.branch[1].block[11].um_I.iw[16] ,
    \top_I.branch[1].block[11].um_I.iw[15] ,
    \top_I.branch[1].block[11].um_I.iw[14] ,
    \top_I.branch[1].block[11].um_I.iw[13] ,
    \top_I.branch[1].block[11].um_I.iw[12] ,
    \top_I.branch[1].block[11].um_I.iw[11] ,
    \top_I.branch[1].block[11].um_I.iw[10] ,
    \top_I.branch[1].block[11].um_I.iw[9] ,
    \top_I.branch[1].block[11].um_I.iw[8] ,
    \top_I.branch[1].block[11].um_I.iw[7] ,
    \top_I.branch[1].block[11].um_I.iw[6] ,
    \top_I.branch[1].block[11].um_I.iw[5] ,
    \top_I.branch[1].block[11].um_I.iw[4] ,
    \top_I.branch[1].block[11].um_I.iw[3] ,
    \top_I.branch[1].block[11].um_I.iw[2] ,
    \top_I.branch[1].block[11].um_I.iw[1] ,
    \top_I.branch[1].block[11].um_I.clk ,
    \top_I.branch[1].block[10].um_I.iw[17] ,
    \top_I.branch[1].block[10].um_I.iw[16] ,
    \top_I.branch[1].block[10].um_I.iw[15] ,
    \top_I.branch[1].block[10].um_I.iw[14] ,
    \top_I.branch[1].block[10].um_I.iw[13] ,
    \top_I.branch[1].block[10].um_I.iw[12] ,
    \top_I.branch[1].block[10].um_I.iw[11] ,
    \top_I.branch[1].block[10].um_I.iw[10] ,
    \top_I.branch[1].block[10].um_I.iw[9] ,
    \top_I.branch[1].block[10].um_I.iw[8] ,
    \top_I.branch[1].block[10].um_I.iw[7] ,
    \top_I.branch[1].block[10].um_I.iw[6] ,
    \top_I.branch[1].block[10].um_I.iw[5] ,
    \top_I.branch[1].block[10].um_I.iw[4] ,
    \top_I.branch[1].block[10].um_I.iw[3] ,
    \top_I.branch[1].block[10].um_I.iw[2] ,
    \top_I.branch[1].block[10].um_I.iw[1] ,
    \top_I.branch[1].block[10].um_I.clk ,
    \top_I.branch[1].block[9].um_I.iw[17] ,
    \top_I.branch[1].block[9].um_I.iw[16] ,
    \top_I.branch[1].block[9].um_I.iw[15] ,
    \top_I.branch[1].block[9].um_I.iw[14] ,
    \top_I.branch[1].block[9].um_I.iw[13] ,
    \top_I.branch[1].block[9].um_I.iw[12] ,
    \top_I.branch[1].block[9].um_I.iw[11] ,
    \top_I.branch[1].block[9].um_I.iw[10] ,
    \top_I.branch[1].block[9].um_I.iw[9] ,
    \top_I.branch[1].block[9].um_I.iw[8] ,
    \top_I.branch[1].block[9].um_I.iw[7] ,
    \top_I.branch[1].block[9].um_I.iw[6] ,
    \top_I.branch[1].block[9].um_I.iw[5] ,
    \top_I.branch[1].block[9].um_I.iw[4] ,
    \top_I.branch[1].block[9].um_I.iw[3] ,
    \top_I.branch[1].block[9].um_I.iw[2] ,
    \top_I.branch[1].block[9].um_I.iw[1] ,
    \top_I.branch[1].block[9].um_I.clk ,
    \top_I.branch[1].block[8].um_I.iw[17] ,
    \top_I.branch[1].block[8].um_I.iw[16] ,
    \top_I.branch[1].block[8].um_I.iw[15] ,
    \top_I.branch[1].block[8].um_I.iw[14] ,
    \top_I.branch[1].block[8].um_I.iw[13] ,
    \top_I.branch[1].block[8].um_I.iw[12] ,
    \top_I.branch[1].block[8].um_I.iw[11] ,
    \top_I.branch[1].block[8].um_I.iw[10] ,
    \top_I.branch[1].block[8].um_I.iw[9] ,
    \top_I.branch[1].block[8].um_I.iw[8] ,
    \top_I.branch[1].block[8].um_I.iw[7] ,
    \top_I.branch[1].block[8].um_I.iw[6] ,
    \top_I.branch[1].block[8].um_I.iw[5] ,
    \top_I.branch[1].block[8].um_I.iw[4] ,
    \top_I.branch[1].block[8].um_I.iw[3] ,
    \top_I.branch[1].block[8].um_I.iw[2] ,
    \top_I.branch[1].block[8].um_I.iw[1] ,
    \top_I.branch[1].block[8].um_I.clk ,
    \top_I.branch[1].block[7].um_I.iw[17] ,
    \top_I.branch[1].block[7].um_I.iw[16] ,
    \top_I.branch[1].block[7].um_I.iw[15] ,
    \top_I.branch[1].block[7].um_I.iw[14] ,
    \top_I.branch[1].block[7].um_I.iw[13] ,
    \top_I.branch[1].block[7].um_I.iw[12] ,
    \top_I.branch[1].block[7].um_I.iw[11] ,
    \top_I.branch[1].block[7].um_I.iw[10] ,
    \top_I.branch[1].block[7].um_I.iw[9] ,
    \top_I.branch[1].block[7].um_I.iw[8] ,
    \top_I.branch[1].block[7].um_I.iw[7] ,
    \top_I.branch[1].block[7].um_I.iw[6] ,
    \top_I.branch[1].block[7].um_I.iw[5] ,
    \top_I.branch[1].block[7].um_I.iw[4] ,
    \top_I.branch[1].block[7].um_I.iw[3] ,
    \top_I.branch[1].block[7].um_I.iw[2] ,
    \top_I.branch[1].block[7].um_I.iw[1] ,
    \top_I.branch[1].block[7].um_I.clk ,
    \top_I.branch[1].block[6].um_I.iw[17] ,
    \top_I.branch[1].block[6].um_I.iw[16] ,
    \top_I.branch[1].block[6].um_I.iw[15] ,
    \top_I.branch[1].block[6].um_I.iw[14] ,
    \top_I.branch[1].block[6].um_I.iw[13] ,
    \top_I.branch[1].block[6].um_I.iw[12] ,
    \top_I.branch[1].block[6].um_I.iw[11] ,
    \top_I.branch[1].block[6].um_I.iw[10] ,
    \top_I.branch[1].block[6].um_I.iw[9] ,
    \top_I.branch[1].block[6].um_I.iw[8] ,
    \top_I.branch[1].block[6].um_I.iw[7] ,
    \top_I.branch[1].block[6].um_I.iw[6] ,
    \top_I.branch[1].block[6].um_I.iw[5] ,
    \top_I.branch[1].block[6].um_I.iw[4] ,
    \top_I.branch[1].block[6].um_I.iw[3] ,
    \top_I.branch[1].block[6].um_I.iw[2] ,
    \top_I.branch[1].block[6].um_I.iw[1] ,
    \top_I.branch[1].block[6].um_I.clk ,
    \top_I.branch[1].block[5].um_I.iw[17] ,
    \top_I.branch[1].block[5].um_I.iw[16] ,
    \top_I.branch[1].block[5].um_I.iw[15] ,
    \top_I.branch[1].block[5].um_I.iw[14] ,
    \top_I.branch[1].block[5].um_I.iw[13] ,
    \top_I.branch[1].block[5].um_I.iw[12] ,
    \top_I.branch[1].block[5].um_I.iw[11] ,
    \top_I.branch[1].block[5].um_I.iw[10] ,
    \top_I.branch[1].block[5].um_I.iw[9] ,
    \top_I.branch[1].block[5].um_I.iw[8] ,
    \top_I.branch[1].block[5].um_I.iw[7] ,
    \top_I.branch[1].block[5].um_I.iw[6] ,
    \top_I.branch[1].block[5].um_I.iw[5] ,
    \top_I.branch[1].block[5].um_I.iw[4] ,
    \top_I.branch[1].block[5].um_I.iw[3] ,
    \top_I.branch[1].block[5].um_I.iw[2] ,
    \top_I.branch[1].block[5].um_I.iw[1] ,
    \top_I.branch[1].block[5].um_I.clk ,
    \top_I.branch[1].block[4].um_I.iw[17] ,
    \top_I.branch[1].block[4].um_I.iw[16] ,
    \top_I.branch[1].block[4].um_I.iw[15] ,
    \top_I.branch[1].block[4].um_I.iw[14] ,
    \top_I.branch[1].block[4].um_I.iw[13] ,
    \top_I.branch[1].block[4].um_I.iw[12] ,
    \top_I.branch[1].block[4].um_I.iw[11] ,
    \top_I.branch[1].block[4].um_I.iw[10] ,
    \top_I.branch[1].block[4].um_I.iw[9] ,
    \top_I.branch[1].block[4].um_I.iw[8] ,
    \top_I.branch[1].block[4].um_I.iw[7] ,
    \top_I.branch[1].block[4].um_I.iw[6] ,
    \top_I.branch[1].block[4].um_I.iw[5] ,
    \top_I.branch[1].block[4].um_I.iw[4] ,
    \top_I.branch[1].block[4].um_I.iw[3] ,
    \top_I.branch[1].block[4].um_I.iw[2] ,
    \top_I.branch[1].block[4].um_I.iw[1] ,
    \top_I.branch[1].block[4].um_I.clk ,
    \top_I.branch[1].block[3].um_I.iw[17] ,
    \top_I.branch[1].block[3].um_I.iw[16] ,
    \top_I.branch[1].block[3].um_I.iw[15] ,
    \top_I.branch[1].block[3].um_I.iw[14] ,
    \top_I.branch[1].block[3].um_I.iw[13] ,
    \top_I.branch[1].block[3].um_I.iw[12] ,
    \top_I.branch[1].block[3].um_I.iw[11] ,
    \top_I.branch[1].block[3].um_I.iw[10] ,
    \top_I.branch[1].block[3].um_I.iw[9] ,
    \top_I.branch[1].block[3].um_I.iw[8] ,
    \top_I.branch[1].block[3].um_I.iw[7] ,
    \top_I.branch[1].block[3].um_I.iw[6] ,
    \top_I.branch[1].block[3].um_I.iw[5] ,
    \top_I.branch[1].block[3].um_I.iw[4] ,
    \top_I.branch[1].block[3].um_I.iw[3] ,
    \top_I.branch[1].block[3].um_I.iw[2] ,
    \top_I.branch[1].block[3].um_I.iw[1] ,
    \top_I.branch[1].block[3].um_I.clk ,
    \top_I.branch[1].block[2].um_I.iw[17] ,
    \top_I.branch[1].block[2].um_I.iw[16] ,
    \top_I.branch[1].block[2].um_I.iw[15] ,
    \top_I.branch[1].block[2].um_I.iw[14] ,
    \top_I.branch[1].block[2].um_I.iw[13] ,
    \top_I.branch[1].block[2].um_I.iw[12] ,
    \top_I.branch[1].block[2].um_I.iw[11] ,
    \top_I.branch[1].block[2].um_I.iw[10] ,
    \top_I.branch[1].block[2].um_I.iw[9] ,
    \top_I.branch[1].block[2].um_I.iw[8] ,
    \top_I.branch[1].block[2].um_I.iw[7] ,
    \top_I.branch[1].block[2].um_I.iw[6] ,
    \top_I.branch[1].block[2].um_I.iw[5] ,
    \top_I.branch[1].block[2].um_I.iw[4] ,
    \top_I.branch[1].block[2].um_I.iw[3] ,
    \top_I.branch[1].block[2].um_I.iw[2] ,
    \top_I.branch[1].block[2].um_I.iw[1] ,
    \top_I.branch[1].block[2].um_I.clk ,
    \top_I.branch[1].block[1].um_I.iw[17] ,
    \top_I.branch[1].block[1].um_I.iw[16] ,
    \top_I.branch[1].block[1].um_I.iw[15] ,
    \top_I.branch[1].block[1].um_I.iw[14] ,
    \top_I.branch[1].block[1].um_I.iw[13] ,
    \top_I.branch[1].block[1].um_I.iw[12] ,
    \top_I.branch[1].block[1].um_I.iw[11] ,
    \top_I.branch[1].block[1].um_I.iw[10] ,
    \top_I.branch[1].block[1].um_I.iw[9] ,
    \top_I.branch[1].block[1].um_I.iw[8] ,
    \top_I.branch[1].block[1].um_I.iw[7] ,
    \top_I.branch[1].block[1].um_I.iw[6] ,
    \top_I.branch[1].block[1].um_I.iw[5] ,
    \top_I.branch[1].block[1].um_I.iw[4] ,
    \top_I.branch[1].block[1].um_I.iw[3] ,
    \top_I.branch[1].block[1].um_I.iw[2] ,
    \top_I.branch[1].block[1].um_I.iw[1] ,
    \top_I.branch[1].block[1].um_I.clk ,
    \top_I.branch[1].block[0].um_I.iw[17] ,
    \top_I.branch[1].block[0].um_I.iw[16] ,
    \top_I.branch[1].block[0].um_I.iw[15] ,
    \top_I.branch[1].block[0].um_I.iw[14] ,
    \top_I.branch[1].block[0].um_I.iw[13] ,
    \top_I.branch[1].block[0].um_I.iw[12] ,
    \top_I.branch[1].block[0].um_I.iw[11] ,
    \top_I.branch[1].block[0].um_I.iw[10] ,
    \top_I.branch[1].block[0].um_I.iw[9] ,
    \top_I.branch[1].block[0].um_I.iw[8] ,
    \top_I.branch[1].block[0].um_I.iw[7] ,
    \top_I.branch[1].block[0].um_I.iw[6] ,
    \top_I.branch[1].block[0].um_I.iw[5] ,
    \top_I.branch[1].block[0].um_I.iw[4] ,
    \top_I.branch[1].block[0].um_I.iw[3] ,
    \top_I.branch[1].block[0].um_I.iw[2] ,
    \top_I.branch[1].block[0].um_I.iw[1] ,
    \top_I.branch[1].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[1].block[15].um_I.pg_vdd ,
    \top_I.branch[1].block[14].um_I.pg_vdd ,
    \top_I.branch[1].block[13].um_I.pg_vdd ,
    \top_I.branch[1].block[12].um_I.pg_vdd ,
    \top_I.branch[1].block[11].um_I.pg_vdd ,
    \top_I.branch[1].block[10].um_I.pg_vdd ,
    \top_I.branch[1].block[9].um_I.pg_vdd ,
    \top_I.branch[1].block[8].um_I.pg_vdd ,
    \top_I.branch[1].block[7].um_I.pg_vdd ,
    \top_I.branch[1].block[6].um_I.pg_vdd ,
    \top_I.branch[1].block[5].um_I.pg_vdd ,
    \top_I.branch[1].block[4].um_I.pg_vdd ,
    \top_I.branch[1].block[3].um_I.pg_vdd ,
    \top_I.branch[1].block[2].um_I.pg_vdd ,
    \top_I.branch[1].block[1].um_I.pg_vdd ,
    \top_I.branch[1].block[0].um_I.pg_vdd }));
 tt_pg_vdd_2 \top_I.branch[20].block[14].um_I.block_20_14.tt_pg_vdd_I  (.ctrl(\top_I.branch[20].block[14].um_I.pg_vdd ));
 tt_um_urish_dffram \top_I.branch[20].block[14].um_I.block_20_14.tt_um_I  (.clk(\top_I.branch[20].block[14].um_I.clk ),
    .ena(\top_I.branch[20].block[14].um_I.ena ),
    .rst_n(\top_I.branch[20].block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[20].block[14].um_I.iw[9] ,
    \top_I.branch[20].block[14].um_I.iw[8] ,
    \top_I.branch[20].block[14].um_I.iw[7] ,
    \top_I.branch[20].block[14].um_I.iw[6] ,
    \top_I.branch[20].block[14].um_I.iw[5] ,
    \top_I.branch[20].block[14].um_I.iw[4] ,
    \top_I.branch[20].block[14].um_I.iw[3] ,
    \top_I.branch[20].block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[20].block[14].um_I.iw[17] ,
    \top_I.branch[20].block[14].um_I.iw[16] ,
    \top_I.branch[20].block[14].um_I.iw[15] ,
    \top_I.branch[20].block[14].um_I.iw[14] ,
    \top_I.branch[20].block[14].um_I.iw[13] ,
    \top_I.branch[20].block[14].um_I.iw[12] ,
    \top_I.branch[20].block[14].um_I.iw[11] ,
    \top_I.branch[20].block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[20].block[14].um_I.ow[23] ,
    \top_I.branch[20].block[14].um_I.ow[22] ,
    \top_I.branch[20].block[14].um_I.ow[21] ,
    \top_I.branch[20].block[14].um_I.ow[20] ,
    \top_I.branch[20].block[14].um_I.ow[19] ,
    \top_I.branch[20].block[14].um_I.ow[18] ,
    \top_I.branch[20].block[14].um_I.ow[17] ,
    \top_I.branch[20].block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[20].block[14].um_I.ow[15] ,
    \top_I.branch[20].block[14].um_I.ow[14] ,
    \top_I.branch[20].block[14].um_I.ow[13] ,
    \top_I.branch[20].block[14].um_I.ow[12] ,
    \top_I.branch[20].block[14].um_I.ow[11] ,
    \top_I.branch[20].block[14].um_I.ow[10] ,
    \top_I.branch[20].block[14].um_I.ow[9] ,
    \top_I.branch[20].block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[20].block[14].um_I.ow[7] ,
    \top_I.branch[20].block[14].um_I.ow[6] ,
    \top_I.branch[20].block[14].um_I.ow[5] ,
    \top_I.branch[20].block[14].um_I.ow[4] ,
    \top_I.branch[20].block[14].um_I.ow[3] ,
    \top_I.branch[20].block[14].um_I.ow[2] ,
    \top_I.branch[20].block[14].um_I.ow[1] ,
    \top_I.branch[20].block[14].um_I.ow[0] }));
 tt_mux \top_I.branch[20].mux_I  (.k_one(\top_I.branch[20].l_addr[1] ),
    .k_zero(\top_I.branch[20].l_addr[0] ),
    .addr({\top_I.branch[20].l_addr[1] ,
    \top_I.branch[20].l_addr[0] ,
    \top_I.branch[20].l_addr[1] ,
    \top_I.branch[20].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[20].block[15].um_I.ena ,
    \top_I.branch[20].block[14].um_I.ena ,
    \top_I.branch[20].block[13].um_I.ena ,
    \top_I.branch[20].block[12].um_I.ena ,
    \top_I.branch[20].block[11].um_I.ena ,
    \top_I.branch[20].block[10].um_I.ena ,
    \top_I.branch[20].block[9].um_I.ena ,
    \top_I.branch[20].block[8].um_I.ena ,
    \top_I.branch[20].block[7].um_I.ena ,
    \top_I.branch[20].block[6].um_I.ena ,
    \top_I.branch[20].block[5].um_I.ena ,
    \top_I.branch[20].block[4].um_I.ena ,
    \top_I.branch[20].block[3].um_I.ena ,
    \top_I.branch[20].block[2].um_I.ena ,
    \top_I.branch[20].block[1].um_I.ena ,
    \top_I.branch[20].block[0].um_I.ena }),
    .um_iw({\top_I.branch[20].block[15].um_I.iw[17] ,
    \top_I.branch[20].block[15].um_I.iw[16] ,
    \top_I.branch[20].block[15].um_I.iw[15] ,
    \top_I.branch[20].block[15].um_I.iw[14] ,
    \top_I.branch[20].block[15].um_I.iw[13] ,
    \top_I.branch[20].block[15].um_I.iw[12] ,
    \top_I.branch[20].block[15].um_I.iw[11] ,
    \top_I.branch[20].block[15].um_I.iw[10] ,
    \top_I.branch[20].block[15].um_I.iw[9] ,
    \top_I.branch[20].block[15].um_I.iw[8] ,
    \top_I.branch[20].block[15].um_I.iw[7] ,
    \top_I.branch[20].block[15].um_I.iw[6] ,
    \top_I.branch[20].block[15].um_I.iw[5] ,
    \top_I.branch[20].block[15].um_I.iw[4] ,
    \top_I.branch[20].block[15].um_I.iw[3] ,
    \top_I.branch[20].block[15].um_I.iw[2] ,
    \top_I.branch[20].block[15].um_I.iw[1] ,
    \top_I.branch[20].block[15].um_I.clk ,
    \top_I.branch[20].block[14].um_I.iw[17] ,
    \top_I.branch[20].block[14].um_I.iw[16] ,
    \top_I.branch[20].block[14].um_I.iw[15] ,
    \top_I.branch[20].block[14].um_I.iw[14] ,
    \top_I.branch[20].block[14].um_I.iw[13] ,
    \top_I.branch[20].block[14].um_I.iw[12] ,
    \top_I.branch[20].block[14].um_I.iw[11] ,
    \top_I.branch[20].block[14].um_I.iw[10] ,
    \top_I.branch[20].block[14].um_I.iw[9] ,
    \top_I.branch[20].block[14].um_I.iw[8] ,
    \top_I.branch[20].block[14].um_I.iw[7] ,
    \top_I.branch[20].block[14].um_I.iw[6] ,
    \top_I.branch[20].block[14].um_I.iw[5] ,
    \top_I.branch[20].block[14].um_I.iw[4] ,
    \top_I.branch[20].block[14].um_I.iw[3] ,
    \top_I.branch[20].block[14].um_I.iw[2] ,
    \top_I.branch[20].block[14].um_I.iw[1] ,
    \top_I.branch[20].block[14].um_I.clk ,
    \top_I.branch[20].block[13].um_I.iw[17] ,
    \top_I.branch[20].block[13].um_I.iw[16] ,
    \top_I.branch[20].block[13].um_I.iw[15] ,
    \top_I.branch[20].block[13].um_I.iw[14] ,
    \top_I.branch[20].block[13].um_I.iw[13] ,
    \top_I.branch[20].block[13].um_I.iw[12] ,
    \top_I.branch[20].block[13].um_I.iw[11] ,
    \top_I.branch[20].block[13].um_I.iw[10] ,
    \top_I.branch[20].block[13].um_I.iw[9] ,
    \top_I.branch[20].block[13].um_I.iw[8] ,
    \top_I.branch[20].block[13].um_I.iw[7] ,
    \top_I.branch[20].block[13].um_I.iw[6] ,
    \top_I.branch[20].block[13].um_I.iw[5] ,
    \top_I.branch[20].block[13].um_I.iw[4] ,
    \top_I.branch[20].block[13].um_I.iw[3] ,
    \top_I.branch[20].block[13].um_I.iw[2] ,
    \top_I.branch[20].block[13].um_I.iw[1] ,
    \top_I.branch[20].block[13].um_I.clk ,
    \top_I.branch[20].block[12].um_I.iw[17] ,
    \top_I.branch[20].block[12].um_I.iw[16] ,
    \top_I.branch[20].block[12].um_I.iw[15] ,
    \top_I.branch[20].block[12].um_I.iw[14] ,
    \top_I.branch[20].block[12].um_I.iw[13] ,
    \top_I.branch[20].block[12].um_I.iw[12] ,
    \top_I.branch[20].block[12].um_I.iw[11] ,
    \top_I.branch[20].block[12].um_I.iw[10] ,
    \top_I.branch[20].block[12].um_I.iw[9] ,
    \top_I.branch[20].block[12].um_I.iw[8] ,
    \top_I.branch[20].block[12].um_I.iw[7] ,
    \top_I.branch[20].block[12].um_I.iw[6] ,
    \top_I.branch[20].block[12].um_I.iw[5] ,
    \top_I.branch[20].block[12].um_I.iw[4] ,
    \top_I.branch[20].block[12].um_I.iw[3] ,
    \top_I.branch[20].block[12].um_I.iw[2] ,
    \top_I.branch[20].block[12].um_I.iw[1] ,
    \top_I.branch[20].block[12].um_I.clk ,
    \top_I.branch[20].block[11].um_I.iw[17] ,
    \top_I.branch[20].block[11].um_I.iw[16] ,
    \top_I.branch[20].block[11].um_I.iw[15] ,
    \top_I.branch[20].block[11].um_I.iw[14] ,
    \top_I.branch[20].block[11].um_I.iw[13] ,
    \top_I.branch[20].block[11].um_I.iw[12] ,
    \top_I.branch[20].block[11].um_I.iw[11] ,
    \top_I.branch[20].block[11].um_I.iw[10] ,
    \top_I.branch[20].block[11].um_I.iw[9] ,
    \top_I.branch[20].block[11].um_I.iw[8] ,
    \top_I.branch[20].block[11].um_I.iw[7] ,
    \top_I.branch[20].block[11].um_I.iw[6] ,
    \top_I.branch[20].block[11].um_I.iw[5] ,
    \top_I.branch[20].block[11].um_I.iw[4] ,
    \top_I.branch[20].block[11].um_I.iw[3] ,
    \top_I.branch[20].block[11].um_I.iw[2] ,
    \top_I.branch[20].block[11].um_I.iw[1] ,
    \top_I.branch[20].block[11].um_I.clk ,
    \top_I.branch[20].block[10].um_I.iw[17] ,
    \top_I.branch[20].block[10].um_I.iw[16] ,
    \top_I.branch[20].block[10].um_I.iw[15] ,
    \top_I.branch[20].block[10].um_I.iw[14] ,
    \top_I.branch[20].block[10].um_I.iw[13] ,
    \top_I.branch[20].block[10].um_I.iw[12] ,
    \top_I.branch[20].block[10].um_I.iw[11] ,
    \top_I.branch[20].block[10].um_I.iw[10] ,
    \top_I.branch[20].block[10].um_I.iw[9] ,
    \top_I.branch[20].block[10].um_I.iw[8] ,
    \top_I.branch[20].block[10].um_I.iw[7] ,
    \top_I.branch[20].block[10].um_I.iw[6] ,
    \top_I.branch[20].block[10].um_I.iw[5] ,
    \top_I.branch[20].block[10].um_I.iw[4] ,
    \top_I.branch[20].block[10].um_I.iw[3] ,
    \top_I.branch[20].block[10].um_I.iw[2] ,
    \top_I.branch[20].block[10].um_I.iw[1] ,
    \top_I.branch[20].block[10].um_I.clk ,
    \top_I.branch[20].block[9].um_I.iw[17] ,
    \top_I.branch[20].block[9].um_I.iw[16] ,
    \top_I.branch[20].block[9].um_I.iw[15] ,
    \top_I.branch[20].block[9].um_I.iw[14] ,
    \top_I.branch[20].block[9].um_I.iw[13] ,
    \top_I.branch[20].block[9].um_I.iw[12] ,
    \top_I.branch[20].block[9].um_I.iw[11] ,
    \top_I.branch[20].block[9].um_I.iw[10] ,
    \top_I.branch[20].block[9].um_I.iw[9] ,
    \top_I.branch[20].block[9].um_I.iw[8] ,
    \top_I.branch[20].block[9].um_I.iw[7] ,
    \top_I.branch[20].block[9].um_I.iw[6] ,
    \top_I.branch[20].block[9].um_I.iw[5] ,
    \top_I.branch[20].block[9].um_I.iw[4] ,
    \top_I.branch[20].block[9].um_I.iw[3] ,
    \top_I.branch[20].block[9].um_I.iw[2] ,
    \top_I.branch[20].block[9].um_I.iw[1] ,
    \top_I.branch[20].block[9].um_I.clk ,
    \top_I.branch[20].block[8].um_I.iw[17] ,
    \top_I.branch[20].block[8].um_I.iw[16] ,
    \top_I.branch[20].block[8].um_I.iw[15] ,
    \top_I.branch[20].block[8].um_I.iw[14] ,
    \top_I.branch[20].block[8].um_I.iw[13] ,
    \top_I.branch[20].block[8].um_I.iw[12] ,
    \top_I.branch[20].block[8].um_I.iw[11] ,
    \top_I.branch[20].block[8].um_I.iw[10] ,
    \top_I.branch[20].block[8].um_I.iw[9] ,
    \top_I.branch[20].block[8].um_I.iw[8] ,
    \top_I.branch[20].block[8].um_I.iw[7] ,
    \top_I.branch[20].block[8].um_I.iw[6] ,
    \top_I.branch[20].block[8].um_I.iw[5] ,
    \top_I.branch[20].block[8].um_I.iw[4] ,
    \top_I.branch[20].block[8].um_I.iw[3] ,
    \top_I.branch[20].block[8].um_I.iw[2] ,
    \top_I.branch[20].block[8].um_I.iw[1] ,
    \top_I.branch[20].block[8].um_I.clk ,
    \top_I.branch[20].block[7].um_I.iw[17] ,
    \top_I.branch[20].block[7].um_I.iw[16] ,
    \top_I.branch[20].block[7].um_I.iw[15] ,
    \top_I.branch[20].block[7].um_I.iw[14] ,
    \top_I.branch[20].block[7].um_I.iw[13] ,
    \top_I.branch[20].block[7].um_I.iw[12] ,
    \top_I.branch[20].block[7].um_I.iw[11] ,
    \top_I.branch[20].block[7].um_I.iw[10] ,
    \top_I.branch[20].block[7].um_I.iw[9] ,
    \top_I.branch[20].block[7].um_I.iw[8] ,
    \top_I.branch[20].block[7].um_I.iw[7] ,
    \top_I.branch[20].block[7].um_I.iw[6] ,
    \top_I.branch[20].block[7].um_I.iw[5] ,
    \top_I.branch[20].block[7].um_I.iw[4] ,
    \top_I.branch[20].block[7].um_I.iw[3] ,
    \top_I.branch[20].block[7].um_I.iw[2] ,
    \top_I.branch[20].block[7].um_I.iw[1] ,
    \top_I.branch[20].block[7].um_I.clk ,
    \top_I.branch[20].block[6].um_I.iw[17] ,
    \top_I.branch[20].block[6].um_I.iw[16] ,
    \top_I.branch[20].block[6].um_I.iw[15] ,
    \top_I.branch[20].block[6].um_I.iw[14] ,
    \top_I.branch[20].block[6].um_I.iw[13] ,
    \top_I.branch[20].block[6].um_I.iw[12] ,
    \top_I.branch[20].block[6].um_I.iw[11] ,
    \top_I.branch[20].block[6].um_I.iw[10] ,
    \top_I.branch[20].block[6].um_I.iw[9] ,
    \top_I.branch[20].block[6].um_I.iw[8] ,
    \top_I.branch[20].block[6].um_I.iw[7] ,
    \top_I.branch[20].block[6].um_I.iw[6] ,
    \top_I.branch[20].block[6].um_I.iw[5] ,
    \top_I.branch[20].block[6].um_I.iw[4] ,
    \top_I.branch[20].block[6].um_I.iw[3] ,
    \top_I.branch[20].block[6].um_I.iw[2] ,
    \top_I.branch[20].block[6].um_I.iw[1] ,
    \top_I.branch[20].block[6].um_I.clk ,
    \top_I.branch[20].block[5].um_I.iw[17] ,
    \top_I.branch[20].block[5].um_I.iw[16] ,
    \top_I.branch[20].block[5].um_I.iw[15] ,
    \top_I.branch[20].block[5].um_I.iw[14] ,
    \top_I.branch[20].block[5].um_I.iw[13] ,
    \top_I.branch[20].block[5].um_I.iw[12] ,
    \top_I.branch[20].block[5].um_I.iw[11] ,
    \top_I.branch[20].block[5].um_I.iw[10] ,
    \top_I.branch[20].block[5].um_I.iw[9] ,
    \top_I.branch[20].block[5].um_I.iw[8] ,
    \top_I.branch[20].block[5].um_I.iw[7] ,
    \top_I.branch[20].block[5].um_I.iw[6] ,
    \top_I.branch[20].block[5].um_I.iw[5] ,
    \top_I.branch[20].block[5].um_I.iw[4] ,
    \top_I.branch[20].block[5].um_I.iw[3] ,
    \top_I.branch[20].block[5].um_I.iw[2] ,
    \top_I.branch[20].block[5].um_I.iw[1] ,
    \top_I.branch[20].block[5].um_I.clk ,
    \top_I.branch[20].block[4].um_I.iw[17] ,
    \top_I.branch[20].block[4].um_I.iw[16] ,
    \top_I.branch[20].block[4].um_I.iw[15] ,
    \top_I.branch[20].block[4].um_I.iw[14] ,
    \top_I.branch[20].block[4].um_I.iw[13] ,
    \top_I.branch[20].block[4].um_I.iw[12] ,
    \top_I.branch[20].block[4].um_I.iw[11] ,
    \top_I.branch[20].block[4].um_I.iw[10] ,
    \top_I.branch[20].block[4].um_I.iw[9] ,
    \top_I.branch[20].block[4].um_I.iw[8] ,
    \top_I.branch[20].block[4].um_I.iw[7] ,
    \top_I.branch[20].block[4].um_I.iw[6] ,
    \top_I.branch[20].block[4].um_I.iw[5] ,
    \top_I.branch[20].block[4].um_I.iw[4] ,
    \top_I.branch[20].block[4].um_I.iw[3] ,
    \top_I.branch[20].block[4].um_I.iw[2] ,
    \top_I.branch[20].block[4].um_I.iw[1] ,
    \top_I.branch[20].block[4].um_I.clk ,
    \top_I.branch[20].block[3].um_I.iw[17] ,
    \top_I.branch[20].block[3].um_I.iw[16] ,
    \top_I.branch[20].block[3].um_I.iw[15] ,
    \top_I.branch[20].block[3].um_I.iw[14] ,
    \top_I.branch[20].block[3].um_I.iw[13] ,
    \top_I.branch[20].block[3].um_I.iw[12] ,
    \top_I.branch[20].block[3].um_I.iw[11] ,
    \top_I.branch[20].block[3].um_I.iw[10] ,
    \top_I.branch[20].block[3].um_I.iw[9] ,
    \top_I.branch[20].block[3].um_I.iw[8] ,
    \top_I.branch[20].block[3].um_I.iw[7] ,
    \top_I.branch[20].block[3].um_I.iw[6] ,
    \top_I.branch[20].block[3].um_I.iw[5] ,
    \top_I.branch[20].block[3].um_I.iw[4] ,
    \top_I.branch[20].block[3].um_I.iw[3] ,
    \top_I.branch[20].block[3].um_I.iw[2] ,
    \top_I.branch[20].block[3].um_I.iw[1] ,
    \top_I.branch[20].block[3].um_I.clk ,
    \top_I.branch[20].block[2].um_I.iw[17] ,
    \top_I.branch[20].block[2].um_I.iw[16] ,
    \top_I.branch[20].block[2].um_I.iw[15] ,
    \top_I.branch[20].block[2].um_I.iw[14] ,
    \top_I.branch[20].block[2].um_I.iw[13] ,
    \top_I.branch[20].block[2].um_I.iw[12] ,
    \top_I.branch[20].block[2].um_I.iw[11] ,
    \top_I.branch[20].block[2].um_I.iw[10] ,
    \top_I.branch[20].block[2].um_I.iw[9] ,
    \top_I.branch[20].block[2].um_I.iw[8] ,
    \top_I.branch[20].block[2].um_I.iw[7] ,
    \top_I.branch[20].block[2].um_I.iw[6] ,
    \top_I.branch[20].block[2].um_I.iw[5] ,
    \top_I.branch[20].block[2].um_I.iw[4] ,
    \top_I.branch[20].block[2].um_I.iw[3] ,
    \top_I.branch[20].block[2].um_I.iw[2] ,
    \top_I.branch[20].block[2].um_I.iw[1] ,
    \top_I.branch[20].block[2].um_I.clk ,
    \top_I.branch[20].block[1].um_I.iw[17] ,
    \top_I.branch[20].block[1].um_I.iw[16] ,
    \top_I.branch[20].block[1].um_I.iw[15] ,
    \top_I.branch[20].block[1].um_I.iw[14] ,
    \top_I.branch[20].block[1].um_I.iw[13] ,
    \top_I.branch[20].block[1].um_I.iw[12] ,
    \top_I.branch[20].block[1].um_I.iw[11] ,
    \top_I.branch[20].block[1].um_I.iw[10] ,
    \top_I.branch[20].block[1].um_I.iw[9] ,
    \top_I.branch[20].block[1].um_I.iw[8] ,
    \top_I.branch[20].block[1].um_I.iw[7] ,
    \top_I.branch[20].block[1].um_I.iw[6] ,
    \top_I.branch[20].block[1].um_I.iw[5] ,
    \top_I.branch[20].block[1].um_I.iw[4] ,
    \top_I.branch[20].block[1].um_I.iw[3] ,
    \top_I.branch[20].block[1].um_I.iw[2] ,
    \top_I.branch[20].block[1].um_I.iw[1] ,
    \top_I.branch[20].block[1].um_I.clk ,
    \top_I.branch[20].block[0].um_I.iw[17] ,
    \top_I.branch[20].block[0].um_I.iw[16] ,
    \top_I.branch[20].block[0].um_I.iw[15] ,
    \top_I.branch[20].block[0].um_I.iw[14] ,
    \top_I.branch[20].block[0].um_I.iw[13] ,
    \top_I.branch[20].block[0].um_I.iw[12] ,
    \top_I.branch[20].block[0].um_I.iw[11] ,
    \top_I.branch[20].block[0].um_I.iw[10] ,
    \top_I.branch[20].block[0].um_I.iw[9] ,
    \top_I.branch[20].block[0].um_I.iw[8] ,
    \top_I.branch[20].block[0].um_I.iw[7] ,
    \top_I.branch[20].block[0].um_I.iw[6] ,
    \top_I.branch[20].block[0].um_I.iw[5] ,
    \top_I.branch[20].block[0].um_I.iw[4] ,
    \top_I.branch[20].block[0].um_I.iw[3] ,
    \top_I.branch[20].block[0].um_I.iw[2] ,
    \top_I.branch[20].block[0].um_I.iw[1] ,
    \top_I.branch[20].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.ow[23] ,
    \top_I.branch[20].block[14].um_I.ow[22] ,
    \top_I.branch[20].block[14].um_I.ow[21] ,
    \top_I.branch[20].block[14].um_I.ow[20] ,
    \top_I.branch[20].block[14].um_I.ow[19] ,
    \top_I.branch[20].block[14].um_I.ow[18] ,
    \top_I.branch[20].block[14].um_I.ow[17] ,
    \top_I.branch[20].block[14].um_I.ow[16] ,
    \top_I.branch[20].block[14].um_I.ow[15] ,
    \top_I.branch[20].block[14].um_I.ow[14] ,
    \top_I.branch[20].block[14].um_I.ow[13] ,
    \top_I.branch[20].block[14].um_I.ow[12] ,
    \top_I.branch[20].block[14].um_I.ow[11] ,
    \top_I.branch[20].block[14].um_I.ow[10] ,
    \top_I.branch[20].block[14].um_I.ow[9] ,
    \top_I.branch[20].block[14].um_I.ow[8] ,
    \top_I.branch[20].block[14].um_I.ow[7] ,
    \top_I.branch[20].block[14].um_I.ow[6] ,
    \top_I.branch[20].block[14].um_I.ow[5] ,
    \top_I.branch[20].block[14].um_I.ow[4] ,
    \top_I.branch[20].block[14].um_I.ow[3] ,
    \top_I.branch[20].block[14].um_I.ow[2] ,
    \top_I.branch[20].block[14].um_I.ow[1] ,
    \top_I.branch[20].block[14].um_I.ow[0] ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[20].block[15].um_I.pg_vdd ,
    \top_I.branch[20].block[14].um_I.pg_vdd ,
    \top_I.branch[20].block[13].um_I.pg_vdd ,
    \top_I.branch[20].block[12].um_I.pg_vdd ,
    \top_I.branch[20].block[11].um_I.pg_vdd ,
    \top_I.branch[20].block[10].um_I.pg_vdd ,
    \top_I.branch[20].block[9].um_I.pg_vdd ,
    \top_I.branch[20].block[8].um_I.pg_vdd ,
    \top_I.branch[20].block[7].um_I.pg_vdd ,
    \top_I.branch[20].block[6].um_I.pg_vdd ,
    \top_I.branch[20].block[5].um_I.pg_vdd ,
    \top_I.branch[20].block[4].um_I.pg_vdd ,
    \top_I.branch[20].block[3].um_I.pg_vdd ,
    \top_I.branch[20].block[2].um_I.pg_vdd ,
    \top_I.branch[20].block[1].um_I.pg_vdd ,
    \top_I.branch[20].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[21].mux_I  (.k_one(\top_I.branch[21].l_addr[1] ),
    .k_zero(\top_I.branch[21].l_addr[0] ),
    .addr({\top_I.branch[21].l_addr[1] ,
    \top_I.branch[21].l_addr[0] ,
    \top_I.branch[21].l_addr[1] ,
    \top_I.branch[21].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[21].block[15].um_I.ena ,
    \top_I.branch[21].block[14].um_I.ena ,
    \top_I.branch[21].block[13].um_I.ena ,
    \top_I.branch[21].block[12].um_I.ena ,
    \top_I.branch[21].block[11].um_I.ena ,
    \top_I.branch[21].block[10].um_I.ena ,
    \top_I.branch[21].block[9].um_I.ena ,
    \top_I.branch[21].block[8].um_I.ena ,
    \top_I.branch[21].block[7].um_I.ena ,
    \top_I.branch[21].block[6].um_I.ena ,
    \top_I.branch[21].block[5].um_I.ena ,
    \top_I.branch[21].block[4].um_I.ena ,
    \top_I.branch[21].block[3].um_I.ena ,
    \top_I.branch[21].block[2].um_I.ena ,
    \top_I.branch[21].block[1].um_I.ena ,
    \top_I.branch[21].block[0].um_I.ena }),
    .um_iw({\top_I.branch[21].block[15].um_I.iw[17] ,
    \top_I.branch[21].block[15].um_I.iw[16] ,
    \top_I.branch[21].block[15].um_I.iw[15] ,
    \top_I.branch[21].block[15].um_I.iw[14] ,
    \top_I.branch[21].block[15].um_I.iw[13] ,
    \top_I.branch[21].block[15].um_I.iw[12] ,
    \top_I.branch[21].block[15].um_I.iw[11] ,
    \top_I.branch[21].block[15].um_I.iw[10] ,
    \top_I.branch[21].block[15].um_I.iw[9] ,
    \top_I.branch[21].block[15].um_I.iw[8] ,
    \top_I.branch[21].block[15].um_I.iw[7] ,
    \top_I.branch[21].block[15].um_I.iw[6] ,
    \top_I.branch[21].block[15].um_I.iw[5] ,
    \top_I.branch[21].block[15].um_I.iw[4] ,
    \top_I.branch[21].block[15].um_I.iw[3] ,
    \top_I.branch[21].block[15].um_I.iw[2] ,
    \top_I.branch[21].block[15].um_I.iw[1] ,
    \top_I.branch[21].block[15].um_I.clk ,
    \top_I.branch[21].block[14].um_I.iw[17] ,
    \top_I.branch[21].block[14].um_I.iw[16] ,
    \top_I.branch[21].block[14].um_I.iw[15] ,
    \top_I.branch[21].block[14].um_I.iw[14] ,
    \top_I.branch[21].block[14].um_I.iw[13] ,
    \top_I.branch[21].block[14].um_I.iw[12] ,
    \top_I.branch[21].block[14].um_I.iw[11] ,
    \top_I.branch[21].block[14].um_I.iw[10] ,
    \top_I.branch[21].block[14].um_I.iw[9] ,
    \top_I.branch[21].block[14].um_I.iw[8] ,
    \top_I.branch[21].block[14].um_I.iw[7] ,
    \top_I.branch[21].block[14].um_I.iw[6] ,
    \top_I.branch[21].block[14].um_I.iw[5] ,
    \top_I.branch[21].block[14].um_I.iw[4] ,
    \top_I.branch[21].block[14].um_I.iw[3] ,
    \top_I.branch[21].block[14].um_I.iw[2] ,
    \top_I.branch[21].block[14].um_I.iw[1] ,
    \top_I.branch[21].block[14].um_I.clk ,
    \top_I.branch[21].block[13].um_I.iw[17] ,
    \top_I.branch[21].block[13].um_I.iw[16] ,
    \top_I.branch[21].block[13].um_I.iw[15] ,
    \top_I.branch[21].block[13].um_I.iw[14] ,
    \top_I.branch[21].block[13].um_I.iw[13] ,
    \top_I.branch[21].block[13].um_I.iw[12] ,
    \top_I.branch[21].block[13].um_I.iw[11] ,
    \top_I.branch[21].block[13].um_I.iw[10] ,
    \top_I.branch[21].block[13].um_I.iw[9] ,
    \top_I.branch[21].block[13].um_I.iw[8] ,
    \top_I.branch[21].block[13].um_I.iw[7] ,
    \top_I.branch[21].block[13].um_I.iw[6] ,
    \top_I.branch[21].block[13].um_I.iw[5] ,
    \top_I.branch[21].block[13].um_I.iw[4] ,
    \top_I.branch[21].block[13].um_I.iw[3] ,
    \top_I.branch[21].block[13].um_I.iw[2] ,
    \top_I.branch[21].block[13].um_I.iw[1] ,
    \top_I.branch[21].block[13].um_I.clk ,
    \top_I.branch[21].block[12].um_I.iw[17] ,
    \top_I.branch[21].block[12].um_I.iw[16] ,
    \top_I.branch[21].block[12].um_I.iw[15] ,
    \top_I.branch[21].block[12].um_I.iw[14] ,
    \top_I.branch[21].block[12].um_I.iw[13] ,
    \top_I.branch[21].block[12].um_I.iw[12] ,
    \top_I.branch[21].block[12].um_I.iw[11] ,
    \top_I.branch[21].block[12].um_I.iw[10] ,
    \top_I.branch[21].block[12].um_I.iw[9] ,
    \top_I.branch[21].block[12].um_I.iw[8] ,
    \top_I.branch[21].block[12].um_I.iw[7] ,
    \top_I.branch[21].block[12].um_I.iw[6] ,
    \top_I.branch[21].block[12].um_I.iw[5] ,
    \top_I.branch[21].block[12].um_I.iw[4] ,
    \top_I.branch[21].block[12].um_I.iw[3] ,
    \top_I.branch[21].block[12].um_I.iw[2] ,
    \top_I.branch[21].block[12].um_I.iw[1] ,
    \top_I.branch[21].block[12].um_I.clk ,
    \top_I.branch[21].block[11].um_I.iw[17] ,
    \top_I.branch[21].block[11].um_I.iw[16] ,
    \top_I.branch[21].block[11].um_I.iw[15] ,
    \top_I.branch[21].block[11].um_I.iw[14] ,
    \top_I.branch[21].block[11].um_I.iw[13] ,
    \top_I.branch[21].block[11].um_I.iw[12] ,
    \top_I.branch[21].block[11].um_I.iw[11] ,
    \top_I.branch[21].block[11].um_I.iw[10] ,
    \top_I.branch[21].block[11].um_I.iw[9] ,
    \top_I.branch[21].block[11].um_I.iw[8] ,
    \top_I.branch[21].block[11].um_I.iw[7] ,
    \top_I.branch[21].block[11].um_I.iw[6] ,
    \top_I.branch[21].block[11].um_I.iw[5] ,
    \top_I.branch[21].block[11].um_I.iw[4] ,
    \top_I.branch[21].block[11].um_I.iw[3] ,
    \top_I.branch[21].block[11].um_I.iw[2] ,
    \top_I.branch[21].block[11].um_I.iw[1] ,
    \top_I.branch[21].block[11].um_I.clk ,
    \top_I.branch[21].block[10].um_I.iw[17] ,
    \top_I.branch[21].block[10].um_I.iw[16] ,
    \top_I.branch[21].block[10].um_I.iw[15] ,
    \top_I.branch[21].block[10].um_I.iw[14] ,
    \top_I.branch[21].block[10].um_I.iw[13] ,
    \top_I.branch[21].block[10].um_I.iw[12] ,
    \top_I.branch[21].block[10].um_I.iw[11] ,
    \top_I.branch[21].block[10].um_I.iw[10] ,
    \top_I.branch[21].block[10].um_I.iw[9] ,
    \top_I.branch[21].block[10].um_I.iw[8] ,
    \top_I.branch[21].block[10].um_I.iw[7] ,
    \top_I.branch[21].block[10].um_I.iw[6] ,
    \top_I.branch[21].block[10].um_I.iw[5] ,
    \top_I.branch[21].block[10].um_I.iw[4] ,
    \top_I.branch[21].block[10].um_I.iw[3] ,
    \top_I.branch[21].block[10].um_I.iw[2] ,
    \top_I.branch[21].block[10].um_I.iw[1] ,
    \top_I.branch[21].block[10].um_I.clk ,
    \top_I.branch[21].block[9].um_I.iw[17] ,
    \top_I.branch[21].block[9].um_I.iw[16] ,
    \top_I.branch[21].block[9].um_I.iw[15] ,
    \top_I.branch[21].block[9].um_I.iw[14] ,
    \top_I.branch[21].block[9].um_I.iw[13] ,
    \top_I.branch[21].block[9].um_I.iw[12] ,
    \top_I.branch[21].block[9].um_I.iw[11] ,
    \top_I.branch[21].block[9].um_I.iw[10] ,
    \top_I.branch[21].block[9].um_I.iw[9] ,
    \top_I.branch[21].block[9].um_I.iw[8] ,
    \top_I.branch[21].block[9].um_I.iw[7] ,
    \top_I.branch[21].block[9].um_I.iw[6] ,
    \top_I.branch[21].block[9].um_I.iw[5] ,
    \top_I.branch[21].block[9].um_I.iw[4] ,
    \top_I.branch[21].block[9].um_I.iw[3] ,
    \top_I.branch[21].block[9].um_I.iw[2] ,
    \top_I.branch[21].block[9].um_I.iw[1] ,
    \top_I.branch[21].block[9].um_I.clk ,
    \top_I.branch[21].block[8].um_I.iw[17] ,
    \top_I.branch[21].block[8].um_I.iw[16] ,
    \top_I.branch[21].block[8].um_I.iw[15] ,
    \top_I.branch[21].block[8].um_I.iw[14] ,
    \top_I.branch[21].block[8].um_I.iw[13] ,
    \top_I.branch[21].block[8].um_I.iw[12] ,
    \top_I.branch[21].block[8].um_I.iw[11] ,
    \top_I.branch[21].block[8].um_I.iw[10] ,
    \top_I.branch[21].block[8].um_I.iw[9] ,
    \top_I.branch[21].block[8].um_I.iw[8] ,
    \top_I.branch[21].block[8].um_I.iw[7] ,
    \top_I.branch[21].block[8].um_I.iw[6] ,
    \top_I.branch[21].block[8].um_I.iw[5] ,
    \top_I.branch[21].block[8].um_I.iw[4] ,
    \top_I.branch[21].block[8].um_I.iw[3] ,
    \top_I.branch[21].block[8].um_I.iw[2] ,
    \top_I.branch[21].block[8].um_I.iw[1] ,
    \top_I.branch[21].block[8].um_I.clk ,
    \top_I.branch[21].block[7].um_I.iw[17] ,
    \top_I.branch[21].block[7].um_I.iw[16] ,
    \top_I.branch[21].block[7].um_I.iw[15] ,
    \top_I.branch[21].block[7].um_I.iw[14] ,
    \top_I.branch[21].block[7].um_I.iw[13] ,
    \top_I.branch[21].block[7].um_I.iw[12] ,
    \top_I.branch[21].block[7].um_I.iw[11] ,
    \top_I.branch[21].block[7].um_I.iw[10] ,
    \top_I.branch[21].block[7].um_I.iw[9] ,
    \top_I.branch[21].block[7].um_I.iw[8] ,
    \top_I.branch[21].block[7].um_I.iw[7] ,
    \top_I.branch[21].block[7].um_I.iw[6] ,
    \top_I.branch[21].block[7].um_I.iw[5] ,
    \top_I.branch[21].block[7].um_I.iw[4] ,
    \top_I.branch[21].block[7].um_I.iw[3] ,
    \top_I.branch[21].block[7].um_I.iw[2] ,
    \top_I.branch[21].block[7].um_I.iw[1] ,
    \top_I.branch[21].block[7].um_I.clk ,
    \top_I.branch[21].block[6].um_I.iw[17] ,
    \top_I.branch[21].block[6].um_I.iw[16] ,
    \top_I.branch[21].block[6].um_I.iw[15] ,
    \top_I.branch[21].block[6].um_I.iw[14] ,
    \top_I.branch[21].block[6].um_I.iw[13] ,
    \top_I.branch[21].block[6].um_I.iw[12] ,
    \top_I.branch[21].block[6].um_I.iw[11] ,
    \top_I.branch[21].block[6].um_I.iw[10] ,
    \top_I.branch[21].block[6].um_I.iw[9] ,
    \top_I.branch[21].block[6].um_I.iw[8] ,
    \top_I.branch[21].block[6].um_I.iw[7] ,
    \top_I.branch[21].block[6].um_I.iw[6] ,
    \top_I.branch[21].block[6].um_I.iw[5] ,
    \top_I.branch[21].block[6].um_I.iw[4] ,
    \top_I.branch[21].block[6].um_I.iw[3] ,
    \top_I.branch[21].block[6].um_I.iw[2] ,
    \top_I.branch[21].block[6].um_I.iw[1] ,
    \top_I.branch[21].block[6].um_I.clk ,
    \top_I.branch[21].block[5].um_I.iw[17] ,
    \top_I.branch[21].block[5].um_I.iw[16] ,
    \top_I.branch[21].block[5].um_I.iw[15] ,
    \top_I.branch[21].block[5].um_I.iw[14] ,
    \top_I.branch[21].block[5].um_I.iw[13] ,
    \top_I.branch[21].block[5].um_I.iw[12] ,
    \top_I.branch[21].block[5].um_I.iw[11] ,
    \top_I.branch[21].block[5].um_I.iw[10] ,
    \top_I.branch[21].block[5].um_I.iw[9] ,
    \top_I.branch[21].block[5].um_I.iw[8] ,
    \top_I.branch[21].block[5].um_I.iw[7] ,
    \top_I.branch[21].block[5].um_I.iw[6] ,
    \top_I.branch[21].block[5].um_I.iw[5] ,
    \top_I.branch[21].block[5].um_I.iw[4] ,
    \top_I.branch[21].block[5].um_I.iw[3] ,
    \top_I.branch[21].block[5].um_I.iw[2] ,
    \top_I.branch[21].block[5].um_I.iw[1] ,
    \top_I.branch[21].block[5].um_I.clk ,
    \top_I.branch[21].block[4].um_I.iw[17] ,
    \top_I.branch[21].block[4].um_I.iw[16] ,
    \top_I.branch[21].block[4].um_I.iw[15] ,
    \top_I.branch[21].block[4].um_I.iw[14] ,
    \top_I.branch[21].block[4].um_I.iw[13] ,
    \top_I.branch[21].block[4].um_I.iw[12] ,
    \top_I.branch[21].block[4].um_I.iw[11] ,
    \top_I.branch[21].block[4].um_I.iw[10] ,
    \top_I.branch[21].block[4].um_I.iw[9] ,
    \top_I.branch[21].block[4].um_I.iw[8] ,
    \top_I.branch[21].block[4].um_I.iw[7] ,
    \top_I.branch[21].block[4].um_I.iw[6] ,
    \top_I.branch[21].block[4].um_I.iw[5] ,
    \top_I.branch[21].block[4].um_I.iw[4] ,
    \top_I.branch[21].block[4].um_I.iw[3] ,
    \top_I.branch[21].block[4].um_I.iw[2] ,
    \top_I.branch[21].block[4].um_I.iw[1] ,
    \top_I.branch[21].block[4].um_I.clk ,
    \top_I.branch[21].block[3].um_I.iw[17] ,
    \top_I.branch[21].block[3].um_I.iw[16] ,
    \top_I.branch[21].block[3].um_I.iw[15] ,
    \top_I.branch[21].block[3].um_I.iw[14] ,
    \top_I.branch[21].block[3].um_I.iw[13] ,
    \top_I.branch[21].block[3].um_I.iw[12] ,
    \top_I.branch[21].block[3].um_I.iw[11] ,
    \top_I.branch[21].block[3].um_I.iw[10] ,
    \top_I.branch[21].block[3].um_I.iw[9] ,
    \top_I.branch[21].block[3].um_I.iw[8] ,
    \top_I.branch[21].block[3].um_I.iw[7] ,
    \top_I.branch[21].block[3].um_I.iw[6] ,
    \top_I.branch[21].block[3].um_I.iw[5] ,
    \top_I.branch[21].block[3].um_I.iw[4] ,
    \top_I.branch[21].block[3].um_I.iw[3] ,
    \top_I.branch[21].block[3].um_I.iw[2] ,
    \top_I.branch[21].block[3].um_I.iw[1] ,
    \top_I.branch[21].block[3].um_I.clk ,
    \top_I.branch[21].block[2].um_I.iw[17] ,
    \top_I.branch[21].block[2].um_I.iw[16] ,
    \top_I.branch[21].block[2].um_I.iw[15] ,
    \top_I.branch[21].block[2].um_I.iw[14] ,
    \top_I.branch[21].block[2].um_I.iw[13] ,
    \top_I.branch[21].block[2].um_I.iw[12] ,
    \top_I.branch[21].block[2].um_I.iw[11] ,
    \top_I.branch[21].block[2].um_I.iw[10] ,
    \top_I.branch[21].block[2].um_I.iw[9] ,
    \top_I.branch[21].block[2].um_I.iw[8] ,
    \top_I.branch[21].block[2].um_I.iw[7] ,
    \top_I.branch[21].block[2].um_I.iw[6] ,
    \top_I.branch[21].block[2].um_I.iw[5] ,
    \top_I.branch[21].block[2].um_I.iw[4] ,
    \top_I.branch[21].block[2].um_I.iw[3] ,
    \top_I.branch[21].block[2].um_I.iw[2] ,
    \top_I.branch[21].block[2].um_I.iw[1] ,
    \top_I.branch[21].block[2].um_I.clk ,
    \top_I.branch[21].block[1].um_I.iw[17] ,
    \top_I.branch[21].block[1].um_I.iw[16] ,
    \top_I.branch[21].block[1].um_I.iw[15] ,
    \top_I.branch[21].block[1].um_I.iw[14] ,
    \top_I.branch[21].block[1].um_I.iw[13] ,
    \top_I.branch[21].block[1].um_I.iw[12] ,
    \top_I.branch[21].block[1].um_I.iw[11] ,
    \top_I.branch[21].block[1].um_I.iw[10] ,
    \top_I.branch[21].block[1].um_I.iw[9] ,
    \top_I.branch[21].block[1].um_I.iw[8] ,
    \top_I.branch[21].block[1].um_I.iw[7] ,
    \top_I.branch[21].block[1].um_I.iw[6] ,
    \top_I.branch[21].block[1].um_I.iw[5] ,
    \top_I.branch[21].block[1].um_I.iw[4] ,
    \top_I.branch[21].block[1].um_I.iw[3] ,
    \top_I.branch[21].block[1].um_I.iw[2] ,
    \top_I.branch[21].block[1].um_I.iw[1] ,
    \top_I.branch[21].block[1].um_I.clk ,
    \top_I.branch[21].block[0].um_I.iw[17] ,
    \top_I.branch[21].block[0].um_I.iw[16] ,
    \top_I.branch[21].block[0].um_I.iw[15] ,
    \top_I.branch[21].block[0].um_I.iw[14] ,
    \top_I.branch[21].block[0].um_I.iw[13] ,
    \top_I.branch[21].block[0].um_I.iw[12] ,
    \top_I.branch[21].block[0].um_I.iw[11] ,
    \top_I.branch[21].block[0].um_I.iw[10] ,
    \top_I.branch[21].block[0].um_I.iw[9] ,
    \top_I.branch[21].block[0].um_I.iw[8] ,
    \top_I.branch[21].block[0].um_I.iw[7] ,
    \top_I.branch[21].block[0].um_I.iw[6] ,
    \top_I.branch[21].block[0].um_I.iw[5] ,
    \top_I.branch[21].block[0].um_I.iw[4] ,
    \top_I.branch[21].block[0].um_I.iw[3] ,
    \top_I.branch[21].block[0].um_I.iw[2] ,
    \top_I.branch[21].block[0].um_I.iw[1] ,
    \top_I.branch[21].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[21].block[15].um_I.pg_vdd ,
    \top_I.branch[21].block[14].um_I.pg_vdd ,
    \top_I.branch[21].block[13].um_I.pg_vdd ,
    \top_I.branch[21].block[12].um_I.pg_vdd ,
    \top_I.branch[21].block[11].um_I.pg_vdd ,
    \top_I.branch[21].block[10].um_I.pg_vdd ,
    \top_I.branch[21].block[9].um_I.pg_vdd ,
    \top_I.branch[21].block[8].um_I.pg_vdd ,
    \top_I.branch[21].block[7].um_I.pg_vdd ,
    \top_I.branch[21].block[6].um_I.pg_vdd ,
    \top_I.branch[21].block[5].um_I.pg_vdd ,
    \top_I.branch[21].block[4].um_I.pg_vdd ,
    \top_I.branch[21].block[3].um_I.pg_vdd ,
    \top_I.branch[21].block[2].um_I.pg_vdd ,
    \top_I.branch[21].block[1].um_I.pg_vdd ,
    \top_I.branch[21].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[22].mux_I  (.k_one(\top_I.branch[22].l_addr[0] ),
    .k_zero(\top_I.branch[22].l_addr[2] ),
    .addr({\top_I.branch[22].l_addr[0] ,
    \top_I.branch[22].l_addr[2] ,
    \top_I.branch[22].l_addr[0] ,
    \top_I.branch[22].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[22].block[15].um_I.ena ,
    \top_I.branch[22].block[14].um_I.ena ,
    \top_I.branch[22].block[13].um_I.ena ,
    \top_I.branch[22].block[12].um_I.ena ,
    \top_I.branch[22].block[11].um_I.ena ,
    \top_I.branch[22].block[10].um_I.ena ,
    \top_I.branch[22].block[9].um_I.ena ,
    \top_I.branch[22].block[8].um_I.ena ,
    \top_I.branch[22].block[7].um_I.ena ,
    \top_I.branch[22].block[6].um_I.ena ,
    \top_I.branch[22].block[5].um_I.ena ,
    \top_I.branch[22].block[4].um_I.ena ,
    \top_I.branch[22].block[3].um_I.ena ,
    \top_I.branch[22].block[2].um_I.ena ,
    \top_I.branch[22].block[1].um_I.ena ,
    \top_I.branch[22].block[0].um_I.ena }),
    .um_iw({\top_I.branch[22].block[15].um_I.iw[17] ,
    \top_I.branch[22].block[15].um_I.iw[16] ,
    \top_I.branch[22].block[15].um_I.iw[15] ,
    \top_I.branch[22].block[15].um_I.iw[14] ,
    \top_I.branch[22].block[15].um_I.iw[13] ,
    \top_I.branch[22].block[15].um_I.iw[12] ,
    \top_I.branch[22].block[15].um_I.iw[11] ,
    \top_I.branch[22].block[15].um_I.iw[10] ,
    \top_I.branch[22].block[15].um_I.iw[9] ,
    \top_I.branch[22].block[15].um_I.iw[8] ,
    \top_I.branch[22].block[15].um_I.iw[7] ,
    \top_I.branch[22].block[15].um_I.iw[6] ,
    \top_I.branch[22].block[15].um_I.iw[5] ,
    \top_I.branch[22].block[15].um_I.iw[4] ,
    \top_I.branch[22].block[15].um_I.iw[3] ,
    \top_I.branch[22].block[15].um_I.iw[2] ,
    \top_I.branch[22].block[15].um_I.iw[1] ,
    \top_I.branch[22].block[15].um_I.clk ,
    \top_I.branch[22].block[14].um_I.iw[17] ,
    \top_I.branch[22].block[14].um_I.iw[16] ,
    \top_I.branch[22].block[14].um_I.iw[15] ,
    \top_I.branch[22].block[14].um_I.iw[14] ,
    \top_I.branch[22].block[14].um_I.iw[13] ,
    \top_I.branch[22].block[14].um_I.iw[12] ,
    \top_I.branch[22].block[14].um_I.iw[11] ,
    \top_I.branch[22].block[14].um_I.iw[10] ,
    \top_I.branch[22].block[14].um_I.iw[9] ,
    \top_I.branch[22].block[14].um_I.iw[8] ,
    \top_I.branch[22].block[14].um_I.iw[7] ,
    \top_I.branch[22].block[14].um_I.iw[6] ,
    \top_I.branch[22].block[14].um_I.iw[5] ,
    \top_I.branch[22].block[14].um_I.iw[4] ,
    \top_I.branch[22].block[14].um_I.iw[3] ,
    \top_I.branch[22].block[14].um_I.iw[2] ,
    \top_I.branch[22].block[14].um_I.iw[1] ,
    \top_I.branch[22].block[14].um_I.clk ,
    \top_I.branch[22].block[13].um_I.iw[17] ,
    \top_I.branch[22].block[13].um_I.iw[16] ,
    \top_I.branch[22].block[13].um_I.iw[15] ,
    \top_I.branch[22].block[13].um_I.iw[14] ,
    \top_I.branch[22].block[13].um_I.iw[13] ,
    \top_I.branch[22].block[13].um_I.iw[12] ,
    \top_I.branch[22].block[13].um_I.iw[11] ,
    \top_I.branch[22].block[13].um_I.iw[10] ,
    \top_I.branch[22].block[13].um_I.iw[9] ,
    \top_I.branch[22].block[13].um_I.iw[8] ,
    \top_I.branch[22].block[13].um_I.iw[7] ,
    \top_I.branch[22].block[13].um_I.iw[6] ,
    \top_I.branch[22].block[13].um_I.iw[5] ,
    \top_I.branch[22].block[13].um_I.iw[4] ,
    \top_I.branch[22].block[13].um_I.iw[3] ,
    \top_I.branch[22].block[13].um_I.iw[2] ,
    \top_I.branch[22].block[13].um_I.iw[1] ,
    \top_I.branch[22].block[13].um_I.clk ,
    \top_I.branch[22].block[12].um_I.iw[17] ,
    \top_I.branch[22].block[12].um_I.iw[16] ,
    \top_I.branch[22].block[12].um_I.iw[15] ,
    \top_I.branch[22].block[12].um_I.iw[14] ,
    \top_I.branch[22].block[12].um_I.iw[13] ,
    \top_I.branch[22].block[12].um_I.iw[12] ,
    \top_I.branch[22].block[12].um_I.iw[11] ,
    \top_I.branch[22].block[12].um_I.iw[10] ,
    \top_I.branch[22].block[12].um_I.iw[9] ,
    \top_I.branch[22].block[12].um_I.iw[8] ,
    \top_I.branch[22].block[12].um_I.iw[7] ,
    \top_I.branch[22].block[12].um_I.iw[6] ,
    \top_I.branch[22].block[12].um_I.iw[5] ,
    \top_I.branch[22].block[12].um_I.iw[4] ,
    \top_I.branch[22].block[12].um_I.iw[3] ,
    \top_I.branch[22].block[12].um_I.iw[2] ,
    \top_I.branch[22].block[12].um_I.iw[1] ,
    \top_I.branch[22].block[12].um_I.clk ,
    \top_I.branch[22].block[11].um_I.iw[17] ,
    \top_I.branch[22].block[11].um_I.iw[16] ,
    \top_I.branch[22].block[11].um_I.iw[15] ,
    \top_I.branch[22].block[11].um_I.iw[14] ,
    \top_I.branch[22].block[11].um_I.iw[13] ,
    \top_I.branch[22].block[11].um_I.iw[12] ,
    \top_I.branch[22].block[11].um_I.iw[11] ,
    \top_I.branch[22].block[11].um_I.iw[10] ,
    \top_I.branch[22].block[11].um_I.iw[9] ,
    \top_I.branch[22].block[11].um_I.iw[8] ,
    \top_I.branch[22].block[11].um_I.iw[7] ,
    \top_I.branch[22].block[11].um_I.iw[6] ,
    \top_I.branch[22].block[11].um_I.iw[5] ,
    \top_I.branch[22].block[11].um_I.iw[4] ,
    \top_I.branch[22].block[11].um_I.iw[3] ,
    \top_I.branch[22].block[11].um_I.iw[2] ,
    \top_I.branch[22].block[11].um_I.iw[1] ,
    \top_I.branch[22].block[11].um_I.clk ,
    \top_I.branch[22].block[10].um_I.iw[17] ,
    \top_I.branch[22].block[10].um_I.iw[16] ,
    \top_I.branch[22].block[10].um_I.iw[15] ,
    \top_I.branch[22].block[10].um_I.iw[14] ,
    \top_I.branch[22].block[10].um_I.iw[13] ,
    \top_I.branch[22].block[10].um_I.iw[12] ,
    \top_I.branch[22].block[10].um_I.iw[11] ,
    \top_I.branch[22].block[10].um_I.iw[10] ,
    \top_I.branch[22].block[10].um_I.iw[9] ,
    \top_I.branch[22].block[10].um_I.iw[8] ,
    \top_I.branch[22].block[10].um_I.iw[7] ,
    \top_I.branch[22].block[10].um_I.iw[6] ,
    \top_I.branch[22].block[10].um_I.iw[5] ,
    \top_I.branch[22].block[10].um_I.iw[4] ,
    \top_I.branch[22].block[10].um_I.iw[3] ,
    \top_I.branch[22].block[10].um_I.iw[2] ,
    \top_I.branch[22].block[10].um_I.iw[1] ,
    \top_I.branch[22].block[10].um_I.clk ,
    \top_I.branch[22].block[9].um_I.iw[17] ,
    \top_I.branch[22].block[9].um_I.iw[16] ,
    \top_I.branch[22].block[9].um_I.iw[15] ,
    \top_I.branch[22].block[9].um_I.iw[14] ,
    \top_I.branch[22].block[9].um_I.iw[13] ,
    \top_I.branch[22].block[9].um_I.iw[12] ,
    \top_I.branch[22].block[9].um_I.iw[11] ,
    \top_I.branch[22].block[9].um_I.iw[10] ,
    \top_I.branch[22].block[9].um_I.iw[9] ,
    \top_I.branch[22].block[9].um_I.iw[8] ,
    \top_I.branch[22].block[9].um_I.iw[7] ,
    \top_I.branch[22].block[9].um_I.iw[6] ,
    \top_I.branch[22].block[9].um_I.iw[5] ,
    \top_I.branch[22].block[9].um_I.iw[4] ,
    \top_I.branch[22].block[9].um_I.iw[3] ,
    \top_I.branch[22].block[9].um_I.iw[2] ,
    \top_I.branch[22].block[9].um_I.iw[1] ,
    \top_I.branch[22].block[9].um_I.clk ,
    \top_I.branch[22].block[8].um_I.iw[17] ,
    \top_I.branch[22].block[8].um_I.iw[16] ,
    \top_I.branch[22].block[8].um_I.iw[15] ,
    \top_I.branch[22].block[8].um_I.iw[14] ,
    \top_I.branch[22].block[8].um_I.iw[13] ,
    \top_I.branch[22].block[8].um_I.iw[12] ,
    \top_I.branch[22].block[8].um_I.iw[11] ,
    \top_I.branch[22].block[8].um_I.iw[10] ,
    \top_I.branch[22].block[8].um_I.iw[9] ,
    \top_I.branch[22].block[8].um_I.iw[8] ,
    \top_I.branch[22].block[8].um_I.iw[7] ,
    \top_I.branch[22].block[8].um_I.iw[6] ,
    \top_I.branch[22].block[8].um_I.iw[5] ,
    \top_I.branch[22].block[8].um_I.iw[4] ,
    \top_I.branch[22].block[8].um_I.iw[3] ,
    \top_I.branch[22].block[8].um_I.iw[2] ,
    \top_I.branch[22].block[8].um_I.iw[1] ,
    \top_I.branch[22].block[8].um_I.clk ,
    \top_I.branch[22].block[7].um_I.iw[17] ,
    \top_I.branch[22].block[7].um_I.iw[16] ,
    \top_I.branch[22].block[7].um_I.iw[15] ,
    \top_I.branch[22].block[7].um_I.iw[14] ,
    \top_I.branch[22].block[7].um_I.iw[13] ,
    \top_I.branch[22].block[7].um_I.iw[12] ,
    \top_I.branch[22].block[7].um_I.iw[11] ,
    \top_I.branch[22].block[7].um_I.iw[10] ,
    \top_I.branch[22].block[7].um_I.iw[9] ,
    \top_I.branch[22].block[7].um_I.iw[8] ,
    \top_I.branch[22].block[7].um_I.iw[7] ,
    \top_I.branch[22].block[7].um_I.iw[6] ,
    \top_I.branch[22].block[7].um_I.iw[5] ,
    \top_I.branch[22].block[7].um_I.iw[4] ,
    \top_I.branch[22].block[7].um_I.iw[3] ,
    \top_I.branch[22].block[7].um_I.iw[2] ,
    \top_I.branch[22].block[7].um_I.iw[1] ,
    \top_I.branch[22].block[7].um_I.clk ,
    \top_I.branch[22].block[6].um_I.iw[17] ,
    \top_I.branch[22].block[6].um_I.iw[16] ,
    \top_I.branch[22].block[6].um_I.iw[15] ,
    \top_I.branch[22].block[6].um_I.iw[14] ,
    \top_I.branch[22].block[6].um_I.iw[13] ,
    \top_I.branch[22].block[6].um_I.iw[12] ,
    \top_I.branch[22].block[6].um_I.iw[11] ,
    \top_I.branch[22].block[6].um_I.iw[10] ,
    \top_I.branch[22].block[6].um_I.iw[9] ,
    \top_I.branch[22].block[6].um_I.iw[8] ,
    \top_I.branch[22].block[6].um_I.iw[7] ,
    \top_I.branch[22].block[6].um_I.iw[6] ,
    \top_I.branch[22].block[6].um_I.iw[5] ,
    \top_I.branch[22].block[6].um_I.iw[4] ,
    \top_I.branch[22].block[6].um_I.iw[3] ,
    \top_I.branch[22].block[6].um_I.iw[2] ,
    \top_I.branch[22].block[6].um_I.iw[1] ,
    \top_I.branch[22].block[6].um_I.clk ,
    \top_I.branch[22].block[5].um_I.iw[17] ,
    \top_I.branch[22].block[5].um_I.iw[16] ,
    \top_I.branch[22].block[5].um_I.iw[15] ,
    \top_I.branch[22].block[5].um_I.iw[14] ,
    \top_I.branch[22].block[5].um_I.iw[13] ,
    \top_I.branch[22].block[5].um_I.iw[12] ,
    \top_I.branch[22].block[5].um_I.iw[11] ,
    \top_I.branch[22].block[5].um_I.iw[10] ,
    \top_I.branch[22].block[5].um_I.iw[9] ,
    \top_I.branch[22].block[5].um_I.iw[8] ,
    \top_I.branch[22].block[5].um_I.iw[7] ,
    \top_I.branch[22].block[5].um_I.iw[6] ,
    \top_I.branch[22].block[5].um_I.iw[5] ,
    \top_I.branch[22].block[5].um_I.iw[4] ,
    \top_I.branch[22].block[5].um_I.iw[3] ,
    \top_I.branch[22].block[5].um_I.iw[2] ,
    \top_I.branch[22].block[5].um_I.iw[1] ,
    \top_I.branch[22].block[5].um_I.clk ,
    \top_I.branch[22].block[4].um_I.iw[17] ,
    \top_I.branch[22].block[4].um_I.iw[16] ,
    \top_I.branch[22].block[4].um_I.iw[15] ,
    \top_I.branch[22].block[4].um_I.iw[14] ,
    \top_I.branch[22].block[4].um_I.iw[13] ,
    \top_I.branch[22].block[4].um_I.iw[12] ,
    \top_I.branch[22].block[4].um_I.iw[11] ,
    \top_I.branch[22].block[4].um_I.iw[10] ,
    \top_I.branch[22].block[4].um_I.iw[9] ,
    \top_I.branch[22].block[4].um_I.iw[8] ,
    \top_I.branch[22].block[4].um_I.iw[7] ,
    \top_I.branch[22].block[4].um_I.iw[6] ,
    \top_I.branch[22].block[4].um_I.iw[5] ,
    \top_I.branch[22].block[4].um_I.iw[4] ,
    \top_I.branch[22].block[4].um_I.iw[3] ,
    \top_I.branch[22].block[4].um_I.iw[2] ,
    \top_I.branch[22].block[4].um_I.iw[1] ,
    \top_I.branch[22].block[4].um_I.clk ,
    \top_I.branch[22].block[3].um_I.iw[17] ,
    \top_I.branch[22].block[3].um_I.iw[16] ,
    \top_I.branch[22].block[3].um_I.iw[15] ,
    \top_I.branch[22].block[3].um_I.iw[14] ,
    \top_I.branch[22].block[3].um_I.iw[13] ,
    \top_I.branch[22].block[3].um_I.iw[12] ,
    \top_I.branch[22].block[3].um_I.iw[11] ,
    \top_I.branch[22].block[3].um_I.iw[10] ,
    \top_I.branch[22].block[3].um_I.iw[9] ,
    \top_I.branch[22].block[3].um_I.iw[8] ,
    \top_I.branch[22].block[3].um_I.iw[7] ,
    \top_I.branch[22].block[3].um_I.iw[6] ,
    \top_I.branch[22].block[3].um_I.iw[5] ,
    \top_I.branch[22].block[3].um_I.iw[4] ,
    \top_I.branch[22].block[3].um_I.iw[3] ,
    \top_I.branch[22].block[3].um_I.iw[2] ,
    \top_I.branch[22].block[3].um_I.iw[1] ,
    \top_I.branch[22].block[3].um_I.clk ,
    \top_I.branch[22].block[2].um_I.iw[17] ,
    \top_I.branch[22].block[2].um_I.iw[16] ,
    \top_I.branch[22].block[2].um_I.iw[15] ,
    \top_I.branch[22].block[2].um_I.iw[14] ,
    \top_I.branch[22].block[2].um_I.iw[13] ,
    \top_I.branch[22].block[2].um_I.iw[12] ,
    \top_I.branch[22].block[2].um_I.iw[11] ,
    \top_I.branch[22].block[2].um_I.iw[10] ,
    \top_I.branch[22].block[2].um_I.iw[9] ,
    \top_I.branch[22].block[2].um_I.iw[8] ,
    \top_I.branch[22].block[2].um_I.iw[7] ,
    \top_I.branch[22].block[2].um_I.iw[6] ,
    \top_I.branch[22].block[2].um_I.iw[5] ,
    \top_I.branch[22].block[2].um_I.iw[4] ,
    \top_I.branch[22].block[2].um_I.iw[3] ,
    \top_I.branch[22].block[2].um_I.iw[2] ,
    \top_I.branch[22].block[2].um_I.iw[1] ,
    \top_I.branch[22].block[2].um_I.clk ,
    \top_I.branch[22].block[1].um_I.iw[17] ,
    \top_I.branch[22].block[1].um_I.iw[16] ,
    \top_I.branch[22].block[1].um_I.iw[15] ,
    \top_I.branch[22].block[1].um_I.iw[14] ,
    \top_I.branch[22].block[1].um_I.iw[13] ,
    \top_I.branch[22].block[1].um_I.iw[12] ,
    \top_I.branch[22].block[1].um_I.iw[11] ,
    \top_I.branch[22].block[1].um_I.iw[10] ,
    \top_I.branch[22].block[1].um_I.iw[9] ,
    \top_I.branch[22].block[1].um_I.iw[8] ,
    \top_I.branch[22].block[1].um_I.iw[7] ,
    \top_I.branch[22].block[1].um_I.iw[6] ,
    \top_I.branch[22].block[1].um_I.iw[5] ,
    \top_I.branch[22].block[1].um_I.iw[4] ,
    \top_I.branch[22].block[1].um_I.iw[3] ,
    \top_I.branch[22].block[1].um_I.iw[2] ,
    \top_I.branch[22].block[1].um_I.iw[1] ,
    \top_I.branch[22].block[1].um_I.clk ,
    \top_I.branch[22].block[0].um_I.iw[17] ,
    \top_I.branch[22].block[0].um_I.iw[16] ,
    \top_I.branch[22].block[0].um_I.iw[15] ,
    \top_I.branch[22].block[0].um_I.iw[14] ,
    \top_I.branch[22].block[0].um_I.iw[13] ,
    \top_I.branch[22].block[0].um_I.iw[12] ,
    \top_I.branch[22].block[0].um_I.iw[11] ,
    \top_I.branch[22].block[0].um_I.iw[10] ,
    \top_I.branch[22].block[0].um_I.iw[9] ,
    \top_I.branch[22].block[0].um_I.iw[8] ,
    \top_I.branch[22].block[0].um_I.iw[7] ,
    \top_I.branch[22].block[0].um_I.iw[6] ,
    \top_I.branch[22].block[0].um_I.iw[5] ,
    \top_I.branch[22].block[0].um_I.iw[4] ,
    \top_I.branch[22].block[0].um_I.iw[3] ,
    \top_I.branch[22].block[0].um_I.iw[2] ,
    \top_I.branch[22].block[0].um_I.iw[1] ,
    \top_I.branch[22].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[22].block[15].um_I.pg_vdd ,
    \top_I.branch[22].block[14].um_I.pg_vdd ,
    \top_I.branch[22].block[13].um_I.pg_vdd ,
    \top_I.branch[22].block[12].um_I.pg_vdd ,
    \top_I.branch[22].block[11].um_I.pg_vdd ,
    \top_I.branch[22].block[10].um_I.pg_vdd ,
    \top_I.branch[22].block[9].um_I.pg_vdd ,
    \top_I.branch[22].block[8].um_I.pg_vdd ,
    \top_I.branch[22].block[7].um_I.pg_vdd ,
    \top_I.branch[22].block[6].um_I.pg_vdd ,
    \top_I.branch[22].block[5].um_I.pg_vdd ,
    \top_I.branch[22].block[4].um_I.pg_vdd ,
    \top_I.branch[22].block[3].um_I.pg_vdd ,
    \top_I.branch[22].block[2].um_I.pg_vdd ,
    \top_I.branch[22].block[1].um_I.pg_vdd ,
    \top_I.branch[22].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[23].mux_I  (.k_one(\top_I.branch[23].l_addr[0] ),
    .k_zero(\top_I.branch[23].l_addr[2] ),
    .addr({\top_I.branch[23].l_addr[0] ,
    \top_I.branch[23].l_addr[2] ,
    \top_I.branch[23].l_addr[0] ,
    \top_I.branch[23].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[23].block[15].um_I.ena ,
    \top_I.branch[23].block[14].um_I.ena ,
    \top_I.branch[23].block[13].um_I.ena ,
    \top_I.branch[23].block[12].um_I.ena ,
    \top_I.branch[23].block[11].um_I.ena ,
    \top_I.branch[23].block[10].um_I.ena ,
    \top_I.branch[23].block[9].um_I.ena ,
    \top_I.branch[23].block[8].um_I.ena ,
    \top_I.branch[23].block[7].um_I.ena ,
    \top_I.branch[23].block[6].um_I.ena ,
    \top_I.branch[23].block[5].um_I.ena ,
    \top_I.branch[23].block[4].um_I.ena ,
    \top_I.branch[23].block[3].um_I.ena ,
    \top_I.branch[23].block[2].um_I.ena ,
    \top_I.branch[23].block[1].um_I.ena ,
    \top_I.branch[23].block[0].um_I.ena }),
    .um_iw({\top_I.branch[23].block[15].um_I.iw[17] ,
    \top_I.branch[23].block[15].um_I.iw[16] ,
    \top_I.branch[23].block[15].um_I.iw[15] ,
    \top_I.branch[23].block[15].um_I.iw[14] ,
    \top_I.branch[23].block[15].um_I.iw[13] ,
    \top_I.branch[23].block[15].um_I.iw[12] ,
    \top_I.branch[23].block[15].um_I.iw[11] ,
    \top_I.branch[23].block[15].um_I.iw[10] ,
    \top_I.branch[23].block[15].um_I.iw[9] ,
    \top_I.branch[23].block[15].um_I.iw[8] ,
    \top_I.branch[23].block[15].um_I.iw[7] ,
    \top_I.branch[23].block[15].um_I.iw[6] ,
    \top_I.branch[23].block[15].um_I.iw[5] ,
    \top_I.branch[23].block[15].um_I.iw[4] ,
    \top_I.branch[23].block[15].um_I.iw[3] ,
    \top_I.branch[23].block[15].um_I.iw[2] ,
    \top_I.branch[23].block[15].um_I.iw[1] ,
    \top_I.branch[23].block[15].um_I.clk ,
    \top_I.branch[23].block[14].um_I.iw[17] ,
    \top_I.branch[23].block[14].um_I.iw[16] ,
    \top_I.branch[23].block[14].um_I.iw[15] ,
    \top_I.branch[23].block[14].um_I.iw[14] ,
    \top_I.branch[23].block[14].um_I.iw[13] ,
    \top_I.branch[23].block[14].um_I.iw[12] ,
    \top_I.branch[23].block[14].um_I.iw[11] ,
    \top_I.branch[23].block[14].um_I.iw[10] ,
    \top_I.branch[23].block[14].um_I.iw[9] ,
    \top_I.branch[23].block[14].um_I.iw[8] ,
    \top_I.branch[23].block[14].um_I.iw[7] ,
    \top_I.branch[23].block[14].um_I.iw[6] ,
    \top_I.branch[23].block[14].um_I.iw[5] ,
    \top_I.branch[23].block[14].um_I.iw[4] ,
    \top_I.branch[23].block[14].um_I.iw[3] ,
    \top_I.branch[23].block[14].um_I.iw[2] ,
    \top_I.branch[23].block[14].um_I.iw[1] ,
    \top_I.branch[23].block[14].um_I.clk ,
    \top_I.branch[23].block[13].um_I.iw[17] ,
    \top_I.branch[23].block[13].um_I.iw[16] ,
    \top_I.branch[23].block[13].um_I.iw[15] ,
    \top_I.branch[23].block[13].um_I.iw[14] ,
    \top_I.branch[23].block[13].um_I.iw[13] ,
    \top_I.branch[23].block[13].um_I.iw[12] ,
    \top_I.branch[23].block[13].um_I.iw[11] ,
    \top_I.branch[23].block[13].um_I.iw[10] ,
    \top_I.branch[23].block[13].um_I.iw[9] ,
    \top_I.branch[23].block[13].um_I.iw[8] ,
    \top_I.branch[23].block[13].um_I.iw[7] ,
    \top_I.branch[23].block[13].um_I.iw[6] ,
    \top_I.branch[23].block[13].um_I.iw[5] ,
    \top_I.branch[23].block[13].um_I.iw[4] ,
    \top_I.branch[23].block[13].um_I.iw[3] ,
    \top_I.branch[23].block[13].um_I.iw[2] ,
    \top_I.branch[23].block[13].um_I.iw[1] ,
    \top_I.branch[23].block[13].um_I.clk ,
    \top_I.branch[23].block[12].um_I.iw[17] ,
    \top_I.branch[23].block[12].um_I.iw[16] ,
    \top_I.branch[23].block[12].um_I.iw[15] ,
    \top_I.branch[23].block[12].um_I.iw[14] ,
    \top_I.branch[23].block[12].um_I.iw[13] ,
    \top_I.branch[23].block[12].um_I.iw[12] ,
    \top_I.branch[23].block[12].um_I.iw[11] ,
    \top_I.branch[23].block[12].um_I.iw[10] ,
    \top_I.branch[23].block[12].um_I.iw[9] ,
    \top_I.branch[23].block[12].um_I.iw[8] ,
    \top_I.branch[23].block[12].um_I.iw[7] ,
    \top_I.branch[23].block[12].um_I.iw[6] ,
    \top_I.branch[23].block[12].um_I.iw[5] ,
    \top_I.branch[23].block[12].um_I.iw[4] ,
    \top_I.branch[23].block[12].um_I.iw[3] ,
    \top_I.branch[23].block[12].um_I.iw[2] ,
    \top_I.branch[23].block[12].um_I.iw[1] ,
    \top_I.branch[23].block[12].um_I.clk ,
    \top_I.branch[23].block[11].um_I.iw[17] ,
    \top_I.branch[23].block[11].um_I.iw[16] ,
    \top_I.branch[23].block[11].um_I.iw[15] ,
    \top_I.branch[23].block[11].um_I.iw[14] ,
    \top_I.branch[23].block[11].um_I.iw[13] ,
    \top_I.branch[23].block[11].um_I.iw[12] ,
    \top_I.branch[23].block[11].um_I.iw[11] ,
    \top_I.branch[23].block[11].um_I.iw[10] ,
    \top_I.branch[23].block[11].um_I.iw[9] ,
    \top_I.branch[23].block[11].um_I.iw[8] ,
    \top_I.branch[23].block[11].um_I.iw[7] ,
    \top_I.branch[23].block[11].um_I.iw[6] ,
    \top_I.branch[23].block[11].um_I.iw[5] ,
    \top_I.branch[23].block[11].um_I.iw[4] ,
    \top_I.branch[23].block[11].um_I.iw[3] ,
    \top_I.branch[23].block[11].um_I.iw[2] ,
    \top_I.branch[23].block[11].um_I.iw[1] ,
    \top_I.branch[23].block[11].um_I.clk ,
    \top_I.branch[23].block[10].um_I.iw[17] ,
    \top_I.branch[23].block[10].um_I.iw[16] ,
    \top_I.branch[23].block[10].um_I.iw[15] ,
    \top_I.branch[23].block[10].um_I.iw[14] ,
    \top_I.branch[23].block[10].um_I.iw[13] ,
    \top_I.branch[23].block[10].um_I.iw[12] ,
    \top_I.branch[23].block[10].um_I.iw[11] ,
    \top_I.branch[23].block[10].um_I.iw[10] ,
    \top_I.branch[23].block[10].um_I.iw[9] ,
    \top_I.branch[23].block[10].um_I.iw[8] ,
    \top_I.branch[23].block[10].um_I.iw[7] ,
    \top_I.branch[23].block[10].um_I.iw[6] ,
    \top_I.branch[23].block[10].um_I.iw[5] ,
    \top_I.branch[23].block[10].um_I.iw[4] ,
    \top_I.branch[23].block[10].um_I.iw[3] ,
    \top_I.branch[23].block[10].um_I.iw[2] ,
    \top_I.branch[23].block[10].um_I.iw[1] ,
    \top_I.branch[23].block[10].um_I.clk ,
    \top_I.branch[23].block[9].um_I.iw[17] ,
    \top_I.branch[23].block[9].um_I.iw[16] ,
    \top_I.branch[23].block[9].um_I.iw[15] ,
    \top_I.branch[23].block[9].um_I.iw[14] ,
    \top_I.branch[23].block[9].um_I.iw[13] ,
    \top_I.branch[23].block[9].um_I.iw[12] ,
    \top_I.branch[23].block[9].um_I.iw[11] ,
    \top_I.branch[23].block[9].um_I.iw[10] ,
    \top_I.branch[23].block[9].um_I.iw[9] ,
    \top_I.branch[23].block[9].um_I.iw[8] ,
    \top_I.branch[23].block[9].um_I.iw[7] ,
    \top_I.branch[23].block[9].um_I.iw[6] ,
    \top_I.branch[23].block[9].um_I.iw[5] ,
    \top_I.branch[23].block[9].um_I.iw[4] ,
    \top_I.branch[23].block[9].um_I.iw[3] ,
    \top_I.branch[23].block[9].um_I.iw[2] ,
    \top_I.branch[23].block[9].um_I.iw[1] ,
    \top_I.branch[23].block[9].um_I.clk ,
    \top_I.branch[23].block[8].um_I.iw[17] ,
    \top_I.branch[23].block[8].um_I.iw[16] ,
    \top_I.branch[23].block[8].um_I.iw[15] ,
    \top_I.branch[23].block[8].um_I.iw[14] ,
    \top_I.branch[23].block[8].um_I.iw[13] ,
    \top_I.branch[23].block[8].um_I.iw[12] ,
    \top_I.branch[23].block[8].um_I.iw[11] ,
    \top_I.branch[23].block[8].um_I.iw[10] ,
    \top_I.branch[23].block[8].um_I.iw[9] ,
    \top_I.branch[23].block[8].um_I.iw[8] ,
    \top_I.branch[23].block[8].um_I.iw[7] ,
    \top_I.branch[23].block[8].um_I.iw[6] ,
    \top_I.branch[23].block[8].um_I.iw[5] ,
    \top_I.branch[23].block[8].um_I.iw[4] ,
    \top_I.branch[23].block[8].um_I.iw[3] ,
    \top_I.branch[23].block[8].um_I.iw[2] ,
    \top_I.branch[23].block[8].um_I.iw[1] ,
    \top_I.branch[23].block[8].um_I.clk ,
    \top_I.branch[23].block[7].um_I.iw[17] ,
    \top_I.branch[23].block[7].um_I.iw[16] ,
    \top_I.branch[23].block[7].um_I.iw[15] ,
    \top_I.branch[23].block[7].um_I.iw[14] ,
    \top_I.branch[23].block[7].um_I.iw[13] ,
    \top_I.branch[23].block[7].um_I.iw[12] ,
    \top_I.branch[23].block[7].um_I.iw[11] ,
    \top_I.branch[23].block[7].um_I.iw[10] ,
    \top_I.branch[23].block[7].um_I.iw[9] ,
    \top_I.branch[23].block[7].um_I.iw[8] ,
    \top_I.branch[23].block[7].um_I.iw[7] ,
    \top_I.branch[23].block[7].um_I.iw[6] ,
    \top_I.branch[23].block[7].um_I.iw[5] ,
    \top_I.branch[23].block[7].um_I.iw[4] ,
    \top_I.branch[23].block[7].um_I.iw[3] ,
    \top_I.branch[23].block[7].um_I.iw[2] ,
    \top_I.branch[23].block[7].um_I.iw[1] ,
    \top_I.branch[23].block[7].um_I.clk ,
    \top_I.branch[23].block[6].um_I.iw[17] ,
    \top_I.branch[23].block[6].um_I.iw[16] ,
    \top_I.branch[23].block[6].um_I.iw[15] ,
    \top_I.branch[23].block[6].um_I.iw[14] ,
    \top_I.branch[23].block[6].um_I.iw[13] ,
    \top_I.branch[23].block[6].um_I.iw[12] ,
    \top_I.branch[23].block[6].um_I.iw[11] ,
    \top_I.branch[23].block[6].um_I.iw[10] ,
    \top_I.branch[23].block[6].um_I.iw[9] ,
    \top_I.branch[23].block[6].um_I.iw[8] ,
    \top_I.branch[23].block[6].um_I.iw[7] ,
    \top_I.branch[23].block[6].um_I.iw[6] ,
    \top_I.branch[23].block[6].um_I.iw[5] ,
    \top_I.branch[23].block[6].um_I.iw[4] ,
    \top_I.branch[23].block[6].um_I.iw[3] ,
    \top_I.branch[23].block[6].um_I.iw[2] ,
    \top_I.branch[23].block[6].um_I.iw[1] ,
    \top_I.branch[23].block[6].um_I.clk ,
    \top_I.branch[23].block[5].um_I.iw[17] ,
    \top_I.branch[23].block[5].um_I.iw[16] ,
    \top_I.branch[23].block[5].um_I.iw[15] ,
    \top_I.branch[23].block[5].um_I.iw[14] ,
    \top_I.branch[23].block[5].um_I.iw[13] ,
    \top_I.branch[23].block[5].um_I.iw[12] ,
    \top_I.branch[23].block[5].um_I.iw[11] ,
    \top_I.branch[23].block[5].um_I.iw[10] ,
    \top_I.branch[23].block[5].um_I.iw[9] ,
    \top_I.branch[23].block[5].um_I.iw[8] ,
    \top_I.branch[23].block[5].um_I.iw[7] ,
    \top_I.branch[23].block[5].um_I.iw[6] ,
    \top_I.branch[23].block[5].um_I.iw[5] ,
    \top_I.branch[23].block[5].um_I.iw[4] ,
    \top_I.branch[23].block[5].um_I.iw[3] ,
    \top_I.branch[23].block[5].um_I.iw[2] ,
    \top_I.branch[23].block[5].um_I.iw[1] ,
    \top_I.branch[23].block[5].um_I.clk ,
    \top_I.branch[23].block[4].um_I.iw[17] ,
    \top_I.branch[23].block[4].um_I.iw[16] ,
    \top_I.branch[23].block[4].um_I.iw[15] ,
    \top_I.branch[23].block[4].um_I.iw[14] ,
    \top_I.branch[23].block[4].um_I.iw[13] ,
    \top_I.branch[23].block[4].um_I.iw[12] ,
    \top_I.branch[23].block[4].um_I.iw[11] ,
    \top_I.branch[23].block[4].um_I.iw[10] ,
    \top_I.branch[23].block[4].um_I.iw[9] ,
    \top_I.branch[23].block[4].um_I.iw[8] ,
    \top_I.branch[23].block[4].um_I.iw[7] ,
    \top_I.branch[23].block[4].um_I.iw[6] ,
    \top_I.branch[23].block[4].um_I.iw[5] ,
    \top_I.branch[23].block[4].um_I.iw[4] ,
    \top_I.branch[23].block[4].um_I.iw[3] ,
    \top_I.branch[23].block[4].um_I.iw[2] ,
    \top_I.branch[23].block[4].um_I.iw[1] ,
    \top_I.branch[23].block[4].um_I.clk ,
    \top_I.branch[23].block[3].um_I.iw[17] ,
    \top_I.branch[23].block[3].um_I.iw[16] ,
    \top_I.branch[23].block[3].um_I.iw[15] ,
    \top_I.branch[23].block[3].um_I.iw[14] ,
    \top_I.branch[23].block[3].um_I.iw[13] ,
    \top_I.branch[23].block[3].um_I.iw[12] ,
    \top_I.branch[23].block[3].um_I.iw[11] ,
    \top_I.branch[23].block[3].um_I.iw[10] ,
    \top_I.branch[23].block[3].um_I.iw[9] ,
    \top_I.branch[23].block[3].um_I.iw[8] ,
    \top_I.branch[23].block[3].um_I.iw[7] ,
    \top_I.branch[23].block[3].um_I.iw[6] ,
    \top_I.branch[23].block[3].um_I.iw[5] ,
    \top_I.branch[23].block[3].um_I.iw[4] ,
    \top_I.branch[23].block[3].um_I.iw[3] ,
    \top_I.branch[23].block[3].um_I.iw[2] ,
    \top_I.branch[23].block[3].um_I.iw[1] ,
    \top_I.branch[23].block[3].um_I.clk ,
    \top_I.branch[23].block[2].um_I.iw[17] ,
    \top_I.branch[23].block[2].um_I.iw[16] ,
    \top_I.branch[23].block[2].um_I.iw[15] ,
    \top_I.branch[23].block[2].um_I.iw[14] ,
    \top_I.branch[23].block[2].um_I.iw[13] ,
    \top_I.branch[23].block[2].um_I.iw[12] ,
    \top_I.branch[23].block[2].um_I.iw[11] ,
    \top_I.branch[23].block[2].um_I.iw[10] ,
    \top_I.branch[23].block[2].um_I.iw[9] ,
    \top_I.branch[23].block[2].um_I.iw[8] ,
    \top_I.branch[23].block[2].um_I.iw[7] ,
    \top_I.branch[23].block[2].um_I.iw[6] ,
    \top_I.branch[23].block[2].um_I.iw[5] ,
    \top_I.branch[23].block[2].um_I.iw[4] ,
    \top_I.branch[23].block[2].um_I.iw[3] ,
    \top_I.branch[23].block[2].um_I.iw[2] ,
    \top_I.branch[23].block[2].um_I.iw[1] ,
    \top_I.branch[23].block[2].um_I.clk ,
    \top_I.branch[23].block[1].um_I.iw[17] ,
    \top_I.branch[23].block[1].um_I.iw[16] ,
    \top_I.branch[23].block[1].um_I.iw[15] ,
    \top_I.branch[23].block[1].um_I.iw[14] ,
    \top_I.branch[23].block[1].um_I.iw[13] ,
    \top_I.branch[23].block[1].um_I.iw[12] ,
    \top_I.branch[23].block[1].um_I.iw[11] ,
    \top_I.branch[23].block[1].um_I.iw[10] ,
    \top_I.branch[23].block[1].um_I.iw[9] ,
    \top_I.branch[23].block[1].um_I.iw[8] ,
    \top_I.branch[23].block[1].um_I.iw[7] ,
    \top_I.branch[23].block[1].um_I.iw[6] ,
    \top_I.branch[23].block[1].um_I.iw[5] ,
    \top_I.branch[23].block[1].um_I.iw[4] ,
    \top_I.branch[23].block[1].um_I.iw[3] ,
    \top_I.branch[23].block[1].um_I.iw[2] ,
    \top_I.branch[23].block[1].um_I.iw[1] ,
    \top_I.branch[23].block[1].um_I.clk ,
    \top_I.branch[23].block[0].um_I.iw[17] ,
    \top_I.branch[23].block[0].um_I.iw[16] ,
    \top_I.branch[23].block[0].um_I.iw[15] ,
    \top_I.branch[23].block[0].um_I.iw[14] ,
    \top_I.branch[23].block[0].um_I.iw[13] ,
    \top_I.branch[23].block[0].um_I.iw[12] ,
    \top_I.branch[23].block[0].um_I.iw[11] ,
    \top_I.branch[23].block[0].um_I.iw[10] ,
    \top_I.branch[23].block[0].um_I.iw[9] ,
    \top_I.branch[23].block[0].um_I.iw[8] ,
    \top_I.branch[23].block[0].um_I.iw[7] ,
    \top_I.branch[23].block[0].um_I.iw[6] ,
    \top_I.branch[23].block[0].um_I.iw[5] ,
    \top_I.branch[23].block[0].um_I.iw[4] ,
    \top_I.branch[23].block[0].um_I.iw[3] ,
    \top_I.branch[23].block[0].um_I.iw[2] ,
    \top_I.branch[23].block[0].um_I.iw[1] ,
    \top_I.branch[23].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[23].block[15].um_I.pg_vdd ,
    \top_I.branch[23].block[14].um_I.pg_vdd ,
    \top_I.branch[23].block[13].um_I.pg_vdd ,
    \top_I.branch[23].block[12].um_I.pg_vdd ,
    \top_I.branch[23].block[11].um_I.pg_vdd ,
    \top_I.branch[23].block[10].um_I.pg_vdd ,
    \top_I.branch[23].block[9].um_I.pg_vdd ,
    \top_I.branch[23].block[8].um_I.pg_vdd ,
    \top_I.branch[23].block[7].um_I.pg_vdd ,
    \top_I.branch[23].block[6].um_I.pg_vdd ,
    \top_I.branch[23].block[5].um_I.pg_vdd ,
    \top_I.branch[23].block[4].um_I.pg_vdd ,
    \top_I.branch[23].block[3].um_I.pg_vdd ,
    \top_I.branch[23].block[2].um_I.pg_vdd ,
    \top_I.branch[23].block[1].um_I.pg_vdd ,
    \top_I.branch[23].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[2].mux_I  (.k_one(\top_I.branch[2].l_addr[0] ),
    .k_zero(\top_I.branch[2].l_addr[1] ),
    .addr({\top_I.branch[2].l_addr[1] ,
    \top_I.branch[2].l_addr[1] ,
    \top_I.branch[2].l_addr[1] ,
    \top_I.branch[2].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[2].block[15].um_I.ena ,
    \top_I.branch[2].block[14].um_I.ena ,
    \top_I.branch[2].block[13].um_I.ena ,
    \top_I.branch[2].block[12].um_I.ena ,
    \top_I.branch[2].block[11].um_I.ena ,
    \top_I.branch[2].block[10].um_I.ena ,
    \top_I.branch[2].block[9].um_I.ena ,
    \top_I.branch[2].block[8].um_I.ena ,
    \top_I.branch[2].block[7].um_I.ena ,
    \top_I.branch[2].block[6].um_I.ena ,
    \top_I.branch[2].block[5].um_I.ena ,
    \top_I.branch[2].block[4].um_I.ena ,
    \top_I.branch[2].block[3].um_I.ena ,
    \top_I.branch[2].block[2].um_I.ena ,
    \top_I.branch[2].block[1].um_I.ena ,
    \top_I.branch[2].block[0].um_I.ena }),
    .um_iw({\top_I.branch[2].block[15].um_I.iw[17] ,
    \top_I.branch[2].block[15].um_I.iw[16] ,
    \top_I.branch[2].block[15].um_I.iw[15] ,
    \top_I.branch[2].block[15].um_I.iw[14] ,
    \top_I.branch[2].block[15].um_I.iw[13] ,
    \top_I.branch[2].block[15].um_I.iw[12] ,
    \top_I.branch[2].block[15].um_I.iw[11] ,
    \top_I.branch[2].block[15].um_I.iw[10] ,
    \top_I.branch[2].block[15].um_I.iw[9] ,
    \top_I.branch[2].block[15].um_I.iw[8] ,
    \top_I.branch[2].block[15].um_I.iw[7] ,
    \top_I.branch[2].block[15].um_I.iw[6] ,
    \top_I.branch[2].block[15].um_I.iw[5] ,
    \top_I.branch[2].block[15].um_I.iw[4] ,
    \top_I.branch[2].block[15].um_I.iw[3] ,
    \top_I.branch[2].block[15].um_I.iw[2] ,
    \top_I.branch[2].block[15].um_I.iw[1] ,
    \top_I.branch[2].block[15].um_I.clk ,
    \top_I.branch[2].block[14].um_I.iw[17] ,
    \top_I.branch[2].block[14].um_I.iw[16] ,
    \top_I.branch[2].block[14].um_I.iw[15] ,
    \top_I.branch[2].block[14].um_I.iw[14] ,
    \top_I.branch[2].block[14].um_I.iw[13] ,
    \top_I.branch[2].block[14].um_I.iw[12] ,
    \top_I.branch[2].block[14].um_I.iw[11] ,
    \top_I.branch[2].block[14].um_I.iw[10] ,
    \top_I.branch[2].block[14].um_I.iw[9] ,
    \top_I.branch[2].block[14].um_I.iw[8] ,
    \top_I.branch[2].block[14].um_I.iw[7] ,
    \top_I.branch[2].block[14].um_I.iw[6] ,
    \top_I.branch[2].block[14].um_I.iw[5] ,
    \top_I.branch[2].block[14].um_I.iw[4] ,
    \top_I.branch[2].block[14].um_I.iw[3] ,
    \top_I.branch[2].block[14].um_I.iw[2] ,
    \top_I.branch[2].block[14].um_I.iw[1] ,
    \top_I.branch[2].block[14].um_I.clk ,
    \top_I.branch[2].block[13].um_I.iw[17] ,
    \top_I.branch[2].block[13].um_I.iw[16] ,
    \top_I.branch[2].block[13].um_I.iw[15] ,
    \top_I.branch[2].block[13].um_I.iw[14] ,
    \top_I.branch[2].block[13].um_I.iw[13] ,
    \top_I.branch[2].block[13].um_I.iw[12] ,
    \top_I.branch[2].block[13].um_I.iw[11] ,
    \top_I.branch[2].block[13].um_I.iw[10] ,
    \top_I.branch[2].block[13].um_I.iw[9] ,
    \top_I.branch[2].block[13].um_I.iw[8] ,
    \top_I.branch[2].block[13].um_I.iw[7] ,
    \top_I.branch[2].block[13].um_I.iw[6] ,
    \top_I.branch[2].block[13].um_I.iw[5] ,
    \top_I.branch[2].block[13].um_I.iw[4] ,
    \top_I.branch[2].block[13].um_I.iw[3] ,
    \top_I.branch[2].block[13].um_I.iw[2] ,
    \top_I.branch[2].block[13].um_I.iw[1] ,
    \top_I.branch[2].block[13].um_I.clk ,
    \top_I.branch[2].block[12].um_I.iw[17] ,
    \top_I.branch[2].block[12].um_I.iw[16] ,
    \top_I.branch[2].block[12].um_I.iw[15] ,
    \top_I.branch[2].block[12].um_I.iw[14] ,
    \top_I.branch[2].block[12].um_I.iw[13] ,
    \top_I.branch[2].block[12].um_I.iw[12] ,
    \top_I.branch[2].block[12].um_I.iw[11] ,
    \top_I.branch[2].block[12].um_I.iw[10] ,
    \top_I.branch[2].block[12].um_I.iw[9] ,
    \top_I.branch[2].block[12].um_I.iw[8] ,
    \top_I.branch[2].block[12].um_I.iw[7] ,
    \top_I.branch[2].block[12].um_I.iw[6] ,
    \top_I.branch[2].block[12].um_I.iw[5] ,
    \top_I.branch[2].block[12].um_I.iw[4] ,
    \top_I.branch[2].block[12].um_I.iw[3] ,
    \top_I.branch[2].block[12].um_I.iw[2] ,
    \top_I.branch[2].block[12].um_I.iw[1] ,
    \top_I.branch[2].block[12].um_I.clk ,
    \top_I.branch[2].block[11].um_I.iw[17] ,
    \top_I.branch[2].block[11].um_I.iw[16] ,
    \top_I.branch[2].block[11].um_I.iw[15] ,
    \top_I.branch[2].block[11].um_I.iw[14] ,
    \top_I.branch[2].block[11].um_I.iw[13] ,
    \top_I.branch[2].block[11].um_I.iw[12] ,
    \top_I.branch[2].block[11].um_I.iw[11] ,
    \top_I.branch[2].block[11].um_I.iw[10] ,
    \top_I.branch[2].block[11].um_I.iw[9] ,
    \top_I.branch[2].block[11].um_I.iw[8] ,
    \top_I.branch[2].block[11].um_I.iw[7] ,
    \top_I.branch[2].block[11].um_I.iw[6] ,
    \top_I.branch[2].block[11].um_I.iw[5] ,
    \top_I.branch[2].block[11].um_I.iw[4] ,
    \top_I.branch[2].block[11].um_I.iw[3] ,
    \top_I.branch[2].block[11].um_I.iw[2] ,
    \top_I.branch[2].block[11].um_I.iw[1] ,
    \top_I.branch[2].block[11].um_I.clk ,
    \top_I.branch[2].block[10].um_I.iw[17] ,
    \top_I.branch[2].block[10].um_I.iw[16] ,
    \top_I.branch[2].block[10].um_I.iw[15] ,
    \top_I.branch[2].block[10].um_I.iw[14] ,
    \top_I.branch[2].block[10].um_I.iw[13] ,
    \top_I.branch[2].block[10].um_I.iw[12] ,
    \top_I.branch[2].block[10].um_I.iw[11] ,
    \top_I.branch[2].block[10].um_I.iw[10] ,
    \top_I.branch[2].block[10].um_I.iw[9] ,
    \top_I.branch[2].block[10].um_I.iw[8] ,
    \top_I.branch[2].block[10].um_I.iw[7] ,
    \top_I.branch[2].block[10].um_I.iw[6] ,
    \top_I.branch[2].block[10].um_I.iw[5] ,
    \top_I.branch[2].block[10].um_I.iw[4] ,
    \top_I.branch[2].block[10].um_I.iw[3] ,
    \top_I.branch[2].block[10].um_I.iw[2] ,
    \top_I.branch[2].block[10].um_I.iw[1] ,
    \top_I.branch[2].block[10].um_I.clk ,
    \top_I.branch[2].block[9].um_I.iw[17] ,
    \top_I.branch[2].block[9].um_I.iw[16] ,
    \top_I.branch[2].block[9].um_I.iw[15] ,
    \top_I.branch[2].block[9].um_I.iw[14] ,
    \top_I.branch[2].block[9].um_I.iw[13] ,
    \top_I.branch[2].block[9].um_I.iw[12] ,
    \top_I.branch[2].block[9].um_I.iw[11] ,
    \top_I.branch[2].block[9].um_I.iw[10] ,
    \top_I.branch[2].block[9].um_I.iw[9] ,
    \top_I.branch[2].block[9].um_I.iw[8] ,
    \top_I.branch[2].block[9].um_I.iw[7] ,
    \top_I.branch[2].block[9].um_I.iw[6] ,
    \top_I.branch[2].block[9].um_I.iw[5] ,
    \top_I.branch[2].block[9].um_I.iw[4] ,
    \top_I.branch[2].block[9].um_I.iw[3] ,
    \top_I.branch[2].block[9].um_I.iw[2] ,
    \top_I.branch[2].block[9].um_I.iw[1] ,
    \top_I.branch[2].block[9].um_I.clk ,
    \top_I.branch[2].block[8].um_I.iw[17] ,
    \top_I.branch[2].block[8].um_I.iw[16] ,
    \top_I.branch[2].block[8].um_I.iw[15] ,
    \top_I.branch[2].block[8].um_I.iw[14] ,
    \top_I.branch[2].block[8].um_I.iw[13] ,
    \top_I.branch[2].block[8].um_I.iw[12] ,
    \top_I.branch[2].block[8].um_I.iw[11] ,
    \top_I.branch[2].block[8].um_I.iw[10] ,
    \top_I.branch[2].block[8].um_I.iw[9] ,
    \top_I.branch[2].block[8].um_I.iw[8] ,
    \top_I.branch[2].block[8].um_I.iw[7] ,
    \top_I.branch[2].block[8].um_I.iw[6] ,
    \top_I.branch[2].block[8].um_I.iw[5] ,
    \top_I.branch[2].block[8].um_I.iw[4] ,
    \top_I.branch[2].block[8].um_I.iw[3] ,
    \top_I.branch[2].block[8].um_I.iw[2] ,
    \top_I.branch[2].block[8].um_I.iw[1] ,
    \top_I.branch[2].block[8].um_I.clk ,
    \top_I.branch[2].block[7].um_I.iw[17] ,
    \top_I.branch[2].block[7].um_I.iw[16] ,
    \top_I.branch[2].block[7].um_I.iw[15] ,
    \top_I.branch[2].block[7].um_I.iw[14] ,
    \top_I.branch[2].block[7].um_I.iw[13] ,
    \top_I.branch[2].block[7].um_I.iw[12] ,
    \top_I.branch[2].block[7].um_I.iw[11] ,
    \top_I.branch[2].block[7].um_I.iw[10] ,
    \top_I.branch[2].block[7].um_I.iw[9] ,
    \top_I.branch[2].block[7].um_I.iw[8] ,
    \top_I.branch[2].block[7].um_I.iw[7] ,
    \top_I.branch[2].block[7].um_I.iw[6] ,
    \top_I.branch[2].block[7].um_I.iw[5] ,
    \top_I.branch[2].block[7].um_I.iw[4] ,
    \top_I.branch[2].block[7].um_I.iw[3] ,
    \top_I.branch[2].block[7].um_I.iw[2] ,
    \top_I.branch[2].block[7].um_I.iw[1] ,
    \top_I.branch[2].block[7].um_I.clk ,
    \top_I.branch[2].block[6].um_I.iw[17] ,
    \top_I.branch[2].block[6].um_I.iw[16] ,
    \top_I.branch[2].block[6].um_I.iw[15] ,
    \top_I.branch[2].block[6].um_I.iw[14] ,
    \top_I.branch[2].block[6].um_I.iw[13] ,
    \top_I.branch[2].block[6].um_I.iw[12] ,
    \top_I.branch[2].block[6].um_I.iw[11] ,
    \top_I.branch[2].block[6].um_I.iw[10] ,
    \top_I.branch[2].block[6].um_I.iw[9] ,
    \top_I.branch[2].block[6].um_I.iw[8] ,
    \top_I.branch[2].block[6].um_I.iw[7] ,
    \top_I.branch[2].block[6].um_I.iw[6] ,
    \top_I.branch[2].block[6].um_I.iw[5] ,
    \top_I.branch[2].block[6].um_I.iw[4] ,
    \top_I.branch[2].block[6].um_I.iw[3] ,
    \top_I.branch[2].block[6].um_I.iw[2] ,
    \top_I.branch[2].block[6].um_I.iw[1] ,
    \top_I.branch[2].block[6].um_I.clk ,
    \top_I.branch[2].block[5].um_I.iw[17] ,
    \top_I.branch[2].block[5].um_I.iw[16] ,
    \top_I.branch[2].block[5].um_I.iw[15] ,
    \top_I.branch[2].block[5].um_I.iw[14] ,
    \top_I.branch[2].block[5].um_I.iw[13] ,
    \top_I.branch[2].block[5].um_I.iw[12] ,
    \top_I.branch[2].block[5].um_I.iw[11] ,
    \top_I.branch[2].block[5].um_I.iw[10] ,
    \top_I.branch[2].block[5].um_I.iw[9] ,
    \top_I.branch[2].block[5].um_I.iw[8] ,
    \top_I.branch[2].block[5].um_I.iw[7] ,
    \top_I.branch[2].block[5].um_I.iw[6] ,
    \top_I.branch[2].block[5].um_I.iw[5] ,
    \top_I.branch[2].block[5].um_I.iw[4] ,
    \top_I.branch[2].block[5].um_I.iw[3] ,
    \top_I.branch[2].block[5].um_I.iw[2] ,
    \top_I.branch[2].block[5].um_I.iw[1] ,
    \top_I.branch[2].block[5].um_I.clk ,
    \top_I.branch[2].block[4].um_I.iw[17] ,
    \top_I.branch[2].block[4].um_I.iw[16] ,
    \top_I.branch[2].block[4].um_I.iw[15] ,
    \top_I.branch[2].block[4].um_I.iw[14] ,
    \top_I.branch[2].block[4].um_I.iw[13] ,
    \top_I.branch[2].block[4].um_I.iw[12] ,
    \top_I.branch[2].block[4].um_I.iw[11] ,
    \top_I.branch[2].block[4].um_I.iw[10] ,
    \top_I.branch[2].block[4].um_I.iw[9] ,
    \top_I.branch[2].block[4].um_I.iw[8] ,
    \top_I.branch[2].block[4].um_I.iw[7] ,
    \top_I.branch[2].block[4].um_I.iw[6] ,
    \top_I.branch[2].block[4].um_I.iw[5] ,
    \top_I.branch[2].block[4].um_I.iw[4] ,
    \top_I.branch[2].block[4].um_I.iw[3] ,
    \top_I.branch[2].block[4].um_I.iw[2] ,
    \top_I.branch[2].block[4].um_I.iw[1] ,
    \top_I.branch[2].block[4].um_I.clk ,
    \top_I.branch[2].block[3].um_I.iw[17] ,
    \top_I.branch[2].block[3].um_I.iw[16] ,
    \top_I.branch[2].block[3].um_I.iw[15] ,
    \top_I.branch[2].block[3].um_I.iw[14] ,
    \top_I.branch[2].block[3].um_I.iw[13] ,
    \top_I.branch[2].block[3].um_I.iw[12] ,
    \top_I.branch[2].block[3].um_I.iw[11] ,
    \top_I.branch[2].block[3].um_I.iw[10] ,
    \top_I.branch[2].block[3].um_I.iw[9] ,
    \top_I.branch[2].block[3].um_I.iw[8] ,
    \top_I.branch[2].block[3].um_I.iw[7] ,
    \top_I.branch[2].block[3].um_I.iw[6] ,
    \top_I.branch[2].block[3].um_I.iw[5] ,
    \top_I.branch[2].block[3].um_I.iw[4] ,
    \top_I.branch[2].block[3].um_I.iw[3] ,
    \top_I.branch[2].block[3].um_I.iw[2] ,
    \top_I.branch[2].block[3].um_I.iw[1] ,
    \top_I.branch[2].block[3].um_I.clk ,
    \top_I.branch[2].block[2].um_I.iw[17] ,
    \top_I.branch[2].block[2].um_I.iw[16] ,
    \top_I.branch[2].block[2].um_I.iw[15] ,
    \top_I.branch[2].block[2].um_I.iw[14] ,
    \top_I.branch[2].block[2].um_I.iw[13] ,
    \top_I.branch[2].block[2].um_I.iw[12] ,
    \top_I.branch[2].block[2].um_I.iw[11] ,
    \top_I.branch[2].block[2].um_I.iw[10] ,
    \top_I.branch[2].block[2].um_I.iw[9] ,
    \top_I.branch[2].block[2].um_I.iw[8] ,
    \top_I.branch[2].block[2].um_I.iw[7] ,
    \top_I.branch[2].block[2].um_I.iw[6] ,
    \top_I.branch[2].block[2].um_I.iw[5] ,
    \top_I.branch[2].block[2].um_I.iw[4] ,
    \top_I.branch[2].block[2].um_I.iw[3] ,
    \top_I.branch[2].block[2].um_I.iw[2] ,
    \top_I.branch[2].block[2].um_I.iw[1] ,
    \top_I.branch[2].block[2].um_I.clk ,
    \top_I.branch[2].block[1].um_I.iw[17] ,
    \top_I.branch[2].block[1].um_I.iw[16] ,
    \top_I.branch[2].block[1].um_I.iw[15] ,
    \top_I.branch[2].block[1].um_I.iw[14] ,
    \top_I.branch[2].block[1].um_I.iw[13] ,
    \top_I.branch[2].block[1].um_I.iw[12] ,
    \top_I.branch[2].block[1].um_I.iw[11] ,
    \top_I.branch[2].block[1].um_I.iw[10] ,
    \top_I.branch[2].block[1].um_I.iw[9] ,
    \top_I.branch[2].block[1].um_I.iw[8] ,
    \top_I.branch[2].block[1].um_I.iw[7] ,
    \top_I.branch[2].block[1].um_I.iw[6] ,
    \top_I.branch[2].block[1].um_I.iw[5] ,
    \top_I.branch[2].block[1].um_I.iw[4] ,
    \top_I.branch[2].block[1].um_I.iw[3] ,
    \top_I.branch[2].block[1].um_I.iw[2] ,
    \top_I.branch[2].block[1].um_I.iw[1] ,
    \top_I.branch[2].block[1].um_I.clk ,
    \top_I.branch[2].block[0].um_I.iw[17] ,
    \top_I.branch[2].block[0].um_I.iw[16] ,
    \top_I.branch[2].block[0].um_I.iw[15] ,
    \top_I.branch[2].block[0].um_I.iw[14] ,
    \top_I.branch[2].block[0].um_I.iw[13] ,
    \top_I.branch[2].block[0].um_I.iw[12] ,
    \top_I.branch[2].block[0].um_I.iw[11] ,
    \top_I.branch[2].block[0].um_I.iw[10] ,
    \top_I.branch[2].block[0].um_I.iw[9] ,
    \top_I.branch[2].block[0].um_I.iw[8] ,
    \top_I.branch[2].block[0].um_I.iw[7] ,
    \top_I.branch[2].block[0].um_I.iw[6] ,
    \top_I.branch[2].block[0].um_I.iw[5] ,
    \top_I.branch[2].block[0].um_I.iw[4] ,
    \top_I.branch[2].block[0].um_I.iw[3] ,
    \top_I.branch[2].block[0].um_I.iw[2] ,
    \top_I.branch[2].block[0].um_I.iw[1] ,
    \top_I.branch[2].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[2].block[15].um_I.pg_vdd ,
    \top_I.branch[2].block[14].um_I.pg_vdd ,
    \top_I.branch[2].block[13].um_I.pg_vdd ,
    \top_I.branch[2].block[12].um_I.pg_vdd ,
    \top_I.branch[2].block[11].um_I.pg_vdd ,
    \top_I.branch[2].block[10].um_I.pg_vdd ,
    \top_I.branch[2].block[9].um_I.pg_vdd ,
    \top_I.branch[2].block[8].um_I.pg_vdd ,
    \top_I.branch[2].block[7].um_I.pg_vdd ,
    \top_I.branch[2].block[6].um_I.pg_vdd ,
    \top_I.branch[2].block[5].um_I.pg_vdd ,
    \top_I.branch[2].block[4].um_I.pg_vdd ,
    \top_I.branch[2].block[3].um_I.pg_vdd ,
    \top_I.branch[2].block[2].um_I.pg_vdd ,
    \top_I.branch[2].block[1].um_I.pg_vdd ,
    \top_I.branch[2].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[3].mux_I  (.k_one(\top_I.branch[3].l_addr[0] ),
    .k_zero(\top_I.branch[3].l_addr[1] ),
    .addr({\top_I.branch[3].l_addr[1] ,
    \top_I.branch[3].l_addr[1] ,
    \top_I.branch[3].l_addr[1] ,
    \top_I.branch[3].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[3].block[15].um_I.ena ,
    \top_I.branch[3].block[14].um_I.ena ,
    \top_I.branch[3].block[13].um_I.ena ,
    \top_I.branch[3].block[12].um_I.ena ,
    \top_I.branch[3].block[11].um_I.ena ,
    \top_I.branch[3].block[10].um_I.ena ,
    \top_I.branch[3].block[9].um_I.ena ,
    \top_I.branch[3].block[8].um_I.ena ,
    \top_I.branch[3].block[7].um_I.ena ,
    \top_I.branch[3].block[6].um_I.ena ,
    \top_I.branch[3].block[5].um_I.ena ,
    \top_I.branch[3].block[4].um_I.ena ,
    \top_I.branch[3].block[3].um_I.ena ,
    \top_I.branch[3].block[2].um_I.ena ,
    \top_I.branch[3].block[1].um_I.ena ,
    \top_I.branch[3].block[0].um_I.ena }),
    .um_iw({\top_I.branch[3].block[15].um_I.iw[17] ,
    \top_I.branch[3].block[15].um_I.iw[16] ,
    \top_I.branch[3].block[15].um_I.iw[15] ,
    \top_I.branch[3].block[15].um_I.iw[14] ,
    \top_I.branch[3].block[15].um_I.iw[13] ,
    \top_I.branch[3].block[15].um_I.iw[12] ,
    \top_I.branch[3].block[15].um_I.iw[11] ,
    \top_I.branch[3].block[15].um_I.iw[10] ,
    \top_I.branch[3].block[15].um_I.iw[9] ,
    \top_I.branch[3].block[15].um_I.iw[8] ,
    \top_I.branch[3].block[15].um_I.iw[7] ,
    \top_I.branch[3].block[15].um_I.iw[6] ,
    \top_I.branch[3].block[15].um_I.iw[5] ,
    \top_I.branch[3].block[15].um_I.iw[4] ,
    \top_I.branch[3].block[15].um_I.iw[3] ,
    \top_I.branch[3].block[15].um_I.iw[2] ,
    \top_I.branch[3].block[15].um_I.iw[1] ,
    \top_I.branch[3].block[15].um_I.clk ,
    \top_I.branch[3].block[14].um_I.iw[17] ,
    \top_I.branch[3].block[14].um_I.iw[16] ,
    \top_I.branch[3].block[14].um_I.iw[15] ,
    \top_I.branch[3].block[14].um_I.iw[14] ,
    \top_I.branch[3].block[14].um_I.iw[13] ,
    \top_I.branch[3].block[14].um_I.iw[12] ,
    \top_I.branch[3].block[14].um_I.iw[11] ,
    \top_I.branch[3].block[14].um_I.iw[10] ,
    \top_I.branch[3].block[14].um_I.iw[9] ,
    \top_I.branch[3].block[14].um_I.iw[8] ,
    \top_I.branch[3].block[14].um_I.iw[7] ,
    \top_I.branch[3].block[14].um_I.iw[6] ,
    \top_I.branch[3].block[14].um_I.iw[5] ,
    \top_I.branch[3].block[14].um_I.iw[4] ,
    \top_I.branch[3].block[14].um_I.iw[3] ,
    \top_I.branch[3].block[14].um_I.iw[2] ,
    \top_I.branch[3].block[14].um_I.iw[1] ,
    \top_I.branch[3].block[14].um_I.clk ,
    \top_I.branch[3].block[13].um_I.iw[17] ,
    \top_I.branch[3].block[13].um_I.iw[16] ,
    \top_I.branch[3].block[13].um_I.iw[15] ,
    \top_I.branch[3].block[13].um_I.iw[14] ,
    \top_I.branch[3].block[13].um_I.iw[13] ,
    \top_I.branch[3].block[13].um_I.iw[12] ,
    \top_I.branch[3].block[13].um_I.iw[11] ,
    \top_I.branch[3].block[13].um_I.iw[10] ,
    \top_I.branch[3].block[13].um_I.iw[9] ,
    \top_I.branch[3].block[13].um_I.iw[8] ,
    \top_I.branch[3].block[13].um_I.iw[7] ,
    \top_I.branch[3].block[13].um_I.iw[6] ,
    \top_I.branch[3].block[13].um_I.iw[5] ,
    \top_I.branch[3].block[13].um_I.iw[4] ,
    \top_I.branch[3].block[13].um_I.iw[3] ,
    \top_I.branch[3].block[13].um_I.iw[2] ,
    \top_I.branch[3].block[13].um_I.iw[1] ,
    \top_I.branch[3].block[13].um_I.clk ,
    \top_I.branch[3].block[12].um_I.iw[17] ,
    \top_I.branch[3].block[12].um_I.iw[16] ,
    \top_I.branch[3].block[12].um_I.iw[15] ,
    \top_I.branch[3].block[12].um_I.iw[14] ,
    \top_I.branch[3].block[12].um_I.iw[13] ,
    \top_I.branch[3].block[12].um_I.iw[12] ,
    \top_I.branch[3].block[12].um_I.iw[11] ,
    \top_I.branch[3].block[12].um_I.iw[10] ,
    \top_I.branch[3].block[12].um_I.iw[9] ,
    \top_I.branch[3].block[12].um_I.iw[8] ,
    \top_I.branch[3].block[12].um_I.iw[7] ,
    \top_I.branch[3].block[12].um_I.iw[6] ,
    \top_I.branch[3].block[12].um_I.iw[5] ,
    \top_I.branch[3].block[12].um_I.iw[4] ,
    \top_I.branch[3].block[12].um_I.iw[3] ,
    \top_I.branch[3].block[12].um_I.iw[2] ,
    \top_I.branch[3].block[12].um_I.iw[1] ,
    \top_I.branch[3].block[12].um_I.clk ,
    \top_I.branch[3].block[11].um_I.iw[17] ,
    \top_I.branch[3].block[11].um_I.iw[16] ,
    \top_I.branch[3].block[11].um_I.iw[15] ,
    \top_I.branch[3].block[11].um_I.iw[14] ,
    \top_I.branch[3].block[11].um_I.iw[13] ,
    \top_I.branch[3].block[11].um_I.iw[12] ,
    \top_I.branch[3].block[11].um_I.iw[11] ,
    \top_I.branch[3].block[11].um_I.iw[10] ,
    \top_I.branch[3].block[11].um_I.iw[9] ,
    \top_I.branch[3].block[11].um_I.iw[8] ,
    \top_I.branch[3].block[11].um_I.iw[7] ,
    \top_I.branch[3].block[11].um_I.iw[6] ,
    \top_I.branch[3].block[11].um_I.iw[5] ,
    \top_I.branch[3].block[11].um_I.iw[4] ,
    \top_I.branch[3].block[11].um_I.iw[3] ,
    \top_I.branch[3].block[11].um_I.iw[2] ,
    \top_I.branch[3].block[11].um_I.iw[1] ,
    \top_I.branch[3].block[11].um_I.clk ,
    \top_I.branch[3].block[10].um_I.iw[17] ,
    \top_I.branch[3].block[10].um_I.iw[16] ,
    \top_I.branch[3].block[10].um_I.iw[15] ,
    \top_I.branch[3].block[10].um_I.iw[14] ,
    \top_I.branch[3].block[10].um_I.iw[13] ,
    \top_I.branch[3].block[10].um_I.iw[12] ,
    \top_I.branch[3].block[10].um_I.iw[11] ,
    \top_I.branch[3].block[10].um_I.iw[10] ,
    \top_I.branch[3].block[10].um_I.iw[9] ,
    \top_I.branch[3].block[10].um_I.iw[8] ,
    \top_I.branch[3].block[10].um_I.iw[7] ,
    \top_I.branch[3].block[10].um_I.iw[6] ,
    \top_I.branch[3].block[10].um_I.iw[5] ,
    \top_I.branch[3].block[10].um_I.iw[4] ,
    \top_I.branch[3].block[10].um_I.iw[3] ,
    \top_I.branch[3].block[10].um_I.iw[2] ,
    \top_I.branch[3].block[10].um_I.iw[1] ,
    \top_I.branch[3].block[10].um_I.clk ,
    \top_I.branch[3].block[9].um_I.iw[17] ,
    \top_I.branch[3].block[9].um_I.iw[16] ,
    \top_I.branch[3].block[9].um_I.iw[15] ,
    \top_I.branch[3].block[9].um_I.iw[14] ,
    \top_I.branch[3].block[9].um_I.iw[13] ,
    \top_I.branch[3].block[9].um_I.iw[12] ,
    \top_I.branch[3].block[9].um_I.iw[11] ,
    \top_I.branch[3].block[9].um_I.iw[10] ,
    \top_I.branch[3].block[9].um_I.iw[9] ,
    \top_I.branch[3].block[9].um_I.iw[8] ,
    \top_I.branch[3].block[9].um_I.iw[7] ,
    \top_I.branch[3].block[9].um_I.iw[6] ,
    \top_I.branch[3].block[9].um_I.iw[5] ,
    \top_I.branch[3].block[9].um_I.iw[4] ,
    \top_I.branch[3].block[9].um_I.iw[3] ,
    \top_I.branch[3].block[9].um_I.iw[2] ,
    \top_I.branch[3].block[9].um_I.iw[1] ,
    \top_I.branch[3].block[9].um_I.clk ,
    \top_I.branch[3].block[8].um_I.iw[17] ,
    \top_I.branch[3].block[8].um_I.iw[16] ,
    \top_I.branch[3].block[8].um_I.iw[15] ,
    \top_I.branch[3].block[8].um_I.iw[14] ,
    \top_I.branch[3].block[8].um_I.iw[13] ,
    \top_I.branch[3].block[8].um_I.iw[12] ,
    \top_I.branch[3].block[8].um_I.iw[11] ,
    \top_I.branch[3].block[8].um_I.iw[10] ,
    \top_I.branch[3].block[8].um_I.iw[9] ,
    \top_I.branch[3].block[8].um_I.iw[8] ,
    \top_I.branch[3].block[8].um_I.iw[7] ,
    \top_I.branch[3].block[8].um_I.iw[6] ,
    \top_I.branch[3].block[8].um_I.iw[5] ,
    \top_I.branch[3].block[8].um_I.iw[4] ,
    \top_I.branch[3].block[8].um_I.iw[3] ,
    \top_I.branch[3].block[8].um_I.iw[2] ,
    \top_I.branch[3].block[8].um_I.iw[1] ,
    \top_I.branch[3].block[8].um_I.clk ,
    \top_I.branch[3].block[7].um_I.iw[17] ,
    \top_I.branch[3].block[7].um_I.iw[16] ,
    \top_I.branch[3].block[7].um_I.iw[15] ,
    \top_I.branch[3].block[7].um_I.iw[14] ,
    \top_I.branch[3].block[7].um_I.iw[13] ,
    \top_I.branch[3].block[7].um_I.iw[12] ,
    \top_I.branch[3].block[7].um_I.iw[11] ,
    \top_I.branch[3].block[7].um_I.iw[10] ,
    \top_I.branch[3].block[7].um_I.iw[9] ,
    \top_I.branch[3].block[7].um_I.iw[8] ,
    \top_I.branch[3].block[7].um_I.iw[7] ,
    \top_I.branch[3].block[7].um_I.iw[6] ,
    \top_I.branch[3].block[7].um_I.iw[5] ,
    \top_I.branch[3].block[7].um_I.iw[4] ,
    \top_I.branch[3].block[7].um_I.iw[3] ,
    \top_I.branch[3].block[7].um_I.iw[2] ,
    \top_I.branch[3].block[7].um_I.iw[1] ,
    \top_I.branch[3].block[7].um_I.clk ,
    \top_I.branch[3].block[6].um_I.iw[17] ,
    \top_I.branch[3].block[6].um_I.iw[16] ,
    \top_I.branch[3].block[6].um_I.iw[15] ,
    \top_I.branch[3].block[6].um_I.iw[14] ,
    \top_I.branch[3].block[6].um_I.iw[13] ,
    \top_I.branch[3].block[6].um_I.iw[12] ,
    \top_I.branch[3].block[6].um_I.iw[11] ,
    \top_I.branch[3].block[6].um_I.iw[10] ,
    \top_I.branch[3].block[6].um_I.iw[9] ,
    \top_I.branch[3].block[6].um_I.iw[8] ,
    \top_I.branch[3].block[6].um_I.iw[7] ,
    \top_I.branch[3].block[6].um_I.iw[6] ,
    \top_I.branch[3].block[6].um_I.iw[5] ,
    \top_I.branch[3].block[6].um_I.iw[4] ,
    \top_I.branch[3].block[6].um_I.iw[3] ,
    \top_I.branch[3].block[6].um_I.iw[2] ,
    \top_I.branch[3].block[6].um_I.iw[1] ,
    \top_I.branch[3].block[6].um_I.clk ,
    \top_I.branch[3].block[5].um_I.iw[17] ,
    \top_I.branch[3].block[5].um_I.iw[16] ,
    \top_I.branch[3].block[5].um_I.iw[15] ,
    \top_I.branch[3].block[5].um_I.iw[14] ,
    \top_I.branch[3].block[5].um_I.iw[13] ,
    \top_I.branch[3].block[5].um_I.iw[12] ,
    \top_I.branch[3].block[5].um_I.iw[11] ,
    \top_I.branch[3].block[5].um_I.iw[10] ,
    \top_I.branch[3].block[5].um_I.iw[9] ,
    \top_I.branch[3].block[5].um_I.iw[8] ,
    \top_I.branch[3].block[5].um_I.iw[7] ,
    \top_I.branch[3].block[5].um_I.iw[6] ,
    \top_I.branch[3].block[5].um_I.iw[5] ,
    \top_I.branch[3].block[5].um_I.iw[4] ,
    \top_I.branch[3].block[5].um_I.iw[3] ,
    \top_I.branch[3].block[5].um_I.iw[2] ,
    \top_I.branch[3].block[5].um_I.iw[1] ,
    \top_I.branch[3].block[5].um_I.clk ,
    \top_I.branch[3].block[4].um_I.iw[17] ,
    \top_I.branch[3].block[4].um_I.iw[16] ,
    \top_I.branch[3].block[4].um_I.iw[15] ,
    \top_I.branch[3].block[4].um_I.iw[14] ,
    \top_I.branch[3].block[4].um_I.iw[13] ,
    \top_I.branch[3].block[4].um_I.iw[12] ,
    \top_I.branch[3].block[4].um_I.iw[11] ,
    \top_I.branch[3].block[4].um_I.iw[10] ,
    \top_I.branch[3].block[4].um_I.iw[9] ,
    \top_I.branch[3].block[4].um_I.iw[8] ,
    \top_I.branch[3].block[4].um_I.iw[7] ,
    \top_I.branch[3].block[4].um_I.iw[6] ,
    \top_I.branch[3].block[4].um_I.iw[5] ,
    \top_I.branch[3].block[4].um_I.iw[4] ,
    \top_I.branch[3].block[4].um_I.iw[3] ,
    \top_I.branch[3].block[4].um_I.iw[2] ,
    \top_I.branch[3].block[4].um_I.iw[1] ,
    \top_I.branch[3].block[4].um_I.clk ,
    \top_I.branch[3].block[3].um_I.iw[17] ,
    \top_I.branch[3].block[3].um_I.iw[16] ,
    \top_I.branch[3].block[3].um_I.iw[15] ,
    \top_I.branch[3].block[3].um_I.iw[14] ,
    \top_I.branch[3].block[3].um_I.iw[13] ,
    \top_I.branch[3].block[3].um_I.iw[12] ,
    \top_I.branch[3].block[3].um_I.iw[11] ,
    \top_I.branch[3].block[3].um_I.iw[10] ,
    \top_I.branch[3].block[3].um_I.iw[9] ,
    \top_I.branch[3].block[3].um_I.iw[8] ,
    \top_I.branch[3].block[3].um_I.iw[7] ,
    \top_I.branch[3].block[3].um_I.iw[6] ,
    \top_I.branch[3].block[3].um_I.iw[5] ,
    \top_I.branch[3].block[3].um_I.iw[4] ,
    \top_I.branch[3].block[3].um_I.iw[3] ,
    \top_I.branch[3].block[3].um_I.iw[2] ,
    \top_I.branch[3].block[3].um_I.iw[1] ,
    \top_I.branch[3].block[3].um_I.clk ,
    \top_I.branch[3].block[2].um_I.iw[17] ,
    \top_I.branch[3].block[2].um_I.iw[16] ,
    \top_I.branch[3].block[2].um_I.iw[15] ,
    \top_I.branch[3].block[2].um_I.iw[14] ,
    \top_I.branch[3].block[2].um_I.iw[13] ,
    \top_I.branch[3].block[2].um_I.iw[12] ,
    \top_I.branch[3].block[2].um_I.iw[11] ,
    \top_I.branch[3].block[2].um_I.iw[10] ,
    \top_I.branch[3].block[2].um_I.iw[9] ,
    \top_I.branch[3].block[2].um_I.iw[8] ,
    \top_I.branch[3].block[2].um_I.iw[7] ,
    \top_I.branch[3].block[2].um_I.iw[6] ,
    \top_I.branch[3].block[2].um_I.iw[5] ,
    \top_I.branch[3].block[2].um_I.iw[4] ,
    \top_I.branch[3].block[2].um_I.iw[3] ,
    \top_I.branch[3].block[2].um_I.iw[2] ,
    \top_I.branch[3].block[2].um_I.iw[1] ,
    \top_I.branch[3].block[2].um_I.clk ,
    \top_I.branch[3].block[1].um_I.iw[17] ,
    \top_I.branch[3].block[1].um_I.iw[16] ,
    \top_I.branch[3].block[1].um_I.iw[15] ,
    \top_I.branch[3].block[1].um_I.iw[14] ,
    \top_I.branch[3].block[1].um_I.iw[13] ,
    \top_I.branch[3].block[1].um_I.iw[12] ,
    \top_I.branch[3].block[1].um_I.iw[11] ,
    \top_I.branch[3].block[1].um_I.iw[10] ,
    \top_I.branch[3].block[1].um_I.iw[9] ,
    \top_I.branch[3].block[1].um_I.iw[8] ,
    \top_I.branch[3].block[1].um_I.iw[7] ,
    \top_I.branch[3].block[1].um_I.iw[6] ,
    \top_I.branch[3].block[1].um_I.iw[5] ,
    \top_I.branch[3].block[1].um_I.iw[4] ,
    \top_I.branch[3].block[1].um_I.iw[3] ,
    \top_I.branch[3].block[1].um_I.iw[2] ,
    \top_I.branch[3].block[1].um_I.iw[1] ,
    \top_I.branch[3].block[1].um_I.clk ,
    \top_I.branch[3].block[0].um_I.iw[17] ,
    \top_I.branch[3].block[0].um_I.iw[16] ,
    \top_I.branch[3].block[0].um_I.iw[15] ,
    \top_I.branch[3].block[0].um_I.iw[14] ,
    \top_I.branch[3].block[0].um_I.iw[13] ,
    \top_I.branch[3].block[0].um_I.iw[12] ,
    \top_I.branch[3].block[0].um_I.iw[11] ,
    \top_I.branch[3].block[0].um_I.iw[10] ,
    \top_I.branch[3].block[0].um_I.iw[9] ,
    \top_I.branch[3].block[0].um_I.iw[8] ,
    \top_I.branch[3].block[0].um_I.iw[7] ,
    \top_I.branch[3].block[0].um_I.iw[6] ,
    \top_I.branch[3].block[0].um_I.iw[5] ,
    \top_I.branch[3].block[0].um_I.iw[4] ,
    \top_I.branch[3].block[0].um_I.iw[3] ,
    \top_I.branch[3].block[0].um_I.iw[2] ,
    \top_I.branch[3].block[0].um_I.iw[1] ,
    \top_I.branch[3].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[3].block[15].um_I.pg_vdd ,
    \top_I.branch[3].block[14].um_I.pg_vdd ,
    \top_I.branch[3].block[13].um_I.pg_vdd ,
    \top_I.branch[3].block[12].um_I.pg_vdd ,
    \top_I.branch[3].block[11].um_I.pg_vdd ,
    \top_I.branch[3].block[10].um_I.pg_vdd ,
    \top_I.branch[3].block[9].um_I.pg_vdd ,
    \top_I.branch[3].block[8].um_I.pg_vdd ,
    \top_I.branch[3].block[7].um_I.pg_vdd ,
    \top_I.branch[3].block[6].um_I.pg_vdd ,
    \top_I.branch[3].block[5].um_I.pg_vdd ,
    \top_I.branch[3].block[4].um_I.pg_vdd ,
    \top_I.branch[3].block[3].um_I.pg_vdd ,
    \top_I.branch[3].block[2].um_I.pg_vdd ,
    \top_I.branch[3].block[1].um_I.pg_vdd ,
    \top_I.branch[3].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[4].mux_I  (.k_one(\top_I.branch[4].l_addr[1] ),
    .k_zero(\top_I.branch[4].l_addr[0] ),
    .addr({\top_I.branch[4].l_addr[0] ,
    \top_I.branch[4].l_addr[0] ,
    \top_I.branch[4].l_addr[1] ,
    \top_I.branch[4].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[4].block[15].um_I.ena ,
    \top_I.branch[4].block[14].um_I.ena ,
    \top_I.branch[4].block[13].um_I.ena ,
    \top_I.branch[4].block[12].um_I.ena ,
    \top_I.branch[4].block[11].um_I.ena ,
    \top_I.branch[4].block[10].um_I.ena ,
    \top_I.branch[4].block[9].um_I.ena ,
    \top_I.branch[4].block[8].um_I.ena ,
    \top_I.branch[4].block[7].um_I.ena ,
    \top_I.branch[4].block[6].um_I.ena ,
    \top_I.branch[4].block[5].um_I.ena ,
    \top_I.branch[4].block[4].um_I.ena ,
    \top_I.branch[4].block[3].um_I.ena ,
    \top_I.branch[4].block[2].um_I.ena ,
    \top_I.branch[4].block[1].um_I.ena ,
    \top_I.branch[4].block[0].um_I.ena }),
    .um_iw({\top_I.branch[4].block[15].um_I.iw[17] ,
    \top_I.branch[4].block[15].um_I.iw[16] ,
    \top_I.branch[4].block[15].um_I.iw[15] ,
    \top_I.branch[4].block[15].um_I.iw[14] ,
    \top_I.branch[4].block[15].um_I.iw[13] ,
    \top_I.branch[4].block[15].um_I.iw[12] ,
    \top_I.branch[4].block[15].um_I.iw[11] ,
    \top_I.branch[4].block[15].um_I.iw[10] ,
    \top_I.branch[4].block[15].um_I.iw[9] ,
    \top_I.branch[4].block[15].um_I.iw[8] ,
    \top_I.branch[4].block[15].um_I.iw[7] ,
    \top_I.branch[4].block[15].um_I.iw[6] ,
    \top_I.branch[4].block[15].um_I.iw[5] ,
    \top_I.branch[4].block[15].um_I.iw[4] ,
    \top_I.branch[4].block[15].um_I.iw[3] ,
    \top_I.branch[4].block[15].um_I.iw[2] ,
    \top_I.branch[4].block[15].um_I.iw[1] ,
    \top_I.branch[4].block[15].um_I.clk ,
    \top_I.branch[4].block[14].um_I.iw[17] ,
    \top_I.branch[4].block[14].um_I.iw[16] ,
    \top_I.branch[4].block[14].um_I.iw[15] ,
    \top_I.branch[4].block[14].um_I.iw[14] ,
    \top_I.branch[4].block[14].um_I.iw[13] ,
    \top_I.branch[4].block[14].um_I.iw[12] ,
    \top_I.branch[4].block[14].um_I.iw[11] ,
    \top_I.branch[4].block[14].um_I.iw[10] ,
    \top_I.branch[4].block[14].um_I.iw[9] ,
    \top_I.branch[4].block[14].um_I.iw[8] ,
    \top_I.branch[4].block[14].um_I.iw[7] ,
    \top_I.branch[4].block[14].um_I.iw[6] ,
    \top_I.branch[4].block[14].um_I.iw[5] ,
    \top_I.branch[4].block[14].um_I.iw[4] ,
    \top_I.branch[4].block[14].um_I.iw[3] ,
    \top_I.branch[4].block[14].um_I.iw[2] ,
    \top_I.branch[4].block[14].um_I.iw[1] ,
    \top_I.branch[4].block[14].um_I.clk ,
    \top_I.branch[4].block[13].um_I.iw[17] ,
    \top_I.branch[4].block[13].um_I.iw[16] ,
    \top_I.branch[4].block[13].um_I.iw[15] ,
    \top_I.branch[4].block[13].um_I.iw[14] ,
    \top_I.branch[4].block[13].um_I.iw[13] ,
    \top_I.branch[4].block[13].um_I.iw[12] ,
    \top_I.branch[4].block[13].um_I.iw[11] ,
    \top_I.branch[4].block[13].um_I.iw[10] ,
    \top_I.branch[4].block[13].um_I.iw[9] ,
    \top_I.branch[4].block[13].um_I.iw[8] ,
    \top_I.branch[4].block[13].um_I.iw[7] ,
    \top_I.branch[4].block[13].um_I.iw[6] ,
    \top_I.branch[4].block[13].um_I.iw[5] ,
    \top_I.branch[4].block[13].um_I.iw[4] ,
    \top_I.branch[4].block[13].um_I.iw[3] ,
    \top_I.branch[4].block[13].um_I.iw[2] ,
    \top_I.branch[4].block[13].um_I.iw[1] ,
    \top_I.branch[4].block[13].um_I.clk ,
    \top_I.branch[4].block[12].um_I.iw[17] ,
    \top_I.branch[4].block[12].um_I.iw[16] ,
    \top_I.branch[4].block[12].um_I.iw[15] ,
    \top_I.branch[4].block[12].um_I.iw[14] ,
    \top_I.branch[4].block[12].um_I.iw[13] ,
    \top_I.branch[4].block[12].um_I.iw[12] ,
    \top_I.branch[4].block[12].um_I.iw[11] ,
    \top_I.branch[4].block[12].um_I.iw[10] ,
    \top_I.branch[4].block[12].um_I.iw[9] ,
    \top_I.branch[4].block[12].um_I.iw[8] ,
    \top_I.branch[4].block[12].um_I.iw[7] ,
    \top_I.branch[4].block[12].um_I.iw[6] ,
    \top_I.branch[4].block[12].um_I.iw[5] ,
    \top_I.branch[4].block[12].um_I.iw[4] ,
    \top_I.branch[4].block[12].um_I.iw[3] ,
    \top_I.branch[4].block[12].um_I.iw[2] ,
    \top_I.branch[4].block[12].um_I.iw[1] ,
    \top_I.branch[4].block[12].um_I.clk ,
    \top_I.branch[4].block[11].um_I.iw[17] ,
    \top_I.branch[4].block[11].um_I.iw[16] ,
    \top_I.branch[4].block[11].um_I.iw[15] ,
    \top_I.branch[4].block[11].um_I.iw[14] ,
    \top_I.branch[4].block[11].um_I.iw[13] ,
    \top_I.branch[4].block[11].um_I.iw[12] ,
    \top_I.branch[4].block[11].um_I.iw[11] ,
    \top_I.branch[4].block[11].um_I.iw[10] ,
    \top_I.branch[4].block[11].um_I.iw[9] ,
    \top_I.branch[4].block[11].um_I.iw[8] ,
    \top_I.branch[4].block[11].um_I.iw[7] ,
    \top_I.branch[4].block[11].um_I.iw[6] ,
    \top_I.branch[4].block[11].um_I.iw[5] ,
    \top_I.branch[4].block[11].um_I.iw[4] ,
    \top_I.branch[4].block[11].um_I.iw[3] ,
    \top_I.branch[4].block[11].um_I.iw[2] ,
    \top_I.branch[4].block[11].um_I.iw[1] ,
    \top_I.branch[4].block[11].um_I.clk ,
    \top_I.branch[4].block[10].um_I.iw[17] ,
    \top_I.branch[4].block[10].um_I.iw[16] ,
    \top_I.branch[4].block[10].um_I.iw[15] ,
    \top_I.branch[4].block[10].um_I.iw[14] ,
    \top_I.branch[4].block[10].um_I.iw[13] ,
    \top_I.branch[4].block[10].um_I.iw[12] ,
    \top_I.branch[4].block[10].um_I.iw[11] ,
    \top_I.branch[4].block[10].um_I.iw[10] ,
    \top_I.branch[4].block[10].um_I.iw[9] ,
    \top_I.branch[4].block[10].um_I.iw[8] ,
    \top_I.branch[4].block[10].um_I.iw[7] ,
    \top_I.branch[4].block[10].um_I.iw[6] ,
    \top_I.branch[4].block[10].um_I.iw[5] ,
    \top_I.branch[4].block[10].um_I.iw[4] ,
    \top_I.branch[4].block[10].um_I.iw[3] ,
    \top_I.branch[4].block[10].um_I.iw[2] ,
    \top_I.branch[4].block[10].um_I.iw[1] ,
    \top_I.branch[4].block[10].um_I.clk ,
    \top_I.branch[4].block[9].um_I.iw[17] ,
    \top_I.branch[4].block[9].um_I.iw[16] ,
    \top_I.branch[4].block[9].um_I.iw[15] ,
    \top_I.branch[4].block[9].um_I.iw[14] ,
    \top_I.branch[4].block[9].um_I.iw[13] ,
    \top_I.branch[4].block[9].um_I.iw[12] ,
    \top_I.branch[4].block[9].um_I.iw[11] ,
    \top_I.branch[4].block[9].um_I.iw[10] ,
    \top_I.branch[4].block[9].um_I.iw[9] ,
    \top_I.branch[4].block[9].um_I.iw[8] ,
    \top_I.branch[4].block[9].um_I.iw[7] ,
    \top_I.branch[4].block[9].um_I.iw[6] ,
    \top_I.branch[4].block[9].um_I.iw[5] ,
    \top_I.branch[4].block[9].um_I.iw[4] ,
    \top_I.branch[4].block[9].um_I.iw[3] ,
    \top_I.branch[4].block[9].um_I.iw[2] ,
    \top_I.branch[4].block[9].um_I.iw[1] ,
    \top_I.branch[4].block[9].um_I.clk ,
    \top_I.branch[4].block[8].um_I.iw[17] ,
    \top_I.branch[4].block[8].um_I.iw[16] ,
    \top_I.branch[4].block[8].um_I.iw[15] ,
    \top_I.branch[4].block[8].um_I.iw[14] ,
    \top_I.branch[4].block[8].um_I.iw[13] ,
    \top_I.branch[4].block[8].um_I.iw[12] ,
    \top_I.branch[4].block[8].um_I.iw[11] ,
    \top_I.branch[4].block[8].um_I.iw[10] ,
    \top_I.branch[4].block[8].um_I.iw[9] ,
    \top_I.branch[4].block[8].um_I.iw[8] ,
    \top_I.branch[4].block[8].um_I.iw[7] ,
    \top_I.branch[4].block[8].um_I.iw[6] ,
    \top_I.branch[4].block[8].um_I.iw[5] ,
    \top_I.branch[4].block[8].um_I.iw[4] ,
    \top_I.branch[4].block[8].um_I.iw[3] ,
    \top_I.branch[4].block[8].um_I.iw[2] ,
    \top_I.branch[4].block[8].um_I.iw[1] ,
    \top_I.branch[4].block[8].um_I.clk ,
    \top_I.branch[4].block[7].um_I.iw[17] ,
    \top_I.branch[4].block[7].um_I.iw[16] ,
    \top_I.branch[4].block[7].um_I.iw[15] ,
    \top_I.branch[4].block[7].um_I.iw[14] ,
    \top_I.branch[4].block[7].um_I.iw[13] ,
    \top_I.branch[4].block[7].um_I.iw[12] ,
    \top_I.branch[4].block[7].um_I.iw[11] ,
    \top_I.branch[4].block[7].um_I.iw[10] ,
    \top_I.branch[4].block[7].um_I.iw[9] ,
    \top_I.branch[4].block[7].um_I.iw[8] ,
    \top_I.branch[4].block[7].um_I.iw[7] ,
    \top_I.branch[4].block[7].um_I.iw[6] ,
    \top_I.branch[4].block[7].um_I.iw[5] ,
    \top_I.branch[4].block[7].um_I.iw[4] ,
    \top_I.branch[4].block[7].um_I.iw[3] ,
    \top_I.branch[4].block[7].um_I.iw[2] ,
    \top_I.branch[4].block[7].um_I.iw[1] ,
    \top_I.branch[4].block[7].um_I.clk ,
    \top_I.branch[4].block[6].um_I.iw[17] ,
    \top_I.branch[4].block[6].um_I.iw[16] ,
    \top_I.branch[4].block[6].um_I.iw[15] ,
    \top_I.branch[4].block[6].um_I.iw[14] ,
    \top_I.branch[4].block[6].um_I.iw[13] ,
    \top_I.branch[4].block[6].um_I.iw[12] ,
    \top_I.branch[4].block[6].um_I.iw[11] ,
    \top_I.branch[4].block[6].um_I.iw[10] ,
    \top_I.branch[4].block[6].um_I.iw[9] ,
    \top_I.branch[4].block[6].um_I.iw[8] ,
    \top_I.branch[4].block[6].um_I.iw[7] ,
    \top_I.branch[4].block[6].um_I.iw[6] ,
    \top_I.branch[4].block[6].um_I.iw[5] ,
    \top_I.branch[4].block[6].um_I.iw[4] ,
    \top_I.branch[4].block[6].um_I.iw[3] ,
    \top_I.branch[4].block[6].um_I.iw[2] ,
    \top_I.branch[4].block[6].um_I.iw[1] ,
    \top_I.branch[4].block[6].um_I.clk ,
    \top_I.branch[4].block[5].um_I.iw[17] ,
    \top_I.branch[4].block[5].um_I.iw[16] ,
    \top_I.branch[4].block[5].um_I.iw[15] ,
    \top_I.branch[4].block[5].um_I.iw[14] ,
    \top_I.branch[4].block[5].um_I.iw[13] ,
    \top_I.branch[4].block[5].um_I.iw[12] ,
    \top_I.branch[4].block[5].um_I.iw[11] ,
    \top_I.branch[4].block[5].um_I.iw[10] ,
    \top_I.branch[4].block[5].um_I.iw[9] ,
    \top_I.branch[4].block[5].um_I.iw[8] ,
    \top_I.branch[4].block[5].um_I.iw[7] ,
    \top_I.branch[4].block[5].um_I.iw[6] ,
    \top_I.branch[4].block[5].um_I.iw[5] ,
    \top_I.branch[4].block[5].um_I.iw[4] ,
    \top_I.branch[4].block[5].um_I.iw[3] ,
    \top_I.branch[4].block[5].um_I.iw[2] ,
    \top_I.branch[4].block[5].um_I.iw[1] ,
    \top_I.branch[4].block[5].um_I.clk ,
    \top_I.branch[4].block[4].um_I.iw[17] ,
    \top_I.branch[4].block[4].um_I.iw[16] ,
    \top_I.branch[4].block[4].um_I.iw[15] ,
    \top_I.branch[4].block[4].um_I.iw[14] ,
    \top_I.branch[4].block[4].um_I.iw[13] ,
    \top_I.branch[4].block[4].um_I.iw[12] ,
    \top_I.branch[4].block[4].um_I.iw[11] ,
    \top_I.branch[4].block[4].um_I.iw[10] ,
    \top_I.branch[4].block[4].um_I.iw[9] ,
    \top_I.branch[4].block[4].um_I.iw[8] ,
    \top_I.branch[4].block[4].um_I.iw[7] ,
    \top_I.branch[4].block[4].um_I.iw[6] ,
    \top_I.branch[4].block[4].um_I.iw[5] ,
    \top_I.branch[4].block[4].um_I.iw[4] ,
    \top_I.branch[4].block[4].um_I.iw[3] ,
    \top_I.branch[4].block[4].um_I.iw[2] ,
    \top_I.branch[4].block[4].um_I.iw[1] ,
    \top_I.branch[4].block[4].um_I.clk ,
    \top_I.branch[4].block[3].um_I.iw[17] ,
    \top_I.branch[4].block[3].um_I.iw[16] ,
    \top_I.branch[4].block[3].um_I.iw[15] ,
    \top_I.branch[4].block[3].um_I.iw[14] ,
    \top_I.branch[4].block[3].um_I.iw[13] ,
    \top_I.branch[4].block[3].um_I.iw[12] ,
    \top_I.branch[4].block[3].um_I.iw[11] ,
    \top_I.branch[4].block[3].um_I.iw[10] ,
    \top_I.branch[4].block[3].um_I.iw[9] ,
    \top_I.branch[4].block[3].um_I.iw[8] ,
    \top_I.branch[4].block[3].um_I.iw[7] ,
    \top_I.branch[4].block[3].um_I.iw[6] ,
    \top_I.branch[4].block[3].um_I.iw[5] ,
    \top_I.branch[4].block[3].um_I.iw[4] ,
    \top_I.branch[4].block[3].um_I.iw[3] ,
    \top_I.branch[4].block[3].um_I.iw[2] ,
    \top_I.branch[4].block[3].um_I.iw[1] ,
    \top_I.branch[4].block[3].um_I.clk ,
    \top_I.branch[4].block[2].um_I.iw[17] ,
    \top_I.branch[4].block[2].um_I.iw[16] ,
    \top_I.branch[4].block[2].um_I.iw[15] ,
    \top_I.branch[4].block[2].um_I.iw[14] ,
    \top_I.branch[4].block[2].um_I.iw[13] ,
    \top_I.branch[4].block[2].um_I.iw[12] ,
    \top_I.branch[4].block[2].um_I.iw[11] ,
    \top_I.branch[4].block[2].um_I.iw[10] ,
    \top_I.branch[4].block[2].um_I.iw[9] ,
    \top_I.branch[4].block[2].um_I.iw[8] ,
    \top_I.branch[4].block[2].um_I.iw[7] ,
    \top_I.branch[4].block[2].um_I.iw[6] ,
    \top_I.branch[4].block[2].um_I.iw[5] ,
    \top_I.branch[4].block[2].um_I.iw[4] ,
    \top_I.branch[4].block[2].um_I.iw[3] ,
    \top_I.branch[4].block[2].um_I.iw[2] ,
    \top_I.branch[4].block[2].um_I.iw[1] ,
    \top_I.branch[4].block[2].um_I.clk ,
    \top_I.branch[4].block[1].um_I.iw[17] ,
    \top_I.branch[4].block[1].um_I.iw[16] ,
    \top_I.branch[4].block[1].um_I.iw[15] ,
    \top_I.branch[4].block[1].um_I.iw[14] ,
    \top_I.branch[4].block[1].um_I.iw[13] ,
    \top_I.branch[4].block[1].um_I.iw[12] ,
    \top_I.branch[4].block[1].um_I.iw[11] ,
    \top_I.branch[4].block[1].um_I.iw[10] ,
    \top_I.branch[4].block[1].um_I.iw[9] ,
    \top_I.branch[4].block[1].um_I.iw[8] ,
    \top_I.branch[4].block[1].um_I.iw[7] ,
    \top_I.branch[4].block[1].um_I.iw[6] ,
    \top_I.branch[4].block[1].um_I.iw[5] ,
    \top_I.branch[4].block[1].um_I.iw[4] ,
    \top_I.branch[4].block[1].um_I.iw[3] ,
    \top_I.branch[4].block[1].um_I.iw[2] ,
    \top_I.branch[4].block[1].um_I.iw[1] ,
    \top_I.branch[4].block[1].um_I.clk ,
    \top_I.branch[4].block[0].um_I.iw[17] ,
    \top_I.branch[4].block[0].um_I.iw[16] ,
    \top_I.branch[4].block[0].um_I.iw[15] ,
    \top_I.branch[4].block[0].um_I.iw[14] ,
    \top_I.branch[4].block[0].um_I.iw[13] ,
    \top_I.branch[4].block[0].um_I.iw[12] ,
    \top_I.branch[4].block[0].um_I.iw[11] ,
    \top_I.branch[4].block[0].um_I.iw[10] ,
    \top_I.branch[4].block[0].um_I.iw[9] ,
    \top_I.branch[4].block[0].um_I.iw[8] ,
    \top_I.branch[4].block[0].um_I.iw[7] ,
    \top_I.branch[4].block[0].um_I.iw[6] ,
    \top_I.branch[4].block[0].um_I.iw[5] ,
    \top_I.branch[4].block[0].um_I.iw[4] ,
    \top_I.branch[4].block[0].um_I.iw[3] ,
    \top_I.branch[4].block[0].um_I.iw[2] ,
    \top_I.branch[4].block[0].um_I.iw[1] ,
    \top_I.branch[4].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[4].block[15].um_I.pg_vdd ,
    \top_I.branch[4].block[14].um_I.pg_vdd ,
    \top_I.branch[4].block[13].um_I.pg_vdd ,
    \top_I.branch[4].block[12].um_I.pg_vdd ,
    \top_I.branch[4].block[11].um_I.pg_vdd ,
    \top_I.branch[4].block[10].um_I.pg_vdd ,
    \top_I.branch[4].block[9].um_I.pg_vdd ,
    \top_I.branch[4].block[8].um_I.pg_vdd ,
    \top_I.branch[4].block[7].um_I.pg_vdd ,
    \top_I.branch[4].block[6].um_I.pg_vdd ,
    \top_I.branch[4].block[5].um_I.pg_vdd ,
    \top_I.branch[4].block[4].um_I.pg_vdd ,
    \top_I.branch[4].block[3].um_I.pg_vdd ,
    \top_I.branch[4].block[2].um_I.pg_vdd ,
    \top_I.branch[4].block[1].um_I.pg_vdd ,
    \top_I.branch[4].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[5].mux_I  (.k_one(\top_I.branch[5].l_addr[1] ),
    .k_zero(\top_I.branch[5].l_addr[0] ),
    .addr({\top_I.branch[5].l_addr[0] ,
    \top_I.branch[5].l_addr[0] ,
    \top_I.branch[5].l_addr[1] ,
    \top_I.branch[5].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[5].block[15].um_I.ena ,
    \top_I.branch[5].block[14].um_I.ena ,
    \top_I.branch[5].block[13].um_I.ena ,
    \top_I.branch[5].block[12].um_I.ena ,
    \top_I.branch[5].block[11].um_I.ena ,
    \top_I.branch[5].block[10].um_I.ena ,
    \top_I.branch[5].block[9].um_I.ena ,
    \top_I.branch[5].block[8].um_I.ena ,
    \top_I.branch[5].block[7].um_I.ena ,
    \top_I.branch[5].block[6].um_I.ena ,
    \top_I.branch[5].block[5].um_I.ena ,
    \top_I.branch[5].block[4].um_I.ena ,
    \top_I.branch[5].block[3].um_I.ena ,
    \top_I.branch[5].block[2].um_I.ena ,
    \top_I.branch[5].block[1].um_I.ena ,
    \top_I.branch[5].block[0].um_I.ena }),
    .um_iw({\top_I.branch[5].block[15].um_I.iw[17] ,
    \top_I.branch[5].block[15].um_I.iw[16] ,
    \top_I.branch[5].block[15].um_I.iw[15] ,
    \top_I.branch[5].block[15].um_I.iw[14] ,
    \top_I.branch[5].block[15].um_I.iw[13] ,
    \top_I.branch[5].block[15].um_I.iw[12] ,
    \top_I.branch[5].block[15].um_I.iw[11] ,
    \top_I.branch[5].block[15].um_I.iw[10] ,
    \top_I.branch[5].block[15].um_I.iw[9] ,
    \top_I.branch[5].block[15].um_I.iw[8] ,
    \top_I.branch[5].block[15].um_I.iw[7] ,
    \top_I.branch[5].block[15].um_I.iw[6] ,
    \top_I.branch[5].block[15].um_I.iw[5] ,
    \top_I.branch[5].block[15].um_I.iw[4] ,
    \top_I.branch[5].block[15].um_I.iw[3] ,
    \top_I.branch[5].block[15].um_I.iw[2] ,
    \top_I.branch[5].block[15].um_I.iw[1] ,
    \top_I.branch[5].block[15].um_I.clk ,
    \top_I.branch[5].block[14].um_I.iw[17] ,
    \top_I.branch[5].block[14].um_I.iw[16] ,
    \top_I.branch[5].block[14].um_I.iw[15] ,
    \top_I.branch[5].block[14].um_I.iw[14] ,
    \top_I.branch[5].block[14].um_I.iw[13] ,
    \top_I.branch[5].block[14].um_I.iw[12] ,
    \top_I.branch[5].block[14].um_I.iw[11] ,
    \top_I.branch[5].block[14].um_I.iw[10] ,
    \top_I.branch[5].block[14].um_I.iw[9] ,
    \top_I.branch[5].block[14].um_I.iw[8] ,
    \top_I.branch[5].block[14].um_I.iw[7] ,
    \top_I.branch[5].block[14].um_I.iw[6] ,
    \top_I.branch[5].block[14].um_I.iw[5] ,
    \top_I.branch[5].block[14].um_I.iw[4] ,
    \top_I.branch[5].block[14].um_I.iw[3] ,
    \top_I.branch[5].block[14].um_I.iw[2] ,
    \top_I.branch[5].block[14].um_I.iw[1] ,
    \top_I.branch[5].block[14].um_I.clk ,
    \top_I.branch[5].block[13].um_I.iw[17] ,
    \top_I.branch[5].block[13].um_I.iw[16] ,
    \top_I.branch[5].block[13].um_I.iw[15] ,
    \top_I.branch[5].block[13].um_I.iw[14] ,
    \top_I.branch[5].block[13].um_I.iw[13] ,
    \top_I.branch[5].block[13].um_I.iw[12] ,
    \top_I.branch[5].block[13].um_I.iw[11] ,
    \top_I.branch[5].block[13].um_I.iw[10] ,
    \top_I.branch[5].block[13].um_I.iw[9] ,
    \top_I.branch[5].block[13].um_I.iw[8] ,
    \top_I.branch[5].block[13].um_I.iw[7] ,
    \top_I.branch[5].block[13].um_I.iw[6] ,
    \top_I.branch[5].block[13].um_I.iw[5] ,
    \top_I.branch[5].block[13].um_I.iw[4] ,
    \top_I.branch[5].block[13].um_I.iw[3] ,
    \top_I.branch[5].block[13].um_I.iw[2] ,
    \top_I.branch[5].block[13].um_I.iw[1] ,
    \top_I.branch[5].block[13].um_I.clk ,
    \top_I.branch[5].block[12].um_I.iw[17] ,
    \top_I.branch[5].block[12].um_I.iw[16] ,
    \top_I.branch[5].block[12].um_I.iw[15] ,
    \top_I.branch[5].block[12].um_I.iw[14] ,
    \top_I.branch[5].block[12].um_I.iw[13] ,
    \top_I.branch[5].block[12].um_I.iw[12] ,
    \top_I.branch[5].block[12].um_I.iw[11] ,
    \top_I.branch[5].block[12].um_I.iw[10] ,
    \top_I.branch[5].block[12].um_I.iw[9] ,
    \top_I.branch[5].block[12].um_I.iw[8] ,
    \top_I.branch[5].block[12].um_I.iw[7] ,
    \top_I.branch[5].block[12].um_I.iw[6] ,
    \top_I.branch[5].block[12].um_I.iw[5] ,
    \top_I.branch[5].block[12].um_I.iw[4] ,
    \top_I.branch[5].block[12].um_I.iw[3] ,
    \top_I.branch[5].block[12].um_I.iw[2] ,
    \top_I.branch[5].block[12].um_I.iw[1] ,
    \top_I.branch[5].block[12].um_I.clk ,
    \top_I.branch[5].block[11].um_I.iw[17] ,
    \top_I.branch[5].block[11].um_I.iw[16] ,
    \top_I.branch[5].block[11].um_I.iw[15] ,
    \top_I.branch[5].block[11].um_I.iw[14] ,
    \top_I.branch[5].block[11].um_I.iw[13] ,
    \top_I.branch[5].block[11].um_I.iw[12] ,
    \top_I.branch[5].block[11].um_I.iw[11] ,
    \top_I.branch[5].block[11].um_I.iw[10] ,
    \top_I.branch[5].block[11].um_I.iw[9] ,
    \top_I.branch[5].block[11].um_I.iw[8] ,
    \top_I.branch[5].block[11].um_I.iw[7] ,
    \top_I.branch[5].block[11].um_I.iw[6] ,
    \top_I.branch[5].block[11].um_I.iw[5] ,
    \top_I.branch[5].block[11].um_I.iw[4] ,
    \top_I.branch[5].block[11].um_I.iw[3] ,
    \top_I.branch[5].block[11].um_I.iw[2] ,
    \top_I.branch[5].block[11].um_I.iw[1] ,
    \top_I.branch[5].block[11].um_I.clk ,
    \top_I.branch[5].block[10].um_I.iw[17] ,
    \top_I.branch[5].block[10].um_I.iw[16] ,
    \top_I.branch[5].block[10].um_I.iw[15] ,
    \top_I.branch[5].block[10].um_I.iw[14] ,
    \top_I.branch[5].block[10].um_I.iw[13] ,
    \top_I.branch[5].block[10].um_I.iw[12] ,
    \top_I.branch[5].block[10].um_I.iw[11] ,
    \top_I.branch[5].block[10].um_I.iw[10] ,
    \top_I.branch[5].block[10].um_I.iw[9] ,
    \top_I.branch[5].block[10].um_I.iw[8] ,
    \top_I.branch[5].block[10].um_I.iw[7] ,
    \top_I.branch[5].block[10].um_I.iw[6] ,
    \top_I.branch[5].block[10].um_I.iw[5] ,
    \top_I.branch[5].block[10].um_I.iw[4] ,
    \top_I.branch[5].block[10].um_I.iw[3] ,
    \top_I.branch[5].block[10].um_I.iw[2] ,
    \top_I.branch[5].block[10].um_I.iw[1] ,
    \top_I.branch[5].block[10].um_I.clk ,
    \top_I.branch[5].block[9].um_I.iw[17] ,
    \top_I.branch[5].block[9].um_I.iw[16] ,
    \top_I.branch[5].block[9].um_I.iw[15] ,
    \top_I.branch[5].block[9].um_I.iw[14] ,
    \top_I.branch[5].block[9].um_I.iw[13] ,
    \top_I.branch[5].block[9].um_I.iw[12] ,
    \top_I.branch[5].block[9].um_I.iw[11] ,
    \top_I.branch[5].block[9].um_I.iw[10] ,
    \top_I.branch[5].block[9].um_I.iw[9] ,
    \top_I.branch[5].block[9].um_I.iw[8] ,
    \top_I.branch[5].block[9].um_I.iw[7] ,
    \top_I.branch[5].block[9].um_I.iw[6] ,
    \top_I.branch[5].block[9].um_I.iw[5] ,
    \top_I.branch[5].block[9].um_I.iw[4] ,
    \top_I.branch[5].block[9].um_I.iw[3] ,
    \top_I.branch[5].block[9].um_I.iw[2] ,
    \top_I.branch[5].block[9].um_I.iw[1] ,
    \top_I.branch[5].block[9].um_I.clk ,
    \top_I.branch[5].block[8].um_I.iw[17] ,
    \top_I.branch[5].block[8].um_I.iw[16] ,
    \top_I.branch[5].block[8].um_I.iw[15] ,
    \top_I.branch[5].block[8].um_I.iw[14] ,
    \top_I.branch[5].block[8].um_I.iw[13] ,
    \top_I.branch[5].block[8].um_I.iw[12] ,
    \top_I.branch[5].block[8].um_I.iw[11] ,
    \top_I.branch[5].block[8].um_I.iw[10] ,
    \top_I.branch[5].block[8].um_I.iw[9] ,
    \top_I.branch[5].block[8].um_I.iw[8] ,
    \top_I.branch[5].block[8].um_I.iw[7] ,
    \top_I.branch[5].block[8].um_I.iw[6] ,
    \top_I.branch[5].block[8].um_I.iw[5] ,
    \top_I.branch[5].block[8].um_I.iw[4] ,
    \top_I.branch[5].block[8].um_I.iw[3] ,
    \top_I.branch[5].block[8].um_I.iw[2] ,
    \top_I.branch[5].block[8].um_I.iw[1] ,
    \top_I.branch[5].block[8].um_I.clk ,
    \top_I.branch[5].block[7].um_I.iw[17] ,
    \top_I.branch[5].block[7].um_I.iw[16] ,
    \top_I.branch[5].block[7].um_I.iw[15] ,
    \top_I.branch[5].block[7].um_I.iw[14] ,
    \top_I.branch[5].block[7].um_I.iw[13] ,
    \top_I.branch[5].block[7].um_I.iw[12] ,
    \top_I.branch[5].block[7].um_I.iw[11] ,
    \top_I.branch[5].block[7].um_I.iw[10] ,
    \top_I.branch[5].block[7].um_I.iw[9] ,
    \top_I.branch[5].block[7].um_I.iw[8] ,
    \top_I.branch[5].block[7].um_I.iw[7] ,
    \top_I.branch[5].block[7].um_I.iw[6] ,
    \top_I.branch[5].block[7].um_I.iw[5] ,
    \top_I.branch[5].block[7].um_I.iw[4] ,
    \top_I.branch[5].block[7].um_I.iw[3] ,
    \top_I.branch[5].block[7].um_I.iw[2] ,
    \top_I.branch[5].block[7].um_I.iw[1] ,
    \top_I.branch[5].block[7].um_I.clk ,
    \top_I.branch[5].block[6].um_I.iw[17] ,
    \top_I.branch[5].block[6].um_I.iw[16] ,
    \top_I.branch[5].block[6].um_I.iw[15] ,
    \top_I.branch[5].block[6].um_I.iw[14] ,
    \top_I.branch[5].block[6].um_I.iw[13] ,
    \top_I.branch[5].block[6].um_I.iw[12] ,
    \top_I.branch[5].block[6].um_I.iw[11] ,
    \top_I.branch[5].block[6].um_I.iw[10] ,
    \top_I.branch[5].block[6].um_I.iw[9] ,
    \top_I.branch[5].block[6].um_I.iw[8] ,
    \top_I.branch[5].block[6].um_I.iw[7] ,
    \top_I.branch[5].block[6].um_I.iw[6] ,
    \top_I.branch[5].block[6].um_I.iw[5] ,
    \top_I.branch[5].block[6].um_I.iw[4] ,
    \top_I.branch[5].block[6].um_I.iw[3] ,
    \top_I.branch[5].block[6].um_I.iw[2] ,
    \top_I.branch[5].block[6].um_I.iw[1] ,
    \top_I.branch[5].block[6].um_I.clk ,
    \top_I.branch[5].block[5].um_I.iw[17] ,
    \top_I.branch[5].block[5].um_I.iw[16] ,
    \top_I.branch[5].block[5].um_I.iw[15] ,
    \top_I.branch[5].block[5].um_I.iw[14] ,
    \top_I.branch[5].block[5].um_I.iw[13] ,
    \top_I.branch[5].block[5].um_I.iw[12] ,
    \top_I.branch[5].block[5].um_I.iw[11] ,
    \top_I.branch[5].block[5].um_I.iw[10] ,
    \top_I.branch[5].block[5].um_I.iw[9] ,
    \top_I.branch[5].block[5].um_I.iw[8] ,
    \top_I.branch[5].block[5].um_I.iw[7] ,
    \top_I.branch[5].block[5].um_I.iw[6] ,
    \top_I.branch[5].block[5].um_I.iw[5] ,
    \top_I.branch[5].block[5].um_I.iw[4] ,
    \top_I.branch[5].block[5].um_I.iw[3] ,
    \top_I.branch[5].block[5].um_I.iw[2] ,
    \top_I.branch[5].block[5].um_I.iw[1] ,
    \top_I.branch[5].block[5].um_I.clk ,
    \top_I.branch[5].block[4].um_I.iw[17] ,
    \top_I.branch[5].block[4].um_I.iw[16] ,
    \top_I.branch[5].block[4].um_I.iw[15] ,
    \top_I.branch[5].block[4].um_I.iw[14] ,
    \top_I.branch[5].block[4].um_I.iw[13] ,
    \top_I.branch[5].block[4].um_I.iw[12] ,
    \top_I.branch[5].block[4].um_I.iw[11] ,
    \top_I.branch[5].block[4].um_I.iw[10] ,
    \top_I.branch[5].block[4].um_I.iw[9] ,
    \top_I.branch[5].block[4].um_I.iw[8] ,
    \top_I.branch[5].block[4].um_I.iw[7] ,
    \top_I.branch[5].block[4].um_I.iw[6] ,
    \top_I.branch[5].block[4].um_I.iw[5] ,
    \top_I.branch[5].block[4].um_I.iw[4] ,
    \top_I.branch[5].block[4].um_I.iw[3] ,
    \top_I.branch[5].block[4].um_I.iw[2] ,
    \top_I.branch[5].block[4].um_I.iw[1] ,
    \top_I.branch[5].block[4].um_I.clk ,
    \top_I.branch[5].block[3].um_I.iw[17] ,
    \top_I.branch[5].block[3].um_I.iw[16] ,
    \top_I.branch[5].block[3].um_I.iw[15] ,
    \top_I.branch[5].block[3].um_I.iw[14] ,
    \top_I.branch[5].block[3].um_I.iw[13] ,
    \top_I.branch[5].block[3].um_I.iw[12] ,
    \top_I.branch[5].block[3].um_I.iw[11] ,
    \top_I.branch[5].block[3].um_I.iw[10] ,
    \top_I.branch[5].block[3].um_I.iw[9] ,
    \top_I.branch[5].block[3].um_I.iw[8] ,
    \top_I.branch[5].block[3].um_I.iw[7] ,
    \top_I.branch[5].block[3].um_I.iw[6] ,
    \top_I.branch[5].block[3].um_I.iw[5] ,
    \top_I.branch[5].block[3].um_I.iw[4] ,
    \top_I.branch[5].block[3].um_I.iw[3] ,
    \top_I.branch[5].block[3].um_I.iw[2] ,
    \top_I.branch[5].block[3].um_I.iw[1] ,
    \top_I.branch[5].block[3].um_I.clk ,
    \top_I.branch[5].block[2].um_I.iw[17] ,
    \top_I.branch[5].block[2].um_I.iw[16] ,
    \top_I.branch[5].block[2].um_I.iw[15] ,
    \top_I.branch[5].block[2].um_I.iw[14] ,
    \top_I.branch[5].block[2].um_I.iw[13] ,
    \top_I.branch[5].block[2].um_I.iw[12] ,
    \top_I.branch[5].block[2].um_I.iw[11] ,
    \top_I.branch[5].block[2].um_I.iw[10] ,
    \top_I.branch[5].block[2].um_I.iw[9] ,
    \top_I.branch[5].block[2].um_I.iw[8] ,
    \top_I.branch[5].block[2].um_I.iw[7] ,
    \top_I.branch[5].block[2].um_I.iw[6] ,
    \top_I.branch[5].block[2].um_I.iw[5] ,
    \top_I.branch[5].block[2].um_I.iw[4] ,
    \top_I.branch[5].block[2].um_I.iw[3] ,
    \top_I.branch[5].block[2].um_I.iw[2] ,
    \top_I.branch[5].block[2].um_I.iw[1] ,
    \top_I.branch[5].block[2].um_I.clk ,
    \top_I.branch[5].block[1].um_I.iw[17] ,
    \top_I.branch[5].block[1].um_I.iw[16] ,
    \top_I.branch[5].block[1].um_I.iw[15] ,
    \top_I.branch[5].block[1].um_I.iw[14] ,
    \top_I.branch[5].block[1].um_I.iw[13] ,
    \top_I.branch[5].block[1].um_I.iw[12] ,
    \top_I.branch[5].block[1].um_I.iw[11] ,
    \top_I.branch[5].block[1].um_I.iw[10] ,
    \top_I.branch[5].block[1].um_I.iw[9] ,
    \top_I.branch[5].block[1].um_I.iw[8] ,
    \top_I.branch[5].block[1].um_I.iw[7] ,
    \top_I.branch[5].block[1].um_I.iw[6] ,
    \top_I.branch[5].block[1].um_I.iw[5] ,
    \top_I.branch[5].block[1].um_I.iw[4] ,
    \top_I.branch[5].block[1].um_I.iw[3] ,
    \top_I.branch[5].block[1].um_I.iw[2] ,
    \top_I.branch[5].block[1].um_I.iw[1] ,
    \top_I.branch[5].block[1].um_I.clk ,
    \top_I.branch[5].block[0].um_I.iw[17] ,
    \top_I.branch[5].block[0].um_I.iw[16] ,
    \top_I.branch[5].block[0].um_I.iw[15] ,
    \top_I.branch[5].block[0].um_I.iw[14] ,
    \top_I.branch[5].block[0].um_I.iw[13] ,
    \top_I.branch[5].block[0].um_I.iw[12] ,
    \top_I.branch[5].block[0].um_I.iw[11] ,
    \top_I.branch[5].block[0].um_I.iw[10] ,
    \top_I.branch[5].block[0].um_I.iw[9] ,
    \top_I.branch[5].block[0].um_I.iw[8] ,
    \top_I.branch[5].block[0].um_I.iw[7] ,
    \top_I.branch[5].block[0].um_I.iw[6] ,
    \top_I.branch[5].block[0].um_I.iw[5] ,
    \top_I.branch[5].block[0].um_I.iw[4] ,
    \top_I.branch[5].block[0].um_I.iw[3] ,
    \top_I.branch[5].block[0].um_I.iw[2] ,
    \top_I.branch[5].block[0].um_I.iw[1] ,
    \top_I.branch[5].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[5].block[15].um_I.pg_vdd ,
    \top_I.branch[5].block[14].um_I.pg_vdd ,
    \top_I.branch[5].block[13].um_I.pg_vdd ,
    \top_I.branch[5].block[12].um_I.pg_vdd ,
    \top_I.branch[5].block[11].um_I.pg_vdd ,
    \top_I.branch[5].block[10].um_I.pg_vdd ,
    \top_I.branch[5].block[9].um_I.pg_vdd ,
    \top_I.branch[5].block[8].um_I.pg_vdd ,
    \top_I.branch[5].block[7].um_I.pg_vdd ,
    \top_I.branch[5].block[6].um_I.pg_vdd ,
    \top_I.branch[5].block[5].um_I.pg_vdd ,
    \top_I.branch[5].block[4].um_I.pg_vdd ,
    \top_I.branch[5].block[3].um_I.pg_vdd ,
    \top_I.branch[5].block[2].um_I.pg_vdd ,
    \top_I.branch[5].block[1].um_I.pg_vdd ,
    \top_I.branch[5].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[6].mux_I  (.k_one(\top_I.branch[6].l_addr[0] ),
    .k_zero(\top_I.branch[6].l_addr[2] ),
    .addr({\top_I.branch[6].l_addr[2] ,
    \top_I.branch[6].l_addr[2] ,
    \top_I.branch[6].l_addr[0] ,
    \top_I.branch[6].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[6].block[15].um_I.ena ,
    \top_I.branch[6].block[14].um_I.ena ,
    \top_I.branch[6].block[13].um_I.ena ,
    \top_I.branch[6].block[12].um_I.ena ,
    \top_I.branch[6].block[11].um_I.ena ,
    \top_I.branch[6].block[10].um_I.ena ,
    \top_I.branch[6].block[9].um_I.ena ,
    \top_I.branch[6].block[8].um_I.ena ,
    \top_I.branch[6].block[7].um_I.ena ,
    \top_I.branch[6].block[6].um_I.ena ,
    \top_I.branch[6].block[5].um_I.ena ,
    \top_I.branch[6].block[4].um_I.ena ,
    \top_I.branch[6].block[3].um_I.ena ,
    \top_I.branch[6].block[2].um_I.ena ,
    \top_I.branch[6].block[1].um_I.ena ,
    \top_I.branch[6].block[0].um_I.ena }),
    .um_iw({\top_I.branch[6].block[15].um_I.iw[17] ,
    \top_I.branch[6].block[15].um_I.iw[16] ,
    \top_I.branch[6].block[15].um_I.iw[15] ,
    \top_I.branch[6].block[15].um_I.iw[14] ,
    \top_I.branch[6].block[15].um_I.iw[13] ,
    \top_I.branch[6].block[15].um_I.iw[12] ,
    \top_I.branch[6].block[15].um_I.iw[11] ,
    \top_I.branch[6].block[15].um_I.iw[10] ,
    \top_I.branch[6].block[15].um_I.iw[9] ,
    \top_I.branch[6].block[15].um_I.iw[8] ,
    \top_I.branch[6].block[15].um_I.iw[7] ,
    \top_I.branch[6].block[15].um_I.iw[6] ,
    \top_I.branch[6].block[15].um_I.iw[5] ,
    \top_I.branch[6].block[15].um_I.iw[4] ,
    \top_I.branch[6].block[15].um_I.iw[3] ,
    \top_I.branch[6].block[15].um_I.iw[2] ,
    \top_I.branch[6].block[15].um_I.iw[1] ,
    \top_I.branch[6].block[15].um_I.clk ,
    \top_I.branch[6].block[14].um_I.iw[17] ,
    \top_I.branch[6].block[14].um_I.iw[16] ,
    \top_I.branch[6].block[14].um_I.iw[15] ,
    \top_I.branch[6].block[14].um_I.iw[14] ,
    \top_I.branch[6].block[14].um_I.iw[13] ,
    \top_I.branch[6].block[14].um_I.iw[12] ,
    \top_I.branch[6].block[14].um_I.iw[11] ,
    \top_I.branch[6].block[14].um_I.iw[10] ,
    \top_I.branch[6].block[14].um_I.iw[9] ,
    \top_I.branch[6].block[14].um_I.iw[8] ,
    \top_I.branch[6].block[14].um_I.iw[7] ,
    \top_I.branch[6].block[14].um_I.iw[6] ,
    \top_I.branch[6].block[14].um_I.iw[5] ,
    \top_I.branch[6].block[14].um_I.iw[4] ,
    \top_I.branch[6].block[14].um_I.iw[3] ,
    \top_I.branch[6].block[14].um_I.iw[2] ,
    \top_I.branch[6].block[14].um_I.iw[1] ,
    \top_I.branch[6].block[14].um_I.clk ,
    \top_I.branch[6].block[13].um_I.iw[17] ,
    \top_I.branch[6].block[13].um_I.iw[16] ,
    \top_I.branch[6].block[13].um_I.iw[15] ,
    \top_I.branch[6].block[13].um_I.iw[14] ,
    \top_I.branch[6].block[13].um_I.iw[13] ,
    \top_I.branch[6].block[13].um_I.iw[12] ,
    \top_I.branch[6].block[13].um_I.iw[11] ,
    \top_I.branch[6].block[13].um_I.iw[10] ,
    \top_I.branch[6].block[13].um_I.iw[9] ,
    \top_I.branch[6].block[13].um_I.iw[8] ,
    \top_I.branch[6].block[13].um_I.iw[7] ,
    \top_I.branch[6].block[13].um_I.iw[6] ,
    \top_I.branch[6].block[13].um_I.iw[5] ,
    \top_I.branch[6].block[13].um_I.iw[4] ,
    \top_I.branch[6].block[13].um_I.iw[3] ,
    \top_I.branch[6].block[13].um_I.iw[2] ,
    \top_I.branch[6].block[13].um_I.iw[1] ,
    \top_I.branch[6].block[13].um_I.clk ,
    \top_I.branch[6].block[12].um_I.iw[17] ,
    \top_I.branch[6].block[12].um_I.iw[16] ,
    \top_I.branch[6].block[12].um_I.iw[15] ,
    \top_I.branch[6].block[12].um_I.iw[14] ,
    \top_I.branch[6].block[12].um_I.iw[13] ,
    \top_I.branch[6].block[12].um_I.iw[12] ,
    \top_I.branch[6].block[12].um_I.iw[11] ,
    \top_I.branch[6].block[12].um_I.iw[10] ,
    \top_I.branch[6].block[12].um_I.iw[9] ,
    \top_I.branch[6].block[12].um_I.iw[8] ,
    \top_I.branch[6].block[12].um_I.iw[7] ,
    \top_I.branch[6].block[12].um_I.iw[6] ,
    \top_I.branch[6].block[12].um_I.iw[5] ,
    \top_I.branch[6].block[12].um_I.iw[4] ,
    \top_I.branch[6].block[12].um_I.iw[3] ,
    \top_I.branch[6].block[12].um_I.iw[2] ,
    \top_I.branch[6].block[12].um_I.iw[1] ,
    \top_I.branch[6].block[12].um_I.clk ,
    \top_I.branch[6].block[11].um_I.iw[17] ,
    \top_I.branch[6].block[11].um_I.iw[16] ,
    \top_I.branch[6].block[11].um_I.iw[15] ,
    \top_I.branch[6].block[11].um_I.iw[14] ,
    \top_I.branch[6].block[11].um_I.iw[13] ,
    \top_I.branch[6].block[11].um_I.iw[12] ,
    \top_I.branch[6].block[11].um_I.iw[11] ,
    \top_I.branch[6].block[11].um_I.iw[10] ,
    \top_I.branch[6].block[11].um_I.iw[9] ,
    \top_I.branch[6].block[11].um_I.iw[8] ,
    \top_I.branch[6].block[11].um_I.iw[7] ,
    \top_I.branch[6].block[11].um_I.iw[6] ,
    \top_I.branch[6].block[11].um_I.iw[5] ,
    \top_I.branch[6].block[11].um_I.iw[4] ,
    \top_I.branch[6].block[11].um_I.iw[3] ,
    \top_I.branch[6].block[11].um_I.iw[2] ,
    \top_I.branch[6].block[11].um_I.iw[1] ,
    \top_I.branch[6].block[11].um_I.clk ,
    \top_I.branch[6].block[10].um_I.iw[17] ,
    \top_I.branch[6].block[10].um_I.iw[16] ,
    \top_I.branch[6].block[10].um_I.iw[15] ,
    \top_I.branch[6].block[10].um_I.iw[14] ,
    \top_I.branch[6].block[10].um_I.iw[13] ,
    \top_I.branch[6].block[10].um_I.iw[12] ,
    \top_I.branch[6].block[10].um_I.iw[11] ,
    \top_I.branch[6].block[10].um_I.iw[10] ,
    \top_I.branch[6].block[10].um_I.iw[9] ,
    \top_I.branch[6].block[10].um_I.iw[8] ,
    \top_I.branch[6].block[10].um_I.iw[7] ,
    \top_I.branch[6].block[10].um_I.iw[6] ,
    \top_I.branch[6].block[10].um_I.iw[5] ,
    \top_I.branch[6].block[10].um_I.iw[4] ,
    \top_I.branch[6].block[10].um_I.iw[3] ,
    \top_I.branch[6].block[10].um_I.iw[2] ,
    \top_I.branch[6].block[10].um_I.iw[1] ,
    \top_I.branch[6].block[10].um_I.clk ,
    \top_I.branch[6].block[9].um_I.iw[17] ,
    \top_I.branch[6].block[9].um_I.iw[16] ,
    \top_I.branch[6].block[9].um_I.iw[15] ,
    \top_I.branch[6].block[9].um_I.iw[14] ,
    \top_I.branch[6].block[9].um_I.iw[13] ,
    \top_I.branch[6].block[9].um_I.iw[12] ,
    \top_I.branch[6].block[9].um_I.iw[11] ,
    \top_I.branch[6].block[9].um_I.iw[10] ,
    \top_I.branch[6].block[9].um_I.iw[9] ,
    \top_I.branch[6].block[9].um_I.iw[8] ,
    \top_I.branch[6].block[9].um_I.iw[7] ,
    \top_I.branch[6].block[9].um_I.iw[6] ,
    \top_I.branch[6].block[9].um_I.iw[5] ,
    \top_I.branch[6].block[9].um_I.iw[4] ,
    \top_I.branch[6].block[9].um_I.iw[3] ,
    \top_I.branch[6].block[9].um_I.iw[2] ,
    \top_I.branch[6].block[9].um_I.iw[1] ,
    \top_I.branch[6].block[9].um_I.clk ,
    \top_I.branch[6].block[8].um_I.iw[17] ,
    \top_I.branch[6].block[8].um_I.iw[16] ,
    \top_I.branch[6].block[8].um_I.iw[15] ,
    \top_I.branch[6].block[8].um_I.iw[14] ,
    \top_I.branch[6].block[8].um_I.iw[13] ,
    \top_I.branch[6].block[8].um_I.iw[12] ,
    \top_I.branch[6].block[8].um_I.iw[11] ,
    \top_I.branch[6].block[8].um_I.iw[10] ,
    \top_I.branch[6].block[8].um_I.iw[9] ,
    \top_I.branch[6].block[8].um_I.iw[8] ,
    \top_I.branch[6].block[8].um_I.iw[7] ,
    \top_I.branch[6].block[8].um_I.iw[6] ,
    \top_I.branch[6].block[8].um_I.iw[5] ,
    \top_I.branch[6].block[8].um_I.iw[4] ,
    \top_I.branch[6].block[8].um_I.iw[3] ,
    \top_I.branch[6].block[8].um_I.iw[2] ,
    \top_I.branch[6].block[8].um_I.iw[1] ,
    \top_I.branch[6].block[8].um_I.clk ,
    \top_I.branch[6].block[7].um_I.iw[17] ,
    \top_I.branch[6].block[7].um_I.iw[16] ,
    \top_I.branch[6].block[7].um_I.iw[15] ,
    \top_I.branch[6].block[7].um_I.iw[14] ,
    \top_I.branch[6].block[7].um_I.iw[13] ,
    \top_I.branch[6].block[7].um_I.iw[12] ,
    \top_I.branch[6].block[7].um_I.iw[11] ,
    \top_I.branch[6].block[7].um_I.iw[10] ,
    \top_I.branch[6].block[7].um_I.iw[9] ,
    \top_I.branch[6].block[7].um_I.iw[8] ,
    \top_I.branch[6].block[7].um_I.iw[7] ,
    \top_I.branch[6].block[7].um_I.iw[6] ,
    \top_I.branch[6].block[7].um_I.iw[5] ,
    \top_I.branch[6].block[7].um_I.iw[4] ,
    \top_I.branch[6].block[7].um_I.iw[3] ,
    \top_I.branch[6].block[7].um_I.iw[2] ,
    \top_I.branch[6].block[7].um_I.iw[1] ,
    \top_I.branch[6].block[7].um_I.clk ,
    \top_I.branch[6].block[6].um_I.iw[17] ,
    \top_I.branch[6].block[6].um_I.iw[16] ,
    \top_I.branch[6].block[6].um_I.iw[15] ,
    \top_I.branch[6].block[6].um_I.iw[14] ,
    \top_I.branch[6].block[6].um_I.iw[13] ,
    \top_I.branch[6].block[6].um_I.iw[12] ,
    \top_I.branch[6].block[6].um_I.iw[11] ,
    \top_I.branch[6].block[6].um_I.iw[10] ,
    \top_I.branch[6].block[6].um_I.iw[9] ,
    \top_I.branch[6].block[6].um_I.iw[8] ,
    \top_I.branch[6].block[6].um_I.iw[7] ,
    \top_I.branch[6].block[6].um_I.iw[6] ,
    \top_I.branch[6].block[6].um_I.iw[5] ,
    \top_I.branch[6].block[6].um_I.iw[4] ,
    \top_I.branch[6].block[6].um_I.iw[3] ,
    \top_I.branch[6].block[6].um_I.iw[2] ,
    \top_I.branch[6].block[6].um_I.iw[1] ,
    \top_I.branch[6].block[6].um_I.clk ,
    \top_I.branch[6].block[5].um_I.iw[17] ,
    \top_I.branch[6].block[5].um_I.iw[16] ,
    \top_I.branch[6].block[5].um_I.iw[15] ,
    \top_I.branch[6].block[5].um_I.iw[14] ,
    \top_I.branch[6].block[5].um_I.iw[13] ,
    \top_I.branch[6].block[5].um_I.iw[12] ,
    \top_I.branch[6].block[5].um_I.iw[11] ,
    \top_I.branch[6].block[5].um_I.iw[10] ,
    \top_I.branch[6].block[5].um_I.iw[9] ,
    \top_I.branch[6].block[5].um_I.iw[8] ,
    \top_I.branch[6].block[5].um_I.iw[7] ,
    \top_I.branch[6].block[5].um_I.iw[6] ,
    \top_I.branch[6].block[5].um_I.iw[5] ,
    \top_I.branch[6].block[5].um_I.iw[4] ,
    \top_I.branch[6].block[5].um_I.iw[3] ,
    \top_I.branch[6].block[5].um_I.iw[2] ,
    \top_I.branch[6].block[5].um_I.iw[1] ,
    \top_I.branch[6].block[5].um_I.clk ,
    \top_I.branch[6].block[4].um_I.iw[17] ,
    \top_I.branch[6].block[4].um_I.iw[16] ,
    \top_I.branch[6].block[4].um_I.iw[15] ,
    \top_I.branch[6].block[4].um_I.iw[14] ,
    \top_I.branch[6].block[4].um_I.iw[13] ,
    \top_I.branch[6].block[4].um_I.iw[12] ,
    \top_I.branch[6].block[4].um_I.iw[11] ,
    \top_I.branch[6].block[4].um_I.iw[10] ,
    \top_I.branch[6].block[4].um_I.iw[9] ,
    \top_I.branch[6].block[4].um_I.iw[8] ,
    \top_I.branch[6].block[4].um_I.iw[7] ,
    \top_I.branch[6].block[4].um_I.iw[6] ,
    \top_I.branch[6].block[4].um_I.iw[5] ,
    \top_I.branch[6].block[4].um_I.iw[4] ,
    \top_I.branch[6].block[4].um_I.iw[3] ,
    \top_I.branch[6].block[4].um_I.iw[2] ,
    \top_I.branch[6].block[4].um_I.iw[1] ,
    \top_I.branch[6].block[4].um_I.clk ,
    \top_I.branch[6].block[3].um_I.iw[17] ,
    \top_I.branch[6].block[3].um_I.iw[16] ,
    \top_I.branch[6].block[3].um_I.iw[15] ,
    \top_I.branch[6].block[3].um_I.iw[14] ,
    \top_I.branch[6].block[3].um_I.iw[13] ,
    \top_I.branch[6].block[3].um_I.iw[12] ,
    \top_I.branch[6].block[3].um_I.iw[11] ,
    \top_I.branch[6].block[3].um_I.iw[10] ,
    \top_I.branch[6].block[3].um_I.iw[9] ,
    \top_I.branch[6].block[3].um_I.iw[8] ,
    \top_I.branch[6].block[3].um_I.iw[7] ,
    \top_I.branch[6].block[3].um_I.iw[6] ,
    \top_I.branch[6].block[3].um_I.iw[5] ,
    \top_I.branch[6].block[3].um_I.iw[4] ,
    \top_I.branch[6].block[3].um_I.iw[3] ,
    \top_I.branch[6].block[3].um_I.iw[2] ,
    \top_I.branch[6].block[3].um_I.iw[1] ,
    \top_I.branch[6].block[3].um_I.clk ,
    \top_I.branch[6].block[2].um_I.iw[17] ,
    \top_I.branch[6].block[2].um_I.iw[16] ,
    \top_I.branch[6].block[2].um_I.iw[15] ,
    \top_I.branch[6].block[2].um_I.iw[14] ,
    \top_I.branch[6].block[2].um_I.iw[13] ,
    \top_I.branch[6].block[2].um_I.iw[12] ,
    \top_I.branch[6].block[2].um_I.iw[11] ,
    \top_I.branch[6].block[2].um_I.iw[10] ,
    \top_I.branch[6].block[2].um_I.iw[9] ,
    \top_I.branch[6].block[2].um_I.iw[8] ,
    \top_I.branch[6].block[2].um_I.iw[7] ,
    \top_I.branch[6].block[2].um_I.iw[6] ,
    \top_I.branch[6].block[2].um_I.iw[5] ,
    \top_I.branch[6].block[2].um_I.iw[4] ,
    \top_I.branch[6].block[2].um_I.iw[3] ,
    \top_I.branch[6].block[2].um_I.iw[2] ,
    \top_I.branch[6].block[2].um_I.iw[1] ,
    \top_I.branch[6].block[2].um_I.clk ,
    \top_I.branch[6].block[1].um_I.iw[17] ,
    \top_I.branch[6].block[1].um_I.iw[16] ,
    \top_I.branch[6].block[1].um_I.iw[15] ,
    \top_I.branch[6].block[1].um_I.iw[14] ,
    \top_I.branch[6].block[1].um_I.iw[13] ,
    \top_I.branch[6].block[1].um_I.iw[12] ,
    \top_I.branch[6].block[1].um_I.iw[11] ,
    \top_I.branch[6].block[1].um_I.iw[10] ,
    \top_I.branch[6].block[1].um_I.iw[9] ,
    \top_I.branch[6].block[1].um_I.iw[8] ,
    \top_I.branch[6].block[1].um_I.iw[7] ,
    \top_I.branch[6].block[1].um_I.iw[6] ,
    \top_I.branch[6].block[1].um_I.iw[5] ,
    \top_I.branch[6].block[1].um_I.iw[4] ,
    \top_I.branch[6].block[1].um_I.iw[3] ,
    \top_I.branch[6].block[1].um_I.iw[2] ,
    \top_I.branch[6].block[1].um_I.iw[1] ,
    \top_I.branch[6].block[1].um_I.clk ,
    \top_I.branch[6].block[0].um_I.iw[17] ,
    \top_I.branch[6].block[0].um_I.iw[16] ,
    \top_I.branch[6].block[0].um_I.iw[15] ,
    \top_I.branch[6].block[0].um_I.iw[14] ,
    \top_I.branch[6].block[0].um_I.iw[13] ,
    \top_I.branch[6].block[0].um_I.iw[12] ,
    \top_I.branch[6].block[0].um_I.iw[11] ,
    \top_I.branch[6].block[0].um_I.iw[10] ,
    \top_I.branch[6].block[0].um_I.iw[9] ,
    \top_I.branch[6].block[0].um_I.iw[8] ,
    \top_I.branch[6].block[0].um_I.iw[7] ,
    \top_I.branch[6].block[0].um_I.iw[6] ,
    \top_I.branch[6].block[0].um_I.iw[5] ,
    \top_I.branch[6].block[0].um_I.iw[4] ,
    \top_I.branch[6].block[0].um_I.iw[3] ,
    \top_I.branch[6].block[0].um_I.iw[2] ,
    \top_I.branch[6].block[0].um_I.iw[1] ,
    \top_I.branch[6].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[6].block[15].um_I.pg_vdd ,
    \top_I.branch[6].block[14].um_I.pg_vdd ,
    \top_I.branch[6].block[13].um_I.pg_vdd ,
    \top_I.branch[6].block[12].um_I.pg_vdd ,
    \top_I.branch[6].block[11].um_I.pg_vdd ,
    \top_I.branch[6].block[10].um_I.pg_vdd ,
    \top_I.branch[6].block[9].um_I.pg_vdd ,
    \top_I.branch[6].block[8].um_I.pg_vdd ,
    \top_I.branch[6].block[7].um_I.pg_vdd ,
    \top_I.branch[6].block[6].um_I.pg_vdd ,
    \top_I.branch[6].block[5].um_I.pg_vdd ,
    \top_I.branch[6].block[4].um_I.pg_vdd ,
    \top_I.branch[6].block[3].um_I.pg_vdd ,
    \top_I.branch[6].block[2].um_I.pg_vdd ,
    \top_I.branch[6].block[1].um_I.pg_vdd ,
    \top_I.branch[6].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[7].mux_I  (.k_one(\top_I.branch[7].l_addr[0] ),
    .k_zero(\top_I.branch[7].l_addr[2] ),
    .addr({\top_I.branch[7].l_addr[2] ,
    \top_I.branch[7].l_addr[2] ,
    \top_I.branch[7].l_addr[0] ,
    \top_I.branch[7].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[7].block[15].um_I.ena ,
    \top_I.branch[7].block[14].um_I.ena ,
    \top_I.branch[7].block[13].um_I.ena ,
    \top_I.branch[7].block[12].um_I.ena ,
    \top_I.branch[7].block[11].um_I.ena ,
    \top_I.branch[7].block[10].um_I.ena ,
    \top_I.branch[7].block[9].um_I.ena ,
    \top_I.branch[7].block[8].um_I.ena ,
    \top_I.branch[7].block[7].um_I.ena ,
    \top_I.branch[7].block[6].um_I.ena ,
    \top_I.branch[7].block[5].um_I.ena ,
    \top_I.branch[7].block[4].um_I.ena ,
    \top_I.branch[7].block[3].um_I.ena ,
    \top_I.branch[7].block[2].um_I.ena ,
    \top_I.branch[7].block[1].um_I.ena ,
    \top_I.branch[7].block[0].um_I.ena }),
    .um_iw({\top_I.branch[7].block[15].um_I.iw[17] ,
    \top_I.branch[7].block[15].um_I.iw[16] ,
    \top_I.branch[7].block[15].um_I.iw[15] ,
    \top_I.branch[7].block[15].um_I.iw[14] ,
    \top_I.branch[7].block[15].um_I.iw[13] ,
    \top_I.branch[7].block[15].um_I.iw[12] ,
    \top_I.branch[7].block[15].um_I.iw[11] ,
    \top_I.branch[7].block[15].um_I.iw[10] ,
    \top_I.branch[7].block[15].um_I.iw[9] ,
    \top_I.branch[7].block[15].um_I.iw[8] ,
    \top_I.branch[7].block[15].um_I.iw[7] ,
    \top_I.branch[7].block[15].um_I.iw[6] ,
    \top_I.branch[7].block[15].um_I.iw[5] ,
    \top_I.branch[7].block[15].um_I.iw[4] ,
    \top_I.branch[7].block[15].um_I.iw[3] ,
    \top_I.branch[7].block[15].um_I.iw[2] ,
    \top_I.branch[7].block[15].um_I.iw[1] ,
    \top_I.branch[7].block[15].um_I.clk ,
    \top_I.branch[7].block[14].um_I.iw[17] ,
    \top_I.branch[7].block[14].um_I.iw[16] ,
    \top_I.branch[7].block[14].um_I.iw[15] ,
    \top_I.branch[7].block[14].um_I.iw[14] ,
    \top_I.branch[7].block[14].um_I.iw[13] ,
    \top_I.branch[7].block[14].um_I.iw[12] ,
    \top_I.branch[7].block[14].um_I.iw[11] ,
    \top_I.branch[7].block[14].um_I.iw[10] ,
    \top_I.branch[7].block[14].um_I.iw[9] ,
    \top_I.branch[7].block[14].um_I.iw[8] ,
    \top_I.branch[7].block[14].um_I.iw[7] ,
    \top_I.branch[7].block[14].um_I.iw[6] ,
    \top_I.branch[7].block[14].um_I.iw[5] ,
    \top_I.branch[7].block[14].um_I.iw[4] ,
    \top_I.branch[7].block[14].um_I.iw[3] ,
    \top_I.branch[7].block[14].um_I.iw[2] ,
    \top_I.branch[7].block[14].um_I.iw[1] ,
    \top_I.branch[7].block[14].um_I.clk ,
    \top_I.branch[7].block[13].um_I.iw[17] ,
    \top_I.branch[7].block[13].um_I.iw[16] ,
    \top_I.branch[7].block[13].um_I.iw[15] ,
    \top_I.branch[7].block[13].um_I.iw[14] ,
    \top_I.branch[7].block[13].um_I.iw[13] ,
    \top_I.branch[7].block[13].um_I.iw[12] ,
    \top_I.branch[7].block[13].um_I.iw[11] ,
    \top_I.branch[7].block[13].um_I.iw[10] ,
    \top_I.branch[7].block[13].um_I.iw[9] ,
    \top_I.branch[7].block[13].um_I.iw[8] ,
    \top_I.branch[7].block[13].um_I.iw[7] ,
    \top_I.branch[7].block[13].um_I.iw[6] ,
    \top_I.branch[7].block[13].um_I.iw[5] ,
    \top_I.branch[7].block[13].um_I.iw[4] ,
    \top_I.branch[7].block[13].um_I.iw[3] ,
    \top_I.branch[7].block[13].um_I.iw[2] ,
    \top_I.branch[7].block[13].um_I.iw[1] ,
    \top_I.branch[7].block[13].um_I.clk ,
    \top_I.branch[7].block[12].um_I.iw[17] ,
    \top_I.branch[7].block[12].um_I.iw[16] ,
    \top_I.branch[7].block[12].um_I.iw[15] ,
    \top_I.branch[7].block[12].um_I.iw[14] ,
    \top_I.branch[7].block[12].um_I.iw[13] ,
    \top_I.branch[7].block[12].um_I.iw[12] ,
    \top_I.branch[7].block[12].um_I.iw[11] ,
    \top_I.branch[7].block[12].um_I.iw[10] ,
    \top_I.branch[7].block[12].um_I.iw[9] ,
    \top_I.branch[7].block[12].um_I.iw[8] ,
    \top_I.branch[7].block[12].um_I.iw[7] ,
    \top_I.branch[7].block[12].um_I.iw[6] ,
    \top_I.branch[7].block[12].um_I.iw[5] ,
    \top_I.branch[7].block[12].um_I.iw[4] ,
    \top_I.branch[7].block[12].um_I.iw[3] ,
    \top_I.branch[7].block[12].um_I.iw[2] ,
    \top_I.branch[7].block[12].um_I.iw[1] ,
    \top_I.branch[7].block[12].um_I.clk ,
    \top_I.branch[7].block[11].um_I.iw[17] ,
    \top_I.branch[7].block[11].um_I.iw[16] ,
    \top_I.branch[7].block[11].um_I.iw[15] ,
    \top_I.branch[7].block[11].um_I.iw[14] ,
    \top_I.branch[7].block[11].um_I.iw[13] ,
    \top_I.branch[7].block[11].um_I.iw[12] ,
    \top_I.branch[7].block[11].um_I.iw[11] ,
    \top_I.branch[7].block[11].um_I.iw[10] ,
    \top_I.branch[7].block[11].um_I.iw[9] ,
    \top_I.branch[7].block[11].um_I.iw[8] ,
    \top_I.branch[7].block[11].um_I.iw[7] ,
    \top_I.branch[7].block[11].um_I.iw[6] ,
    \top_I.branch[7].block[11].um_I.iw[5] ,
    \top_I.branch[7].block[11].um_I.iw[4] ,
    \top_I.branch[7].block[11].um_I.iw[3] ,
    \top_I.branch[7].block[11].um_I.iw[2] ,
    \top_I.branch[7].block[11].um_I.iw[1] ,
    \top_I.branch[7].block[11].um_I.clk ,
    \top_I.branch[7].block[10].um_I.iw[17] ,
    \top_I.branch[7].block[10].um_I.iw[16] ,
    \top_I.branch[7].block[10].um_I.iw[15] ,
    \top_I.branch[7].block[10].um_I.iw[14] ,
    \top_I.branch[7].block[10].um_I.iw[13] ,
    \top_I.branch[7].block[10].um_I.iw[12] ,
    \top_I.branch[7].block[10].um_I.iw[11] ,
    \top_I.branch[7].block[10].um_I.iw[10] ,
    \top_I.branch[7].block[10].um_I.iw[9] ,
    \top_I.branch[7].block[10].um_I.iw[8] ,
    \top_I.branch[7].block[10].um_I.iw[7] ,
    \top_I.branch[7].block[10].um_I.iw[6] ,
    \top_I.branch[7].block[10].um_I.iw[5] ,
    \top_I.branch[7].block[10].um_I.iw[4] ,
    \top_I.branch[7].block[10].um_I.iw[3] ,
    \top_I.branch[7].block[10].um_I.iw[2] ,
    \top_I.branch[7].block[10].um_I.iw[1] ,
    \top_I.branch[7].block[10].um_I.clk ,
    \top_I.branch[7].block[9].um_I.iw[17] ,
    \top_I.branch[7].block[9].um_I.iw[16] ,
    \top_I.branch[7].block[9].um_I.iw[15] ,
    \top_I.branch[7].block[9].um_I.iw[14] ,
    \top_I.branch[7].block[9].um_I.iw[13] ,
    \top_I.branch[7].block[9].um_I.iw[12] ,
    \top_I.branch[7].block[9].um_I.iw[11] ,
    \top_I.branch[7].block[9].um_I.iw[10] ,
    \top_I.branch[7].block[9].um_I.iw[9] ,
    \top_I.branch[7].block[9].um_I.iw[8] ,
    \top_I.branch[7].block[9].um_I.iw[7] ,
    \top_I.branch[7].block[9].um_I.iw[6] ,
    \top_I.branch[7].block[9].um_I.iw[5] ,
    \top_I.branch[7].block[9].um_I.iw[4] ,
    \top_I.branch[7].block[9].um_I.iw[3] ,
    \top_I.branch[7].block[9].um_I.iw[2] ,
    \top_I.branch[7].block[9].um_I.iw[1] ,
    \top_I.branch[7].block[9].um_I.clk ,
    \top_I.branch[7].block[8].um_I.iw[17] ,
    \top_I.branch[7].block[8].um_I.iw[16] ,
    \top_I.branch[7].block[8].um_I.iw[15] ,
    \top_I.branch[7].block[8].um_I.iw[14] ,
    \top_I.branch[7].block[8].um_I.iw[13] ,
    \top_I.branch[7].block[8].um_I.iw[12] ,
    \top_I.branch[7].block[8].um_I.iw[11] ,
    \top_I.branch[7].block[8].um_I.iw[10] ,
    \top_I.branch[7].block[8].um_I.iw[9] ,
    \top_I.branch[7].block[8].um_I.iw[8] ,
    \top_I.branch[7].block[8].um_I.iw[7] ,
    \top_I.branch[7].block[8].um_I.iw[6] ,
    \top_I.branch[7].block[8].um_I.iw[5] ,
    \top_I.branch[7].block[8].um_I.iw[4] ,
    \top_I.branch[7].block[8].um_I.iw[3] ,
    \top_I.branch[7].block[8].um_I.iw[2] ,
    \top_I.branch[7].block[8].um_I.iw[1] ,
    \top_I.branch[7].block[8].um_I.clk ,
    \top_I.branch[7].block[7].um_I.iw[17] ,
    \top_I.branch[7].block[7].um_I.iw[16] ,
    \top_I.branch[7].block[7].um_I.iw[15] ,
    \top_I.branch[7].block[7].um_I.iw[14] ,
    \top_I.branch[7].block[7].um_I.iw[13] ,
    \top_I.branch[7].block[7].um_I.iw[12] ,
    \top_I.branch[7].block[7].um_I.iw[11] ,
    \top_I.branch[7].block[7].um_I.iw[10] ,
    \top_I.branch[7].block[7].um_I.iw[9] ,
    \top_I.branch[7].block[7].um_I.iw[8] ,
    \top_I.branch[7].block[7].um_I.iw[7] ,
    \top_I.branch[7].block[7].um_I.iw[6] ,
    \top_I.branch[7].block[7].um_I.iw[5] ,
    \top_I.branch[7].block[7].um_I.iw[4] ,
    \top_I.branch[7].block[7].um_I.iw[3] ,
    \top_I.branch[7].block[7].um_I.iw[2] ,
    \top_I.branch[7].block[7].um_I.iw[1] ,
    \top_I.branch[7].block[7].um_I.clk ,
    \top_I.branch[7].block[6].um_I.iw[17] ,
    \top_I.branch[7].block[6].um_I.iw[16] ,
    \top_I.branch[7].block[6].um_I.iw[15] ,
    \top_I.branch[7].block[6].um_I.iw[14] ,
    \top_I.branch[7].block[6].um_I.iw[13] ,
    \top_I.branch[7].block[6].um_I.iw[12] ,
    \top_I.branch[7].block[6].um_I.iw[11] ,
    \top_I.branch[7].block[6].um_I.iw[10] ,
    \top_I.branch[7].block[6].um_I.iw[9] ,
    \top_I.branch[7].block[6].um_I.iw[8] ,
    \top_I.branch[7].block[6].um_I.iw[7] ,
    \top_I.branch[7].block[6].um_I.iw[6] ,
    \top_I.branch[7].block[6].um_I.iw[5] ,
    \top_I.branch[7].block[6].um_I.iw[4] ,
    \top_I.branch[7].block[6].um_I.iw[3] ,
    \top_I.branch[7].block[6].um_I.iw[2] ,
    \top_I.branch[7].block[6].um_I.iw[1] ,
    \top_I.branch[7].block[6].um_I.clk ,
    \top_I.branch[7].block[5].um_I.iw[17] ,
    \top_I.branch[7].block[5].um_I.iw[16] ,
    \top_I.branch[7].block[5].um_I.iw[15] ,
    \top_I.branch[7].block[5].um_I.iw[14] ,
    \top_I.branch[7].block[5].um_I.iw[13] ,
    \top_I.branch[7].block[5].um_I.iw[12] ,
    \top_I.branch[7].block[5].um_I.iw[11] ,
    \top_I.branch[7].block[5].um_I.iw[10] ,
    \top_I.branch[7].block[5].um_I.iw[9] ,
    \top_I.branch[7].block[5].um_I.iw[8] ,
    \top_I.branch[7].block[5].um_I.iw[7] ,
    \top_I.branch[7].block[5].um_I.iw[6] ,
    \top_I.branch[7].block[5].um_I.iw[5] ,
    \top_I.branch[7].block[5].um_I.iw[4] ,
    \top_I.branch[7].block[5].um_I.iw[3] ,
    \top_I.branch[7].block[5].um_I.iw[2] ,
    \top_I.branch[7].block[5].um_I.iw[1] ,
    \top_I.branch[7].block[5].um_I.clk ,
    \top_I.branch[7].block[4].um_I.iw[17] ,
    \top_I.branch[7].block[4].um_I.iw[16] ,
    \top_I.branch[7].block[4].um_I.iw[15] ,
    \top_I.branch[7].block[4].um_I.iw[14] ,
    \top_I.branch[7].block[4].um_I.iw[13] ,
    \top_I.branch[7].block[4].um_I.iw[12] ,
    \top_I.branch[7].block[4].um_I.iw[11] ,
    \top_I.branch[7].block[4].um_I.iw[10] ,
    \top_I.branch[7].block[4].um_I.iw[9] ,
    \top_I.branch[7].block[4].um_I.iw[8] ,
    \top_I.branch[7].block[4].um_I.iw[7] ,
    \top_I.branch[7].block[4].um_I.iw[6] ,
    \top_I.branch[7].block[4].um_I.iw[5] ,
    \top_I.branch[7].block[4].um_I.iw[4] ,
    \top_I.branch[7].block[4].um_I.iw[3] ,
    \top_I.branch[7].block[4].um_I.iw[2] ,
    \top_I.branch[7].block[4].um_I.iw[1] ,
    \top_I.branch[7].block[4].um_I.clk ,
    \top_I.branch[7].block[3].um_I.iw[17] ,
    \top_I.branch[7].block[3].um_I.iw[16] ,
    \top_I.branch[7].block[3].um_I.iw[15] ,
    \top_I.branch[7].block[3].um_I.iw[14] ,
    \top_I.branch[7].block[3].um_I.iw[13] ,
    \top_I.branch[7].block[3].um_I.iw[12] ,
    \top_I.branch[7].block[3].um_I.iw[11] ,
    \top_I.branch[7].block[3].um_I.iw[10] ,
    \top_I.branch[7].block[3].um_I.iw[9] ,
    \top_I.branch[7].block[3].um_I.iw[8] ,
    \top_I.branch[7].block[3].um_I.iw[7] ,
    \top_I.branch[7].block[3].um_I.iw[6] ,
    \top_I.branch[7].block[3].um_I.iw[5] ,
    \top_I.branch[7].block[3].um_I.iw[4] ,
    \top_I.branch[7].block[3].um_I.iw[3] ,
    \top_I.branch[7].block[3].um_I.iw[2] ,
    \top_I.branch[7].block[3].um_I.iw[1] ,
    \top_I.branch[7].block[3].um_I.clk ,
    \top_I.branch[7].block[2].um_I.iw[17] ,
    \top_I.branch[7].block[2].um_I.iw[16] ,
    \top_I.branch[7].block[2].um_I.iw[15] ,
    \top_I.branch[7].block[2].um_I.iw[14] ,
    \top_I.branch[7].block[2].um_I.iw[13] ,
    \top_I.branch[7].block[2].um_I.iw[12] ,
    \top_I.branch[7].block[2].um_I.iw[11] ,
    \top_I.branch[7].block[2].um_I.iw[10] ,
    \top_I.branch[7].block[2].um_I.iw[9] ,
    \top_I.branch[7].block[2].um_I.iw[8] ,
    \top_I.branch[7].block[2].um_I.iw[7] ,
    \top_I.branch[7].block[2].um_I.iw[6] ,
    \top_I.branch[7].block[2].um_I.iw[5] ,
    \top_I.branch[7].block[2].um_I.iw[4] ,
    \top_I.branch[7].block[2].um_I.iw[3] ,
    \top_I.branch[7].block[2].um_I.iw[2] ,
    \top_I.branch[7].block[2].um_I.iw[1] ,
    \top_I.branch[7].block[2].um_I.clk ,
    \top_I.branch[7].block[1].um_I.iw[17] ,
    \top_I.branch[7].block[1].um_I.iw[16] ,
    \top_I.branch[7].block[1].um_I.iw[15] ,
    \top_I.branch[7].block[1].um_I.iw[14] ,
    \top_I.branch[7].block[1].um_I.iw[13] ,
    \top_I.branch[7].block[1].um_I.iw[12] ,
    \top_I.branch[7].block[1].um_I.iw[11] ,
    \top_I.branch[7].block[1].um_I.iw[10] ,
    \top_I.branch[7].block[1].um_I.iw[9] ,
    \top_I.branch[7].block[1].um_I.iw[8] ,
    \top_I.branch[7].block[1].um_I.iw[7] ,
    \top_I.branch[7].block[1].um_I.iw[6] ,
    \top_I.branch[7].block[1].um_I.iw[5] ,
    \top_I.branch[7].block[1].um_I.iw[4] ,
    \top_I.branch[7].block[1].um_I.iw[3] ,
    \top_I.branch[7].block[1].um_I.iw[2] ,
    \top_I.branch[7].block[1].um_I.iw[1] ,
    \top_I.branch[7].block[1].um_I.clk ,
    \top_I.branch[7].block[0].um_I.iw[17] ,
    \top_I.branch[7].block[0].um_I.iw[16] ,
    \top_I.branch[7].block[0].um_I.iw[15] ,
    \top_I.branch[7].block[0].um_I.iw[14] ,
    \top_I.branch[7].block[0].um_I.iw[13] ,
    \top_I.branch[7].block[0].um_I.iw[12] ,
    \top_I.branch[7].block[0].um_I.iw[11] ,
    \top_I.branch[7].block[0].um_I.iw[10] ,
    \top_I.branch[7].block[0].um_I.iw[9] ,
    \top_I.branch[7].block[0].um_I.iw[8] ,
    \top_I.branch[7].block[0].um_I.iw[7] ,
    \top_I.branch[7].block[0].um_I.iw[6] ,
    \top_I.branch[7].block[0].um_I.iw[5] ,
    \top_I.branch[7].block[0].um_I.iw[4] ,
    \top_I.branch[7].block[0].um_I.iw[3] ,
    \top_I.branch[7].block[0].um_I.iw[2] ,
    \top_I.branch[7].block[0].um_I.iw[1] ,
    \top_I.branch[7].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[7].block[15].um_I.pg_vdd ,
    \top_I.branch[7].block[14].um_I.pg_vdd ,
    \top_I.branch[7].block[13].um_I.pg_vdd ,
    \top_I.branch[7].block[12].um_I.pg_vdd ,
    \top_I.branch[7].block[11].um_I.pg_vdd ,
    \top_I.branch[7].block[10].um_I.pg_vdd ,
    \top_I.branch[7].block[9].um_I.pg_vdd ,
    \top_I.branch[7].block[8].um_I.pg_vdd ,
    \top_I.branch[7].block[7].um_I.pg_vdd ,
    \top_I.branch[7].block[6].um_I.pg_vdd ,
    \top_I.branch[7].block[5].um_I.pg_vdd ,
    \top_I.branch[7].block[4].um_I.pg_vdd ,
    \top_I.branch[7].block[3].um_I.pg_vdd ,
    \top_I.branch[7].block[2].um_I.pg_vdd ,
    \top_I.branch[7].block[1].um_I.pg_vdd ,
    \top_I.branch[7].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[8].mux_I  (.k_one(\top_I.branch[8].l_addr[2] ),
    .k_zero(\top_I.branch[8].l_addr[0] ),
    .addr({\top_I.branch[8].l_addr[0] ,
    \top_I.branch[8].l_addr[2] ,
    \top_I.branch[8].l_addr[0] ,
    \top_I.branch[8].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[8].block[15].um_I.ena ,
    \top_I.branch[8].block[14].um_I.ena ,
    \top_I.branch[8].block[13].um_I.ena ,
    \top_I.branch[8].block[12].um_I.ena ,
    \top_I.branch[8].block[11].um_I.ena ,
    \top_I.branch[8].block[10].um_I.ena ,
    \top_I.branch[8].block[9].um_I.ena ,
    \top_I.branch[8].block[8].um_I.ena ,
    \top_I.branch[8].block[7].um_I.ena ,
    \top_I.branch[8].block[6].um_I.ena ,
    \top_I.branch[8].block[5].um_I.ena ,
    \top_I.branch[8].block[4].um_I.ena ,
    \top_I.branch[8].block[3].um_I.ena ,
    \top_I.branch[8].block[2].um_I.ena ,
    \top_I.branch[8].block[1].um_I.ena ,
    \top_I.branch[8].block[0].um_I.ena }),
    .um_iw({\top_I.branch[8].block[15].um_I.iw[17] ,
    \top_I.branch[8].block[15].um_I.iw[16] ,
    \top_I.branch[8].block[15].um_I.iw[15] ,
    \top_I.branch[8].block[15].um_I.iw[14] ,
    \top_I.branch[8].block[15].um_I.iw[13] ,
    \top_I.branch[8].block[15].um_I.iw[12] ,
    \top_I.branch[8].block[15].um_I.iw[11] ,
    \top_I.branch[8].block[15].um_I.iw[10] ,
    \top_I.branch[8].block[15].um_I.iw[9] ,
    \top_I.branch[8].block[15].um_I.iw[8] ,
    \top_I.branch[8].block[15].um_I.iw[7] ,
    \top_I.branch[8].block[15].um_I.iw[6] ,
    \top_I.branch[8].block[15].um_I.iw[5] ,
    \top_I.branch[8].block[15].um_I.iw[4] ,
    \top_I.branch[8].block[15].um_I.iw[3] ,
    \top_I.branch[8].block[15].um_I.iw[2] ,
    \top_I.branch[8].block[15].um_I.iw[1] ,
    \top_I.branch[8].block[15].um_I.clk ,
    \top_I.branch[8].block[14].um_I.iw[17] ,
    \top_I.branch[8].block[14].um_I.iw[16] ,
    \top_I.branch[8].block[14].um_I.iw[15] ,
    \top_I.branch[8].block[14].um_I.iw[14] ,
    \top_I.branch[8].block[14].um_I.iw[13] ,
    \top_I.branch[8].block[14].um_I.iw[12] ,
    \top_I.branch[8].block[14].um_I.iw[11] ,
    \top_I.branch[8].block[14].um_I.iw[10] ,
    \top_I.branch[8].block[14].um_I.iw[9] ,
    \top_I.branch[8].block[14].um_I.iw[8] ,
    \top_I.branch[8].block[14].um_I.iw[7] ,
    \top_I.branch[8].block[14].um_I.iw[6] ,
    \top_I.branch[8].block[14].um_I.iw[5] ,
    \top_I.branch[8].block[14].um_I.iw[4] ,
    \top_I.branch[8].block[14].um_I.iw[3] ,
    \top_I.branch[8].block[14].um_I.iw[2] ,
    \top_I.branch[8].block[14].um_I.iw[1] ,
    \top_I.branch[8].block[14].um_I.clk ,
    \top_I.branch[8].block[13].um_I.iw[17] ,
    \top_I.branch[8].block[13].um_I.iw[16] ,
    \top_I.branch[8].block[13].um_I.iw[15] ,
    \top_I.branch[8].block[13].um_I.iw[14] ,
    \top_I.branch[8].block[13].um_I.iw[13] ,
    \top_I.branch[8].block[13].um_I.iw[12] ,
    \top_I.branch[8].block[13].um_I.iw[11] ,
    \top_I.branch[8].block[13].um_I.iw[10] ,
    \top_I.branch[8].block[13].um_I.iw[9] ,
    \top_I.branch[8].block[13].um_I.iw[8] ,
    \top_I.branch[8].block[13].um_I.iw[7] ,
    \top_I.branch[8].block[13].um_I.iw[6] ,
    \top_I.branch[8].block[13].um_I.iw[5] ,
    \top_I.branch[8].block[13].um_I.iw[4] ,
    \top_I.branch[8].block[13].um_I.iw[3] ,
    \top_I.branch[8].block[13].um_I.iw[2] ,
    \top_I.branch[8].block[13].um_I.iw[1] ,
    \top_I.branch[8].block[13].um_I.clk ,
    \top_I.branch[8].block[12].um_I.iw[17] ,
    \top_I.branch[8].block[12].um_I.iw[16] ,
    \top_I.branch[8].block[12].um_I.iw[15] ,
    \top_I.branch[8].block[12].um_I.iw[14] ,
    \top_I.branch[8].block[12].um_I.iw[13] ,
    \top_I.branch[8].block[12].um_I.iw[12] ,
    \top_I.branch[8].block[12].um_I.iw[11] ,
    \top_I.branch[8].block[12].um_I.iw[10] ,
    \top_I.branch[8].block[12].um_I.iw[9] ,
    \top_I.branch[8].block[12].um_I.iw[8] ,
    \top_I.branch[8].block[12].um_I.iw[7] ,
    \top_I.branch[8].block[12].um_I.iw[6] ,
    \top_I.branch[8].block[12].um_I.iw[5] ,
    \top_I.branch[8].block[12].um_I.iw[4] ,
    \top_I.branch[8].block[12].um_I.iw[3] ,
    \top_I.branch[8].block[12].um_I.iw[2] ,
    \top_I.branch[8].block[12].um_I.iw[1] ,
    \top_I.branch[8].block[12].um_I.clk ,
    \top_I.branch[8].block[11].um_I.iw[17] ,
    \top_I.branch[8].block[11].um_I.iw[16] ,
    \top_I.branch[8].block[11].um_I.iw[15] ,
    \top_I.branch[8].block[11].um_I.iw[14] ,
    \top_I.branch[8].block[11].um_I.iw[13] ,
    \top_I.branch[8].block[11].um_I.iw[12] ,
    \top_I.branch[8].block[11].um_I.iw[11] ,
    \top_I.branch[8].block[11].um_I.iw[10] ,
    \top_I.branch[8].block[11].um_I.iw[9] ,
    \top_I.branch[8].block[11].um_I.iw[8] ,
    \top_I.branch[8].block[11].um_I.iw[7] ,
    \top_I.branch[8].block[11].um_I.iw[6] ,
    \top_I.branch[8].block[11].um_I.iw[5] ,
    \top_I.branch[8].block[11].um_I.iw[4] ,
    \top_I.branch[8].block[11].um_I.iw[3] ,
    \top_I.branch[8].block[11].um_I.iw[2] ,
    \top_I.branch[8].block[11].um_I.iw[1] ,
    \top_I.branch[8].block[11].um_I.clk ,
    \top_I.branch[8].block[10].um_I.iw[17] ,
    \top_I.branch[8].block[10].um_I.iw[16] ,
    \top_I.branch[8].block[10].um_I.iw[15] ,
    \top_I.branch[8].block[10].um_I.iw[14] ,
    \top_I.branch[8].block[10].um_I.iw[13] ,
    \top_I.branch[8].block[10].um_I.iw[12] ,
    \top_I.branch[8].block[10].um_I.iw[11] ,
    \top_I.branch[8].block[10].um_I.iw[10] ,
    \top_I.branch[8].block[10].um_I.iw[9] ,
    \top_I.branch[8].block[10].um_I.iw[8] ,
    \top_I.branch[8].block[10].um_I.iw[7] ,
    \top_I.branch[8].block[10].um_I.iw[6] ,
    \top_I.branch[8].block[10].um_I.iw[5] ,
    \top_I.branch[8].block[10].um_I.iw[4] ,
    \top_I.branch[8].block[10].um_I.iw[3] ,
    \top_I.branch[8].block[10].um_I.iw[2] ,
    \top_I.branch[8].block[10].um_I.iw[1] ,
    \top_I.branch[8].block[10].um_I.clk ,
    \top_I.branch[8].block[9].um_I.iw[17] ,
    \top_I.branch[8].block[9].um_I.iw[16] ,
    \top_I.branch[8].block[9].um_I.iw[15] ,
    \top_I.branch[8].block[9].um_I.iw[14] ,
    \top_I.branch[8].block[9].um_I.iw[13] ,
    \top_I.branch[8].block[9].um_I.iw[12] ,
    \top_I.branch[8].block[9].um_I.iw[11] ,
    \top_I.branch[8].block[9].um_I.iw[10] ,
    \top_I.branch[8].block[9].um_I.iw[9] ,
    \top_I.branch[8].block[9].um_I.iw[8] ,
    \top_I.branch[8].block[9].um_I.iw[7] ,
    \top_I.branch[8].block[9].um_I.iw[6] ,
    \top_I.branch[8].block[9].um_I.iw[5] ,
    \top_I.branch[8].block[9].um_I.iw[4] ,
    \top_I.branch[8].block[9].um_I.iw[3] ,
    \top_I.branch[8].block[9].um_I.iw[2] ,
    \top_I.branch[8].block[9].um_I.iw[1] ,
    \top_I.branch[8].block[9].um_I.clk ,
    \top_I.branch[8].block[8].um_I.iw[17] ,
    \top_I.branch[8].block[8].um_I.iw[16] ,
    \top_I.branch[8].block[8].um_I.iw[15] ,
    \top_I.branch[8].block[8].um_I.iw[14] ,
    \top_I.branch[8].block[8].um_I.iw[13] ,
    \top_I.branch[8].block[8].um_I.iw[12] ,
    \top_I.branch[8].block[8].um_I.iw[11] ,
    \top_I.branch[8].block[8].um_I.iw[10] ,
    \top_I.branch[8].block[8].um_I.iw[9] ,
    \top_I.branch[8].block[8].um_I.iw[8] ,
    \top_I.branch[8].block[8].um_I.iw[7] ,
    \top_I.branch[8].block[8].um_I.iw[6] ,
    \top_I.branch[8].block[8].um_I.iw[5] ,
    \top_I.branch[8].block[8].um_I.iw[4] ,
    \top_I.branch[8].block[8].um_I.iw[3] ,
    \top_I.branch[8].block[8].um_I.iw[2] ,
    \top_I.branch[8].block[8].um_I.iw[1] ,
    \top_I.branch[8].block[8].um_I.clk ,
    \top_I.branch[8].block[7].um_I.iw[17] ,
    \top_I.branch[8].block[7].um_I.iw[16] ,
    \top_I.branch[8].block[7].um_I.iw[15] ,
    \top_I.branch[8].block[7].um_I.iw[14] ,
    \top_I.branch[8].block[7].um_I.iw[13] ,
    \top_I.branch[8].block[7].um_I.iw[12] ,
    \top_I.branch[8].block[7].um_I.iw[11] ,
    \top_I.branch[8].block[7].um_I.iw[10] ,
    \top_I.branch[8].block[7].um_I.iw[9] ,
    \top_I.branch[8].block[7].um_I.iw[8] ,
    \top_I.branch[8].block[7].um_I.iw[7] ,
    \top_I.branch[8].block[7].um_I.iw[6] ,
    \top_I.branch[8].block[7].um_I.iw[5] ,
    \top_I.branch[8].block[7].um_I.iw[4] ,
    \top_I.branch[8].block[7].um_I.iw[3] ,
    \top_I.branch[8].block[7].um_I.iw[2] ,
    \top_I.branch[8].block[7].um_I.iw[1] ,
    \top_I.branch[8].block[7].um_I.clk ,
    \top_I.branch[8].block[6].um_I.iw[17] ,
    \top_I.branch[8].block[6].um_I.iw[16] ,
    \top_I.branch[8].block[6].um_I.iw[15] ,
    \top_I.branch[8].block[6].um_I.iw[14] ,
    \top_I.branch[8].block[6].um_I.iw[13] ,
    \top_I.branch[8].block[6].um_I.iw[12] ,
    \top_I.branch[8].block[6].um_I.iw[11] ,
    \top_I.branch[8].block[6].um_I.iw[10] ,
    \top_I.branch[8].block[6].um_I.iw[9] ,
    \top_I.branch[8].block[6].um_I.iw[8] ,
    \top_I.branch[8].block[6].um_I.iw[7] ,
    \top_I.branch[8].block[6].um_I.iw[6] ,
    \top_I.branch[8].block[6].um_I.iw[5] ,
    \top_I.branch[8].block[6].um_I.iw[4] ,
    \top_I.branch[8].block[6].um_I.iw[3] ,
    \top_I.branch[8].block[6].um_I.iw[2] ,
    \top_I.branch[8].block[6].um_I.iw[1] ,
    \top_I.branch[8].block[6].um_I.clk ,
    \top_I.branch[8].block[5].um_I.iw[17] ,
    \top_I.branch[8].block[5].um_I.iw[16] ,
    \top_I.branch[8].block[5].um_I.iw[15] ,
    \top_I.branch[8].block[5].um_I.iw[14] ,
    \top_I.branch[8].block[5].um_I.iw[13] ,
    \top_I.branch[8].block[5].um_I.iw[12] ,
    \top_I.branch[8].block[5].um_I.iw[11] ,
    \top_I.branch[8].block[5].um_I.iw[10] ,
    \top_I.branch[8].block[5].um_I.iw[9] ,
    \top_I.branch[8].block[5].um_I.iw[8] ,
    \top_I.branch[8].block[5].um_I.iw[7] ,
    \top_I.branch[8].block[5].um_I.iw[6] ,
    \top_I.branch[8].block[5].um_I.iw[5] ,
    \top_I.branch[8].block[5].um_I.iw[4] ,
    \top_I.branch[8].block[5].um_I.iw[3] ,
    \top_I.branch[8].block[5].um_I.iw[2] ,
    \top_I.branch[8].block[5].um_I.iw[1] ,
    \top_I.branch[8].block[5].um_I.clk ,
    \top_I.branch[8].block[4].um_I.iw[17] ,
    \top_I.branch[8].block[4].um_I.iw[16] ,
    \top_I.branch[8].block[4].um_I.iw[15] ,
    \top_I.branch[8].block[4].um_I.iw[14] ,
    \top_I.branch[8].block[4].um_I.iw[13] ,
    \top_I.branch[8].block[4].um_I.iw[12] ,
    \top_I.branch[8].block[4].um_I.iw[11] ,
    \top_I.branch[8].block[4].um_I.iw[10] ,
    \top_I.branch[8].block[4].um_I.iw[9] ,
    \top_I.branch[8].block[4].um_I.iw[8] ,
    \top_I.branch[8].block[4].um_I.iw[7] ,
    \top_I.branch[8].block[4].um_I.iw[6] ,
    \top_I.branch[8].block[4].um_I.iw[5] ,
    \top_I.branch[8].block[4].um_I.iw[4] ,
    \top_I.branch[8].block[4].um_I.iw[3] ,
    \top_I.branch[8].block[4].um_I.iw[2] ,
    \top_I.branch[8].block[4].um_I.iw[1] ,
    \top_I.branch[8].block[4].um_I.clk ,
    \top_I.branch[8].block[3].um_I.iw[17] ,
    \top_I.branch[8].block[3].um_I.iw[16] ,
    \top_I.branch[8].block[3].um_I.iw[15] ,
    \top_I.branch[8].block[3].um_I.iw[14] ,
    \top_I.branch[8].block[3].um_I.iw[13] ,
    \top_I.branch[8].block[3].um_I.iw[12] ,
    \top_I.branch[8].block[3].um_I.iw[11] ,
    \top_I.branch[8].block[3].um_I.iw[10] ,
    \top_I.branch[8].block[3].um_I.iw[9] ,
    \top_I.branch[8].block[3].um_I.iw[8] ,
    \top_I.branch[8].block[3].um_I.iw[7] ,
    \top_I.branch[8].block[3].um_I.iw[6] ,
    \top_I.branch[8].block[3].um_I.iw[5] ,
    \top_I.branch[8].block[3].um_I.iw[4] ,
    \top_I.branch[8].block[3].um_I.iw[3] ,
    \top_I.branch[8].block[3].um_I.iw[2] ,
    \top_I.branch[8].block[3].um_I.iw[1] ,
    \top_I.branch[8].block[3].um_I.clk ,
    \top_I.branch[8].block[2].um_I.iw[17] ,
    \top_I.branch[8].block[2].um_I.iw[16] ,
    \top_I.branch[8].block[2].um_I.iw[15] ,
    \top_I.branch[8].block[2].um_I.iw[14] ,
    \top_I.branch[8].block[2].um_I.iw[13] ,
    \top_I.branch[8].block[2].um_I.iw[12] ,
    \top_I.branch[8].block[2].um_I.iw[11] ,
    \top_I.branch[8].block[2].um_I.iw[10] ,
    \top_I.branch[8].block[2].um_I.iw[9] ,
    \top_I.branch[8].block[2].um_I.iw[8] ,
    \top_I.branch[8].block[2].um_I.iw[7] ,
    \top_I.branch[8].block[2].um_I.iw[6] ,
    \top_I.branch[8].block[2].um_I.iw[5] ,
    \top_I.branch[8].block[2].um_I.iw[4] ,
    \top_I.branch[8].block[2].um_I.iw[3] ,
    \top_I.branch[8].block[2].um_I.iw[2] ,
    \top_I.branch[8].block[2].um_I.iw[1] ,
    \top_I.branch[8].block[2].um_I.clk ,
    \top_I.branch[8].block[1].um_I.iw[17] ,
    \top_I.branch[8].block[1].um_I.iw[16] ,
    \top_I.branch[8].block[1].um_I.iw[15] ,
    \top_I.branch[8].block[1].um_I.iw[14] ,
    \top_I.branch[8].block[1].um_I.iw[13] ,
    \top_I.branch[8].block[1].um_I.iw[12] ,
    \top_I.branch[8].block[1].um_I.iw[11] ,
    \top_I.branch[8].block[1].um_I.iw[10] ,
    \top_I.branch[8].block[1].um_I.iw[9] ,
    \top_I.branch[8].block[1].um_I.iw[8] ,
    \top_I.branch[8].block[1].um_I.iw[7] ,
    \top_I.branch[8].block[1].um_I.iw[6] ,
    \top_I.branch[8].block[1].um_I.iw[5] ,
    \top_I.branch[8].block[1].um_I.iw[4] ,
    \top_I.branch[8].block[1].um_I.iw[3] ,
    \top_I.branch[8].block[1].um_I.iw[2] ,
    \top_I.branch[8].block[1].um_I.iw[1] ,
    \top_I.branch[8].block[1].um_I.clk ,
    \top_I.branch[8].block[0].um_I.iw[17] ,
    \top_I.branch[8].block[0].um_I.iw[16] ,
    \top_I.branch[8].block[0].um_I.iw[15] ,
    \top_I.branch[8].block[0].um_I.iw[14] ,
    \top_I.branch[8].block[0].um_I.iw[13] ,
    \top_I.branch[8].block[0].um_I.iw[12] ,
    \top_I.branch[8].block[0].um_I.iw[11] ,
    \top_I.branch[8].block[0].um_I.iw[10] ,
    \top_I.branch[8].block[0].um_I.iw[9] ,
    \top_I.branch[8].block[0].um_I.iw[8] ,
    \top_I.branch[8].block[0].um_I.iw[7] ,
    \top_I.branch[8].block[0].um_I.iw[6] ,
    \top_I.branch[8].block[0].um_I.iw[5] ,
    \top_I.branch[8].block[0].um_I.iw[4] ,
    \top_I.branch[8].block[0].um_I.iw[3] ,
    \top_I.branch[8].block[0].um_I.iw[2] ,
    \top_I.branch[8].block[0].um_I.iw[1] ,
    \top_I.branch[8].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[8].block[15].um_I.pg_vdd ,
    \top_I.branch[8].block[14].um_I.pg_vdd ,
    \top_I.branch[8].block[13].um_I.pg_vdd ,
    \top_I.branch[8].block[12].um_I.pg_vdd ,
    \top_I.branch[8].block[11].um_I.pg_vdd ,
    \top_I.branch[8].block[10].um_I.pg_vdd ,
    \top_I.branch[8].block[9].um_I.pg_vdd ,
    \top_I.branch[8].block[8].um_I.pg_vdd ,
    \top_I.branch[8].block[7].um_I.pg_vdd ,
    \top_I.branch[8].block[6].um_I.pg_vdd ,
    \top_I.branch[8].block[5].um_I.pg_vdd ,
    \top_I.branch[8].block[4].um_I.pg_vdd ,
    \top_I.branch[8].block[3].um_I.pg_vdd ,
    \top_I.branch[8].block[2].um_I.pg_vdd ,
    \top_I.branch[8].block[1].um_I.pg_vdd ,
    \top_I.branch[8].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[9].mux_I  (.k_one(\top_I.branch[9].l_addr[2] ),
    .k_zero(\top_I.branch[9].l_addr[0] ),
    .addr({\top_I.branch[9].l_addr[0] ,
    \top_I.branch[9].l_addr[2] ,
    \top_I.branch[9].l_addr[0] ,
    \top_I.branch[9].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[9].block[15].um_I.ena ,
    \top_I.branch[9].block[14].um_I.ena ,
    \top_I.branch[9].block[13].um_I.ena ,
    \top_I.branch[9].block[12].um_I.ena ,
    \top_I.branch[9].block[11].um_I.ena ,
    \top_I.branch[9].block[10].um_I.ena ,
    \top_I.branch[9].block[9].um_I.ena ,
    \top_I.branch[9].block[8].um_I.ena ,
    \top_I.branch[9].block[7].um_I.ena ,
    \top_I.branch[9].block[6].um_I.ena ,
    \top_I.branch[9].block[5].um_I.ena ,
    \top_I.branch[9].block[4].um_I.ena ,
    \top_I.branch[9].block[3].um_I.ena ,
    \top_I.branch[9].block[2].um_I.ena ,
    \top_I.branch[9].block[1].um_I.ena ,
    \top_I.branch[9].block[0].um_I.ena }),
    .um_iw({\top_I.branch[9].block[15].um_I.iw[17] ,
    \top_I.branch[9].block[15].um_I.iw[16] ,
    \top_I.branch[9].block[15].um_I.iw[15] ,
    \top_I.branch[9].block[15].um_I.iw[14] ,
    \top_I.branch[9].block[15].um_I.iw[13] ,
    \top_I.branch[9].block[15].um_I.iw[12] ,
    \top_I.branch[9].block[15].um_I.iw[11] ,
    \top_I.branch[9].block[15].um_I.iw[10] ,
    \top_I.branch[9].block[15].um_I.iw[9] ,
    \top_I.branch[9].block[15].um_I.iw[8] ,
    \top_I.branch[9].block[15].um_I.iw[7] ,
    \top_I.branch[9].block[15].um_I.iw[6] ,
    \top_I.branch[9].block[15].um_I.iw[5] ,
    \top_I.branch[9].block[15].um_I.iw[4] ,
    \top_I.branch[9].block[15].um_I.iw[3] ,
    \top_I.branch[9].block[15].um_I.iw[2] ,
    \top_I.branch[9].block[15].um_I.iw[1] ,
    \top_I.branch[9].block[15].um_I.clk ,
    \top_I.branch[9].block[14].um_I.iw[17] ,
    \top_I.branch[9].block[14].um_I.iw[16] ,
    \top_I.branch[9].block[14].um_I.iw[15] ,
    \top_I.branch[9].block[14].um_I.iw[14] ,
    \top_I.branch[9].block[14].um_I.iw[13] ,
    \top_I.branch[9].block[14].um_I.iw[12] ,
    \top_I.branch[9].block[14].um_I.iw[11] ,
    \top_I.branch[9].block[14].um_I.iw[10] ,
    \top_I.branch[9].block[14].um_I.iw[9] ,
    \top_I.branch[9].block[14].um_I.iw[8] ,
    \top_I.branch[9].block[14].um_I.iw[7] ,
    \top_I.branch[9].block[14].um_I.iw[6] ,
    \top_I.branch[9].block[14].um_I.iw[5] ,
    \top_I.branch[9].block[14].um_I.iw[4] ,
    \top_I.branch[9].block[14].um_I.iw[3] ,
    \top_I.branch[9].block[14].um_I.iw[2] ,
    \top_I.branch[9].block[14].um_I.iw[1] ,
    \top_I.branch[9].block[14].um_I.clk ,
    \top_I.branch[9].block[13].um_I.iw[17] ,
    \top_I.branch[9].block[13].um_I.iw[16] ,
    \top_I.branch[9].block[13].um_I.iw[15] ,
    \top_I.branch[9].block[13].um_I.iw[14] ,
    \top_I.branch[9].block[13].um_I.iw[13] ,
    \top_I.branch[9].block[13].um_I.iw[12] ,
    \top_I.branch[9].block[13].um_I.iw[11] ,
    \top_I.branch[9].block[13].um_I.iw[10] ,
    \top_I.branch[9].block[13].um_I.iw[9] ,
    \top_I.branch[9].block[13].um_I.iw[8] ,
    \top_I.branch[9].block[13].um_I.iw[7] ,
    \top_I.branch[9].block[13].um_I.iw[6] ,
    \top_I.branch[9].block[13].um_I.iw[5] ,
    \top_I.branch[9].block[13].um_I.iw[4] ,
    \top_I.branch[9].block[13].um_I.iw[3] ,
    \top_I.branch[9].block[13].um_I.iw[2] ,
    \top_I.branch[9].block[13].um_I.iw[1] ,
    \top_I.branch[9].block[13].um_I.clk ,
    \top_I.branch[9].block[12].um_I.iw[17] ,
    \top_I.branch[9].block[12].um_I.iw[16] ,
    \top_I.branch[9].block[12].um_I.iw[15] ,
    \top_I.branch[9].block[12].um_I.iw[14] ,
    \top_I.branch[9].block[12].um_I.iw[13] ,
    \top_I.branch[9].block[12].um_I.iw[12] ,
    \top_I.branch[9].block[12].um_I.iw[11] ,
    \top_I.branch[9].block[12].um_I.iw[10] ,
    \top_I.branch[9].block[12].um_I.iw[9] ,
    \top_I.branch[9].block[12].um_I.iw[8] ,
    \top_I.branch[9].block[12].um_I.iw[7] ,
    \top_I.branch[9].block[12].um_I.iw[6] ,
    \top_I.branch[9].block[12].um_I.iw[5] ,
    \top_I.branch[9].block[12].um_I.iw[4] ,
    \top_I.branch[9].block[12].um_I.iw[3] ,
    \top_I.branch[9].block[12].um_I.iw[2] ,
    \top_I.branch[9].block[12].um_I.iw[1] ,
    \top_I.branch[9].block[12].um_I.clk ,
    \top_I.branch[9].block[11].um_I.iw[17] ,
    \top_I.branch[9].block[11].um_I.iw[16] ,
    \top_I.branch[9].block[11].um_I.iw[15] ,
    \top_I.branch[9].block[11].um_I.iw[14] ,
    \top_I.branch[9].block[11].um_I.iw[13] ,
    \top_I.branch[9].block[11].um_I.iw[12] ,
    \top_I.branch[9].block[11].um_I.iw[11] ,
    \top_I.branch[9].block[11].um_I.iw[10] ,
    \top_I.branch[9].block[11].um_I.iw[9] ,
    \top_I.branch[9].block[11].um_I.iw[8] ,
    \top_I.branch[9].block[11].um_I.iw[7] ,
    \top_I.branch[9].block[11].um_I.iw[6] ,
    \top_I.branch[9].block[11].um_I.iw[5] ,
    \top_I.branch[9].block[11].um_I.iw[4] ,
    \top_I.branch[9].block[11].um_I.iw[3] ,
    \top_I.branch[9].block[11].um_I.iw[2] ,
    \top_I.branch[9].block[11].um_I.iw[1] ,
    \top_I.branch[9].block[11].um_I.clk ,
    \top_I.branch[9].block[10].um_I.iw[17] ,
    \top_I.branch[9].block[10].um_I.iw[16] ,
    \top_I.branch[9].block[10].um_I.iw[15] ,
    \top_I.branch[9].block[10].um_I.iw[14] ,
    \top_I.branch[9].block[10].um_I.iw[13] ,
    \top_I.branch[9].block[10].um_I.iw[12] ,
    \top_I.branch[9].block[10].um_I.iw[11] ,
    \top_I.branch[9].block[10].um_I.iw[10] ,
    \top_I.branch[9].block[10].um_I.iw[9] ,
    \top_I.branch[9].block[10].um_I.iw[8] ,
    \top_I.branch[9].block[10].um_I.iw[7] ,
    \top_I.branch[9].block[10].um_I.iw[6] ,
    \top_I.branch[9].block[10].um_I.iw[5] ,
    \top_I.branch[9].block[10].um_I.iw[4] ,
    \top_I.branch[9].block[10].um_I.iw[3] ,
    \top_I.branch[9].block[10].um_I.iw[2] ,
    \top_I.branch[9].block[10].um_I.iw[1] ,
    \top_I.branch[9].block[10].um_I.clk ,
    \top_I.branch[9].block[9].um_I.iw[17] ,
    \top_I.branch[9].block[9].um_I.iw[16] ,
    \top_I.branch[9].block[9].um_I.iw[15] ,
    \top_I.branch[9].block[9].um_I.iw[14] ,
    \top_I.branch[9].block[9].um_I.iw[13] ,
    \top_I.branch[9].block[9].um_I.iw[12] ,
    \top_I.branch[9].block[9].um_I.iw[11] ,
    \top_I.branch[9].block[9].um_I.iw[10] ,
    \top_I.branch[9].block[9].um_I.iw[9] ,
    \top_I.branch[9].block[9].um_I.iw[8] ,
    \top_I.branch[9].block[9].um_I.iw[7] ,
    \top_I.branch[9].block[9].um_I.iw[6] ,
    \top_I.branch[9].block[9].um_I.iw[5] ,
    \top_I.branch[9].block[9].um_I.iw[4] ,
    \top_I.branch[9].block[9].um_I.iw[3] ,
    \top_I.branch[9].block[9].um_I.iw[2] ,
    \top_I.branch[9].block[9].um_I.iw[1] ,
    \top_I.branch[9].block[9].um_I.clk ,
    \top_I.branch[9].block[8].um_I.iw[17] ,
    \top_I.branch[9].block[8].um_I.iw[16] ,
    \top_I.branch[9].block[8].um_I.iw[15] ,
    \top_I.branch[9].block[8].um_I.iw[14] ,
    \top_I.branch[9].block[8].um_I.iw[13] ,
    \top_I.branch[9].block[8].um_I.iw[12] ,
    \top_I.branch[9].block[8].um_I.iw[11] ,
    \top_I.branch[9].block[8].um_I.iw[10] ,
    \top_I.branch[9].block[8].um_I.iw[9] ,
    \top_I.branch[9].block[8].um_I.iw[8] ,
    \top_I.branch[9].block[8].um_I.iw[7] ,
    \top_I.branch[9].block[8].um_I.iw[6] ,
    \top_I.branch[9].block[8].um_I.iw[5] ,
    \top_I.branch[9].block[8].um_I.iw[4] ,
    \top_I.branch[9].block[8].um_I.iw[3] ,
    \top_I.branch[9].block[8].um_I.iw[2] ,
    \top_I.branch[9].block[8].um_I.iw[1] ,
    \top_I.branch[9].block[8].um_I.clk ,
    \top_I.branch[9].block[7].um_I.iw[17] ,
    \top_I.branch[9].block[7].um_I.iw[16] ,
    \top_I.branch[9].block[7].um_I.iw[15] ,
    \top_I.branch[9].block[7].um_I.iw[14] ,
    \top_I.branch[9].block[7].um_I.iw[13] ,
    \top_I.branch[9].block[7].um_I.iw[12] ,
    \top_I.branch[9].block[7].um_I.iw[11] ,
    \top_I.branch[9].block[7].um_I.iw[10] ,
    \top_I.branch[9].block[7].um_I.iw[9] ,
    \top_I.branch[9].block[7].um_I.iw[8] ,
    \top_I.branch[9].block[7].um_I.iw[7] ,
    \top_I.branch[9].block[7].um_I.iw[6] ,
    \top_I.branch[9].block[7].um_I.iw[5] ,
    \top_I.branch[9].block[7].um_I.iw[4] ,
    \top_I.branch[9].block[7].um_I.iw[3] ,
    \top_I.branch[9].block[7].um_I.iw[2] ,
    \top_I.branch[9].block[7].um_I.iw[1] ,
    \top_I.branch[9].block[7].um_I.clk ,
    \top_I.branch[9].block[6].um_I.iw[17] ,
    \top_I.branch[9].block[6].um_I.iw[16] ,
    \top_I.branch[9].block[6].um_I.iw[15] ,
    \top_I.branch[9].block[6].um_I.iw[14] ,
    \top_I.branch[9].block[6].um_I.iw[13] ,
    \top_I.branch[9].block[6].um_I.iw[12] ,
    \top_I.branch[9].block[6].um_I.iw[11] ,
    \top_I.branch[9].block[6].um_I.iw[10] ,
    \top_I.branch[9].block[6].um_I.iw[9] ,
    \top_I.branch[9].block[6].um_I.iw[8] ,
    \top_I.branch[9].block[6].um_I.iw[7] ,
    \top_I.branch[9].block[6].um_I.iw[6] ,
    \top_I.branch[9].block[6].um_I.iw[5] ,
    \top_I.branch[9].block[6].um_I.iw[4] ,
    \top_I.branch[9].block[6].um_I.iw[3] ,
    \top_I.branch[9].block[6].um_I.iw[2] ,
    \top_I.branch[9].block[6].um_I.iw[1] ,
    \top_I.branch[9].block[6].um_I.clk ,
    \top_I.branch[9].block[5].um_I.iw[17] ,
    \top_I.branch[9].block[5].um_I.iw[16] ,
    \top_I.branch[9].block[5].um_I.iw[15] ,
    \top_I.branch[9].block[5].um_I.iw[14] ,
    \top_I.branch[9].block[5].um_I.iw[13] ,
    \top_I.branch[9].block[5].um_I.iw[12] ,
    \top_I.branch[9].block[5].um_I.iw[11] ,
    \top_I.branch[9].block[5].um_I.iw[10] ,
    \top_I.branch[9].block[5].um_I.iw[9] ,
    \top_I.branch[9].block[5].um_I.iw[8] ,
    \top_I.branch[9].block[5].um_I.iw[7] ,
    \top_I.branch[9].block[5].um_I.iw[6] ,
    \top_I.branch[9].block[5].um_I.iw[5] ,
    \top_I.branch[9].block[5].um_I.iw[4] ,
    \top_I.branch[9].block[5].um_I.iw[3] ,
    \top_I.branch[9].block[5].um_I.iw[2] ,
    \top_I.branch[9].block[5].um_I.iw[1] ,
    \top_I.branch[9].block[5].um_I.clk ,
    \top_I.branch[9].block[4].um_I.iw[17] ,
    \top_I.branch[9].block[4].um_I.iw[16] ,
    \top_I.branch[9].block[4].um_I.iw[15] ,
    \top_I.branch[9].block[4].um_I.iw[14] ,
    \top_I.branch[9].block[4].um_I.iw[13] ,
    \top_I.branch[9].block[4].um_I.iw[12] ,
    \top_I.branch[9].block[4].um_I.iw[11] ,
    \top_I.branch[9].block[4].um_I.iw[10] ,
    \top_I.branch[9].block[4].um_I.iw[9] ,
    \top_I.branch[9].block[4].um_I.iw[8] ,
    \top_I.branch[9].block[4].um_I.iw[7] ,
    \top_I.branch[9].block[4].um_I.iw[6] ,
    \top_I.branch[9].block[4].um_I.iw[5] ,
    \top_I.branch[9].block[4].um_I.iw[4] ,
    \top_I.branch[9].block[4].um_I.iw[3] ,
    \top_I.branch[9].block[4].um_I.iw[2] ,
    \top_I.branch[9].block[4].um_I.iw[1] ,
    \top_I.branch[9].block[4].um_I.clk ,
    \top_I.branch[9].block[3].um_I.iw[17] ,
    \top_I.branch[9].block[3].um_I.iw[16] ,
    \top_I.branch[9].block[3].um_I.iw[15] ,
    \top_I.branch[9].block[3].um_I.iw[14] ,
    \top_I.branch[9].block[3].um_I.iw[13] ,
    \top_I.branch[9].block[3].um_I.iw[12] ,
    \top_I.branch[9].block[3].um_I.iw[11] ,
    \top_I.branch[9].block[3].um_I.iw[10] ,
    \top_I.branch[9].block[3].um_I.iw[9] ,
    \top_I.branch[9].block[3].um_I.iw[8] ,
    \top_I.branch[9].block[3].um_I.iw[7] ,
    \top_I.branch[9].block[3].um_I.iw[6] ,
    \top_I.branch[9].block[3].um_I.iw[5] ,
    \top_I.branch[9].block[3].um_I.iw[4] ,
    \top_I.branch[9].block[3].um_I.iw[3] ,
    \top_I.branch[9].block[3].um_I.iw[2] ,
    \top_I.branch[9].block[3].um_I.iw[1] ,
    \top_I.branch[9].block[3].um_I.clk ,
    \top_I.branch[9].block[2].um_I.iw[17] ,
    \top_I.branch[9].block[2].um_I.iw[16] ,
    \top_I.branch[9].block[2].um_I.iw[15] ,
    \top_I.branch[9].block[2].um_I.iw[14] ,
    \top_I.branch[9].block[2].um_I.iw[13] ,
    \top_I.branch[9].block[2].um_I.iw[12] ,
    \top_I.branch[9].block[2].um_I.iw[11] ,
    \top_I.branch[9].block[2].um_I.iw[10] ,
    \top_I.branch[9].block[2].um_I.iw[9] ,
    \top_I.branch[9].block[2].um_I.iw[8] ,
    \top_I.branch[9].block[2].um_I.iw[7] ,
    \top_I.branch[9].block[2].um_I.iw[6] ,
    \top_I.branch[9].block[2].um_I.iw[5] ,
    \top_I.branch[9].block[2].um_I.iw[4] ,
    \top_I.branch[9].block[2].um_I.iw[3] ,
    \top_I.branch[9].block[2].um_I.iw[2] ,
    \top_I.branch[9].block[2].um_I.iw[1] ,
    \top_I.branch[9].block[2].um_I.clk ,
    \top_I.branch[9].block[1].um_I.iw[17] ,
    \top_I.branch[9].block[1].um_I.iw[16] ,
    \top_I.branch[9].block[1].um_I.iw[15] ,
    \top_I.branch[9].block[1].um_I.iw[14] ,
    \top_I.branch[9].block[1].um_I.iw[13] ,
    \top_I.branch[9].block[1].um_I.iw[12] ,
    \top_I.branch[9].block[1].um_I.iw[11] ,
    \top_I.branch[9].block[1].um_I.iw[10] ,
    \top_I.branch[9].block[1].um_I.iw[9] ,
    \top_I.branch[9].block[1].um_I.iw[8] ,
    \top_I.branch[9].block[1].um_I.iw[7] ,
    \top_I.branch[9].block[1].um_I.iw[6] ,
    \top_I.branch[9].block[1].um_I.iw[5] ,
    \top_I.branch[9].block[1].um_I.iw[4] ,
    \top_I.branch[9].block[1].um_I.iw[3] ,
    \top_I.branch[9].block[1].um_I.iw[2] ,
    \top_I.branch[9].block[1].um_I.iw[1] ,
    \top_I.branch[9].block[1].um_I.clk ,
    \top_I.branch[9].block[0].um_I.iw[17] ,
    \top_I.branch[9].block[0].um_I.iw[16] ,
    \top_I.branch[9].block[0].um_I.iw[15] ,
    \top_I.branch[9].block[0].um_I.iw[14] ,
    \top_I.branch[9].block[0].um_I.iw[13] ,
    \top_I.branch[9].block[0].um_I.iw[12] ,
    \top_I.branch[9].block[0].um_I.iw[11] ,
    \top_I.branch[9].block[0].um_I.iw[10] ,
    \top_I.branch[9].block[0].um_I.iw[9] ,
    \top_I.branch[9].block[0].um_I.iw[8] ,
    \top_I.branch[9].block[0].um_I.iw[7] ,
    \top_I.branch[9].block[0].um_I.iw[6] ,
    \top_I.branch[9].block[0].um_I.iw[5] ,
    \top_I.branch[9].block[0].um_I.iw[4] ,
    \top_I.branch[9].block[0].um_I.iw[3] ,
    \top_I.branch[9].block[0].um_I.iw[2] ,
    \top_I.branch[9].block[0].um_I.iw[1] ,
    \top_I.branch[9].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[9].block[15].um_I.pg_vdd ,
    \top_I.branch[9].block[14].um_I.pg_vdd ,
    \top_I.branch[9].block[13].um_I.pg_vdd ,
    \top_I.branch[9].block[12].um_I.pg_vdd ,
    \top_I.branch[9].block[11].um_I.pg_vdd ,
    \top_I.branch[9].block[10].um_I.pg_vdd ,
    \top_I.branch[9].block[9].um_I.pg_vdd ,
    \top_I.branch[9].block[8].um_I.pg_vdd ,
    \top_I.branch[9].block[7].um_I.pg_vdd ,
    \top_I.branch[9].block[6].um_I.pg_vdd ,
    \top_I.branch[9].block[5].um_I.pg_vdd ,
    \top_I.branch[9].block[4].um_I.pg_vdd ,
    \top_I.branch[9].block[3].um_I.pg_vdd ,
    \top_I.branch[9].block[2].um_I.pg_vdd ,
    \top_I.branch[9].block[1].um_I.pg_vdd ,
    \top_I.branch[9].block[0].um_I.pg_vdd }));
 tt_ctrl \top_I.ctrl_I  (.ctrl_ena(io_in[32]),
    .ctrl_sel_inc(io_in[34]),
    .ctrl_sel_rst_n(io_in[36]),
    .k_one(\top_I.io_oeb[0] ),
    .k_zero(wbs_ack_o),
    .pad_ui_in({io_in[15],
    io_in[14],
    io_in[13],
    io_in[12],
    io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6]}),
    .pad_uio_in({io_in[31],
    io_in[30],
    io_in[29],
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24]}),
    .pad_uio_oe_n({io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24]}),
    .pad_uio_out({io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24]}),
    .pad_uo_out({io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16]}),
    .spine_bot_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_bot_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .spine_top_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_top_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }));
 assign io_oeb[0] = \top_I.io_oeb[0] ;
 assign io_oeb[10] = \top_I.io_oeb[0] ;
 assign io_oeb[11] = \top_I.io_oeb[0] ;
 assign io_oeb[12] = \top_I.io_oeb[0] ;
 assign io_oeb[13] = \top_I.io_oeb[0] ;
 assign io_oeb[14] = \top_I.io_oeb[0] ;
 assign io_oeb[15] = \top_I.io_oeb[0] ;
 assign io_oeb[1] = \top_I.io_oeb[0] ;
 assign io_oeb[2] = \top_I.io_oeb[0] ;
 assign io_oeb[32] = \top_I.io_oeb[0] ;
 assign io_oeb[34] = \top_I.io_oeb[0] ;
 assign io_oeb[36] = \top_I.io_oeb[0] ;
 assign io_oeb[3] = \top_I.io_oeb[0] ;
 assign io_oeb[6] = \top_I.io_oeb[0] ;
 assign io_oeb[7] = \top_I.io_oeb[0] ;
 assign io_oeb[8] = \top_I.io_oeb[0] ;
 assign io_oeb[9] = \top_I.io_oeb[0] ;
 assign io_out[0] = \top_I.io_oeb[0] ;
 assign io_out[10] = \top_I.io_oeb[0] ;
 assign io_out[11] = \top_I.io_oeb[0] ;
 assign io_out[12] = \top_I.io_oeb[0] ;
 assign io_out[13] = \top_I.io_oeb[0] ;
 assign io_out[14] = \top_I.io_oeb[0] ;
 assign io_out[15] = \top_I.io_oeb[0] ;
 assign io_out[1] = \top_I.io_oeb[0] ;
 assign io_out[2] = \top_I.io_oeb[0] ;
 assign io_out[3] = \top_I.io_oeb[0] ;
 assign io_out[6] = \top_I.io_oeb[0] ;
 assign io_out[7] = \top_I.io_oeb[0] ;
 assign io_out[8] = \top_I.io_oeb[0] ;
 assign io_out[9] = \top_I.io_oeb[0] ;
 assign io_out[5] = user_clock2;
 assign io_oeb[16] = wbs_ack_o;
 assign io_oeb[17] = wbs_ack_o;
 assign io_oeb[18] = wbs_ack_o;
 assign io_oeb[19] = wbs_ack_o;
 assign io_oeb[20] = wbs_ack_o;
 assign io_oeb[21] = wbs_ack_o;
 assign io_oeb[22] = wbs_ack_o;
 assign io_oeb[23] = wbs_ack_o;
 assign io_oeb[33] = wbs_ack_o;
 assign io_oeb[35] = wbs_ack_o;
 assign io_oeb[37] = wbs_ack_o;
 assign io_oeb[4] = wbs_ack_o;
 assign io_oeb[5] = wbs_ack_o;
 assign io_out[32] = wbs_ack_o;
 assign io_out[33] = wbs_ack_o;
 assign io_out[34] = wbs_ack_o;
 assign io_out[35] = wbs_ack_o;
 assign io_out[36] = wbs_ack_o;
 assign io_out[37] = wbs_ack_o;
 assign io_out[4] = wbs_ack_o;
 assign la_data_out[0] = wbs_ack_o;
 assign la_data_out[100] = wbs_ack_o;
 assign la_data_out[101] = wbs_ack_o;
 assign la_data_out[102] = wbs_ack_o;
 assign la_data_out[103] = wbs_ack_o;
 assign la_data_out[104] = wbs_ack_o;
 assign la_data_out[105] = wbs_ack_o;
 assign la_data_out[106] = wbs_ack_o;
 assign la_data_out[107] = wbs_ack_o;
 assign la_data_out[108] = wbs_ack_o;
 assign la_data_out[109] = wbs_ack_o;
 assign la_data_out[10] = wbs_ack_o;
 assign la_data_out[110] = wbs_ack_o;
 assign la_data_out[111] = wbs_ack_o;
 assign la_data_out[112] = wbs_ack_o;
 assign la_data_out[113] = wbs_ack_o;
 assign la_data_out[114] = wbs_ack_o;
 assign la_data_out[115] = wbs_ack_o;
 assign la_data_out[116] = wbs_ack_o;
 assign la_data_out[117] = wbs_ack_o;
 assign la_data_out[118] = wbs_ack_o;
 assign la_data_out[119] = wbs_ack_o;
 assign la_data_out[11] = wbs_ack_o;
 assign la_data_out[120] = wbs_ack_o;
 assign la_data_out[121] = wbs_ack_o;
 assign la_data_out[122] = wbs_ack_o;
 assign la_data_out[123] = wbs_ack_o;
 assign la_data_out[124] = wbs_ack_o;
 assign la_data_out[125] = wbs_ack_o;
 assign la_data_out[126] = wbs_ack_o;
 assign la_data_out[127] = wbs_ack_o;
 assign la_data_out[12] = wbs_ack_o;
 assign la_data_out[13] = wbs_ack_o;
 assign la_data_out[14] = wbs_ack_o;
 assign la_data_out[15] = wbs_ack_o;
 assign la_data_out[16] = wbs_ack_o;
 assign la_data_out[17] = wbs_ack_o;
 assign la_data_out[18] = wbs_ack_o;
 assign la_data_out[19] = wbs_ack_o;
 assign la_data_out[1] = wbs_ack_o;
 assign la_data_out[20] = wbs_ack_o;
 assign la_data_out[21] = wbs_ack_o;
 assign la_data_out[22] = wbs_ack_o;
 assign la_data_out[23] = wbs_ack_o;
 assign la_data_out[24] = wbs_ack_o;
 assign la_data_out[25] = wbs_ack_o;
 assign la_data_out[26] = wbs_ack_o;
 assign la_data_out[27] = wbs_ack_o;
 assign la_data_out[28] = wbs_ack_o;
 assign la_data_out[29] = wbs_ack_o;
 assign la_data_out[2] = wbs_ack_o;
 assign la_data_out[30] = wbs_ack_o;
 assign la_data_out[31] = wbs_ack_o;
 assign la_data_out[32] = wbs_ack_o;
 assign la_data_out[33] = wbs_ack_o;
 assign la_data_out[34] = wbs_ack_o;
 assign la_data_out[35] = wbs_ack_o;
 assign la_data_out[36] = wbs_ack_o;
 assign la_data_out[37] = wbs_ack_o;
 assign la_data_out[38] = wbs_ack_o;
 assign la_data_out[39] = wbs_ack_o;
 assign la_data_out[3] = wbs_ack_o;
 assign la_data_out[40] = wbs_ack_o;
 assign la_data_out[41] = wbs_ack_o;
 assign la_data_out[42] = wbs_ack_o;
 assign la_data_out[43] = wbs_ack_o;
 assign la_data_out[44] = wbs_ack_o;
 assign la_data_out[45] = wbs_ack_o;
 assign la_data_out[46] = wbs_ack_o;
 assign la_data_out[47] = wbs_ack_o;
 assign la_data_out[48] = wbs_ack_o;
 assign la_data_out[49] = wbs_ack_o;
 assign la_data_out[4] = wbs_ack_o;
 assign la_data_out[50] = wbs_ack_o;
 assign la_data_out[51] = wbs_ack_o;
 assign la_data_out[52] = wbs_ack_o;
 assign la_data_out[53] = wbs_ack_o;
 assign la_data_out[54] = wbs_ack_o;
 assign la_data_out[55] = wbs_ack_o;
 assign la_data_out[56] = wbs_ack_o;
 assign la_data_out[57] = wbs_ack_o;
 assign la_data_out[58] = wbs_ack_o;
 assign la_data_out[59] = wbs_ack_o;
 assign la_data_out[5] = wbs_ack_o;
 assign la_data_out[60] = wbs_ack_o;
 assign la_data_out[61] = wbs_ack_o;
 assign la_data_out[62] = wbs_ack_o;
 assign la_data_out[63] = wbs_ack_o;
 assign la_data_out[64] = wbs_ack_o;
 assign la_data_out[65] = wbs_ack_o;
 assign la_data_out[66] = wbs_ack_o;
 assign la_data_out[67] = wbs_ack_o;
 assign la_data_out[68] = wbs_ack_o;
 assign la_data_out[69] = wbs_ack_o;
 assign la_data_out[6] = wbs_ack_o;
 assign la_data_out[70] = wbs_ack_o;
 assign la_data_out[71] = wbs_ack_o;
 assign la_data_out[72] = wbs_ack_o;
 assign la_data_out[73] = wbs_ack_o;
 assign la_data_out[74] = wbs_ack_o;
 assign la_data_out[75] = wbs_ack_o;
 assign la_data_out[76] = wbs_ack_o;
 assign la_data_out[77] = wbs_ack_o;
 assign la_data_out[78] = wbs_ack_o;
 assign la_data_out[79] = wbs_ack_o;
 assign la_data_out[7] = wbs_ack_o;
 assign la_data_out[80] = wbs_ack_o;
 assign la_data_out[81] = wbs_ack_o;
 assign la_data_out[82] = wbs_ack_o;
 assign la_data_out[83] = wbs_ack_o;
 assign la_data_out[84] = wbs_ack_o;
 assign la_data_out[85] = wbs_ack_o;
 assign la_data_out[86] = wbs_ack_o;
 assign la_data_out[87] = wbs_ack_o;
 assign la_data_out[88] = wbs_ack_o;
 assign la_data_out[89] = wbs_ack_o;
 assign la_data_out[8] = wbs_ack_o;
 assign la_data_out[90] = wbs_ack_o;
 assign la_data_out[91] = wbs_ack_o;
 assign la_data_out[92] = wbs_ack_o;
 assign la_data_out[93] = wbs_ack_o;
 assign la_data_out[94] = wbs_ack_o;
 assign la_data_out[95] = wbs_ack_o;
 assign la_data_out[96] = wbs_ack_o;
 assign la_data_out[97] = wbs_ack_o;
 assign la_data_out[98] = wbs_ack_o;
 assign la_data_out[99] = wbs_ack_o;
 assign la_data_out[9] = wbs_ack_o;
 assign user_irq[0] = wbs_ack_o;
 assign user_irq[1] = wbs_ack_o;
 assign user_irq[2] = wbs_ack_o;
 assign wbs_dat_o[0] = wbs_ack_o;
 assign wbs_dat_o[10] = wbs_ack_o;
 assign wbs_dat_o[11] = wbs_ack_o;
 assign wbs_dat_o[12] = wbs_ack_o;
 assign wbs_dat_o[13] = wbs_ack_o;
 assign wbs_dat_o[14] = wbs_ack_o;
 assign wbs_dat_o[15] = wbs_ack_o;
 assign wbs_dat_o[16] = wbs_ack_o;
 assign wbs_dat_o[17] = wbs_ack_o;
 assign wbs_dat_o[18] = wbs_ack_o;
 assign wbs_dat_o[19] = wbs_ack_o;
 assign wbs_dat_o[1] = wbs_ack_o;
 assign wbs_dat_o[20] = wbs_ack_o;
 assign wbs_dat_o[21] = wbs_ack_o;
 assign wbs_dat_o[22] = wbs_ack_o;
 assign wbs_dat_o[23] = wbs_ack_o;
 assign wbs_dat_o[24] = wbs_ack_o;
 assign wbs_dat_o[25] = wbs_ack_o;
 assign wbs_dat_o[26] = wbs_ack_o;
 assign wbs_dat_o[27] = wbs_ack_o;
 assign wbs_dat_o[28] = wbs_ack_o;
 assign wbs_dat_o[29] = wbs_ack_o;
 assign wbs_dat_o[2] = wbs_ack_o;
 assign wbs_dat_o[30] = wbs_ack_o;
 assign wbs_dat_o[31] = wbs_ack_o;
 assign wbs_dat_o[3] = wbs_ack_o;
 assign wbs_dat_o[4] = wbs_ack_o;
 assign wbs_dat_o[5] = wbs_ack_o;
 assign wbs_dat_o[6] = wbs_ack_o;
 assign wbs_dat_o[7] = wbs_ack_o;
 assign wbs_dat_o[8] = wbs_ack_o;
 assign wbs_dat_o[9] = wbs_ack_o;
endmodule
