module tt_um_delay_line_tmng (VGND,
    VPWR,
    clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input VGND;
 input VPWR;
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire net1;
 wire net2;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net5;
 wire net6;
 wire \tmng_0._e_621 ;
 wire \tmng_0._e_630 ;
 wire \tmng_0._e_642 ;
 wire \tmng_0._e_647 ;
 wire \tmng_0._e_650 ;
 wire \tmng_0._e_662 ;
 wire \tmng_0.opa ;
 wire \tmng_0.opb ;
 wire \tmng_0.shift_reg_0.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_9.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_9.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_9.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.s1_val ;
 wire \tmng_0.shift_reg_0.shift_reg100_0.val ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_9.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_9.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_9.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_1.s1_val ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_9.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_9.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_9.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_2.s1_val ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_9.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_9.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_9.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_3.s1_val ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_4.s1_val ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_9.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_9.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_9.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_5.s1_val ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_9.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_9.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_9.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_6.s1_val ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_9.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_9.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_9.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg100_7.s1_val ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_0.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_39.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_39.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_39.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.dlygate_1.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.output__ ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_9.dlygate_0.X_mut ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_9.dlygate_1.A ;
 wire \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_9.dlygate_1.X_mut ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_179 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_41_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_279 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_291 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_177 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_189 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_201 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_48_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_322 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_182 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_124 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_177 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_79_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__mux2_1 _022_ (.A0(\tmng_0.shift_reg_0.output__ ),
    .A1(\tmng_0._e_650 ),
    .S(\tmng_0._e_647 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_010_));
 sky130_fd_sc_hd__and3_1 _023_ (.A(\tmng_0.opb ),
    .B(\tmng_0.opa ),
    .C(\tmng_0._e_642 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_011_));
 sky130_fd_sc_hd__o21ba_1 _024_ (.A1(net38),
    .A2(_010_),
    .B1_N(_011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.val ));
 sky130_fd_sc_hd__mux2_1 _025_ (.A0(net41),
    .A1(\tmng_0.shift_reg_0.output__ ),
    .S(\tmng_0._e_621 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_012_));
 sky130_fd_sc_hd__clkbuf_1 _026_ (.A(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _027_ (.A0(uo_out[0]),
    .A1(\tmng_0.shift_reg_0.output__ ),
    .S(\tmng_0._e_662 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_013_));
 sky130_fd_sc_hd__clkbuf_1 _028_ (.A(_013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _029_ (.A0(uo_out[1]),
    .A1(uo_out[0]),
    .S(\tmng_0._e_662 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_014_));
 sky130_fd_sc_hd__clkbuf_1 _030_ (.A(_014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _031_ (.A0(uo_out[2]),
    .A1(uo_out[1]),
    .S(\tmng_0._e_662 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_015_));
 sky130_fd_sc_hd__clkbuf_1 _032_ (.A(_015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _033_ (.A0(uo_out[3]),
    .A1(uo_out[2]),
    .S(\tmng_0._e_662 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_016_));
 sky130_fd_sc_hd__clkbuf_1 _034_ (.A(_016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _035_ (.A0(uo_out[4]),
    .A1(uo_out[3]),
    .S(\tmng_0._e_662 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_017_));
 sky130_fd_sc_hd__clkbuf_1 _036_ (.A(_017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _037_ (.A0(uo_out[5]),
    .A1(uo_out[4]),
    .S(\tmng_0._e_662 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_018_));
 sky130_fd_sc_hd__clkbuf_1 _038_ (.A(_018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _039_ (.A0(uo_out[6]),
    .A1(uo_out[5]),
    .S(\tmng_0._e_662 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_019_));
 sky130_fd_sc_hd__clkbuf_1 _040_ (.A(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _041_ (.A0(uo_out[7]),
    .A1(uo_out[6]),
    .S(\tmng_0._e_662 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_020_));
 sky130_fd_sc_hd__clkbuf_1 _042_ (.A(_020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _043_ (.A0(net39),
    .A1(\tmng_0.shift_reg_0.output__ ),
    .S(\tmng_0._e_630 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_021_));
 sky130_fd_sc_hd__clkbuf_1 _044_ (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_009_));
 sky130_fd_sc_hd__dfxtp_1 _045_ (.CLK(clknet_leaf_17_clk),
    .D(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0._e_642 ));
 sky130_fd_sc_hd__dfxtp_1 _046_ (.CLK(clknet_leaf_17_clk),
    .D(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0._e_647 ));
 sky130_fd_sc_hd__dfxtp_1 _047_ (.CLK(clknet_leaf_17_clk),
    .D(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0._e_650 ));
 sky130_fd_sc_hd__dfxtp_1 _048_ (.CLK(clknet_leaf_17_clk),
    .D(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0._e_621 ));
 sky130_fd_sc_hd__dfxtp_1 _049_ (.CLK(clknet_leaf_17_clk),
    .D(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0._e_630 ));
 sky130_fd_sc_hd__dfxtp_2 _050_ (.CLK(clknet_leaf_17_clk),
    .D(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0._e_662 ));
 sky130_fd_sc_hd__dfxtp_1 _051_ (.CLK(clknet_leaf_17_clk),
    .D(_000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.opa ));
 sky130_fd_sc_hd__dfxtp_1 _052_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _053_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _054_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _055_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _056_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _057_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _058_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _059_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _060_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _061_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _062_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _063_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _064_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _065_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _066_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _067_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _068_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _069_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _070_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _071_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _072_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _073_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _074_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _075_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _076_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _077_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _078_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _079_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _080_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _081_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _082_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _083_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _084_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _085_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _086_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _087_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _088_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _089_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _090_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _091_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _092_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _093_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _094_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _095_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _096_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _097_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _098_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _099_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _100_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _101_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _102_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _103_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _104_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _105_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _106_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _107_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _108_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _109_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _110_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _111_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _112_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _113_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _114_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _115_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _116_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _117_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _118_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _119_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _120_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _121_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _122_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _123_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _124_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _125_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _126_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _127_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _128_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _129_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _130_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_9.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _131_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_9.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_9.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _132_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _133_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _134_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _135_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _136_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _137_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _138_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _139_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _140_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _141_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _142_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _143_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _144_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _145_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _146_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _147_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _148_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _149_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _150_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_0.val ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.s1_val ));
 sky130_fd_sc_hd__dfxtp_1 _151_ (.CLK(clknet_leaf_17_clk),
    .D(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _152_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _153_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _154_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _155_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _156_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _157_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _158_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _159_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _160_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _161_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _162_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _163_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _164_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _165_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _166_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _167_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _168_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _169_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _170_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _171_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _172_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _173_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _174_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _175_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _176_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _177_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _178_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _179_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _180_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _181_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _182_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _183_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _184_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _185_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _186_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _187_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _188_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _189_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _190_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _191_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _192_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _193_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _194_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _195_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _196_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _197_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _198_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _199_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _200_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _201_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _202_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _203_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _204_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _205_ (.CLK(clknet_leaf_6_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _206_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _207_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _208_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _209_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _210_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _211_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _212_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _213_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _214_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _215_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _216_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _217_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _218_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _219_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _220_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _221_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _222_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _223_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _224_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _225_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _226_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _227_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _228_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _229_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _230_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_9.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _231_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_9.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_9.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _232_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _233_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _234_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _235_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _236_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _237_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _238_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _239_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _240_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _241_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _242_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _243_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _244_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _245_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _246_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _247_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _248_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _249_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _250_ (.CLK(clknet_leaf_7_clk),
    .D(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.s1_val ));
 sky130_fd_sc_hd__dfxtp_1 _251_ (.CLK(clknet_leaf_7_clk),
    .D(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _252_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _253_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _254_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _255_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _256_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _257_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _258_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _259_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _260_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _261_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _262_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _263_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _264_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _265_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _266_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _267_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _268_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _269_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _270_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _271_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _272_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _273_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _274_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _275_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _276_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _277_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _278_ (.CLK(clknet_leaf_37_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _279_ (.CLK(clknet_leaf_37_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _280_ (.CLK(clknet_leaf_37_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _281_ (.CLK(clknet_leaf_37_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _282_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _283_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _284_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _285_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _286_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _287_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _288_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _289_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _290_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _291_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _292_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _293_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _294_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _295_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _296_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _297_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _298_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _299_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _300_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _301_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _302_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _303_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _304_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _305_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _306_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _307_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _308_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _309_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _310_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _311_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _312_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _313_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _314_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _315_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _316_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _317_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _318_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _319_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _320_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _321_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _322_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _323_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _324_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _325_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _326_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _327_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _328_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _329_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _330_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_9.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _331_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_9.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_9.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _332_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _333_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _334_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _335_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _336_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _337_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _338_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _339_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _340_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _341_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _342_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _343_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _344_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _345_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _346_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _347_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _348_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _349_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _350_ (.CLK(clknet_leaf_4_clk),
    .D(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.s1_val ));
 sky130_fd_sc_hd__dfxtp_1 _351_ (.CLK(clknet_leaf_3_clk),
    .D(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _352_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _353_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _354_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _355_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _356_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _357_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _358_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _359_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _360_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _361_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _362_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _363_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _364_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _365_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _366_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _367_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _368_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _369_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _370_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _371_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _372_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _373_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _374_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _375_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _376_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _377_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _378_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _379_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _380_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _381_ (.CLK(clknet_leaf_37_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _382_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _383_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _384_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _385_ (.CLK(clknet_leaf_37_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _386_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _387_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _388_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _389_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _390_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _391_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _392_ (.CLK(clknet_leaf_0_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _393_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _394_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _395_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _396_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _397_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _398_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _399_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _400_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _401_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _402_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _403_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _404_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _405_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _406_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _407_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _408_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _409_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _410_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _411_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _412_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _413_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _414_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _415_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _416_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _417_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _418_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _419_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _420_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _421_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _422_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _423_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _424_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _425_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _426_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _427_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _428_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _429_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _430_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_9.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _431_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_9.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_9.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _432_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _433_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _434_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _435_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _436_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _437_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _438_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _439_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _440_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _441_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _442_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _443_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _444_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _445_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _446_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _447_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _448_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _449_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _450_ (.CLK(clknet_leaf_32_clk),
    .D(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.s1_val ));
 sky130_fd_sc_hd__dfxtp_1 _451_ (.CLK(clknet_leaf_32_clk),
    .D(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _452_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _453_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _454_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _455_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _456_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _457_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _458_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _459_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _460_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _461_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _462_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _463_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _464_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _465_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _466_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _467_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _468_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _469_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _470_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _471_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _472_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _473_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _474_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _475_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _476_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _477_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _478_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _479_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _480_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _481_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _482_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _483_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _484_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _485_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _486_ (.CLK(clknet_leaf_36_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _487_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _488_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _489_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _490_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _491_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _492_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _493_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _494_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _495_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _496_ (.CLK(clknet_leaf_35_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _497_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _498_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _499_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _500_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _501_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _502_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _503_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _504_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _505_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _506_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _507_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _508_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _509_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _510_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _511_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _512_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _513_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _514_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _515_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _516_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _517_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _518_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _519_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _520_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _521_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _522_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _523_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _524_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _525_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _526_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _527_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _528_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _529_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _530_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _531_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _532_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _533_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _534_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _535_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _536_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _537_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _538_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _539_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _540_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _541_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _542_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _543_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _544_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _545_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _546_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _547_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _548_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _549_ (.CLK(clknet_leaf_34_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _550_ (.CLK(clknet_leaf_34_clk),
    .D(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.s1_val ));
 sky130_fd_sc_hd__dfxtp_1 _551_ (.CLK(clknet_leaf_34_clk),
    .D(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _552_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _553_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _554_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _555_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _556_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _557_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _558_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _559_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _560_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _561_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _562_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _563_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _564_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _565_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _566_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _567_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _568_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _569_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _570_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _571_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _572_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _573_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _574_ (.CLK(clknet_leaf_32_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _575_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _576_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _577_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _578_ (.CLK(clknet_leaf_33_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _579_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _580_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _581_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _582_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _583_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _584_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _585_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _586_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _587_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _588_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _589_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _590_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _591_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _592_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _593_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _594_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _595_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _596_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _597_ (.CLK(clknet_leaf_30_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _598_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _599_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _600_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _601_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _602_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _603_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _604_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _605_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _606_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _607_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _608_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _609_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _610_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _611_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _612_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _613_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _614_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _615_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _616_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _617_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _618_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _619_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _620_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _621_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _622_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _623_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _624_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _625_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _626_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _627_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _628_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _629_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _630_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_9.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _631_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_9.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_9.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _632_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _633_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _634_ (.CLK(clknet_leaf_27_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _635_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _636_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _637_ (.CLK(clknet_leaf_26_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _638_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _639_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _640_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _641_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _642_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _643_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _644_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _645_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _646_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _647_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _648_ (.CLK(clknet_leaf_29_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _649_ (.CLK(clknet_leaf_28_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _650_ (.CLK(clknet_leaf_29_clk),
    .D(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.s1_val ));
 sky130_fd_sc_hd__dfxtp_1 _651_ (.CLK(clknet_leaf_29_clk),
    .D(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _652_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _653_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _654_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _655_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _656_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _657_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _658_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _659_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _660_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _661_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _662_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _663_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _664_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _665_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _666_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _667_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _668_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _669_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _670_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _671_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _672_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _673_ (.CLK(clknet_leaf_1_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _674_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _675_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _676_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _677_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _678_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _679_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _680_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _681_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _682_ (.CLK(clknet_leaf_2_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _683_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _684_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _685_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _686_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _687_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _688_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _689_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _690_ (.CLK(clknet_leaf_3_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _691_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _692_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _693_ (.CLK(clknet_leaf_31_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _694_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _695_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _696_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _697_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _698_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _699_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _700_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _701_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _702_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _703_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _704_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _705_ (.CLK(clknet_leaf_22_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _706_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _707_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _708_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _709_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _710_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _711_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _712_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _713_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _714_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _715_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _716_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _717_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _718_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _719_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _720_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _721_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _722_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _723_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _724_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _725_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _726_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _727_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _728_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _729_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _730_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_9.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _731_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_9.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_9.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _732_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _733_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _734_ (.CLK(clknet_leaf_25_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _735_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _736_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _737_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _738_ (.CLK(clknet_leaf_23_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _739_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _740_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _741_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _742_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _743_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _744_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _745_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _746_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _747_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _748_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _749_ (.CLK(clknet_leaf_24_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _750_ (.CLK(clknet_leaf_24_clk),
    .D(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.s1_val ));
 sky130_fd_sc_hd__dfxtp_1 _751_ (.CLK(clknet_leaf_24_clk),
    .D(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _752_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _753_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _754_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _755_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _756_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _757_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _758_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _759_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _760_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _761_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _762_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _763_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _764_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _765_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _766_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _767_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _768_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _769_ (.CLK(clknet_leaf_9_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _770_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _771_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _772_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _773_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _774_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _775_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _776_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _777_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _778_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _779_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _780_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _781_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _782_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _783_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _784_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _785_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _786_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _787_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _788_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _789_ (.CLK(clknet_leaf_8_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _790_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _791_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _792_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _793_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _794_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _795_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _796_ (.CLK(clknet_leaf_5_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _797_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _798_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _799_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _800_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _801_ (.CLK(clknet_leaf_7_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _802_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _803_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _804_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _805_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _806_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _807_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _808_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _809_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _810_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _811_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _812_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _813_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _814_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _815_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _816_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _817_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _818_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _819_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _820_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _821_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _822_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _823_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _824_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _825_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _826_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _827_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _828_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _829_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _830_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_9.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _831_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_9.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_9.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _832_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _833_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _834_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _835_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _836_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _837_ (.CLK(clknet_leaf_13_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _838_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _839_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _840_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _841_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _842_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _843_ (.CLK(clknet_leaf_12_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _844_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _845_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _846_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _847_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _848_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _849_ (.CLK(clknet_leaf_4_clk),
    .D(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _850_ (.CLK(clknet_leaf_5_clk),
    .D(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.s1_val ));
 sky130_fd_sc_hd__dfxtp_1 _851_ (.CLK(clknet_leaf_4_clk),
    .D(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _852_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_39.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _853_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_39.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_39.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _854_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _855_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _856_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _857_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _858_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _859_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _860_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _861_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _862_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _863_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _864_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _865_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _866_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _867_ (.CLK(clknet_leaf_18_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _868_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _869_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _870_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _871_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _872_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _873_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _874_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _875_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _876_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _877_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _878_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _879_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _880_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _881_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _882_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _883_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _884_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _885_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _886_ (.CLK(clknet_leaf_20_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _887_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _888_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _889_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _890_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _891_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _892_ (.CLK(clknet_leaf_19_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _893_ (.CLK(clknet_leaf_21_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _894_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _895_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _896_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _897_ (.CLK(clknet_leaf_14_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _898_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _899_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _900_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _901_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _902_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _903_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _904_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _905_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _906_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _907_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _908_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _909_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _910_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _911_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _912_ (.CLK(clknet_leaf_17_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_9.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_0.A ));
 sky130_fd_sc_hd__dfxtp_1 _913_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_9.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_9.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _914_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _915_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _916_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _917_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _918_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _919_ (.CLK(clknet_leaf_16_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _920_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _921_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _922_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _923_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _924_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _925_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _926_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _927_ (.CLK(clknet_leaf_15_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _928_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _929_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_1 _930_ (.CLK(clknet_leaf_11_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.dlygate_1.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.output__ ));
 sky130_fd_sc_hd__dfxtp_1 _931_ (.CLK(clknet_leaf_10_clk),
    .D(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.dlygate_0.X_mut ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.dlygate_1.A ));
 sky130_fd_sc_hd__dfxtp_2 _932_ (.CLK(clknet_leaf_15_clk),
    .D(_001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__dfxtp_2 _933_ (.CLK(clknet_leaf_10_clk),
    .D(_002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__dfxtp_2 _934_ (.CLK(clknet_leaf_10_clk),
    .D(_003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__dfxtp_2 _935_ (.CLK(clknet_leaf_10_clk),
    .D(_004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[3]));
 sky130_fd_sc_hd__dfxtp_2 _936_ (.CLK(clknet_leaf_10_clk),
    .D(_005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__dfxtp_2 _937_ (.CLK(clknet_leaf_10_clk),
    .D(_006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfxtp_2 _938_ (.CLK(clknet_leaf_10_clk),
    .D(_007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfxtp_2 _939_ (.CLK(clknet_leaf_10_clk),
    .D(_008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(uo_out[7]));
 sky130_fd_sc_hd__dfxtp_1 _940_ (.CLK(clknet_leaf_17_clk),
    .D(_009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tmng_0.opb ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_2_2__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\tmng_0.shift_reg_0.shift_reg100_2.s1_val ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\tmng_0.shift_reg_0.shift_reg100_0.s1_val ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\tmng_0.shift_reg_0.shift_reg100_4.s1_val ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\tmng_0.shift_reg_0.shift_reg100_1.s1_val ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\tmng_0.shift_reg_0.shift_reg100_5.s1_val ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\tmng_0._e_642 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\tmng_0.opb ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\tmng_0.opa ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\tmng_0.shift_reg_0.shift_reg100_7.s1_val ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\tmng_0.shift_reg_0.shift_reg100_3.s1_val ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\tmng_0.shift_reg_0.shift_reg100_6.s1_val ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_0.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_10.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_11.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_12.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_13.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_14.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_15.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_16.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_17.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_18.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_1.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_19.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_20.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_21.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_22.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_23.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_24.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_25.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_26.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_27.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_28.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_2.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_29.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_30.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_31.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_32.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_33.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_34.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_35.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_36.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_37.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_38.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_3.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_39.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_40.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_41.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_42.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_43.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_44.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_45.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_46.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_47.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_48.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_4.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_5.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_6.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_7.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_9.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_8.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_9.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_0.inv_reg_9.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_9.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_0.inv_reg_9.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_0.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_10.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_11.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_12.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_13.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_14.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_15.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_16.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_17.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_18.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_1.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_19.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_20.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_21.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_22.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_23.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_24.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_25.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_26.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_27.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_28.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_2.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_29.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_30.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_31.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_32.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_33.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_34.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_35.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_36.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_37.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_38.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_3.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_39.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_40.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_41.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_42.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_43.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_44.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_45.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_46.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_47.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_48.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_4.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_5.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_6.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_7.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_9.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_8.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_9.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_1.inv_reg_9.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_9.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_1.inv_reg_9.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_0.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_10.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_11.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_12.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_13.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_14.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_15.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_16.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_17.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_18.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_1.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_19.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_20.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_21.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_22.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_23.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_24.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_25.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_26.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_27.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_28.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_2.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_29.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_30.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_31.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_32.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_33.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_34.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_35.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_36.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_37.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_38.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_3.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_39.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_40.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_41.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_42.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_43.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_44.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_45.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_46.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_47.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_48.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_4.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_5.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_6.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_7.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_9.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_8.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_9.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_2.inv_reg_9.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_9.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_2.inv_reg_9.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_0.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_10.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_11.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_12.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_13.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_14.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_15.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_16.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_17.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_18.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_1.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_19.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_20.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_21.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_22.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_23.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_24.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_25.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_26.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_27.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_28.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_2.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_29.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_30.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_31.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_32.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_33.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_34.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_35.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_36.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_37.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_38.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_3.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_39.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_40.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_41.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_42.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_43.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_44.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_45.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_46.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_47.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_48.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_4.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_5.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_6.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_7.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_9.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_8.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_9.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_3.inv_reg_9.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_9.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_3.inv_reg_9.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_0.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_10.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_11.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_12.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_13.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_14.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_15.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_16.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_17.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_18.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_1.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_19.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_20.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_21.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_22.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_23.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_24.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_25.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_26.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_27.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_28.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_2.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_29.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_30.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_31.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_32.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_33.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_34.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_35.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_36.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_37.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_38.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_3.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_39.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_40.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_41.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_42.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_43.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_44.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_45.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_46.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_47.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_48.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_4.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_5.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_6.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_7.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_8.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_4.inv_reg_9.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_0.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_10.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_11.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_12.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_13.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_14.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_15.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_16.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_17.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_18.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_1.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_19.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_20.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_21.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_22.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_23.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_24.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_25.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_26.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_27.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_28.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_2.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_29.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_30.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_31.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_32.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_33.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_34.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_35.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_36.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_37.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_38.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_3.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_39.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_40.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_41.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_42.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_43.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_44.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_45.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_46.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_47.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_48.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_4.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_5.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_6.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_7.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_9.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_8.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_9.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_5.inv_reg_9.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_9.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_5.inv_reg_9.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_0.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_10.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_11.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_12.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_13.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_14.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_15.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_16.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_17.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_18.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_1.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_19.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_20.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_21.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_22.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_23.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_24.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_25.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_26.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_27.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_28.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_2.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_29.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_30.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_31.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_32.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_33.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_34.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_35.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_36.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_37.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_38.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_3.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_39.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_40.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_41.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_42.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_43.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_44.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_45.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_46.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_47.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_48.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_4.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_5.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_6.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_7.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_9.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_8.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_9.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_6.inv_reg_9.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_9.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_6.inv_reg_9.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_0.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_10.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_11.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_12.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_13.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_14.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_15.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_16.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_17.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_18.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_1.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_19.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_20.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_21.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_22.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_23.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_24.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_25.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_26.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_27.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_28.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_2.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_29.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_30.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_31.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_32.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_33.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_34.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_35.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_36.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_37.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_38.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_3.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_39.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_40.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_41.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_42.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_43.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_44.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_45.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_46.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_47.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_4.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_5.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_6.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_7.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_9.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_8.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_9.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg100_7.inv_reg_9.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_9.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_9.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg100_7.inv_reg_48.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_0.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_10.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_11.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_12.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_13.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_14.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_15.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_16.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_17.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_18.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_1.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_19.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_20.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_21.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_22.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_23.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_24.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_25.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_26.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_27.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_28.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_2.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_29.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_30.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_31.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_32.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_33.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_34.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_35.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_36.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_37.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_39.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_38.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_39.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_39.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_39.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_39.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_3.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_4.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_5.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_6.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_7.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.dlygate_1.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_9.dlygate_0.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_8.output__ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_9.dlygate_0.X_mut ));
 sky130_fd_sc_hd__dlygate4sd3_1 \tmng_0.shift_reg_0.shift_reg80_0.inv_reg_9.dlygate_1.sky130_fd_sc_hd__dlygate4sd3_1_0  (.A(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_9.dlygate_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\tmng_0.shift_reg_0.shift_reg80_0.inv_reg_9.dlygate_1.X_mut ));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net10));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net11));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net12));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net13));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net14));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net15));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net16));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net17));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net18));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net19));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net20));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net21));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net22));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net7));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net8));
 sky130_fd_sc_hd__conb_1 tt_um_delay_line_tmng_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net9));
 assign uio_oe[0] = net7;
 assign uio_oe[1] = net8;
 assign uio_oe[2] = net9;
 assign uio_oe[3] = net10;
 assign uio_oe[4] = net11;
 assign uio_oe[5] = net12;
 assign uio_oe[6] = net13;
 assign uio_oe[7] = net14;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[4] = net19;
 assign uio_out[5] = net20;
 assign uio_out[6] = net21;
 assign uio_out[7] = net22;
endmodule
