module tt_um_litneet64_ro_puf (VGND,
    VPWR,
    clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input VGND;
 input VPWR;
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[0] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[10] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[11] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[12] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[13] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[14] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[15] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[1] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[2] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[3] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[4] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[5] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[6] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[7] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[8] ;
 wire \genblk1[0].puf_buffer.cnt_1.ctr[9] ;
 wire \genblk1[0].puf_buffer.cnt_1.finish ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[0] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[10] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[11] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[12] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[13] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[14] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[15] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[1] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[2] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[3] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[4] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[5] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[6] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[7] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[8] ;
 wire \genblk1[0].puf_buffer.cnt_2.ctr[9] ;
 wire \genblk1[0].puf_buffer.cnt_2.finish ;
 wire \genblk1[0].puf_buffer.race_arb.marked_1 ;
 wire \genblk1[0].puf_buffer.race_arb.marked_2 ;
 wire \genblk1[0].puf_buffer.race_arb.resp ;
 wire \genblk1[0].puf_buffer.race_arb.win_1 ;
 wire \genblk1[0].puf_buffer.ro_array_1[0].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[0].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[0].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[0].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[0].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[0].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[0].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[0].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[10].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[10].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[10].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[10].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[10].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[10].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[10].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[10].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[11].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[11].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[11].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[11].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[11].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[11].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[11].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[11].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[12].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[12].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[12].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[12].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[12].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[12].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[12].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[12].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[13].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[13].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[13].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[13].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[13].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[13].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[13].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[13].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[14].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[14].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[14].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[14].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[14].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[14].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[14].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[14].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[15].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[15].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[15].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[15].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[15].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[15].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[15].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[15].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[1].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[1].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[1].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[1].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[1].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[1].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[1].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[1].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[2].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[2].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[2].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[2].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[2].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[2].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[2].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[2].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[3].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[3].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[3].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[3].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[3].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[3].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[3].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[3].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[4].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[4].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[4].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[4].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[4].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[4].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[4].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[4].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[5].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[5].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[5].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[5].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[5].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[5].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[5].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[5].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[6].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[6].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[6].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[6].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[6].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[6].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[6].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[6].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[7].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[7].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[7].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[7].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[7].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[7].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[7].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[7].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[8].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[8].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[8].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[8].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[8].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[8].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[8].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[8].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_1[9].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_1[9].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_1[9].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_1[9].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_1[9].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_1[9].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_1[9].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_1[9].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[0].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[0].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[0].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[0].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[0].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[0].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[0].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[0].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[10].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[10].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[10].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[10].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[10].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[10].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[10].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[10].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[11].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[11].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[11].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[11].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[11].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[11].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[11].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[11].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[12].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[12].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[12].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[12].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[12].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[12].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[12].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[12].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[13].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[13].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[13].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[13].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[13].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[13].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[13].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[13].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[14].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[14].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[14].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[14].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[14].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[14].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[14].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[14].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[15].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[15].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[15].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[15].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[15].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[15].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[15].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[15].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[1].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[1].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[1].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[1].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[1].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[1].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[1].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[1].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[2].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[2].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[2].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[2].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[2].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[2].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[2].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[2].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[3].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[3].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[3].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[3].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[3].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[3].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[3].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[3].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[4].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[4].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[4].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[4].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[4].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[4].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[4].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[4].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[5].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[5].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[5].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[5].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[5].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[5].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[5].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[5].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[6].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[6].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[6].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[6].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[6].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[6].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[6].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[6].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[7].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[7].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[7].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[7].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[7].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[7].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[7].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[7].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[8].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[8].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[8].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[8].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[8].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[8].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[8].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[8].inter_wire[7] ;
 wire \genblk1[0].puf_buffer.ro_array_2[9].inter_wire[0] ;
 wire \genblk1[0].puf_buffer.ro_array_2[9].inter_wire[1] ;
 wire \genblk1[0].puf_buffer.ro_array_2[9].inter_wire[2] ;
 wire \genblk1[0].puf_buffer.ro_array_2[9].inter_wire[3] ;
 wire \genblk1[0].puf_buffer.ro_array_2[9].inter_wire[4] ;
 wire \genblk1[0].puf_buffer.ro_array_2[9].inter_wire[5] ;
 wire \genblk1[0].puf_buffer.ro_array_2[9].inter_wire[6] ;
 wire \genblk1[0].puf_buffer.ro_array_2[9].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[0] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[10] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[11] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[12] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[13] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[14] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[15] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[1] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[2] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[3] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[4] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[5] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[6] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[7] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[8] ;
 wire \genblk1[1].puf_buffer.cnt_1.ctr[9] ;
 wire \genblk1[1].puf_buffer.cnt_1.finish ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[0] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[10] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[11] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[12] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[13] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[14] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[15] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[1] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[2] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[3] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[4] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[5] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[6] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[7] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[8] ;
 wire \genblk1[1].puf_buffer.cnt_2.ctr[9] ;
 wire \genblk1[1].puf_buffer.cnt_2.finish ;
 wire \genblk1[1].puf_buffer.race_arb.marked_1 ;
 wire \genblk1[1].puf_buffer.race_arb.marked_2 ;
 wire \genblk1[1].puf_buffer.race_arb.resp ;
 wire \genblk1[1].puf_buffer.race_arb.win_1 ;
 wire \genblk1[1].puf_buffer.ro_array_1[0].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[0].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[0].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[0].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[0].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[0].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[0].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[0].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[10].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[10].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[10].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[10].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[10].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[10].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[10].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[10].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[11].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[11].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[11].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[11].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[11].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[11].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[11].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[11].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[12].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[12].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[12].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[12].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[12].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[12].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[12].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[12].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[13].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[13].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[13].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[13].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[13].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[13].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[13].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[13].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[14].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[14].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[14].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[14].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[14].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[14].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[14].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[14].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[15].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[15].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[15].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[15].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[15].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[15].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[15].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[15].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[1].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[1].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[1].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[1].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[1].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[1].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[1].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[1].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[2].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[2].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[2].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[2].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[2].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[2].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[2].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[2].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[3].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[3].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[3].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[3].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[3].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[3].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[3].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[3].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[4].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[4].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[4].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[4].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[4].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[4].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[4].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[4].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[5].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[5].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[5].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[5].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[5].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[5].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[5].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[5].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[6].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[6].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[6].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[6].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[6].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[6].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[6].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[6].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[7].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[7].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[7].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[7].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[7].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[7].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[7].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[7].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[8].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[8].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[8].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[8].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[8].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[8].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[8].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[8].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_1[9].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_1[9].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_1[9].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_1[9].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_1[9].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_1[9].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_1[9].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_1[9].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[0].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[0].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[0].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[0].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[0].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[0].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[0].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[0].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[10].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[10].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[10].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[10].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[10].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[10].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[10].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[10].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[11].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[11].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[11].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[11].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[11].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[11].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[11].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[11].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[12].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[12].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[12].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[12].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[12].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[12].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[12].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[12].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[13].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[13].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[13].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[13].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[13].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[13].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[13].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[13].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[14].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[14].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[14].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[14].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[14].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[14].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[14].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[14].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[15].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[15].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[15].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[15].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[15].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[15].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[15].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[15].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[1].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[1].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[1].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[1].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[1].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[1].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[1].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[1].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[2].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[2].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[2].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[2].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[2].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[2].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[2].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[2].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[3].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[3].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[3].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[3].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[3].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[3].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[3].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[3].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[4].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[4].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[4].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[4].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[4].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[4].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[4].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[4].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[5].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[5].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[5].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[5].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[5].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[5].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[5].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[5].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[6].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[6].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[6].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[6].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[6].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[6].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[6].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[6].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[7].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[7].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[7].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[7].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[7].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[7].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[7].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[7].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[8].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[8].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[8].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[8].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[8].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[8].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[8].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[8].inter_wire[7] ;
 wire \genblk1[1].puf_buffer.ro_array_2[9].inter_wire[0] ;
 wire \genblk1[1].puf_buffer.ro_array_2[9].inter_wire[1] ;
 wire \genblk1[1].puf_buffer.ro_array_2[9].inter_wire[2] ;
 wire \genblk1[1].puf_buffer.ro_array_2[9].inter_wire[3] ;
 wire \genblk1[1].puf_buffer.ro_array_2[9].inter_wire[4] ;
 wire \genblk1[1].puf_buffer.ro_array_2[9].inter_wire[5] ;
 wire \genblk1[1].puf_buffer.ro_array_2[9].inter_wire[6] ;
 wire \genblk1[1].puf_buffer.ro_array_2[9].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[0] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[10] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[11] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[12] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[13] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[14] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[15] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[1] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[2] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[3] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[4] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[5] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[6] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[7] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[8] ;
 wire \genblk1[2].puf_buffer.cnt_1.ctr[9] ;
 wire \genblk1[2].puf_buffer.cnt_1.finish ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[0] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[10] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[11] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[12] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[13] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[14] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[15] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[1] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[2] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[3] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[4] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[5] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[6] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[7] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[8] ;
 wire \genblk1[2].puf_buffer.cnt_2.ctr[9] ;
 wire \genblk1[2].puf_buffer.cnt_2.finish ;
 wire \genblk1[2].puf_buffer.race_arb.marked_1 ;
 wire \genblk1[2].puf_buffer.race_arb.marked_2 ;
 wire \genblk1[2].puf_buffer.race_arb.resp ;
 wire \genblk1[2].puf_buffer.race_arb.win_1 ;
 wire \genblk1[2].puf_buffer.ro_array_1[0].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[0].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[0].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[0].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[0].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[0].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[0].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[0].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[10].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[10].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[10].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[10].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[10].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[10].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[10].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[10].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[11].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[11].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[11].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[11].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[11].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[11].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[11].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[11].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[12].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[12].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[12].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[12].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[12].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[12].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[12].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[12].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[13].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[13].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[13].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[13].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[13].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[13].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[13].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[13].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[14].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[14].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[14].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[14].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[14].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[14].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[14].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[14].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[15].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[15].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[15].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[15].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[15].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[15].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[15].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[15].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[1].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[1].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[1].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[1].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[1].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[1].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[1].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[1].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[2].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[2].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[2].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[2].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[2].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[2].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[2].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[2].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[3].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[3].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[3].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[3].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[3].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[3].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[3].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[3].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[4].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[4].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[4].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[4].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[4].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[4].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[4].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[4].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[5].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[5].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[5].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[5].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[5].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[5].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[5].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[5].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[6].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[6].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[6].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[6].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[6].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[6].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[6].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[6].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[7].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[7].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[7].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[7].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[7].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[7].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[7].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[7].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[8].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[8].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[8].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[8].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[8].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[8].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[8].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[8].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_1[9].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_1[9].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_1[9].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_1[9].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_1[9].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_1[9].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_1[9].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_1[9].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[0].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[0].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[0].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[0].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[0].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[0].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[0].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[0].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[10].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[10].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[10].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[10].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[10].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[10].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[10].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[10].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[11].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[11].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[11].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[11].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[11].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[11].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[11].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[11].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[12].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[12].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[12].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[12].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[12].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[12].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[12].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[12].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[13].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[13].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[13].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[13].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[13].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[13].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[13].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[13].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[14].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[14].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[14].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[14].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[14].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[14].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[14].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[14].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[15].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[15].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[15].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[15].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[15].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[15].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[15].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[15].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[1].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[1].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[1].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[1].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[1].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[1].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[1].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[1].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[2].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[2].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[2].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[2].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[2].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[2].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[2].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[2].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[3].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[3].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[3].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[3].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[3].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[3].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[3].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[3].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[4].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[4].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[4].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[4].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[4].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[4].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[4].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[4].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[5].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[5].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[5].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[5].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[5].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[5].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[5].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[5].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[6].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[6].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[6].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[6].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[6].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[6].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[6].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[6].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[7].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[7].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[7].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[7].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[7].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[7].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[7].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[7].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[8].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[8].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[8].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[8].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[8].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[8].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[8].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[8].inter_wire[7] ;
 wire \genblk1[2].puf_buffer.ro_array_2[9].inter_wire[0] ;
 wire \genblk1[2].puf_buffer.ro_array_2[9].inter_wire[1] ;
 wire \genblk1[2].puf_buffer.ro_array_2[9].inter_wire[2] ;
 wire \genblk1[2].puf_buffer.ro_array_2[9].inter_wire[3] ;
 wire \genblk1[2].puf_buffer.ro_array_2[9].inter_wire[4] ;
 wire \genblk1[2].puf_buffer.ro_array_2[9].inter_wire[5] ;
 wire \genblk1[2].puf_buffer.ro_array_2[9].inter_wire[6] ;
 wire \genblk1[2].puf_buffer.ro_array_2[9].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[0] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[10] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[11] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[12] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[13] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[14] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[15] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[1] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[2] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[3] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[4] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[5] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[6] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[7] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[8] ;
 wire \genblk1[3].puf_buffer.cnt_1.ctr[9] ;
 wire \genblk1[3].puf_buffer.cnt_1.finish ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[0] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[10] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[11] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[12] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[13] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[14] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[15] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[1] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[2] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[3] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[4] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[5] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[6] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[7] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[8] ;
 wire \genblk1[3].puf_buffer.cnt_2.ctr[9] ;
 wire \genblk1[3].puf_buffer.cnt_2.finish ;
 wire \genblk1[3].puf_buffer.race_arb.marked_1 ;
 wire \genblk1[3].puf_buffer.race_arb.marked_2 ;
 wire \genblk1[3].puf_buffer.race_arb.resp ;
 wire \genblk1[3].puf_buffer.race_arb.win_1 ;
 wire \genblk1[3].puf_buffer.ro_array_1[0].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[0].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[0].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[0].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[0].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[0].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[0].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[0].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[10].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[10].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[10].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[10].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[10].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[10].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[10].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[10].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[11].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[11].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[11].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[11].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[11].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[11].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[11].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[11].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[12].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[12].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[12].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[12].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[12].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[12].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[12].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[12].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[13].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[13].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[13].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[13].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[13].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[13].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[13].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[13].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[14].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[14].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[14].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[14].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[14].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[14].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[14].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[14].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[15].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[15].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[15].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[15].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[15].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[15].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[15].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[15].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[1].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[1].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[1].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[1].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[1].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[1].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[1].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[1].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[2].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[2].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[2].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[2].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[2].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[2].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[2].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[2].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[3].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[3].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[3].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[3].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[3].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[3].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[3].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[3].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[4].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[4].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[4].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[4].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[4].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[4].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[4].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[4].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[5].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[5].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[5].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[5].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[5].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[5].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[5].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[5].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[6].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[6].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[6].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[6].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[6].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[6].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[6].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[6].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[7].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[7].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[7].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[7].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[7].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[7].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[7].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[7].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[8].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[8].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[8].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[8].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[8].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[8].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[8].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[8].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_1[9].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_1[9].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_1[9].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_1[9].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_1[9].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_1[9].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_1[9].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_1[9].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[0].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[0].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[0].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[0].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[0].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[0].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[0].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[0].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[10].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[10].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[10].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[10].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[10].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[10].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[10].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[10].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[11].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[11].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[11].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[11].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[11].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[11].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[11].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[11].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[12].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[12].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[12].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[12].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[12].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[12].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[12].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[12].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[13].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[13].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[13].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[13].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[13].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[13].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[13].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[13].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[14].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[14].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[14].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[14].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[14].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[14].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[14].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[14].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[15].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[15].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[15].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[15].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[15].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[15].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[15].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[15].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[1].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[1].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[1].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[1].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[1].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[1].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[1].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[1].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[2].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[2].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[2].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[2].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[2].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[2].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[2].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[2].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[3].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[3].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[3].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[3].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[3].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[3].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[3].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[3].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[4].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[4].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[4].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[4].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[4].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[4].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[4].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[4].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[5].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[5].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[5].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[5].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[5].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[5].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[5].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[5].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[6].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[6].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[6].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[6].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[6].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[6].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[6].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[6].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[7].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[7].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[7].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[7].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[7].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[7].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[7].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[7].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[8].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[8].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[8].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[8].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[8].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[8].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[8].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[8].inter_wire[7] ;
 wire \genblk1[3].puf_buffer.ro_array_2[9].inter_wire[0] ;
 wire \genblk1[3].puf_buffer.ro_array_2[9].inter_wire[1] ;
 wire \genblk1[3].puf_buffer.ro_array_2[9].inter_wire[2] ;
 wire \genblk1[3].puf_buffer.ro_array_2[9].inter_wire[3] ;
 wire \genblk1[3].puf_buffer.ro_array_2[9].inter_wire[4] ;
 wire \genblk1[3].puf_buffer.ro_array_2[9].inter_wire[5] ;
 wire \genblk1[3].puf_buffer.ro_array_2[9].inter_wire[6] ;
 wire \genblk1[3].puf_buffer.ro_array_2[9].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[0] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[10] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[11] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[12] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[13] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[14] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[15] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[1] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[2] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[3] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[4] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[5] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[6] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[7] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[8] ;
 wire \genblk1[4].puf_buffer.cnt_1.ctr[9] ;
 wire \genblk1[4].puf_buffer.cnt_1.finish ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[0] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[10] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[11] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[12] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[13] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[14] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[15] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[1] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[2] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[3] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[4] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[5] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[6] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[7] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[8] ;
 wire \genblk1[4].puf_buffer.cnt_2.ctr[9] ;
 wire \genblk1[4].puf_buffer.cnt_2.finish ;
 wire \genblk1[4].puf_buffer.race_arb.marked_1 ;
 wire \genblk1[4].puf_buffer.race_arb.marked_2 ;
 wire \genblk1[4].puf_buffer.race_arb.resp ;
 wire \genblk1[4].puf_buffer.race_arb.win_1 ;
 wire \genblk1[4].puf_buffer.ro_array_1[0].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[0].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[0].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[0].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[0].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[0].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[0].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[0].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[10].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[10].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[10].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[10].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[10].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[10].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[10].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[10].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[11].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[11].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[11].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[11].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[11].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[11].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[11].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[11].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[12].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[12].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[12].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[12].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[12].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[12].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[12].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[12].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[13].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[13].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[13].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[13].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[13].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[13].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[13].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[13].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[14].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[14].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[14].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[14].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[14].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[14].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[14].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[14].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[15].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[15].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[15].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[15].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[15].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[15].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[15].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[15].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[1].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[1].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[1].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[1].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[1].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[1].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[1].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[1].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[2].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[2].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[2].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[2].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[2].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[2].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[2].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[2].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[3].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[3].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[3].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[3].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[3].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[3].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[3].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[3].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[4].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[4].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[4].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[4].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[4].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[4].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[4].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[4].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[5].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[5].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[5].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[5].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[5].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[5].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[5].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[5].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[6].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[6].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[6].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[6].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[6].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[6].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[6].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[6].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[7].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[7].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[7].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[7].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[7].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[7].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[7].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[7].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[8].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[8].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[8].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[8].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[8].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[8].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[8].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[8].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_1[9].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_1[9].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_1[9].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_1[9].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_1[9].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_1[9].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_1[9].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_1[9].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[0].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[0].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[0].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[0].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[0].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[0].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[0].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[0].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[10].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[10].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[10].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[10].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[10].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[10].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[10].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[10].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[11].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[11].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[11].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[11].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[11].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[11].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[11].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[11].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[12].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[12].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[12].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[12].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[12].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[12].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[12].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[12].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[13].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[13].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[13].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[13].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[13].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[13].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[13].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[13].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[14].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[14].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[14].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[14].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[14].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[14].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[14].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[14].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[15].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[15].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[15].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[15].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[15].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[15].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[15].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[15].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[1].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[1].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[1].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[1].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[1].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[1].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[1].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[1].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[2].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[2].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[2].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[2].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[2].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[2].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[2].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[2].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[3].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[3].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[3].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[3].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[3].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[3].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[3].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[3].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[4].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[4].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[4].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[4].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[4].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[4].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[4].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[4].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[5].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[5].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[5].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[5].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[5].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[5].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[5].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[5].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[6].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[6].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[6].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[6].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[6].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[6].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[6].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[6].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[7].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[7].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[7].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[7].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[7].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[7].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[7].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[7].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[8].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[8].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[8].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[8].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[8].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[8].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[8].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[8].inter_wire[7] ;
 wire \genblk1[4].puf_buffer.ro_array_2[9].inter_wire[0] ;
 wire \genblk1[4].puf_buffer.ro_array_2[9].inter_wire[1] ;
 wire \genblk1[4].puf_buffer.ro_array_2[9].inter_wire[2] ;
 wire \genblk1[4].puf_buffer.ro_array_2[9].inter_wire[3] ;
 wire \genblk1[4].puf_buffer.ro_array_2[9].inter_wire[4] ;
 wire \genblk1[4].puf_buffer.ro_array_2[9].inter_wire[5] ;
 wire \genblk1[4].puf_buffer.ro_array_2[9].inter_wire[6] ;
 wire \genblk1[4].puf_buffer.ro_array_2[9].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[0] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[10] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[11] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[12] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[13] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[14] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[15] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[1] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[2] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[3] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[4] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[5] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[6] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[7] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[8] ;
 wire \genblk1[5].puf_buffer.cnt_1.ctr[9] ;
 wire \genblk1[5].puf_buffer.cnt_1.finish ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[0] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[10] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[11] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[12] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[13] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[14] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[15] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[1] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[2] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[3] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[4] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[5] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[6] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[7] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[8] ;
 wire \genblk1[5].puf_buffer.cnt_2.ctr[9] ;
 wire \genblk1[5].puf_buffer.cnt_2.finish ;
 wire \genblk1[5].puf_buffer.race_arb.marked_1 ;
 wire \genblk1[5].puf_buffer.race_arb.marked_2 ;
 wire \genblk1[5].puf_buffer.race_arb.resp ;
 wire \genblk1[5].puf_buffer.race_arb.win_1 ;
 wire \genblk1[5].puf_buffer.ro_array_1[0].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[0].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[0].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[0].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[0].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[0].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[0].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[0].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[10].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[10].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[10].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[10].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[10].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[10].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[10].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[10].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[11].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[11].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[11].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[11].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[11].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[11].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[11].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[11].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[12].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[12].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[12].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[12].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[12].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[12].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[12].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[12].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[13].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[13].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[13].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[13].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[13].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[13].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[13].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[13].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[14].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[14].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[14].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[14].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[14].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[14].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[14].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[14].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[15].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[15].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[15].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[15].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[15].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[15].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[15].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[15].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[1].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[1].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[1].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[1].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[1].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[1].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[1].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[1].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[2].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[2].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[2].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[2].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[2].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[2].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[2].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[2].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[3].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[3].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[3].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[3].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[3].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[3].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[3].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[3].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[4].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[4].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[4].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[4].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[4].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[4].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[4].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[4].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[5].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[5].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[5].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[5].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[5].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[5].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[5].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[5].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[6].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[6].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[6].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[6].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[6].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[6].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[6].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[6].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[7].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[7].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[7].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[7].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[7].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[7].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[7].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[7].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[8].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[8].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[8].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[8].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[8].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[8].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[8].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[8].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_1[9].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_1[9].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_1[9].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_1[9].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_1[9].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_1[9].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_1[9].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_1[9].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[0].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[0].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[0].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[0].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[0].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[0].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[0].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[0].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[10].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[10].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[10].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[10].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[10].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[10].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[10].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[10].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[11].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[11].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[11].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[11].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[11].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[11].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[11].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[11].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[12].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[12].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[12].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[12].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[12].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[12].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[12].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[12].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[13].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[13].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[13].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[13].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[13].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[13].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[13].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[13].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[14].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[14].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[14].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[14].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[14].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[14].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[14].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[14].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[15].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[15].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[15].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[15].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[15].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[15].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[15].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[15].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[1].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[1].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[1].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[1].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[1].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[1].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[1].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[1].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[2].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[2].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[2].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[2].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[2].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[2].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[2].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[2].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[3].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[3].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[3].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[3].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[3].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[3].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[3].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[3].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[4].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[4].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[4].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[4].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[4].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[4].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[4].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[4].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[5].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[5].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[5].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[5].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[5].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[5].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[5].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[5].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[6].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[6].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[6].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[6].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[6].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[6].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[6].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[6].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[7].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[7].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[7].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[7].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[7].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[7].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[7].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[7].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[8].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[8].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[8].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[8].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[8].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[8].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[8].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[8].inter_wire[7] ;
 wire \genblk1[5].puf_buffer.ro_array_2[9].inter_wire[0] ;
 wire \genblk1[5].puf_buffer.ro_array_2[9].inter_wire[1] ;
 wire \genblk1[5].puf_buffer.ro_array_2[9].inter_wire[2] ;
 wire \genblk1[5].puf_buffer.ro_array_2[9].inter_wire[3] ;
 wire \genblk1[5].puf_buffer.ro_array_2[9].inter_wire[4] ;
 wire \genblk1[5].puf_buffer.ro_array_2[9].inter_wire[5] ;
 wire \genblk1[5].puf_buffer.ro_array_2[9].inter_wire[6] ;
 wire \genblk1[5].puf_buffer.ro_array_2[9].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[0] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[10] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[11] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[12] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[13] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[14] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[15] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[1] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[2] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[3] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[4] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[5] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[6] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[7] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[8] ;
 wire \genblk1[6].puf_buffer.cnt_1.ctr[9] ;
 wire \genblk1[6].puf_buffer.cnt_1.finish ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[0] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[10] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[11] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[12] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[13] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[14] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[15] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[1] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[2] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[3] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[4] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[5] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[6] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[7] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[8] ;
 wire \genblk1[6].puf_buffer.cnt_2.ctr[9] ;
 wire \genblk1[6].puf_buffer.cnt_2.finish ;
 wire \genblk1[6].puf_buffer.race_arb.marked_1 ;
 wire \genblk1[6].puf_buffer.race_arb.marked_2 ;
 wire \genblk1[6].puf_buffer.race_arb.resp ;
 wire \genblk1[6].puf_buffer.race_arb.win_1 ;
 wire \genblk1[6].puf_buffer.ro_array_1[0].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[0].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[0].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[0].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[0].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[0].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[0].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[0].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[10].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[10].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[10].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[10].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[10].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[10].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[10].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[10].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[11].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[11].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[11].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[11].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[11].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[11].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[11].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[11].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[12].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[12].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[12].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[12].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[12].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[12].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[12].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[12].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[13].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[13].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[13].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[13].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[13].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[13].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[13].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[13].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[14].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[14].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[14].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[14].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[14].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[14].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[14].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[14].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[15].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[15].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[15].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[15].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[15].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[15].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[15].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[15].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[1].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[1].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[1].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[1].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[1].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[1].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[1].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[1].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[2].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[2].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[2].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[2].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[2].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[2].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[2].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[2].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[3].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[3].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[3].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[3].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[3].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[3].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[3].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[3].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[4].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[4].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[4].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[4].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[4].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[4].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[4].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[4].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[5].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[5].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[5].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[5].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[5].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[5].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[5].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[5].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[6].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[6].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[6].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[6].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[6].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[6].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[6].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[6].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[7].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[7].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[7].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[7].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[7].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[7].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[7].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[7].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[8].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[8].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[8].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[8].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[8].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[8].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[8].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[8].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_1[9].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_1[9].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_1[9].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_1[9].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_1[9].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_1[9].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_1[9].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_1[9].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[0].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[0].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[0].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[0].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[0].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[0].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[0].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[0].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[10].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[10].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[10].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[10].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[10].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[10].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[10].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[10].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[11].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[11].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[11].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[11].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[11].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[11].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[11].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[11].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[12].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[12].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[12].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[12].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[12].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[12].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[12].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[12].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[13].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[13].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[13].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[13].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[13].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[13].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[13].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[13].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[14].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[14].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[14].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[14].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[14].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[14].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[14].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[14].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[15].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[15].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[15].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[15].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[15].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[15].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[15].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[15].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[1].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[1].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[1].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[1].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[1].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[1].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[1].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[1].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[2].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[2].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[2].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[2].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[2].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[2].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[2].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[2].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[3].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[3].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[3].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[3].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[3].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[3].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[3].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[3].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[4].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[4].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[4].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[4].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[4].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[4].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[4].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[4].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[5].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[5].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[5].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[5].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[5].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[5].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[5].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[5].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[6].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[6].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[6].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[6].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[6].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[6].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[6].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[6].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[7].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[7].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[7].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[7].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[7].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[7].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[7].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[7].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[8].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[8].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[8].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[8].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[8].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[8].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[8].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[8].inter_wire[7] ;
 wire \genblk1[6].puf_buffer.ro_array_2[9].inter_wire[0] ;
 wire \genblk1[6].puf_buffer.ro_array_2[9].inter_wire[1] ;
 wire \genblk1[6].puf_buffer.ro_array_2[9].inter_wire[2] ;
 wire \genblk1[6].puf_buffer.ro_array_2[9].inter_wire[3] ;
 wire \genblk1[6].puf_buffer.ro_array_2[9].inter_wire[4] ;
 wire \genblk1[6].puf_buffer.ro_array_2[9].inter_wire[5] ;
 wire \genblk1[6].puf_buffer.ro_array_2[9].inter_wire[6] ;
 wire \genblk1[6].puf_buffer.ro_array_2[9].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[0] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[10] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[11] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[12] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[13] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[14] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[15] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[1] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[2] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[3] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[4] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[5] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[6] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[7] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[8] ;
 wire \genblk1[7].puf_buffer.cnt_1.ctr[9] ;
 wire \genblk1[7].puf_buffer.cnt_1.finish ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[0] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[10] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[11] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[12] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[13] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[14] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[15] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[1] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[2] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[3] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[4] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[5] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[6] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[7] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[8] ;
 wire \genblk1[7].puf_buffer.cnt_2.ctr[9] ;
 wire \genblk1[7].puf_buffer.cnt_2.finish ;
 wire \genblk1[7].puf_buffer.race_arb.marked_1 ;
 wire \genblk1[7].puf_buffer.race_arb.marked_2 ;
 wire \genblk1[7].puf_buffer.race_arb.resp ;
 wire \genblk1[7].puf_buffer.race_arb.win_1 ;
 wire \genblk1[7].puf_buffer.ro_array_1[0].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[0].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[0].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[0].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[0].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[0].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[0].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[0].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[10].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[10].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[10].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[10].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[10].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[10].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[10].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[10].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[11].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[11].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[11].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[11].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[11].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[11].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[11].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[11].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[12].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[12].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[12].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[12].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[12].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[12].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[12].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[12].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[13].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[13].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[13].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[13].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[13].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[13].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[13].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[13].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[14].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[14].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[14].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[14].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[14].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[14].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[14].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[14].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[15].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[15].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[15].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[15].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[15].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[15].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[15].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[15].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[1].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[1].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[1].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[1].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[1].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[1].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[1].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[1].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[2].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[2].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[2].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[2].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[2].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[2].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[2].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[2].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[3].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[3].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[3].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[3].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[3].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[3].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[3].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[3].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[4].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[4].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[4].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[4].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[4].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[4].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[4].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[4].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[5].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[5].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[5].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[5].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[5].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[5].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[5].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[5].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[6].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[6].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[6].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[6].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[6].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[6].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[6].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[6].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[7].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[7].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[7].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[7].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[7].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[7].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[7].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[7].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[8].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[8].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[8].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[8].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[8].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[8].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[8].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[8].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_1[9].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_1[9].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_1[9].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_1[9].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_1[9].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_1[9].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_1[9].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_1[9].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[0].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[0].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[0].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[0].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[0].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[0].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[0].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[0].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[10].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[10].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[10].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[10].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[10].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[10].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[10].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[10].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[11].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[11].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[11].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[11].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[11].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[11].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[11].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[11].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[12].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[12].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[12].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[12].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[12].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[12].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[12].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[12].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[13].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[13].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[13].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[13].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[13].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[13].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[13].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[13].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[14].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[14].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[14].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[14].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[14].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[14].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[14].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[14].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[15].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[15].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[15].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[15].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[15].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[15].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[15].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[15].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[1].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[1].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[1].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[1].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[1].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[1].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[1].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[1].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[2].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[2].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[2].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[2].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[2].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[2].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[2].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[2].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[3].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[3].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[3].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[3].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[3].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[3].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[3].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[3].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[4].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[4].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[4].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[4].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[4].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[4].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[4].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[4].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[5].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[5].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[5].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[5].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[5].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[5].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[5].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[5].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[6].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[6].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[6].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[6].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[6].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[6].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[6].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[6].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[7].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[7].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[7].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[7].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[7].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[7].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[7].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[7].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[8].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[8].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[8].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[8].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[8].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[8].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[8].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[8].inter_wire[7] ;
 wire \genblk1[7].puf_buffer.ro_array_2[9].inter_wire[0] ;
 wire \genblk1[7].puf_buffer.ro_array_2[9].inter_wire[1] ;
 wire \genblk1[7].puf_buffer.ro_array_2[9].inter_wire[2] ;
 wire \genblk1[7].puf_buffer.ro_array_2[9].inter_wire[3] ;
 wire \genblk1[7].puf_buffer.ro_array_2[9].inter_wire[4] ;
 wire \genblk1[7].puf_buffer.ro_array_2[9].inter_wire[5] ;
 wire \genblk1[7].puf_buffer.ro_array_2[9].inter_wire[6] ;
 wire \genblk1[7].puf_buffer.ro_array_2[9].inter_wire[7] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net24;
 wire net25;
 wire net26;
 wire net3;
 wire net4;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__decap_4 FILLER_0_0_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_240 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_10 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_183 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_252 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_222 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_175 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_158 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_170 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_245 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_248 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_213 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_173 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_158 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_170 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_204 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_206 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_48_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_48 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_60 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_143 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_288 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_184 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_126 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_138 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_60_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_175 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_74_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_76_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_76_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_78_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_78_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_78_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_78_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_78_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_79_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_79_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_79_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_79_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_79_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_285 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_80_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_80_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_80_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_80_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_80_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__and3b_1 _1618_ (.A_N(_1227_),
    .B(_1164_),
    .C(_1228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _1619_ (.A(_1229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0166_));
 sky130_fd_sc_hd__and3_1 _1620_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[5].puf_buffer.cnt_1.ctr[4] ),
    .C(_1196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1230_));
 sky130_fd_sc_hd__inv_2 _1621_ (.A(_1230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1231_));
 sky130_fd_sc_hd__o221a_1 _1622_ (.A1(_1231_),
    .A2(_1220_),
    .B1(_1227_),
    .B2(net174),
    .C1(_1221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0167_));
 sky130_fd_sc_hd__and4_1 _1623_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[6] ),
    .B(_1230_),
    .C(_1203_),
    .D(_1213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1232_));
 sky130_fd_sc_hd__a31o_1 _1624_ (.A1(_1230_),
    .A2(_1215_),
    .A3(_1216_),
    .B1(\genblk1[5].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1233_));
 sky130_fd_sc_hd__and3b_1 _1625_ (.A_N(_1232_),
    .B(_1164_),
    .C(_1233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _1626_ (.A(_1234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0168_));
 sky130_fd_sc_hd__inv_2 _1627_ (.A(_1198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1235_));
 sky130_fd_sc_hd__o221a_1 _1628_ (.A1(_1235_),
    .A2(_1220_),
    .B1(_1232_),
    .B2(net160),
    .C1(_1221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0169_));
 sky130_fd_sc_hd__and4_1 _1629_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[8] ),
    .B(_1198_),
    .C(_1203_),
    .D(_1213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1236_));
 sky130_fd_sc_hd__clkbuf_2 _1630_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1237_));
 sky130_fd_sc_hd__a31o_1 _1631_ (.A1(_1198_),
    .A2(_1215_),
    .A3(_1216_),
    .B1(\genblk1[5].puf_buffer.cnt_1.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1238_));
 sky130_fd_sc_hd__and3b_1 _1632_ (.A_N(_1236_),
    .B(_1237_),
    .C(_1238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1239_));
 sky130_fd_sc_hd__clkbuf_1 _1633_ (.A(_1239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0170_));
 sky130_fd_sc_hd__nand3_1 _1634_ (.A(_1199_),
    .B(_1215_),
    .C(_1216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1240_));
 sky130_fd_sc_hd__o211a_1 _1635_ (.A1(net152),
    .A2(_1236_),
    .B1(_1240_),
    .C1(_1007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0171_));
 sky130_fd_sc_hd__and4_1 _1636_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[10] ),
    .B(_1199_),
    .C(_1203_),
    .D(_1213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1241_));
 sky130_fd_sc_hd__a31o_1 _1637_ (.A1(_1199_),
    .A2(_1215_),
    .A3(_1216_),
    .B1(\genblk1[5].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1242_));
 sky130_fd_sc_hd__and3b_1 _1638_ (.A_N(_1241_),
    .B(_1237_),
    .C(_1242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1243_));
 sky130_fd_sc_hd__clkbuf_1 _1639_ (.A(_1243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0172_));
 sky130_fd_sc_hd__nand2_1 _1640_ (.A(net189),
    .B(\genblk1[5].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1244_));
 sky130_fd_sc_hd__o221a_1 _1641_ (.A1(_1244_),
    .A2(_1240_),
    .B1(_1241_),
    .B2(net189),
    .C1(_1221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0173_));
 sky130_fd_sc_hd__inv_2 _1642_ (.A(_1200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1245_));
 sky130_fd_sc_hd__and2_1 _1643_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[11] ),
    .B(\genblk1[5].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1246_));
 sky130_fd_sc_hd__a41o_1 _1644_ (.A1(_1199_),
    .A2(_1246_),
    .A3(_1215_),
    .A4(_1216_),
    .B1(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1247_));
 sky130_fd_sc_hd__o211a_1 _1645_ (.A1(_1245_),
    .A2(_1240_),
    .B1(_1247_),
    .C1(_1007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0174_));
 sky130_fd_sc_hd__and4_1 _1646_ (.A(_1199_),
    .B(_1201_),
    .C(_1203_),
    .D(_1213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1248_));
 sky130_fd_sc_hd__a41o_1 _1647_ (.A1(_1199_),
    .A2(_1200_),
    .A3(_1203_),
    .A4(_1213_),
    .B1(\genblk1[5].puf_buffer.cnt_1.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1249_));
 sky130_fd_sc_hd__and3b_1 _1648_ (.A_N(_1248_),
    .B(_1237_),
    .C(_1249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1250_));
 sky130_fd_sc_hd__clkbuf_1 _1649_ (.A(_1250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0175_));
 sky130_fd_sc_hd__inv_2 _1650_ (.A(_1202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1251_));
 sky130_fd_sc_hd__o221a_1 _1651_ (.A1(_1251_),
    .A2(_1220_),
    .B1(_1248_),
    .B2(net103),
    .C1(_1221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0176_));
 sky130_fd_sc_hd__nand4_1 _1652_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[15] ),
    .B(_1202_),
    .C(_1215_),
    .D(_1216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1252_));
 sky130_fd_sc_hd__a31o_1 _1653_ (.A1(_1202_),
    .A2(_1215_),
    .A3(_1216_),
    .B1(\genblk1[5].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1253_));
 sky130_fd_sc_hd__and3_1 _1654_ (.A(_1129_),
    .B(_1252_),
    .C(_1253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1254_));
 sky130_fd_sc_hd__clkbuf_1 _1655_ (.A(_1254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0177_));
 sky130_fd_sc_hd__inv_2 _1656_ (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1255_));
 sky130_fd_sc_hd__and3b_1 _1657_ (.A_N(\genblk1[6].puf_buffer.cnt_1.finish ),
    .B(\genblk1[6].puf_buffer.cnt_2.finish ),
    .C(_0475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_1 _1658_ (.A(_1256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0215_));
 sky130_fd_sc_hd__o21bai_1 _1659_ (.A1(_1255_),
    .A2(_0215_),
    .B1_N(\genblk1[6].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0178_));
 sky130_fd_sc_hd__and4_1 _1660_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[3] ),
    .B(\genblk1[6].puf_buffer.cnt_2.ctr[2] ),
    .C(\genblk1[6].puf_buffer.cnt_2.ctr[1] ),
    .D(\genblk1[6].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1257_));
 sky130_fd_sc_hd__and2_1 _1661_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[6].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1258_));
 sky130_fd_sc_hd__and4_1 _1662_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[6].puf_buffer.cnt_2.ctr[4] ),
    .C(_1257_),
    .D(_1258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1259_));
 sky130_fd_sc_hd__and3_1 _1663_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[9] ),
    .B(\genblk1[6].puf_buffer.cnt_2.ctr[8] ),
    .C(_1259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1260_));
 sky130_fd_sc_hd__and3_1 _1664_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[12] ),
    .B(\genblk1[6].puf_buffer.cnt_2.ctr[11] ),
    .C(\genblk1[6].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1261_));
 sky130_fd_sc_hd__and2_1 _1665_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[13] ),
    .B(_1261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1262_));
 sky130_fd_sc_hd__and3_1 _1666_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[14] ),
    .B(_1260_),
    .C(_1262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1263_));
 sky130_fd_sc_hd__a22o_1 _1667_ (.A1(_0670_),
    .A2(\genblk1[6].puf_buffer.cnt_2.finish ),
    .B1(_1263_),
    .B2(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0180_));
 sky130_fd_sc_hd__or2_2 _1668_ (.A(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1264_));
 sky130_fd_sc_hd__a22o_1 _1669_ (.A1(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .A2(_0621_),
    .B1(_0603_),
    .B2(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1265_));
 sky130_fd_sc_hd__a221o_1 _1670_ (.A1(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .A2(_0605_),
    .B1(_0625_),
    .B2(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .C1(_1265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1266_));
 sky130_fd_sc_hd__a22o_1 _1671_ (.A1(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .A2(_0611_),
    .B1(_0618_),
    .B2(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1267_));
 sky130_fd_sc_hd__a211o_1 _1672_ (.A1(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .A2(_0615_),
    .B1(_1267_),
    .C1(_0613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1268_));
 sky130_fd_sc_hd__a22o_1 _1673_ (.A1(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .A2(_0606_),
    .B1(_0619_),
    .B2(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1269_));
 sky130_fd_sc_hd__a22o_1 _1674_ (.A1(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .A2(net232),
    .B1(_0604_),
    .B2(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1270_));
 sky130_fd_sc_hd__a22o_1 _1675_ (.A1(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .A2(_0610_),
    .B1(_0616_),
    .B2(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1271_));
 sky130_fd_sc_hd__a22o_1 _1676_ (.A1(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .A2(_0624_),
    .B1(_0622_),
    .B2(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1272_));
 sky130_fd_sc_hd__or4_1 _1677_ (.A(_1269_),
    .B(_1270_),
    .C(_1271_),
    .D(_1272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1273_));
 sky130_fd_sc_hd__or3_4 _1678_ (.A(_1266_),
    .B(_1268_),
    .C(_1273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1274_));
 sky130_fd_sc_hd__and3_1 _1679_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[0] ),
    .B(_1264_),
    .C(_1274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1275_));
 sky130_fd_sc_hd__buf_2 _1680_ (.A(_1264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1276_));
 sky130_fd_sc_hd__buf_2 _1681_ (.A(_1274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1277_));
 sky130_fd_sc_hd__a21o_1 _1682_ (.A1(_1276_),
    .A2(_1277_),
    .B1(\genblk1[6].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1278_));
 sky130_fd_sc_hd__and3b_1 _1683_ (.A_N(_1275_),
    .B(_1237_),
    .C(_1278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1279_));
 sky130_fd_sc_hd__clkbuf_1 _1684_ (.A(_1279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_1 _1685_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[1] ),
    .B(\genblk1[6].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1280_));
 sky130_fd_sc_hd__nand2_2 _1686_ (.A(_1276_),
    .B(_1277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1281_));
 sky130_fd_sc_hd__o221a_1 _1687_ (.A1(_1280_),
    .A2(_1281_),
    .B1(_1275_),
    .B2(net218),
    .C1(_1221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0182_));
 sky130_fd_sc_hd__inv_2 _1688_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1282_));
 sky130_fd_sc_hd__and4bb_1 _1689_ (.A_N(_1282_),
    .B_N(_1280_),
    .C(_1264_),
    .D(_1274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1283_));
 sky130_fd_sc_hd__a41o_1 _1690_ (.A1(\genblk1[6].puf_buffer.cnt_2.ctr[1] ),
    .A2(\genblk1[6].puf_buffer.cnt_2.ctr[0] ),
    .A3(_1264_),
    .A4(_1274_),
    .B1(\genblk1[6].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1284_));
 sky130_fd_sc_hd__and3b_1 _1691_ (.A_N(_1283_),
    .B(_1237_),
    .C(_1284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1285_));
 sky130_fd_sc_hd__clkbuf_1 _1692_ (.A(_1285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0183_));
 sky130_fd_sc_hd__inv_2 _1693_ (.A(_1257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1286_));
 sky130_fd_sc_hd__o221a_1 _1694_ (.A1(_1286_),
    .A2(_1281_),
    .B1(_1283_),
    .B2(net100),
    .C1(_1221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0184_));
 sky130_fd_sc_hd__and4_1 _1695_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[4] ),
    .B(_1257_),
    .C(_1264_),
    .D(_1274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1287_));
 sky130_fd_sc_hd__a31o_1 _1696_ (.A1(_1257_),
    .A2(_1276_),
    .A3(_1277_),
    .B1(\genblk1[6].puf_buffer.cnt_2.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1288_));
 sky130_fd_sc_hd__and3b_1 _1697_ (.A_N(_1287_),
    .B(_1237_),
    .C(_1288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _1698_ (.A(_1289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0185_));
 sky130_fd_sc_hd__and3_1 _1699_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[6].puf_buffer.cnt_2.ctr[4] ),
    .C(_1257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1290_));
 sky130_fd_sc_hd__inv_2 _1700_ (.A(_1290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1291_));
 sky130_fd_sc_hd__o221a_1 _1701_ (.A1(_1291_),
    .A2(_1281_),
    .B1(_1287_),
    .B2(net176),
    .C1(_1221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0186_));
 sky130_fd_sc_hd__and4_1 _1702_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[6] ),
    .B(_1290_),
    .C(_1264_),
    .D(_1274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1292_));
 sky130_fd_sc_hd__a31o_1 _1703_ (.A1(_1290_),
    .A2(_1276_),
    .A3(_1277_),
    .B1(\genblk1[6].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1293_));
 sky130_fd_sc_hd__and3b_1 _1704_ (.A_N(_1292_),
    .B(_1237_),
    .C(_1293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _1705_ (.A(_1294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0187_));
 sky130_fd_sc_hd__inv_2 _1706_ (.A(_1259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1295_));
 sky130_fd_sc_hd__o221a_1 _1707_ (.A1(_1295_),
    .A2(_1281_),
    .B1(_1292_),
    .B2(net118),
    .C1(_1221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0188_));
 sky130_fd_sc_hd__and4_1 _1708_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[8] ),
    .B(_1259_),
    .C(_1264_),
    .D(_1274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1296_));
 sky130_fd_sc_hd__a31o_1 _1709_ (.A1(_1259_),
    .A2(_1276_),
    .A3(_1277_),
    .B1(\genblk1[6].puf_buffer.cnt_2.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1297_));
 sky130_fd_sc_hd__and3b_1 _1710_ (.A_N(_1296_),
    .B(_1237_),
    .C(_1297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_1 _1711_ (.A(_1298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0189_));
 sky130_fd_sc_hd__nand3_1 _1712_ (.A(_1260_),
    .B(_1276_),
    .C(_1277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1299_));
 sky130_fd_sc_hd__o211a_1 _1713_ (.A1(net155),
    .A2(_1296_),
    .B1(_1299_),
    .C1(_1007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0190_));
 sky130_fd_sc_hd__and4_1 _1714_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[10] ),
    .B(_1260_),
    .C(_1264_),
    .D(_1274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1300_));
 sky130_fd_sc_hd__a31o_1 _1715_ (.A1(_1260_),
    .A2(_1276_),
    .A3(_1277_),
    .B1(\genblk1[6].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1301_));
 sky130_fd_sc_hd__and3b_1 _1716_ (.A_N(_1300_),
    .B(_1237_),
    .C(_1301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _1717_ (.A(_1302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0191_));
 sky130_fd_sc_hd__nand2_1 _1718_ (.A(net199),
    .B(\genblk1[6].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1303_));
 sky130_fd_sc_hd__clkbuf_4 _1719_ (.A(_0638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1304_));
 sky130_fd_sc_hd__o221a_1 _1720_ (.A1(_1303_),
    .A2(_1299_),
    .B1(_1300_),
    .B2(net199),
    .C1(_1304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0192_));
 sky130_fd_sc_hd__inv_2 _1721_ (.A(_1261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1305_));
 sky130_fd_sc_hd__and2_1 _1722_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[11] ),
    .B(\genblk1[6].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1306_));
 sky130_fd_sc_hd__a41o_1 _1723_ (.A1(_1260_),
    .A2(_1306_),
    .A3(_1276_),
    .A4(_1277_),
    .B1(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_4 _1724_ (.A(_0631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1308_));
 sky130_fd_sc_hd__o211a_1 _1725_ (.A1(_1305_),
    .A2(_1299_),
    .B1(_1307_),
    .C1(_1308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0193_));
 sky130_fd_sc_hd__and4_1 _1726_ (.A(_1260_),
    .B(_1262_),
    .C(_1264_),
    .D(_1274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1309_));
 sky130_fd_sc_hd__a41o_1 _1727_ (.A1(_1260_),
    .A2(_1261_),
    .A3(_1264_),
    .A4(_1274_),
    .B1(\genblk1[6].puf_buffer.cnt_2.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1310_));
 sky130_fd_sc_hd__and3b_1 _1728_ (.A_N(_1309_),
    .B(_1237_),
    .C(_1310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1311_));
 sky130_fd_sc_hd__clkbuf_1 _1729_ (.A(_1311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0194_));
 sky130_fd_sc_hd__inv_2 _1730_ (.A(_1263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1312_));
 sky130_fd_sc_hd__o221a_1 _1731_ (.A1(_1312_),
    .A2(_1281_),
    .B1(_1309_),
    .B2(net82),
    .C1(_1304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0195_));
 sky130_fd_sc_hd__nand4_1 _1732_ (.A(\genblk1[6].puf_buffer.cnt_2.ctr[15] ),
    .B(_1263_),
    .C(_1276_),
    .D(_1277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1313_));
 sky130_fd_sc_hd__a31o_1 _1733_ (.A1(_1263_),
    .A2(_1276_),
    .A3(_1277_),
    .B1(\genblk1[6].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1314_));
 sky130_fd_sc_hd__and3_1 _1734_ (.A(_1129_),
    .B(_1313_),
    .C(_1314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1315_));
 sky130_fd_sc_hd__clkbuf_1 _1735_ (.A(_1315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0196_));
 sky130_fd_sc_hd__and4_1 _1736_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[3] ),
    .B(\genblk1[6].puf_buffer.cnt_1.ctr[2] ),
    .C(\genblk1[6].puf_buffer.cnt_1.ctr[1] ),
    .D(\genblk1[6].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1316_));
 sky130_fd_sc_hd__and2_1 _1737_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[6].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1317_));
 sky130_fd_sc_hd__and4_1 _1738_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[6].puf_buffer.cnt_1.ctr[4] ),
    .C(_1316_),
    .D(_1317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1318_));
 sky130_fd_sc_hd__and3_1 _1739_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[9] ),
    .B(\genblk1[6].puf_buffer.cnt_1.ctr[8] ),
    .C(_1318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1319_));
 sky130_fd_sc_hd__and3_1 _1740_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[12] ),
    .B(\genblk1[6].puf_buffer.cnt_1.ctr[11] ),
    .C(\genblk1[6].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1320_));
 sky130_fd_sc_hd__and2_1 _1741_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[13] ),
    .B(_1320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1321_));
 sky130_fd_sc_hd__and3_1 _1742_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[14] ),
    .B(_1319_),
    .C(_1321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1322_));
 sky130_fd_sc_hd__a22o_1 _1743_ (.A1(_0670_),
    .A2(\genblk1[6].puf_buffer.cnt_1.finish ),
    .B1(_1322_),
    .B2(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0197_));
 sky130_fd_sc_hd__or2_2 _1744_ (.A(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1323_));
 sky130_fd_sc_hd__a22o_1 _1745_ (.A1(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .A2(_0706_),
    .B1(_0709_),
    .B2(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1324_));
 sky130_fd_sc_hd__a22o_1 _1746_ (.A1(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .A2(_0700_),
    .B1(_0702_),
    .B2(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1325_));
 sky130_fd_sc_hd__a211o_1 _1747_ (.A1(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .A2(_0688_),
    .B1(_1324_),
    .C1(_1325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1326_));
 sky130_fd_sc_hd__a22o_1 _1748_ (.A1(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .A2(net24),
    .B1(_0693_),
    .B2(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1327_));
 sky130_fd_sc_hd__a221o_1 _1749_ (.A1(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .A2(_0705_),
    .B1(_0689_),
    .B2(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .C1(_1327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1328_));
 sky130_fd_sc_hd__a22o_1 _1750_ (.A1(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .A2(_0699_),
    .B1(_0695_),
    .B2(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1329_));
 sky130_fd_sc_hd__a221o_1 _1751_ (.A1(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .A2(_0694_),
    .B1(_0687_),
    .B2(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .C1(_0697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1330_));
 sky130_fd_sc_hd__a22o_1 _1752_ (.A1(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .A2(_0690_),
    .B1(net229),
    .B2(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1331_));
 sky130_fd_sc_hd__or3_1 _1753_ (.A(_1329_),
    .B(_1330_),
    .C(_1331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1332_));
 sky130_fd_sc_hd__or3_4 _1754_ (.A(_1326_),
    .B(_1328_),
    .C(_1332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1333_));
 sky130_fd_sc_hd__and3_1 _1755_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[0] ),
    .B(_1323_),
    .C(_1333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1334_));
 sky130_fd_sc_hd__clkbuf_2 _1756_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1335_));
 sky130_fd_sc_hd__buf_2 _1757_ (.A(_1323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1336_));
 sky130_fd_sc_hd__buf_2 _1758_ (.A(_1333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1337_));
 sky130_fd_sc_hd__a21o_1 _1759_ (.A1(_1336_),
    .A2(_1337_),
    .B1(\genblk1[6].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1338_));
 sky130_fd_sc_hd__and3b_1 _1760_ (.A_N(_1334_),
    .B(_1335_),
    .C(_1338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1339_));
 sky130_fd_sc_hd__clkbuf_1 _1761_ (.A(_1339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0198_));
 sky130_fd_sc_hd__nand2_1 _1762_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[1] ),
    .B(\genblk1[6].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1340_));
 sky130_fd_sc_hd__nand2_2 _1763_ (.A(_1336_),
    .B(_1337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1341_));
 sky130_fd_sc_hd__o221a_1 _1764_ (.A1(_1340_),
    .A2(_1341_),
    .B1(_1334_),
    .B2(net210),
    .C1(_1304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0199_));
 sky130_fd_sc_hd__inv_2 _1765_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1342_));
 sky130_fd_sc_hd__and4bb_1 _1766_ (.A_N(_1342_),
    .B_N(_1340_),
    .C(_1323_),
    .D(_1333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1343_));
 sky130_fd_sc_hd__a41o_1 _1767_ (.A1(\genblk1[6].puf_buffer.cnt_1.ctr[1] ),
    .A2(\genblk1[6].puf_buffer.cnt_1.ctr[0] ),
    .A3(_1323_),
    .A4(_1333_),
    .B1(\genblk1[6].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1344_));
 sky130_fd_sc_hd__and3b_1 _1768_ (.A_N(_1343_),
    .B(_1335_),
    .C(_1344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1345_));
 sky130_fd_sc_hd__clkbuf_1 _1769_ (.A(_1345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0200_));
 sky130_fd_sc_hd__inv_2 _1770_ (.A(_1316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1346_));
 sky130_fd_sc_hd__o221a_1 _1771_ (.A1(_1346_),
    .A2(_1341_),
    .B1(_1343_),
    .B2(net92),
    .C1(_1304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0201_));
 sky130_fd_sc_hd__and4_1 _1772_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[4] ),
    .B(_1316_),
    .C(_1323_),
    .D(_1333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1347_));
 sky130_fd_sc_hd__a31o_1 _1773_ (.A1(_1316_),
    .A2(_1336_),
    .A3(_1337_),
    .B1(\genblk1[6].puf_buffer.cnt_1.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1348_));
 sky130_fd_sc_hd__and3b_1 _1774_ (.A_N(_1347_),
    .B(_1335_),
    .C(_1348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1349_));
 sky130_fd_sc_hd__clkbuf_1 _1775_ (.A(_1349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0202_));
 sky130_fd_sc_hd__and3_1 _1776_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[6].puf_buffer.cnt_1.ctr[4] ),
    .C(_1316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1350_));
 sky130_fd_sc_hd__inv_2 _1777_ (.A(_1350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1351_));
 sky130_fd_sc_hd__o221a_1 _1778_ (.A1(_1351_),
    .A2(_1341_),
    .B1(_1347_),
    .B2(net172),
    .C1(_1304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0203_));
 sky130_fd_sc_hd__and4_1 _1779_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[6] ),
    .B(_1350_),
    .C(_1323_),
    .D(_1333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1352_));
 sky130_fd_sc_hd__a31o_1 _1780_ (.A1(_1350_),
    .A2(_1336_),
    .A3(_1337_),
    .B1(\genblk1[6].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1353_));
 sky130_fd_sc_hd__and3b_1 _1781_ (.A_N(_1352_),
    .B(_1335_),
    .C(_1353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1354_));
 sky130_fd_sc_hd__clkbuf_1 _1782_ (.A(_1354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0204_));
 sky130_fd_sc_hd__inv_2 _1783_ (.A(_1318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1355_));
 sky130_fd_sc_hd__o221a_1 _1784_ (.A1(_1355_),
    .A2(_1341_),
    .B1(_1352_),
    .B2(net81),
    .C1(_1304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0205_));
 sky130_fd_sc_hd__and4_1 _1785_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[8] ),
    .B(_1318_),
    .C(_1323_),
    .D(_1333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1356_));
 sky130_fd_sc_hd__a31o_1 _1786_ (.A1(_1318_),
    .A2(_1336_),
    .A3(_1337_),
    .B1(\genblk1[6].puf_buffer.cnt_1.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1357_));
 sky130_fd_sc_hd__and3b_1 _1787_ (.A_N(_1356_),
    .B(_1335_),
    .C(_1357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1358_));
 sky130_fd_sc_hd__clkbuf_1 _1788_ (.A(_1358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0206_));
 sky130_fd_sc_hd__nand3_1 _1789_ (.A(_1319_),
    .B(_1336_),
    .C(_1337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1359_));
 sky130_fd_sc_hd__o211a_1 _1790_ (.A1(net106),
    .A2(_1356_),
    .B1(_1359_),
    .C1(_1308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0207_));
 sky130_fd_sc_hd__and4_1 _1791_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[10] ),
    .B(_1319_),
    .C(_1323_),
    .D(_1333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1360_));
 sky130_fd_sc_hd__a31o_1 _1792_ (.A1(_1319_),
    .A2(_1336_),
    .A3(_1337_),
    .B1(\genblk1[6].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1361_));
 sky130_fd_sc_hd__and3b_1 _1793_ (.A_N(_1360_),
    .B(_1335_),
    .C(_1361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_1 _1794_ (.A(_1362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0208_));
 sky130_fd_sc_hd__nand2_1 _1795_ (.A(net192),
    .B(\genblk1[6].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1363_));
 sky130_fd_sc_hd__o221a_1 _1796_ (.A1(_1363_),
    .A2(_1359_),
    .B1(_1360_),
    .B2(net192),
    .C1(_1304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0209_));
 sky130_fd_sc_hd__inv_2 _1797_ (.A(_1320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1364_));
 sky130_fd_sc_hd__and2_1 _1798_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[11] ),
    .B(\genblk1[6].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1365_));
 sky130_fd_sc_hd__a41o_1 _1799_ (.A1(_1319_),
    .A2(_1365_),
    .A3(_1336_),
    .A4(_1337_),
    .B1(net226),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1366_));
 sky130_fd_sc_hd__o211a_1 _1800_ (.A1(_1364_),
    .A2(_1359_),
    .B1(_1366_),
    .C1(_1308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0210_));
 sky130_fd_sc_hd__and4_1 _1801_ (.A(_1319_),
    .B(_1321_),
    .C(_1323_),
    .D(_1333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1367_));
 sky130_fd_sc_hd__a41o_1 _1802_ (.A1(_1319_),
    .A2(_1320_),
    .A3(_1323_),
    .A4(_1333_),
    .B1(\genblk1[6].puf_buffer.cnt_1.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1368_));
 sky130_fd_sc_hd__and3b_1 _1803_ (.A_N(_1367_),
    .B(_1335_),
    .C(_1368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1369_));
 sky130_fd_sc_hd__clkbuf_1 _1804_ (.A(_1369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0211_));
 sky130_fd_sc_hd__inv_2 _1805_ (.A(_1322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1370_));
 sky130_fd_sc_hd__o221a_1 _1806_ (.A1(_1370_),
    .A2(_1341_),
    .B1(_1367_),
    .B2(net83),
    .C1(_1304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0212_));
 sky130_fd_sc_hd__nand4_1 _1807_ (.A(\genblk1[6].puf_buffer.cnt_1.ctr[15] ),
    .B(_1322_),
    .C(_1336_),
    .D(_1337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1371_));
 sky130_fd_sc_hd__a31o_1 _1808_ (.A1(_1322_),
    .A2(_1336_),
    .A3(_1337_),
    .B1(\genblk1[6].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1372_));
 sky130_fd_sc_hd__and3_1 _1809_ (.A(_1129_),
    .B(_1371_),
    .C(_1372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1373_));
 sky130_fd_sc_hd__clkbuf_1 _1810_ (.A(_1373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0213_));
 sky130_fd_sc_hd__inv_2 _1811_ (.A(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1374_));
 sky130_fd_sc_hd__and3b_1 _1812_ (.A_N(\genblk1[7].puf_buffer.cnt_1.finish ),
    .B(\genblk1[7].puf_buffer.cnt_2.finish ),
    .C(_0513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1375_));
 sky130_fd_sc_hd__clkbuf_1 _1813_ (.A(_1375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0250_));
 sky130_fd_sc_hd__o21bai_1 _1814_ (.A1(_1374_),
    .A2(_0250_),
    .B1_N(\genblk1[7].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0214_));
 sky130_fd_sc_hd__and3_1 _1815_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[12] ),
    .B(\genblk1[7].puf_buffer.cnt_2.ctr[11] ),
    .C(\genblk1[7].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1376_));
 sky130_fd_sc_hd__and2_1 _1816_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[13] ),
    .B(_1376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1377_));
 sky130_fd_sc_hd__and2_1 _1817_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[9] ),
    .B(\genblk1[7].puf_buffer.cnt_2.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1378_));
 sky130_fd_sc_hd__and4_1 _1818_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[3] ),
    .B(\genblk1[7].puf_buffer.cnt_2.ctr[2] ),
    .C(\genblk1[7].puf_buffer.cnt_2.ctr[1] ),
    .D(\genblk1[7].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1379_));
 sky130_fd_sc_hd__and3_1 _1819_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[7].puf_buffer.cnt_2.ctr[4] ),
    .C(_1379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1380_));
 sky130_fd_sc_hd__and4_1 _1820_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[7].puf_buffer.cnt_2.ctr[6] ),
    .C(_1378_),
    .D(_1380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1381_));
 sky130_fd_sc_hd__and3_1 _1821_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[14] ),
    .B(_1377_),
    .C(_1381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1382_));
 sky130_fd_sc_hd__a22o_1 _1822_ (.A1(_0670_),
    .A2(\genblk1[7].puf_buffer.cnt_2.finish ),
    .B1(_1382_),
    .B2(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0216_));
 sky130_fd_sc_hd__or2_1 _1823_ (.A(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1383_));
 sky130_fd_sc_hd__buf_2 _1824_ (.A(_1383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1384_));
 sky130_fd_sc_hd__a22o_1 _1825_ (.A1(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .A2(_0606_),
    .B1(_0619_),
    .B2(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1385_));
 sky130_fd_sc_hd__a221o_1 _1826_ (.A1(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .A2(_0603_),
    .B1(_0604_),
    .B2(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .C1(_1385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1386_));
 sky130_fd_sc_hd__a22o_1 _1827_ (.A1(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .A2(_0610_),
    .B1(_0622_),
    .B2(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1387_));
 sky130_fd_sc_hd__a211o_1 _1828_ (.A1(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .A2(net26),
    .B1(_1387_),
    .C1(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1388_));
 sky130_fd_sc_hd__a22o_1 _1829_ (.A1(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .A2(_0611_),
    .B1(_0621_),
    .B2(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1389_));
 sky130_fd_sc_hd__a22o_1 _1830_ (.A1(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .A2(_0624_),
    .B1(_0625_),
    .B2(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1390_));
 sky130_fd_sc_hd__a22o_1 _1831_ (.A1(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .A2(_0615_),
    .B1(_0618_),
    .B2(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1391_));
 sky130_fd_sc_hd__a22o_1 _1832_ (.A1(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .A2(_0616_),
    .B1(_0605_),
    .B2(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1392_));
 sky130_fd_sc_hd__or4_1 _1833_ (.A(_1389_),
    .B(_1390_),
    .C(_1391_),
    .D(_1392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1393_));
 sky130_fd_sc_hd__or3_1 _1834_ (.A(_1386_),
    .B(_1388_),
    .C(_1393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1394_));
 sky130_fd_sc_hd__buf_2 _1835_ (.A(_1394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1395_));
 sky130_fd_sc_hd__and3_1 _1836_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[0] ),
    .B(_1384_),
    .C(_1395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1396_));
 sky130_fd_sc_hd__a21o_1 _1837_ (.A1(_1384_),
    .A2(_1395_),
    .B1(\genblk1[7].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1397_));
 sky130_fd_sc_hd__and3b_1 _1838_ (.A_N(_1396_),
    .B(_1335_),
    .C(_1397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1398_));
 sky130_fd_sc_hd__clkbuf_1 _1839_ (.A(_1398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0217_));
 sky130_fd_sc_hd__nand2_1 _1840_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[1] ),
    .B(\genblk1[7].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1399_));
 sky130_fd_sc_hd__clkbuf_2 _1841_ (.A(_1383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_2 _1842_ (.A(_1394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1401_));
 sky130_fd_sc_hd__nand2_1 _1843_ (.A(_1400_),
    .B(_1401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1402_));
 sky130_fd_sc_hd__o221a_1 _1844_ (.A1(_1399_),
    .A2(_1402_),
    .B1(_1396_),
    .B2(net193),
    .C1(_1304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0218_));
 sky130_fd_sc_hd__inv_2 _1845_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1403_));
 sky130_fd_sc_hd__and4bb_1 _1846_ (.A_N(_1403_),
    .B_N(_1399_),
    .C(_1383_),
    .D(_1394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1404_));
 sky130_fd_sc_hd__a41o_1 _1847_ (.A1(\genblk1[7].puf_buffer.cnt_2.ctr[1] ),
    .A2(\genblk1[7].puf_buffer.cnt_2.ctr[0] ),
    .A3(_1384_),
    .A4(_1395_),
    .B1(\genblk1[7].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1405_));
 sky130_fd_sc_hd__and3b_1 _1848_ (.A_N(_1404_),
    .B(_1335_),
    .C(_1405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1406_));
 sky130_fd_sc_hd__clkbuf_1 _1849_ (.A(_1406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0219_));
 sky130_fd_sc_hd__inv_2 _1850_ (.A(_1379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1407_));
 sky130_fd_sc_hd__o221a_1 _1851_ (.A1(_1407_),
    .A2(_1402_),
    .B1(_1404_),
    .B2(net145),
    .C1(_1304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0220_));
 sky130_fd_sc_hd__and4_1 _1852_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[4] ),
    .B(_1379_),
    .C(_1383_),
    .D(_1394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1408_));
 sky130_fd_sc_hd__a31o_1 _1853_ (.A1(_1379_),
    .A2(_1384_),
    .A3(_1395_),
    .B1(\genblk1[7].puf_buffer.cnt_2.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1409_));
 sky130_fd_sc_hd__and3b_1 _1854_ (.A_N(_1408_),
    .B(_1335_),
    .C(_1409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1410_));
 sky130_fd_sc_hd__clkbuf_1 _1855_ (.A(_1410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0221_));
 sky130_fd_sc_hd__inv_2 _1856_ (.A(_1380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1411_));
 sky130_fd_sc_hd__buf_2 _1857_ (.A(_0638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1412_));
 sky130_fd_sc_hd__o221a_1 _1858_ (.A1(_1411_),
    .A2(_1402_),
    .B1(_1408_),
    .B2(net98),
    .C1(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0222_));
 sky130_fd_sc_hd__and4_1 _1859_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[6] ),
    .B(_1380_),
    .C(_1384_),
    .D(_1395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1413_));
 sky130_fd_sc_hd__clkbuf_2 _1860_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1414_));
 sky130_fd_sc_hd__a31o_1 _1861_ (.A1(_1380_),
    .A2(_1384_),
    .A3(_1395_),
    .B1(\genblk1[7].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1415_));
 sky130_fd_sc_hd__and3b_1 _1862_ (.A_N(_1413_),
    .B(_1414_),
    .C(_1415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1416_));
 sky130_fd_sc_hd__clkbuf_1 _1863_ (.A(_1416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0223_));
 sky130_fd_sc_hd__and3_1 _1864_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[7].puf_buffer.cnt_2.ctr[6] ),
    .C(_1380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1417_));
 sky130_fd_sc_hd__nand3_1 _1865_ (.A(_1417_),
    .B(_1400_),
    .C(_1401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1418_));
 sky130_fd_sc_hd__o211a_1 _1866_ (.A1(net184),
    .A2(_1413_),
    .B1(_1418_),
    .C1(_1308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0224_));
 sky130_fd_sc_hd__and4_1 _1867_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[8] ),
    .B(_1417_),
    .C(_1384_),
    .D(_1395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1419_));
 sky130_fd_sc_hd__a31o_1 _1868_ (.A1(_1417_),
    .A2(_1384_),
    .A3(_1395_),
    .B1(\genblk1[7].puf_buffer.cnt_2.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1420_));
 sky130_fd_sc_hd__and3b_1 _1869_ (.A_N(_1419_),
    .B(_1414_),
    .C(_1420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1421_));
 sky130_fd_sc_hd__clkbuf_1 _1870_ (.A(_1421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0225_));
 sky130_fd_sc_hd__and4_2 _1871_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[7].puf_buffer.cnt_2.ctr[6] ),
    .C(_1378_),
    .D(_1380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1422_));
 sky130_fd_sc_hd__a31o_1 _1872_ (.A1(_1422_),
    .A2(_1400_),
    .A3(_1401_),
    .B1(_0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1423_));
 sky130_fd_sc_hd__o21ba_1 _1873_ (.A1(net60),
    .A2(_1419_),
    .B1_N(_1423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0226_));
 sky130_fd_sc_hd__a31o_1 _1874_ (.A1(_1422_),
    .A2(_1384_),
    .A3(_1395_),
    .B1(\genblk1[7].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1424_));
 sky130_fd_sc_hd__nand4_1 _1875_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[10] ),
    .B(_1422_),
    .C(_1400_),
    .D(_1401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1425_));
 sky130_fd_sc_hd__and3_1 _1876_ (.A(_1129_),
    .B(_1424_),
    .C(_1425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1426_));
 sky130_fd_sc_hd__clkbuf_1 _1877_ (.A(_1426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0227_));
 sky130_fd_sc_hd__inv_2 _1878_ (.A(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1427_));
 sky130_fd_sc_hd__and2_1 _1879_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[11] ),
    .B(\genblk1[7].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1428_));
 sky130_fd_sc_hd__and4_1 _1880_ (.A(_1428_),
    .B(_1422_),
    .C(_1400_),
    .D(_1401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1429_));
 sky130_fd_sc_hd__a211oi_1 _1881_ (.A1(_1427_),
    .A2(_1425_),
    .B1(_1429_),
    .C1(_0814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0228_));
 sky130_fd_sc_hd__a41o_1 _1882_ (.A1(_1376_),
    .A2(_1422_),
    .A3(_1400_),
    .A4(_1401_),
    .B1(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1430_));
 sky130_fd_sc_hd__o21ba_1 _1883_ (.A1(net69),
    .A2(_1429_),
    .B1_N(_1430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0229_));
 sky130_fd_sc_hd__and4_1 _1884_ (.A(_1376_),
    .B(_1422_),
    .C(_1400_),
    .D(_1401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1431_));
 sky130_fd_sc_hd__nand4_1 _1885_ (.A(_1377_),
    .B(_1422_),
    .C(_1400_),
    .D(_1401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1432_));
 sky130_fd_sc_hd__o211a_1 _1886_ (.A1(net142),
    .A2(_1431_),
    .B1(_1432_),
    .C1(_1308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0230_));
 sky130_fd_sc_hd__inv_2 _1887_ (.A(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1433_));
 sky130_fd_sc_hd__and3_1 _1888_ (.A(_1382_),
    .B(_1400_),
    .C(_1401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1434_));
 sky130_fd_sc_hd__a211oi_1 _1889_ (.A1(_1433_),
    .A2(_1432_),
    .B1(_1434_),
    .C1(_0814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0231_));
 sky130_fd_sc_hd__a31o_1 _1890_ (.A1(_1382_),
    .A2(_1384_),
    .A3(_1395_),
    .B1(\genblk1[7].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1435_));
 sky130_fd_sc_hd__nand4_1 _1891_ (.A(\genblk1[7].puf_buffer.cnt_2.ctr[15] ),
    .B(_1382_),
    .C(_1400_),
    .D(_1401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1436_));
 sky130_fd_sc_hd__and3_1 _1892_ (.A(_1129_),
    .B(_1435_),
    .C(_1436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1437_));
 sky130_fd_sc_hd__clkbuf_1 _1893_ (.A(_1437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0232_));
 sky130_fd_sc_hd__and3_1 _1894_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[12] ),
    .B(\genblk1[7].puf_buffer.cnt_1.ctr[11] ),
    .C(\genblk1[7].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1438_));
 sky130_fd_sc_hd__and2_1 _1895_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[13] ),
    .B(_1438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1439_));
 sky130_fd_sc_hd__and2_1 _1896_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[9] ),
    .B(\genblk1[7].puf_buffer.cnt_1.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1440_));
 sky130_fd_sc_hd__and4_1 _1897_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[3] ),
    .B(\genblk1[7].puf_buffer.cnt_1.ctr[2] ),
    .C(\genblk1[7].puf_buffer.cnt_1.ctr[1] ),
    .D(\genblk1[7].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1441_));
 sky130_fd_sc_hd__and3_1 _1898_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[7].puf_buffer.cnt_1.ctr[4] ),
    .C(_1441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1442_));
 sky130_fd_sc_hd__and4_1 _1899_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[7].puf_buffer.cnt_1.ctr[6] ),
    .C(_1440_),
    .D(_1442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1443_));
 sky130_fd_sc_hd__and3_1 _1900_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[14] ),
    .B(_1439_),
    .C(_1443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1444_));
 sky130_fd_sc_hd__a22o_1 _1901_ (.A1(_0670_),
    .A2(\genblk1[7].puf_buffer.cnt_1.finish ),
    .B1(_1444_),
    .B2(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0233_));
 sky130_fd_sc_hd__or2_1 _1902_ (.A(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1445_));
 sky130_fd_sc_hd__buf_2 _1903_ (.A(_1445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1446_));
 sky130_fd_sc_hd__a22o_1 _1904_ (.A1(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .A2(_0700_),
    .B1(_0695_),
    .B2(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1447_));
 sky130_fd_sc_hd__a221o_1 _1905_ (.A1(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .A2(_0699_),
    .B1(net11),
    .B2(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .C1(_1447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1448_));
 sky130_fd_sc_hd__a22o_1 _1906_ (.A1(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .A2(_0687_),
    .B1(_0706_),
    .B2(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1449_));
 sky130_fd_sc_hd__a22o_1 _1907_ (.A1(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .A2(_0705_),
    .B1(_0702_),
    .B2(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1450_));
 sky130_fd_sc_hd__a211o_1 _1908_ (.A1(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .A2(_0688_),
    .B1(_1449_),
    .C1(_1450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1451_));
 sky130_fd_sc_hd__a221o_1 _1909_ (.A1(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .A2(_0690_),
    .B1(_0709_),
    .B2(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .C1(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1452_));
 sky130_fd_sc_hd__a22o_1 _1910_ (.A1(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .A2(_0689_),
    .B1(net24),
    .B2(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1453_));
 sky130_fd_sc_hd__a22o_1 _1911_ (.A1(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .A2(_0694_),
    .B1(net14),
    .B2(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1454_));
 sky130_fd_sc_hd__or3_1 _1912_ (.A(_1452_),
    .B(_1453_),
    .C(_1454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1455_));
 sky130_fd_sc_hd__or3_2 _1913_ (.A(_1448_),
    .B(_1451_),
    .C(_1455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1456_));
 sky130_fd_sc_hd__buf_2 _1914_ (.A(_1456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1457_));
 sky130_fd_sc_hd__and3_1 _1915_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[0] ),
    .B(_1446_),
    .C(_1457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1458_));
 sky130_fd_sc_hd__a21o_1 _1916_ (.A1(_1446_),
    .A2(_1457_),
    .B1(\genblk1[7].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1459_));
 sky130_fd_sc_hd__and3b_1 _1917_ (.A_N(_1458_),
    .B(_1414_),
    .C(_1459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1460_));
 sky130_fd_sc_hd__clkbuf_1 _1918_ (.A(_1460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0234_));
 sky130_fd_sc_hd__nand2_1 _1919_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[1] ),
    .B(\genblk1[7].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1461_));
 sky130_fd_sc_hd__buf_2 _1920_ (.A(_1445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1462_));
 sky130_fd_sc_hd__buf_2 _1921_ (.A(_1456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1463_));
 sky130_fd_sc_hd__nand2_1 _1922_ (.A(_1462_),
    .B(_1463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1464_));
 sky130_fd_sc_hd__o221a_1 _1923_ (.A1(_1461_),
    .A2(_1464_),
    .B1(_1458_),
    .B2(net205),
    .C1(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0235_));
 sky130_fd_sc_hd__inv_2 _1924_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1465_));
 sky130_fd_sc_hd__and4bb_1 _1925_ (.A_N(_1465_),
    .B_N(_1461_),
    .C(_1445_),
    .D(_1456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1466_));
 sky130_fd_sc_hd__a41o_1 _1926_ (.A1(\genblk1[7].puf_buffer.cnt_1.ctr[1] ),
    .A2(\genblk1[7].puf_buffer.cnt_1.ctr[0] ),
    .A3(_1446_),
    .A4(_1457_),
    .B1(\genblk1[7].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1467_));
 sky130_fd_sc_hd__and3b_1 _1927_ (.A_N(_1466_),
    .B(_1414_),
    .C(_1467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1468_));
 sky130_fd_sc_hd__clkbuf_1 _1928_ (.A(_1468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0236_));
 sky130_fd_sc_hd__inv_2 _1929_ (.A(_1441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1469_));
 sky130_fd_sc_hd__o221a_1 _1930_ (.A1(_1469_),
    .A2(_1464_),
    .B1(_1466_),
    .B2(net115),
    .C1(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0237_));
 sky130_fd_sc_hd__and4_1 _1931_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[4] ),
    .B(_1441_),
    .C(_1445_),
    .D(_1456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1470_));
 sky130_fd_sc_hd__a31o_1 _1932_ (.A1(_1441_),
    .A2(_1446_),
    .A3(_1457_),
    .B1(\genblk1[7].puf_buffer.cnt_1.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1471_));
 sky130_fd_sc_hd__and3b_1 _1933_ (.A_N(_1470_),
    .B(_1414_),
    .C(_1471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1472_));
 sky130_fd_sc_hd__clkbuf_1 _1934_ (.A(_1472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0238_));
 sky130_fd_sc_hd__inv_2 _1935_ (.A(_1442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1473_));
 sky130_fd_sc_hd__o221a_1 _1936_ (.A1(_1473_),
    .A2(_1464_),
    .B1(_1470_),
    .B2(net126),
    .C1(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0239_));
 sky130_fd_sc_hd__and4_1 _1937_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[6] ),
    .B(_1442_),
    .C(_1446_),
    .D(_1457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1474_));
 sky130_fd_sc_hd__a31o_1 _1938_ (.A1(_1442_),
    .A2(_1446_),
    .A3(_1457_),
    .B1(\genblk1[7].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1475_));
 sky130_fd_sc_hd__and3b_1 _1939_ (.A_N(_1474_),
    .B(_1414_),
    .C(_1475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1476_));
 sky130_fd_sc_hd__clkbuf_1 _1940_ (.A(_1476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0240_));
 sky130_fd_sc_hd__and3_1 _1941_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[7].puf_buffer.cnt_1.ctr[6] ),
    .C(_1442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1477_));
 sky130_fd_sc_hd__nand3_1 _1942_ (.A(_1477_),
    .B(_1462_),
    .C(_1463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1478_));
 sky130_fd_sc_hd__o211a_1 _1943_ (.A1(net180),
    .A2(_1474_),
    .B1(_1478_),
    .C1(_1308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0241_));
 sky130_fd_sc_hd__and4_1 _1944_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[8] ),
    .B(_1477_),
    .C(_1446_),
    .D(_1457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1479_));
 sky130_fd_sc_hd__a31o_1 _1945_ (.A1(_1477_),
    .A2(_1446_),
    .A3(_1457_),
    .B1(\genblk1[7].puf_buffer.cnt_1.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1480_));
 sky130_fd_sc_hd__and3b_1 _1946_ (.A_N(_1479_),
    .B(_1414_),
    .C(_1480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1481_));
 sky130_fd_sc_hd__clkbuf_1 _1947_ (.A(_1481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0242_));
 sky130_fd_sc_hd__and4_2 _1948_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[7].puf_buffer.cnt_1.ctr[6] ),
    .C(_1440_),
    .D(_1442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1482_));
 sky130_fd_sc_hd__a31o_1 _1949_ (.A1(_1482_),
    .A2(_1462_),
    .A3(_1463_),
    .B1(_0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1483_));
 sky130_fd_sc_hd__o21ba_1 _1950_ (.A1(net67),
    .A2(_1479_),
    .B1_N(_1483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0243_));
 sky130_fd_sc_hd__a31o_1 _1951_ (.A1(_1482_),
    .A2(_1446_),
    .A3(_1457_),
    .B1(\genblk1[7].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1484_));
 sky130_fd_sc_hd__nand4_1 _1952_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[10] ),
    .B(_1482_),
    .C(_1462_),
    .D(_1463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1485_));
 sky130_fd_sc_hd__and3_1 _1953_ (.A(_1129_),
    .B(_1484_),
    .C(_1485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1486_));
 sky130_fd_sc_hd__clkbuf_1 _1954_ (.A(_1486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0244_));
 sky130_fd_sc_hd__inv_2 _1955_ (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1487_));
 sky130_fd_sc_hd__and2_1 _1956_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[11] ),
    .B(\genblk1[7].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1488_));
 sky130_fd_sc_hd__and4_1 _1957_ (.A(_1488_),
    .B(_1482_),
    .C(_1462_),
    .D(_1463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1489_));
 sky130_fd_sc_hd__a211oi_1 _1958_ (.A1(_1487_),
    .A2(_1485_),
    .B1(_1489_),
    .C1(_0814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0245_));
 sky130_fd_sc_hd__a41o_1 _1959_ (.A1(_1438_),
    .A2(_1482_),
    .A3(_1462_),
    .A4(_1463_),
    .B1(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1490_));
 sky130_fd_sc_hd__o21ba_1 _1960_ (.A1(net51),
    .A2(_1489_),
    .B1_N(_1490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0246_));
 sky130_fd_sc_hd__and4_1 _1961_ (.A(_1438_),
    .B(_1482_),
    .C(_1462_),
    .D(_1463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1491_));
 sky130_fd_sc_hd__nand4_1 _1962_ (.A(_1439_),
    .B(_1482_),
    .C(_1462_),
    .D(_1463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1492_));
 sky130_fd_sc_hd__o211a_1 _1963_ (.A1(net119),
    .A2(_1491_),
    .B1(_1492_),
    .C1(_1308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0247_));
 sky130_fd_sc_hd__inv_2 _1964_ (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1493_));
 sky130_fd_sc_hd__and3_1 _1965_ (.A(_1444_),
    .B(_1462_),
    .C(_1463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1494_));
 sky130_fd_sc_hd__a211oi_1 _1966_ (.A1(_1493_),
    .A2(_1492_),
    .B1(_1494_),
    .C1(_0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0248_));
 sky130_fd_sc_hd__a31o_1 _1967_ (.A1(_1444_),
    .A2(_1446_),
    .A3(_1457_),
    .B1(\genblk1[7].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1495_));
 sky130_fd_sc_hd__nand4_1 _1968_ (.A(\genblk1[7].puf_buffer.cnt_1.ctr[15] ),
    .B(_1444_),
    .C(_1462_),
    .D(_1463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1496_));
 sky130_fd_sc_hd__and3_1 _1969_ (.A(_1129_),
    .B(_1495_),
    .C(_1496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1497_));
 sky130_fd_sc_hd__clkbuf_1 _1970_ (.A(_1497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0249_));
 sky130_fd_sc_hd__inv_2 _1971_ (.A(net161),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1498_));
 sky130_fd_sc_hd__and3b_1 _1972_ (.A_N(\genblk1[0].puf_buffer.cnt_1.finish ),
    .B(\genblk1[0].puf_buffer.cnt_2.finish ),
    .C(_0550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1499_));
 sky130_fd_sc_hd__clkbuf_1 _1973_ (.A(_1499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0287_));
 sky130_fd_sc_hd__o21bai_1 _1974_ (.A1(_1498_),
    .A2(_0287_),
    .B1_N(\genblk1[0].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0251_));
 sky130_fd_sc_hd__and4_1 _1975_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[3] ),
    .B(\genblk1[0].puf_buffer.cnt_2.ctr[2] ),
    .C(\genblk1[0].puf_buffer.cnt_2.ctr[1] ),
    .D(\genblk1[0].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1500_));
 sky130_fd_sc_hd__and2_1 _1976_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[0].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1501_));
 sky130_fd_sc_hd__and4_1 _1977_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[0].puf_buffer.cnt_2.ctr[4] ),
    .C(_1500_),
    .D(_1501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1502_));
 sky130_fd_sc_hd__and3_1 _1978_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[9] ),
    .B(\genblk1[0].puf_buffer.cnt_2.ctr[8] ),
    .C(_1502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1503_));
 sky130_fd_sc_hd__and3_1 _1979_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[12] ),
    .B(\genblk1[0].puf_buffer.cnt_2.ctr[11] ),
    .C(\genblk1[0].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1504_));
 sky130_fd_sc_hd__and2_1 _1980_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[13] ),
    .B(_1504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1505_));
 sky130_fd_sc_hd__and3_1 _1981_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[14] ),
    .B(_1503_),
    .C(_1505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1506_));
 sky130_fd_sc_hd__a22o_1 _1982_ (.A1(_0670_),
    .A2(net127),
    .B1(_1506_),
    .B2(\genblk1[0].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0252_));
 sky130_fd_sc_hd__or2_2 _1983_ (.A(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1507_));
 sky130_fd_sc_hd__a22o_1 _1984_ (.A1(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .A2(_0603_),
    .B1(_0604_),
    .B2(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1508_));
 sky130_fd_sc_hd__a221o_1 _1985_ (.A1(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .A2(_0624_),
    .B1(_0605_),
    .B2(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .C1(_1508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1509_));
 sky130_fd_sc_hd__a22o_1 _1986_ (.A1(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .A2(_0615_),
    .B1(net19),
    .B2(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1510_));
 sky130_fd_sc_hd__a211o_1 _1987_ (.A1(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .A2(_0610_),
    .B1(_1510_),
    .C1(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1511_));
 sky130_fd_sc_hd__a22o_1 _1988_ (.A1(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .A2(_0606_),
    .B1(net17),
    .B2(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1512_));
 sky130_fd_sc_hd__a22o_1 _1989_ (.A1(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .A2(net26),
    .B1(_0625_),
    .B2(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1513_));
 sky130_fd_sc_hd__a22o_1 _1990_ (.A1(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .A2(_0611_),
    .B1(_0618_),
    .B2(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1514_));
 sky130_fd_sc_hd__a22o_1 _1991_ (.A1(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .A2(_0621_),
    .B1(_0622_),
    .B2(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1515_));
 sky130_fd_sc_hd__or4_1 _1992_ (.A(_1512_),
    .B(_1513_),
    .C(_1514_),
    .D(_1515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1516_));
 sky130_fd_sc_hd__or3_4 _1993_ (.A(_1509_),
    .B(_1511_),
    .C(_1516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1517_));
 sky130_fd_sc_hd__and3_1 _1994_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[0] ),
    .B(_1507_),
    .C(_1517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1518_));
 sky130_fd_sc_hd__buf_2 _1995_ (.A(_1507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1519_));
 sky130_fd_sc_hd__buf_2 _1996_ (.A(_1517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1520_));
 sky130_fd_sc_hd__a21o_1 _1997_ (.A1(_1519_),
    .A2(_1520_),
    .B1(\genblk1[0].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1521_));
 sky130_fd_sc_hd__and3b_1 _1998_ (.A_N(_1518_),
    .B(_1414_),
    .C(_1521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1522_));
 sky130_fd_sc_hd__clkbuf_1 _1999_ (.A(_1522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0253_));
 sky130_fd_sc_hd__nand2_1 _2000_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[1] ),
    .B(\genblk1[0].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1523_));
 sky130_fd_sc_hd__nand2_2 _2001_ (.A(_1519_),
    .B(_1520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1524_));
 sky130_fd_sc_hd__o221a_1 _2002_ (.A1(_1523_),
    .A2(_1524_),
    .B1(_1518_),
    .B2(net187),
    .C1(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0254_));
 sky130_fd_sc_hd__inv_2 _2003_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1525_));
 sky130_fd_sc_hd__and4bb_1 _2004_ (.A_N(_1525_),
    .B_N(_1523_),
    .C(_1507_),
    .D(_1517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1526_));
 sky130_fd_sc_hd__a41o_1 _2005_ (.A1(\genblk1[0].puf_buffer.cnt_2.ctr[1] ),
    .A2(\genblk1[0].puf_buffer.cnt_2.ctr[0] ),
    .A3(_1507_),
    .A4(_1517_),
    .B1(\genblk1[0].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1527_));
 sky130_fd_sc_hd__and3b_1 _2006_ (.A_N(_1526_),
    .B(_1414_),
    .C(_1527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1528_));
 sky130_fd_sc_hd__clkbuf_1 _2007_ (.A(_1528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0255_));
 sky130_fd_sc_hd__inv_2 _2008_ (.A(_1500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1529_));
 sky130_fd_sc_hd__o221a_1 _2009_ (.A1(_1529_),
    .A2(_1524_),
    .B1(_1526_),
    .B2(net64),
    .C1(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0256_));
 sky130_fd_sc_hd__and4_1 _2010_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[4] ),
    .B(_1500_),
    .C(_1507_),
    .D(_1517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1530_));
 sky130_fd_sc_hd__a31o_1 _2011_ (.A1(_1500_),
    .A2(_1519_),
    .A3(_1520_),
    .B1(\genblk1[0].puf_buffer.cnt_2.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1531_));
 sky130_fd_sc_hd__and3b_1 _2012_ (.A_N(_1530_),
    .B(_1414_),
    .C(_1531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1532_));
 sky130_fd_sc_hd__clkbuf_1 _2013_ (.A(_1532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0257_));
 sky130_fd_sc_hd__and3_1 _2014_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[0].puf_buffer.cnt_2.ctr[4] ),
    .C(_1500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1533_));
 sky130_fd_sc_hd__inv_2 _2015_ (.A(_1533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1534_));
 sky130_fd_sc_hd__o221a_1 _2016_ (.A1(_1534_),
    .A2(_1524_),
    .B1(_1530_),
    .B2(net162),
    .C1(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0258_));
 sky130_fd_sc_hd__and4_1 _2017_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[6] ),
    .B(_1533_),
    .C(_1507_),
    .D(_1517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1535_));
 sky130_fd_sc_hd__a31o_1 _2018_ (.A1(_1533_),
    .A2(_1519_),
    .A3(_1520_),
    .B1(\genblk1[0].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1536_));
 sky130_fd_sc_hd__and3b_1 _2019_ (.A_N(_1535_),
    .B(_0588_),
    .C(_1536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1537_));
 sky130_fd_sc_hd__clkbuf_1 _2020_ (.A(_1537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0259_));
 sky130_fd_sc_hd__inv_2 _2021_ (.A(_1502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1538_));
 sky130_fd_sc_hd__o221a_1 _2022_ (.A1(_1538_),
    .A2(_1524_),
    .B1(_1535_),
    .B2(net68),
    .C1(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0260_));
 sky130_fd_sc_hd__and4_1 _2023_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[8] ),
    .B(_1502_),
    .C(_1507_),
    .D(_1517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1539_));
 sky130_fd_sc_hd__a31o_1 _2024_ (.A1(_1502_),
    .A2(_1519_),
    .A3(_1520_),
    .B1(\genblk1[0].puf_buffer.cnt_2.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1540_));
 sky130_fd_sc_hd__and3b_1 _2025_ (.A_N(_1539_),
    .B(_0588_),
    .C(_1540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _2026_ (.A(_1541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0261_));
 sky130_fd_sc_hd__nand3_1 _2027_ (.A(_1503_),
    .B(_1519_),
    .C(_1520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1542_));
 sky130_fd_sc_hd__o211a_1 _2028_ (.A1(net88),
    .A2(_1539_),
    .B1(_1542_),
    .C1(_1308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0262_));
 sky130_fd_sc_hd__and4_1 _2029_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[10] ),
    .B(_1503_),
    .C(_1507_),
    .D(_1517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1543_));
 sky130_fd_sc_hd__a31o_1 _2030_ (.A1(_1503_),
    .A2(_1519_),
    .A3(_1520_),
    .B1(\genblk1[0].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1544_));
 sky130_fd_sc_hd__and3b_1 _2031_ (.A_N(_1543_),
    .B(_0588_),
    .C(_1544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1545_));
 sky130_fd_sc_hd__clkbuf_1 _2032_ (.A(_1545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0263_));
 sky130_fd_sc_hd__nand2_1 _2033_ (.A(net190),
    .B(\genblk1[0].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1546_));
 sky130_fd_sc_hd__o221a_1 _2034_ (.A1(_1546_),
    .A2(_1542_),
    .B1(_1543_),
    .B2(net190),
    .C1(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0264_));
 sky130_fd_sc_hd__inv_2 _2035_ (.A(_1504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1547_));
 sky130_fd_sc_hd__and2_1 _2036_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[11] ),
    .B(\genblk1[0].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1548_));
 sky130_fd_sc_hd__a41o_1 _2037_ (.A1(_1503_),
    .A2(_1548_),
    .A3(_1519_),
    .A4(_1520_),
    .B1(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1549_));
 sky130_fd_sc_hd__o211a_1 _2038_ (.A1(_1547_),
    .A2(_1542_),
    .B1(_1549_),
    .C1(_1308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0265_));
 sky130_fd_sc_hd__and4_1 _2039_ (.A(_1503_),
    .B(_1505_),
    .C(_1507_),
    .D(_1517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1550_));
 sky130_fd_sc_hd__a41o_1 _2040_ (.A1(_1503_),
    .A2(_1504_),
    .A3(_1507_),
    .A4(_1517_),
    .B1(\genblk1[0].puf_buffer.cnt_2.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1551_));
 sky130_fd_sc_hd__and3b_1 _2041_ (.A_N(_1550_),
    .B(_0588_),
    .C(_1551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1552_));
 sky130_fd_sc_hd__clkbuf_1 _2042_ (.A(_1552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0266_));
 sky130_fd_sc_hd__inv_2 _2043_ (.A(_1506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1553_));
 sky130_fd_sc_hd__o221a_1 _2044_ (.A1(_1553_),
    .A2(_1524_),
    .B1(_1550_),
    .B2(net72),
    .C1(_1412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0267_));
 sky130_fd_sc_hd__nand4_1 _2045_ (.A(\genblk1[0].puf_buffer.cnt_2.ctr[15] ),
    .B(_1506_),
    .C(_1519_),
    .D(_1520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1554_));
 sky130_fd_sc_hd__a31o_1 _2046_ (.A1(_1506_),
    .A2(_1519_),
    .A3(_1520_),
    .B1(\genblk1[0].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1555_));
 sky130_fd_sc_hd__and3_1 _2047_ (.A(_1129_),
    .B(_1554_),
    .C(_1555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1556_));
 sky130_fd_sc_hd__clkbuf_1 _2048_ (.A(_1556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0268_));
 sky130_fd_sc_hd__and3_1 _2049_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[12] ),
    .B(\genblk1[0].puf_buffer.cnt_1.ctr[11] ),
    .C(\genblk1[0].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1557_));
 sky130_fd_sc_hd__and2_1 _2050_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[13] ),
    .B(_1557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1558_));
 sky130_fd_sc_hd__and2_1 _2051_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[9] ),
    .B(\genblk1[0].puf_buffer.cnt_1.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1559_));
 sky130_fd_sc_hd__and4_1 _2052_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[3] ),
    .B(\genblk1[0].puf_buffer.cnt_1.ctr[2] ),
    .C(\genblk1[0].puf_buffer.cnt_1.ctr[1] ),
    .D(\genblk1[0].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1560_));
 sky130_fd_sc_hd__and3_1 _2053_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[0].puf_buffer.cnt_1.ctr[4] ),
    .C(_1560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1561_));
 sky130_fd_sc_hd__and4_1 _2054_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[0].puf_buffer.cnt_1.ctr[6] ),
    .C(_1559_),
    .D(_1561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1562_));
 sky130_fd_sc_hd__and3_1 _2055_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[14] ),
    .B(_1558_),
    .C(_1562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1563_));
 sky130_fd_sc_hd__a22o_1 _2056_ (.A1(\genblk1[0].puf_buffer.cnt_1.finish ),
    .A2(_0670_),
    .B1(_1563_),
    .B2(net167),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0269_));
 sky130_fd_sc_hd__or2_1 _2057_ (.A(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1564_));
 sky130_fd_sc_hd__buf_2 _2058_ (.A(_1564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1565_));
 sky130_fd_sc_hd__a22o_1 _2059_ (.A1(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .A2(_0687_),
    .B1(_0706_),
    .B2(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1566_));
 sky130_fd_sc_hd__a22o_1 _2060_ (.A1(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .A2(net23),
    .B1(net13),
    .B2(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1567_));
 sky130_fd_sc_hd__a211o_1 _2061_ (.A1(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .A2(_0709_),
    .B1(_1566_),
    .C1(_1567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1568_));
 sky130_fd_sc_hd__a22o_1 _2062_ (.A1(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .A2(_0705_),
    .B1(_0690_),
    .B2(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1569_));
 sky130_fd_sc_hd__a221o_1 _2063_ (.A1(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .A2(_0699_),
    .B1(net10),
    .B2(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .C1(_1569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1570_));
 sky130_fd_sc_hd__a22o_1 _2064_ (.A1(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .A2(_0700_),
    .B1(_0694_),
    .B2(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1571_));
 sky130_fd_sc_hd__a221o_1 _2065_ (.A1(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .A2(_0689_),
    .B1(net15),
    .B2(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .C1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1572_));
 sky130_fd_sc_hd__a22o_1 _2066_ (.A1(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .A2(_0695_),
    .B1(_0702_),
    .B2(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1573_));
 sky130_fd_sc_hd__or3_1 _2067_ (.A(_1571_),
    .B(_1572_),
    .C(_1573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1574_));
 sky130_fd_sc_hd__or3_2 _2068_ (.A(_1568_),
    .B(_1570_),
    .C(_1574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1575_));
 sky130_fd_sc_hd__buf_2 _2069_ (.A(_1575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1576_));
 sky130_fd_sc_hd__and3_1 _2070_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[0] ),
    .B(_1565_),
    .C(_1576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1577_));
 sky130_fd_sc_hd__a21o_1 _2071_ (.A1(_1565_),
    .A2(_1576_),
    .B1(\genblk1[0].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1578_));
 sky130_fd_sc_hd__and3b_1 _2072_ (.A_N(_1577_),
    .B(_0588_),
    .C(_1578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1579_));
 sky130_fd_sc_hd__clkbuf_1 _2073_ (.A(_1579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0270_));
 sky130_fd_sc_hd__nand2_1 _2074_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[1] ),
    .B(\genblk1[0].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1580_));
 sky130_fd_sc_hd__clkbuf_2 _2075_ (.A(_1564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1581_));
 sky130_fd_sc_hd__clkbuf_2 _2076_ (.A(_1575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1582_));
 sky130_fd_sc_hd__nand2_1 _2077_ (.A(_1581_),
    .B(_1582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1583_));
 sky130_fd_sc_hd__o221a_1 _2078_ (.A1(_1580_),
    .A2(_1583_),
    .B1(_1577_),
    .B2(net202),
    .C1(_0589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0271_));
 sky130_fd_sc_hd__inv_2 _2079_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1584_));
 sky130_fd_sc_hd__and4bb_1 _2080_ (.A_N(_1584_),
    .B_N(_1580_),
    .C(_1564_),
    .D(_1575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1585_));
 sky130_fd_sc_hd__a41o_1 _2081_ (.A1(\genblk1[0].puf_buffer.cnt_1.ctr[1] ),
    .A2(\genblk1[0].puf_buffer.cnt_1.ctr[0] ),
    .A3(_1565_),
    .A4(_1576_),
    .B1(\genblk1[0].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1586_));
 sky130_fd_sc_hd__and3b_1 _2082_ (.A_N(_1585_),
    .B(_0588_),
    .C(_1586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1587_));
 sky130_fd_sc_hd__clkbuf_1 _2083_ (.A(_1587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0272_));
 sky130_fd_sc_hd__inv_2 _2084_ (.A(_1560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1588_));
 sky130_fd_sc_hd__o221a_1 _2085_ (.A1(_1588_),
    .A2(_1583_),
    .B1(_1585_),
    .B2(net132),
    .C1(_0589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0273_));
 sky130_fd_sc_hd__and4_1 _2086_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[4] ),
    .B(_1560_),
    .C(_1564_),
    .D(_1575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1589_));
 sky130_fd_sc_hd__a31o_1 _2087_ (.A1(_1560_),
    .A2(_1565_),
    .A3(_1576_),
    .B1(\genblk1[0].puf_buffer.cnt_1.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1590_));
 sky130_fd_sc_hd__and3b_1 _2088_ (.A_N(_1589_),
    .B(_0588_),
    .C(_1590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1591_));
 sky130_fd_sc_hd__clkbuf_1 _2089_ (.A(_1591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0274_));
 sky130_fd_sc_hd__inv_2 _2090_ (.A(_1561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1592_));
 sky130_fd_sc_hd__o221a_1 _2091_ (.A1(_1592_),
    .A2(_1583_),
    .B1(_1589_),
    .B2(net91),
    .C1(_0589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0275_));
 sky130_fd_sc_hd__and4_1 _2092_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[6] ),
    .B(_1561_),
    .C(_1565_),
    .D(_1576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1593_));
 sky130_fd_sc_hd__a31o_1 _2093_ (.A1(_1561_),
    .A2(_1565_),
    .A3(_1576_),
    .B1(\genblk1[0].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1594_));
 sky130_fd_sc_hd__and3b_1 _2094_ (.A_N(_1593_),
    .B(_0588_),
    .C(_1594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1595_));
 sky130_fd_sc_hd__clkbuf_1 _2095_ (.A(_1595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0276_));
 sky130_fd_sc_hd__and3_1 _2096_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[0].puf_buffer.cnt_1.ctr[6] ),
    .C(_1561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1596_));
 sky130_fd_sc_hd__nand3_1 _2097_ (.A(_1596_),
    .B(_1581_),
    .C(_1582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1597_));
 sky130_fd_sc_hd__o211a_1 _2098_ (.A1(net181),
    .A2(_1593_),
    .B1(_1597_),
    .C1(_1308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0277_));
 sky130_fd_sc_hd__and4_1 _2099_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[8] ),
    .B(_1596_),
    .C(_1565_),
    .D(_1576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1598_));
 sky130_fd_sc_hd__a31o_1 _2100_ (.A1(_1596_),
    .A2(_1565_),
    .A3(_1576_),
    .B1(\genblk1[0].puf_buffer.cnt_1.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1599_));
 sky130_fd_sc_hd__and3b_1 _2101_ (.A_N(_1598_),
    .B(_0588_),
    .C(_1599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1600_));
 sky130_fd_sc_hd__clkbuf_1 _2102_ (.A(_1600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0278_));
 sky130_fd_sc_hd__and4_2 _2103_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[0].puf_buffer.cnt_1.ctr[6] ),
    .C(_1559_),
    .D(_1561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1601_));
 sky130_fd_sc_hd__a31o_1 _2104_ (.A1(_1601_),
    .A2(_1581_),
    .A3(_1582_),
    .B1(_0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1602_));
 sky130_fd_sc_hd__o21ba_1 _2105_ (.A1(net44),
    .A2(_1598_),
    .B1_N(_1602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0279_));
 sky130_fd_sc_hd__a31o_1 _2106_ (.A1(_1601_),
    .A2(_1565_),
    .A3(_1576_),
    .B1(\genblk1[0].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1603_));
 sky130_fd_sc_hd__nand4_1 _2107_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[10] ),
    .B(_1601_),
    .C(_1581_),
    .D(_1582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1604_));
 sky130_fd_sc_hd__and3_1 _2108_ (.A(_0638_),
    .B(_1603_),
    .C(_1604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1605_));
 sky130_fd_sc_hd__clkbuf_1 _2109_ (.A(_1605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0280_));
 sky130_fd_sc_hd__inv_2 _2110_ (.A(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1606_));
 sky130_fd_sc_hd__and2_1 _2111_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[11] ),
    .B(\genblk1[0].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1607_));
 sky130_fd_sc_hd__and4_1 _2112_ (.A(_1607_),
    .B(_1601_),
    .C(_1581_),
    .D(_1582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1608_));
 sky130_fd_sc_hd__a211oi_1 _2113_ (.A1(_1606_),
    .A2(_1604_),
    .B1(_1608_),
    .C1(_0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0281_));
 sky130_fd_sc_hd__a41o_1 _2114_ (.A1(_1557_),
    .A2(_1601_),
    .A3(_1581_),
    .A4(_1582_),
    .B1(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1609_));
 sky130_fd_sc_hd__o21ba_1 _2115_ (.A1(net61),
    .A2(_1608_),
    .B1_N(_1609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0282_));
 sky130_fd_sc_hd__and4_1 _2116_ (.A(_1557_),
    .B(_1601_),
    .C(_1581_),
    .D(_1582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1610_));
 sky130_fd_sc_hd__nand4_1 _2117_ (.A(_1558_),
    .B(_1601_),
    .C(_1581_),
    .D(_1582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1611_));
 sky130_fd_sc_hd__o211a_1 _2118_ (.A1(net135),
    .A2(_1610_),
    .B1(_1611_),
    .C1(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0283_));
 sky130_fd_sc_hd__inv_2 _2119_ (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1612_));
 sky130_fd_sc_hd__and3_1 _2120_ (.A(_1563_),
    .B(_1581_),
    .C(_1582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1613_));
 sky130_fd_sc_hd__a211oi_1 _2121_ (.A1(_1612_),
    .A2(_1611_),
    .B1(_1613_),
    .C1(_0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0284_));
 sky130_fd_sc_hd__a31o_1 _2122_ (.A1(_1563_),
    .A2(_1565_),
    .A3(_1576_),
    .B1(\genblk1[0].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1614_));
 sky130_fd_sc_hd__nand4_1 _2123_ (.A(\genblk1[0].puf_buffer.cnt_1.ctr[15] ),
    .B(_1563_),
    .C(_1581_),
    .D(_1582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1615_));
 sky130_fd_sc_hd__and3_1 _2124_ (.A(_0638_),
    .B(_1614_),
    .C(_1615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1616_));
 sky130_fd_sc_hd__clkbuf_1 _2125_ (.A(_1616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0285_));
 sky130_fd_sc_hd__inv_2 _2126_ (.A(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1617_));
 sky130_fd_sc_hd__o21bai_1 _2127_ (.A1(_1617_),
    .A2(_0035_),
    .B1_N(\genblk1[1].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0286_));
 sky130_fd_sc_hd__buf_2 _2128_ (.A(ena),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0288_));
 sky130_fd_sc_hd__clkbuf_2 _2129_ (.A(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0289_));
 sky130_fd_sc_hd__and2_1 _2130_ (.A(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0290_));
 sky130_fd_sc_hd__clkbuf_1 _2131_ (.A(_0290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2132_ (.A(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _2133_ (.A(_0291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2134_ (.A(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_1 _2135_ (.A(_0292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2136_ (.A(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0293_));
 sky130_fd_sc_hd__clkbuf_1 _2137_ (.A(_0293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2138_ (.A(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_1 _2139_ (.A(_0294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2140_ (.A(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_1 _2141_ (.A(_0295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2142_ (.A(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0296_));
 sky130_fd_sc_hd__clkbuf_1 _2143_ (.A(_0296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2144_ (.A(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0297_));
 sky130_fd_sc_hd__clkbuf_1 _2145_ (.A(_0297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2146_ (.A(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_1 _2147_ (.A(_0298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2148_ (.A(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .B(_0289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _2149_ (.A(_0299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2150_ (.A(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0300_));
 sky130_fd_sc_hd__and2_1 _2151_ (.A(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _2152_ (.A(_0301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2153_ (.A(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0302_));
 sky130_fd_sc_hd__clkbuf_1 _2154_ (.A(_0302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2155_ (.A(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_1 _2156_ (.A(_0303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2157_ (.A(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_1 _2158_ (.A(_0304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2159_ (.A(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_1 _2160_ (.A(_0305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2161_ (.A(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_1 _2162_ (.A(_0306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2163_ (.A(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0307_));
 sky130_fd_sc_hd__clkbuf_1 _2164_ (.A(_0307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2165_ (.A(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_1 _2166_ (.A(_0308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2167_ (.A(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_1 _2168_ (.A(_0309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2169_ (.A(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .B(_0300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _2170_ (.A(_0310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2171_ (.A(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0311_));
 sky130_fd_sc_hd__and2_1 _2172_ (.A(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _2173_ (.A(_0312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2174_ (.A(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _2175_ (.A(_0313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2176_ (.A(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _2177_ (.A(_0314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2178_ (.A(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_1 _2179_ (.A(_0315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2180_ (.A(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_1 _2181_ (.A(_0316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2182_ (.A(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0317_));
 sky130_fd_sc_hd__clkbuf_1 _2183_ (.A(_0317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2184_ (.A(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0318_));
 sky130_fd_sc_hd__clkbuf_1 _2185_ (.A(_0318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2186_ (.A(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_1 _2187_ (.A(_0319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2188_ (.A(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_1 _2189_ (.A(_0320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2190_ (.A(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .B(_0311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _2191_ (.A(_0321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2192_ (.A(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0322_));
 sky130_fd_sc_hd__and2_1 _2193_ (.A(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_1 _2194_ (.A(_0323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2195_ (.A(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_1 _2196_ (.A(_0324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[0] ));
 sky130_fd_sc_hd__nor2_1 _2197_ (.A(\genblk1[2].puf_buffer.race_arb.marked_2 ),
    .B(\genblk1[2].puf_buffer.race_arb.marked_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0325_));
 sky130_fd_sc_hd__and3b_1 _2198_ (.A_N(\genblk1[2].puf_buffer.cnt_2.finish ),
    .B(_0325_),
    .C(\genblk1[2].puf_buffer.cnt_1.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _2199_ (.A(_0326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[2].puf_buffer.race_arb.win_1 ));
 sky130_fd_sc_hd__and2_1 _2200_ (.A(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_1 _2201_ (.A(_0327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2202_ (.A(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_1 _2203_ (.A(_0328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2204_ (.A(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _2205_ (.A(_0329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2206_ (.A(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_1 _2207_ (.A(_0330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2208_ (.A(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_1 _2209_ (.A(_0331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2210_ (.A(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_1 _2211_ (.A(_0332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2212_ (.A(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_1 _2213_ (.A(_0333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2214_ (.A(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .B(_0322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0334_));
 sky130_fd_sc_hd__clkbuf_1 _2215_ (.A(_0334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_4 _2216_ (.A(ena),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_2 _2217_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0336_));
 sky130_fd_sc_hd__and2_1 _2218_ (.A(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_1 _2219_ (.A(_0337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2220_ (.A(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_1 _2221_ (.A(_0338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2222_ (.A(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_1 _2223_ (.A(_0339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2224_ (.A(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _2225_ (.A(_0340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2226_ (.A(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _2227_ (.A(_0341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2228_ (.A(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0342_));
 sky130_fd_sc_hd__clkbuf_1 _2229_ (.A(_0342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2230_ (.A(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_1 _2231_ (.A(_0343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2232_ (.A(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _2233_ (.A(_0344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2234_ (.A(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _2235_ (.A(_0345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2236_ (.A(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .B(_0336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_1 _2237_ (.A(_0346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2238_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0347_));
 sky130_fd_sc_hd__and2_1 _2239_ (.A(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0348_));
 sky130_fd_sc_hd__clkbuf_1 _2240_ (.A(_0348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2241_ (.A(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0349_));
 sky130_fd_sc_hd__clkbuf_1 _2242_ (.A(_0349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2243_ (.A(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0350_));
 sky130_fd_sc_hd__clkbuf_1 _2244_ (.A(_0350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2245_ (.A(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _2246_ (.A(_0351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2247_ (.A(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_1 _2248_ (.A(_0352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2249_ (.A(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_1 _2250_ (.A(_0353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2251_ (.A(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _2252_ (.A(_0354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2253_ (.A(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _2254_ (.A(_0355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2255_ (.A(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_1 _2256_ (.A(_0356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2257_ (.A(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .B(_0347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _2258_ (.A(_0357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[0] ));
 sky130_fd_sc_hd__buf_2 _2259_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0358_));
 sky130_fd_sc_hd__and2_1 _2260_ (.A(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .B(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _2261_ (.A(_0359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2262_ (.A(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .B(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _2263_ (.A(_0360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2264_ (.A(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .B(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_1 _2265_ (.A(_0361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2266_ (.A(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _2267_ (.A(_0362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[0] ));
 sky130_fd_sc_hd__nor2_1 _2268_ (.A(\genblk1[3].puf_buffer.race_arb.marked_2 ),
    .B(\genblk1[3].puf_buffer.race_arb.marked_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0363_));
 sky130_fd_sc_hd__and3b_1 _2269_ (.A_N(\genblk1[3].puf_buffer.cnt_2.finish ),
    .B(_0363_),
    .C(\genblk1[3].puf_buffer.cnt_1.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_1 _2270_ (.A(_0364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[3].puf_buffer.race_arb.win_1 ));
 sky130_fd_sc_hd__and2_1 _2271_ (.A(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .B(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _2272_ (.A(_0365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2273_ (.A(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .B(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _2274_ (.A(_0366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2275_ (.A(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .B(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0367_));
 sky130_fd_sc_hd__clkbuf_1 _2276_ (.A(_0367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2277_ (.A(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .B(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_1 _2278_ (.A(_0368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2279_ (.A(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .B(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _2280_ (.A(_0369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2281_ (.A(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .B(_0358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_1 _2282_ (.A(_0370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2283_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0371_));
 sky130_fd_sc_hd__and2_1 _2284_ (.A(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0372_));
 sky130_fd_sc_hd__clkbuf_1 _2285_ (.A(_0372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2286_ (.A(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0373_));
 sky130_fd_sc_hd__clkbuf_1 _2287_ (.A(_0373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2288_ (.A(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _2289_ (.A(_0374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2290_ (.A(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _2291_ (.A(_0375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2292_ (.A(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _2293_ (.A(_0376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2294_ (.A(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _2295_ (.A(_0377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2296_ (.A(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _2297_ (.A(_0378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2298_ (.A(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_1 _2299_ (.A(_0379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2300_ (.A(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _2301_ (.A(_0380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2302_ (.A(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_1 _2303_ (.A(_0381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2304_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0382_));
 sky130_fd_sc_hd__and2_1 _2305_ (.A(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .B(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_1 _2306_ (.A(_0383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2307_ (.A(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .B(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_1 _2308_ (.A(_0384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2309_ (.A(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .B(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_1 _2310_ (.A(_0385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2311_ (.A(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .B(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_1 _2312_ (.A(_0386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2313_ (.A(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .B(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_1 _2314_ (.A(_0387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2315_ (.A(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .B(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_1 _2316_ (.A(_0388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2317_ (.A(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .B(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_1 _2318_ (.A(_0389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2319_ (.A(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .B(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _2320_ (.A(_0390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2321_ (.A(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .B(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_1 _2322_ (.A(_0391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2323_ (.A(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .B(_0382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_1 _2324_ (.A(_0392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2325_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0393_));
 sky130_fd_sc_hd__and2_1 _2326_ (.A(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .B(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _2327_ (.A(_0394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2328_ (.A(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .B(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _2329_ (.A(_0395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2330_ (.A(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .B(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _2331_ (.A(_0396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2332_ (.A(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .B(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_1 _2333_ (.A(_0397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2334_ (.A(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .B(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_1 _2335_ (.A(_0398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2336_ (.A(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_1 _2337_ (.A(_0399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[0] ));
 sky130_fd_sc_hd__nor2_1 _2338_ (.A(\genblk1[4].puf_buffer.race_arb.marked_2 ),
    .B(\genblk1[4].puf_buffer.race_arb.marked_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0400_));
 sky130_fd_sc_hd__and3b_1 _2339_ (.A_N(\genblk1[4].puf_buffer.cnt_2.finish ),
    .B(_0400_),
    .C(\genblk1[4].puf_buffer.cnt_1.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _2340_ (.A(_0401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[4].puf_buffer.race_arb.win_1 ));
 sky130_fd_sc_hd__and2_1 _2341_ (.A(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .B(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_1 _2342_ (.A(_0402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2343_ (.A(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .B(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_1 _2344_ (.A(_0403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2345_ (.A(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .B(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_1 _2346_ (.A(_0404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2347_ (.A(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .B(_0393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _2348_ (.A(_0405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2349_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0406_));
 sky130_fd_sc_hd__and2_1 _2350_ (.A(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .B(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_1 _2351_ (.A(_0407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2352_ (.A(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .B(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0408_));
 sky130_fd_sc_hd__clkbuf_1 _2353_ (.A(_0408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2354_ (.A(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .B(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_1 _2355_ (.A(_0409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2356_ (.A(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .B(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_1 _2357_ (.A(_0410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2358_ (.A(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .B(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _2359_ (.A(_0411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2360_ (.A(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .B(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_1 _2361_ (.A(_0412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2362_ (.A(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .B(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_1 _2363_ (.A(_0413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2364_ (.A(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .B(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _2365_ (.A(_0414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2366_ (.A(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .B(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _2367_ (.A(_0415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2368_ (.A(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .B(_0406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _2369_ (.A(_0416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2370_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0417_));
 sky130_fd_sc_hd__and2_1 _2371_ (.A(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _2372_ (.A(_0418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2373_ (.A(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_1 _2374_ (.A(_0419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2375_ (.A(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_1 _2376_ (.A(_0420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2377_ (.A(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _2378_ (.A(_0421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2379_ (.A(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _2380_ (.A(_0422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2381_ (.A(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _2382_ (.A(_0423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2383_ (.A(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_1 _2384_ (.A(_0424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2385_ (.A(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_1 _2386_ (.A(_0425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2387_ (.A(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_1 _2388_ (.A(_0426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2389_ (.A(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .B(_0417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_1 _2390_ (.A(_0427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2391_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0428_));
 sky130_fd_sc_hd__and2_1 _2392_ (.A(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0429_));
 sky130_fd_sc_hd__clkbuf_1 _2393_ (.A(_0429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2394_ (.A(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0430_));
 sky130_fd_sc_hd__clkbuf_1 _2395_ (.A(_0430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2396_ (.A(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _2397_ (.A(_0431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2398_ (.A(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _2399_ (.A(_0432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2400_ (.A(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _2401_ (.A(_0433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2402_ (.A(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_1 _2403_ (.A(_0434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2404_ (.A(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_1 _2405_ (.A(_0435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2406_ (.A(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _2407_ (.A(_0436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[0] ));
 sky130_fd_sc_hd__nor2_1 _2408_ (.A(\genblk1[5].puf_buffer.race_arb.marked_2 ),
    .B(\genblk1[5].puf_buffer.race_arb.marked_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0437_));
 sky130_fd_sc_hd__and3b_1 _2409_ (.A_N(\genblk1[5].puf_buffer.cnt_2.finish ),
    .B(_0437_),
    .C(\genblk1[5].puf_buffer.cnt_1.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _2410_ (.A(_0438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[5].puf_buffer.race_arb.win_1 ));
 sky130_fd_sc_hd__and2_1 _2411_ (.A(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_1 _2412_ (.A(_0439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2413_ (.A(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .B(_0428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_1 _2414_ (.A(_0440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2415_ (.A(_0335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0441_));
 sky130_fd_sc_hd__and2_1 _2416_ (.A(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .B(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _2417_ (.A(_0442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2418_ (.A(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .B(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _2419_ (.A(_0443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2420_ (.A(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .B(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_1 _2421_ (.A(_0444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2422_ (.A(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .B(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _2423_ (.A(_0445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2424_ (.A(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .B(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _2425_ (.A(_0446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2426_ (.A(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .B(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _2427_ (.A(_0447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2428_ (.A(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .B(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _2429_ (.A(_0448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2430_ (.A(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .B(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _2431_ (.A(_0449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2432_ (.A(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .B(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _2433_ (.A(_0450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2434_ (.A(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .B(_0441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _2435_ (.A(_0451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[0] ));
 sky130_fd_sc_hd__buf_2 _2436_ (.A(ena),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0452_));
 sky130_fd_sc_hd__buf_2 _2437_ (.A(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0453_));
 sky130_fd_sc_hd__and2_1 _2438_ (.A(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _2439_ (.A(_0454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2440_ (.A(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_1 _2441_ (.A(_0455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2442_ (.A(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _2443_ (.A(_0456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2444_ (.A(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _2445_ (.A(_0457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2446_ (.A(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _2447_ (.A(_0458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2448_ (.A(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0459_));
 sky130_fd_sc_hd__clkbuf_1 _2449_ (.A(_0459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2450_ (.A(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _2451_ (.A(_0460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2452_ (.A(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _2453_ (.A(_0461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2454_ (.A(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_1 _2455_ (.A(_0462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2456_ (.A(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .B(_0453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_1 _2457_ (.A(_0463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2458_ (.A(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0464_));
 sky130_fd_sc_hd__and2_1 _2459_ (.A(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .B(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _2460_ (.A(_0465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2461_ (.A(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .B(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _2462_ (.A(_0466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2463_ (.A(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .B(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_1 _2464_ (.A(_0467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2465_ (.A(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .B(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_1 _2466_ (.A(_0468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2467_ (.A(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .B(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_1 _2468_ (.A(_0469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2469_ (.A(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .B(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0470_));
 sky130_fd_sc_hd__clkbuf_1 _2470_ (.A(_0470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2471_ (.A(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .B(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_1 _2472_ (.A(_0471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2473_ (.A(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .B(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _2474_ (.A(_0472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2475_ (.A(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .B(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_1 _2476_ (.A(_0473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2477_ (.A(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_1 _2478_ (.A(_0474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[0] ));
 sky130_fd_sc_hd__nor2_1 _2479_ (.A(\genblk1[6].puf_buffer.race_arb.marked_2 ),
    .B(\genblk1[6].puf_buffer.race_arb.marked_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0475_));
 sky130_fd_sc_hd__and3b_1 _2480_ (.A_N(\genblk1[6].puf_buffer.cnt_2.finish ),
    .B(_0475_),
    .C(\genblk1[6].puf_buffer.cnt_1.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_1 _2481_ (.A(_0476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[6].puf_buffer.race_arb.win_1 ));
 sky130_fd_sc_hd__clkbuf_2 _2482_ (.A(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0477_));
 sky130_fd_sc_hd__and2_1 _2483_ (.A(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .B(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _2484_ (.A(_0478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2485_ (.A(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .B(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_1 _2486_ (.A(_0479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2487_ (.A(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .B(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0480_));
 sky130_fd_sc_hd__clkbuf_1 _2488_ (.A(_0480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2489_ (.A(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .B(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0481_));
 sky130_fd_sc_hd__clkbuf_1 _2490_ (.A(_0481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2491_ (.A(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .B(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0482_));
 sky130_fd_sc_hd__clkbuf_1 _2492_ (.A(_0482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2493_ (.A(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .B(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0483_));
 sky130_fd_sc_hd__clkbuf_1 _2494_ (.A(_0483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2495_ (.A(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .B(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0484_));
 sky130_fd_sc_hd__clkbuf_1 _2496_ (.A(_0484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2497_ (.A(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .B(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_1 _2498_ (.A(_0485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2499_ (.A(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .B(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_1 _2500_ (.A(_0486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2501_ (.A(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .B(_0477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_1 _2502_ (.A(_0487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2503_ (.A(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0488_));
 sky130_fd_sc_hd__and2_1 _2504_ (.A(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .B(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0489_));
 sky130_fd_sc_hd__clkbuf_1 _2505_ (.A(_0489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2506_ (.A(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .B(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_1 _2507_ (.A(_0490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2508_ (.A(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .B(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0491_));
 sky130_fd_sc_hd__clkbuf_1 _2509_ (.A(_0491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2510_ (.A(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .B(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0492_));
 sky130_fd_sc_hd__clkbuf_1 _2511_ (.A(_0492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2512_ (.A(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .B(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0493_));
 sky130_fd_sc_hd__clkbuf_1 _2513_ (.A(_0493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2514_ (.A(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0494_));
 sky130_fd_sc_hd__clkbuf_1 _2515_ (.A(_0494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2516_ (.A(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .B(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _2517_ (.A(_0495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2518_ (.A(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .B(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0496_));
 sky130_fd_sc_hd__clkbuf_1 _2519_ (.A(_0496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2520_ (.A(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .B(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0497_));
 sky130_fd_sc_hd__clkbuf_1 _2521_ (.A(_0497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2522_ (.A(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .B(_0488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0498_));
 sky130_fd_sc_hd__clkbuf_1 _2523_ (.A(_0498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2524_ (.A(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0499_));
 sky130_fd_sc_hd__and2_1 _2525_ (.A(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .B(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0500_));
 sky130_fd_sc_hd__clkbuf_1 _2526_ (.A(_0500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2527_ (.A(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .B(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_1 _2528_ (.A(_0501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2529_ (.A(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .B(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0502_));
 sky130_fd_sc_hd__clkbuf_1 _2530_ (.A(_0502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2531_ (.A(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .B(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0503_));
 sky130_fd_sc_hd__clkbuf_1 _2532_ (.A(_0503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2533_ (.A(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .B(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0504_));
 sky130_fd_sc_hd__clkbuf_1 _2534_ (.A(_0504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2535_ (.A(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .B(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_1 _2536_ (.A(_0505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2537_ (.A(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .B(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0506_));
 sky130_fd_sc_hd__clkbuf_1 _2538_ (.A(_0506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2539_ (.A(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .B(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0507_));
 sky130_fd_sc_hd__clkbuf_1 _2540_ (.A(_0507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2541_ (.A(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .B(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0508_));
 sky130_fd_sc_hd__clkbuf_1 _2542_ (.A(_0508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2543_ (.A(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .B(_0499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_1 _2544_ (.A(_0509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2545_ (.A(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0510_));
 sky130_fd_sc_hd__and2_1 _2546_ (.A(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .B(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0511_));
 sky130_fd_sc_hd__clkbuf_1 _2547_ (.A(_0511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2548_ (.A(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_1 _2549_ (.A(_0512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[0] ));
 sky130_fd_sc_hd__nor2_1 _2550_ (.A(\genblk1[7].puf_buffer.race_arb.marked_2 ),
    .B(\genblk1[7].puf_buffer.race_arb.marked_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0513_));
 sky130_fd_sc_hd__and3b_1 _2551_ (.A_N(\genblk1[7].puf_buffer.cnt_2.finish ),
    .B(_0513_),
    .C(\genblk1[7].puf_buffer.cnt_1.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_1 _2552_ (.A(_0514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[7].puf_buffer.race_arb.win_1 ));
 sky130_fd_sc_hd__and2_1 _2553_ (.A(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .B(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0515_));
 sky130_fd_sc_hd__clkbuf_1 _2554_ (.A(_0515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2555_ (.A(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .B(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_1 _2556_ (.A(_0516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2557_ (.A(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .B(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0517_));
 sky130_fd_sc_hd__clkbuf_1 _2558_ (.A(_0517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2559_ (.A(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .B(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _2560_ (.A(_0518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2561_ (.A(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .B(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0519_));
 sky130_fd_sc_hd__clkbuf_1 _2562_ (.A(_0519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2563_ (.A(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .B(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0520_));
 sky130_fd_sc_hd__clkbuf_1 _2564_ (.A(_0520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2565_ (.A(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .B(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0521_));
 sky130_fd_sc_hd__clkbuf_1 _2566_ (.A(_0521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2567_ (.A(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .B(_0510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0522_));
 sky130_fd_sc_hd__clkbuf_1 _2568_ (.A(_0522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2569_ (.A(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0523_));
 sky130_fd_sc_hd__and2_1 _2570_ (.A(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .B(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0524_));
 sky130_fd_sc_hd__clkbuf_1 _2571_ (.A(_0524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2572_ (.A(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .B(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0525_));
 sky130_fd_sc_hd__clkbuf_1 _2573_ (.A(_0525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2574_ (.A(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .B(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_1 _2575_ (.A(_0526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2576_ (.A(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .B(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_1 _2577_ (.A(_0527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2578_ (.A(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .B(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0528_));
 sky130_fd_sc_hd__clkbuf_1 _2579_ (.A(_0528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2580_ (.A(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .B(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0529_));
 sky130_fd_sc_hd__clkbuf_1 _2581_ (.A(_0529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2582_ (.A(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .B(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_1 _2583_ (.A(_0530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2584_ (.A(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0531_));
 sky130_fd_sc_hd__clkbuf_1 _2585_ (.A(_0531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2586_ (.A(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .B(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_1 _2587_ (.A(_0532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2588_ (.A(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .B(_0523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0533_));
 sky130_fd_sc_hd__clkbuf_1 _2589_ (.A(_0533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2590_ (.A(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0534_));
 sky130_fd_sc_hd__and2_1 _2591_ (.A(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .B(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0535_));
 sky130_fd_sc_hd__clkbuf_1 _2592_ (.A(_0535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2593_ (.A(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .B(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_1 _2594_ (.A(_0536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2595_ (.A(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .B(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0537_));
 sky130_fd_sc_hd__clkbuf_1 _2596_ (.A(_0537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2597_ (.A(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .B(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0538_));
 sky130_fd_sc_hd__clkbuf_1 _2598_ (.A(_0538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2599_ (.A(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .B(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_1 _2600_ (.A(_0539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2601_ (.A(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .B(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0540_));
 sky130_fd_sc_hd__clkbuf_1 _2602_ (.A(_0540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2603_ (.A(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .B(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0541_));
 sky130_fd_sc_hd__clkbuf_1 _2604_ (.A(_0541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2605_ (.A(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .B(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0542_));
 sky130_fd_sc_hd__clkbuf_1 _2606_ (.A(_0542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2607_ (.A(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .B(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0543_));
 sky130_fd_sc_hd__clkbuf_1 _2608_ (.A(_0543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2609_ (.A(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .B(_0534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0544_));
 sky130_fd_sc_hd__clkbuf_1 _2610_ (.A(_0544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2611_ (.A(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0545_));
 sky130_fd_sc_hd__and2_1 _2612_ (.A(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .B(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0546_));
 sky130_fd_sc_hd__clkbuf_1 _2613_ (.A(_0546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2614_ (.A(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .B(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0547_));
 sky130_fd_sc_hd__clkbuf_1 _2615_ (.A(_0547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2616_ (.A(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .B(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0548_));
 sky130_fd_sc_hd__clkbuf_1 _2617_ (.A(_0548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2618_ (.A(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0549_));
 sky130_fd_sc_hd__clkbuf_1 _2619_ (.A(_0549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[0] ));
 sky130_fd_sc_hd__nor2_1 _2620_ (.A(\genblk1[0].puf_buffer.race_arb.marked_2 ),
    .B(\genblk1[0].puf_buffer.race_arb.marked_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0550_));
 sky130_fd_sc_hd__and3b_1 _2621_ (.A_N(\genblk1[0].puf_buffer.cnt_2.finish ),
    .B(_0550_),
    .C(\genblk1[0].puf_buffer.cnt_1.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0551_));
 sky130_fd_sc_hd__clkbuf_1 _2622_ (.A(_0551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[0].puf_buffer.race_arb.win_1 ));
 sky130_fd_sc_hd__and2_1 _2623_ (.A(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .B(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0552_));
 sky130_fd_sc_hd__clkbuf_1 _2624_ (.A(_0552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2625_ (.A(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .B(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0553_));
 sky130_fd_sc_hd__clkbuf_1 _2626_ (.A(_0553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2627_ (.A(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .B(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_1 _2628_ (.A(_0554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2629_ (.A(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .B(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0555_));
 sky130_fd_sc_hd__clkbuf_1 _2630_ (.A(_0555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2631_ (.A(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .B(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0556_));
 sky130_fd_sc_hd__clkbuf_1 _2632_ (.A(_0556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2633_ (.A(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .B(_0545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0557_));
 sky130_fd_sc_hd__clkbuf_1 _2634_ (.A(_0557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2635_ (.A(_0452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0558_));
 sky130_fd_sc_hd__and2_1 _2636_ (.A(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .B(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0559_));
 sky130_fd_sc_hd__clkbuf_1 _2637_ (.A(_0559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2638_ (.A(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .B(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0560_));
 sky130_fd_sc_hd__clkbuf_1 _2639_ (.A(_0560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2640_ (.A(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .B(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0561_));
 sky130_fd_sc_hd__clkbuf_1 _2641_ (.A(_0561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2642_ (.A(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .B(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0562_));
 sky130_fd_sc_hd__clkbuf_1 _2643_ (.A(_0562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2644_ (.A(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .B(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0563_));
 sky130_fd_sc_hd__clkbuf_1 _2645_ (.A(_0563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2646_ (.A(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .B(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0564_));
 sky130_fd_sc_hd__clkbuf_1 _2647_ (.A(_0564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2648_ (.A(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .B(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_1 _2649_ (.A(_0565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2650_ (.A(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .B(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0566_));
 sky130_fd_sc_hd__clkbuf_1 _2651_ (.A(_0566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2652_ (.A(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .B(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0567_));
 sky130_fd_sc_hd__clkbuf_1 _2653_ (.A(_0567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2654_ (.A(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0568_));
 sky130_fd_sc_hd__clkbuf_1 _2655_ (.A(_0568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[0] ));
 sky130_fd_sc_hd__clkbuf_2 _2656_ (.A(ena),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0569_));
 sky130_fd_sc_hd__and2_1 _2657_ (.A(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .B(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0570_));
 sky130_fd_sc_hd__clkbuf_1 _2658_ (.A(_0570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2659_ (.A(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .B(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_1 _2660_ (.A(_0571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2661_ (.A(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .B(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_1 _2662_ (.A(_0572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2663_ (.A(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .B(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0573_));
 sky130_fd_sc_hd__clkbuf_1 _2664_ (.A(_0573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2665_ (.A(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .B(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0574_));
 sky130_fd_sc_hd__clkbuf_1 _2666_ (.A(_0574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2667_ (.A(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .B(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0575_));
 sky130_fd_sc_hd__clkbuf_1 _2668_ (.A(_0575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2669_ (.A(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .B(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0576_));
 sky130_fd_sc_hd__clkbuf_1 _2670_ (.A(_0576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2671_ (.A(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .B(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_1 _2672_ (.A(_0577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2673_ (.A(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .B(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0578_));
 sky130_fd_sc_hd__clkbuf_1 _2674_ (.A(_0578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2675_ (.A(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .B(_0569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0579_));
 sky130_fd_sc_hd__clkbuf_1 _2676_ (.A(_0579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2677_ (.A(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .B(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0580_));
 sky130_fd_sc_hd__clkbuf_1 _2678_ (.A(_0580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2679_ (.A(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .B(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0581_));
 sky130_fd_sc_hd__clkbuf_1 _2680_ (.A(_0581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2681_ (.A(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .B(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0582_));
 sky130_fd_sc_hd__clkbuf_1 _2682_ (.A(_0582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2683_ (.A(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .B(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0583_));
 sky130_fd_sc_hd__clkbuf_1 _2684_ (.A(_0583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2685_ (.A(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .B(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0584_));
 sky130_fd_sc_hd__clkbuf_1 _2686_ (.A(_0584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[0] ));
 sky130_fd_sc_hd__and2_1 _2687_ (.A(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0585_));
 sky130_fd_sc_hd__clkbuf_1 _2688_ (.A(_0585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[0] ));
 sky130_fd_sc_hd__nor2_1 _2689_ (.A(\genblk1[1].puf_buffer.race_arb.marked_2 ),
    .B(\genblk1[1].puf_buffer.race_arb.marked_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0586_));
 sky130_fd_sc_hd__and3b_1 _2690_ (.A_N(\genblk1[1].puf_buffer.cnt_2.finish ),
    .B(_0586_),
    .C(\genblk1[1].puf_buffer.cnt_1.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_1 _2691_ (.A(_0587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\genblk1[1].puf_buffer.race_arb.win_1 ));
 sky130_fd_sc_hd__clkbuf_2 _2692_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0588_));
 sky130_fd_sc_hd__clkbuf_4 _2693_ (.A(_0588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0589_));
 sky130_fd_sc_hd__and4_1 _2694_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[3] ),
    .B(\genblk1[1].puf_buffer.cnt_2.ctr[2] ),
    .C(\genblk1[1].puf_buffer.cnt_2.ctr[1] ),
    .D(\genblk1[1].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0590_));
 sky130_fd_sc_hd__and2_1 _2695_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[1].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0591_));
 sky130_fd_sc_hd__and4_1 _2696_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[1].puf_buffer.cnt_2.ctr[4] ),
    .C(_0590_),
    .D(_0591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0592_));
 sky130_fd_sc_hd__and3_1 _2697_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[9] ),
    .B(\genblk1[1].puf_buffer.cnt_2.ctr[8] ),
    .C(_0592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0593_));
 sky130_fd_sc_hd__and3_1 _2698_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[12] ),
    .B(\genblk1[1].puf_buffer.cnt_2.ctr[11] ),
    .C(\genblk1[1].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0594_));
 sky130_fd_sc_hd__and2_1 _2699_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[13] ),
    .B(_0594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0595_));
 sky130_fd_sc_hd__and3_1 _2700_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[14] ),
    .B(_0593_),
    .C(_0595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0596_));
 sky130_fd_sc_hd__a22o_1 _2701_ (.A1(_0589_),
    .A2(\genblk1[1].puf_buffer.cnt_2.finish ),
    .B1(_0596_),
    .B2(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0000_));
 sky130_fd_sc_hd__clkbuf_2 _2702_ (.A(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0597_));
 sky130_fd_sc_hd__buf_2 _2703_ (.A(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0598_));
 sky130_fd_sc_hd__buf_2 _2704_ (.A(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0599_));
 sky130_fd_sc_hd__buf_2 _2705_ (.A(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0600_));
 sky130_fd_sc_hd__or4_4 _2706_ (.A(_0597_),
    .B(_0598_),
    .C(_0599_),
    .D(_0600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0601_));
 sky130_fd_sc_hd__or2_2 _2707_ (.A(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0602_));
 sky130_fd_sc_hd__and4bb_4 _2708_ (.A_N(_0599_),
    .B_N(_0600_),
    .C(_0597_),
    .D(_0598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0603_));
 sky130_fd_sc_hd__and4b_4 _2709_ (.A_N(_0599_),
    .B(_0600_),
    .C(_0597_),
    .D(_0598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0604_));
 sky130_fd_sc_hd__and4bb_4 _2710_ (.A_N(_0597_),
    .B_N(_0599_),
    .C(net6),
    .D(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0605_));
 sky130_fd_sc_hd__nor4b_4 _2711_ (.A(_0598_),
    .B(_0599_),
    .C(_0600_),
    .D_N(_0597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0606_));
 sky130_fd_sc_hd__a22o_1 _2712_ (.A1(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .A2(_0605_),
    .B1(net22),
    .B2(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0607_));
 sky130_fd_sc_hd__a221o_1 _2713_ (.A1(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .A2(_0603_),
    .B1(_0604_),
    .B2(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .C1(_0607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0608_));
 sky130_fd_sc_hd__nor4b_1 _2714_ (.A(net8),
    .B(net9),
    .C(net7),
    .D_N(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0609_));
 sky130_fd_sc_hd__and4bb_4 _2715_ (.A_N(net8),
    .B_N(net9),
    .C(net7),
    .D(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0610_));
 sky130_fd_sc_hd__and4b_4 _2716_ (.A_N(net9),
    .B(net7),
    .C(net6),
    .D(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0611_));
 sky130_fd_sc_hd__a22o_1 _2717_ (.A1(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .A2(_0610_),
    .B1(_0611_),
    .B2(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0612_));
 sky130_fd_sc_hd__nor4_1 _2718_ (.A(_0597_),
    .B(_0598_),
    .C(_0599_),
    .D(_0600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0613_));
 sky130_fd_sc_hd__a211o_1 _2719_ (.A1(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .A2(net25),
    .B1(_0612_),
    .C1(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0614_));
 sky130_fd_sc_hd__and4b_4 _2720_ (.A_N(net6),
    .B(net7),
    .C(net9),
    .D(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0615_));
 sky130_fd_sc_hd__nor4b_2 _2721_ (.A(_0597_),
    .B(_0598_),
    .C(_0600_),
    .D_N(net7),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0616_));
 sky130_fd_sc_hd__a22o_1 _2722_ (.A1(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .A2(_0615_),
    .B1(net18),
    .B2(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0617_));
 sky130_fd_sc_hd__and4_4 _2723_ (.A(_0597_),
    .B(_0598_),
    .C(_0599_),
    .D(_0600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0618_));
 sky130_fd_sc_hd__nor4b_2 _2724_ (.A(_0597_),
    .B(_0599_),
    .C(_0600_),
    .D_N(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0619_));
 sky130_fd_sc_hd__a22o_1 _2725_ (.A1(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .A2(_0618_),
    .B1(net16),
    .B2(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0620_));
 sky130_fd_sc_hd__and4b_4 _2726_ (.A_N(_0597_),
    .B(_0598_),
    .C(_0599_),
    .D(_0600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0621_));
 sky130_fd_sc_hd__and4bb_4 _2727_ (.A_N(_0598_),
    .B_N(_0600_),
    .C(net7),
    .D(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0622_));
 sky130_fd_sc_hd__a22o_1 _2728_ (.A1(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .A2(_0621_),
    .B1(_0622_),
    .B2(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0623_));
 sky130_fd_sc_hd__and4bb_4 _2729_ (.A_N(net8),
    .B_N(net6),
    .C(net7),
    .D(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0624_));
 sky130_fd_sc_hd__and4bb_4 _2730_ (.A_N(_0598_),
    .B_N(_0599_),
    .C(net6),
    .D(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0625_));
 sky130_fd_sc_hd__a22o_1 _2731_ (.A1(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .A2(_0624_),
    .B1(_0625_),
    .B2(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0626_));
 sky130_fd_sc_hd__or4_1 _2732_ (.A(_0617_),
    .B(_0620_),
    .C(_0623_),
    .D(_0626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0627_));
 sky130_fd_sc_hd__or3_4 _2733_ (.A(_0608_),
    .B(_0614_),
    .C(_0627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0628_));
 sky130_fd_sc_hd__and3_1 _2734_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[0] ),
    .B(_0602_),
    .C(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0629_));
 sky130_fd_sc_hd__clkbuf_4 _2735_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0630_));
 sky130_fd_sc_hd__buf_2 _2736_ (.A(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0631_));
 sky130_fd_sc_hd__buf_2 _2737_ (.A(_0602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0632_));
 sky130_fd_sc_hd__buf_2 _2738_ (.A(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0633_));
 sky130_fd_sc_hd__a21o_1 _2739_ (.A1(_0632_),
    .A2(_0633_),
    .B1(\genblk1[1].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0634_));
 sky130_fd_sc_hd__and3b_1 _2740_ (.A_N(_0629_),
    .B(_0631_),
    .C(_0634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0635_));
 sky130_fd_sc_hd__clkbuf_1 _2741_ (.A(_0635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0001_));
 sky130_fd_sc_hd__nand2_1 _2742_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[1] ),
    .B(\genblk1[1].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0636_));
 sky130_fd_sc_hd__nand2_2 _2743_ (.A(_0632_),
    .B(_0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0637_));
 sky130_fd_sc_hd__clkbuf_4 _2744_ (.A(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0638_));
 sky130_fd_sc_hd__clkbuf_4 _2745_ (.A(_0638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0639_));
 sky130_fd_sc_hd__o221a_1 _2746_ (.A1(_0636_),
    .A2(_0637_),
    .B1(_0629_),
    .B2(net203),
    .C1(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0002_));
 sky130_fd_sc_hd__inv_2 _2747_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0640_));
 sky130_fd_sc_hd__and4bb_1 _2748_ (.A_N(_0640_),
    .B_N(_0636_),
    .C(_0602_),
    .D(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0641_));
 sky130_fd_sc_hd__a41o_1 _2749_ (.A1(\genblk1[1].puf_buffer.cnt_2.ctr[1] ),
    .A2(\genblk1[1].puf_buffer.cnt_2.ctr[0] ),
    .A3(_0602_),
    .A4(_0628_),
    .B1(\genblk1[1].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0642_));
 sky130_fd_sc_hd__and3b_1 _2750_ (.A_N(_0641_),
    .B(_0631_),
    .C(_0642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0643_));
 sky130_fd_sc_hd__clkbuf_1 _2751_ (.A(_0643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0003_));
 sky130_fd_sc_hd__inv_2 _2752_ (.A(_0590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0644_));
 sky130_fd_sc_hd__o221a_1 _2753_ (.A1(_0644_),
    .A2(_0637_),
    .B1(_0641_),
    .B2(net123),
    .C1(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0004_));
 sky130_fd_sc_hd__and4_1 _2754_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[4] ),
    .B(_0590_),
    .C(_0602_),
    .D(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0645_));
 sky130_fd_sc_hd__a31o_1 _2755_ (.A1(_0590_),
    .A2(_0632_),
    .A3(_0633_),
    .B1(\genblk1[1].puf_buffer.cnt_2.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0646_));
 sky130_fd_sc_hd__and3b_1 _2756_ (.A_N(_0645_),
    .B(_0631_),
    .C(_0646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0647_));
 sky130_fd_sc_hd__clkbuf_1 _2757_ (.A(_0647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0005_));
 sky130_fd_sc_hd__and3_1 _2758_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[1].puf_buffer.cnt_2.ctr[4] ),
    .C(_0590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0648_));
 sky130_fd_sc_hd__inv_2 _2759_ (.A(_0648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0649_));
 sky130_fd_sc_hd__o221a_1 _2760_ (.A1(_0649_),
    .A2(_0637_),
    .B1(_0645_),
    .B2(net171),
    .C1(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0006_));
 sky130_fd_sc_hd__and4_1 _2761_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[6] ),
    .B(_0648_),
    .C(_0602_),
    .D(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0650_));
 sky130_fd_sc_hd__a31o_1 _2762_ (.A1(_0648_),
    .A2(_0632_),
    .A3(_0633_),
    .B1(\genblk1[1].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0651_));
 sky130_fd_sc_hd__and3b_1 _2763_ (.A_N(_0650_),
    .B(_0631_),
    .C(_0651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0652_));
 sky130_fd_sc_hd__clkbuf_1 _2764_ (.A(_0652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0007_));
 sky130_fd_sc_hd__inv_2 _2765_ (.A(_0592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0653_));
 sky130_fd_sc_hd__o221a_1 _2766_ (.A1(_0653_),
    .A2(_0637_),
    .B1(_0650_),
    .B2(net90),
    .C1(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0008_));
 sky130_fd_sc_hd__and4_1 _2767_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[8] ),
    .B(_0592_),
    .C(_0602_),
    .D(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0654_));
 sky130_fd_sc_hd__a31o_1 _2768_ (.A1(_0592_),
    .A2(_0632_),
    .A3(_0633_),
    .B1(\genblk1[1].puf_buffer.cnt_2.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0655_));
 sky130_fd_sc_hd__and3b_1 _2769_ (.A_N(_0654_),
    .B(_0631_),
    .C(_0655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0656_));
 sky130_fd_sc_hd__clkbuf_1 _2770_ (.A(_0656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0009_));
 sky130_fd_sc_hd__nand3_1 _2771_ (.A(_0593_),
    .B(_0632_),
    .C(_0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0657_));
 sky130_fd_sc_hd__clkbuf_4 _2772_ (.A(_0638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0658_));
 sky130_fd_sc_hd__o211a_1 _2773_ (.A1(net101),
    .A2(_0654_),
    .B1(_0657_),
    .C1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0010_));
 sky130_fd_sc_hd__and4_1 _2774_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[10] ),
    .B(_0593_),
    .C(_0602_),
    .D(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0659_));
 sky130_fd_sc_hd__a31o_1 _2775_ (.A1(_0593_),
    .A2(_0632_),
    .A3(_0633_),
    .B1(\genblk1[1].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0660_));
 sky130_fd_sc_hd__and3b_1 _2776_ (.A_N(_0659_),
    .B(_0631_),
    .C(_0660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0661_));
 sky130_fd_sc_hd__clkbuf_1 _2777_ (.A(_0661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0011_));
 sky130_fd_sc_hd__nand2_1 _2778_ (.A(net198),
    .B(\genblk1[1].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0662_));
 sky130_fd_sc_hd__o221a_1 _2779_ (.A1(_0662_),
    .A2(_0657_),
    .B1(_0659_),
    .B2(net198),
    .C1(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0012_));
 sky130_fd_sc_hd__inv_2 _2780_ (.A(_0594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0663_));
 sky130_fd_sc_hd__and2_1 _2781_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[11] ),
    .B(\genblk1[1].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0664_));
 sky130_fd_sc_hd__a41o_1 _2782_ (.A1(_0593_),
    .A2(_0664_),
    .A3(_0632_),
    .A4(_0633_),
    .B1(net209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0665_));
 sky130_fd_sc_hd__o211a_1 _2783_ (.A1(_0663_),
    .A2(_0657_),
    .B1(_0665_),
    .C1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0013_));
 sky130_fd_sc_hd__and4_1 _2784_ (.A(_0593_),
    .B(_0595_),
    .C(_0602_),
    .D(_0628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0666_));
 sky130_fd_sc_hd__a41o_1 _2785_ (.A1(_0593_),
    .A2(_0594_),
    .A3(_0602_),
    .A4(_0628_),
    .B1(\genblk1[1].puf_buffer.cnt_2.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0667_));
 sky130_fd_sc_hd__and3b_1 _2786_ (.A_N(_0666_),
    .B(_0631_),
    .C(_0667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0668_));
 sky130_fd_sc_hd__clkbuf_1 _2787_ (.A(_0668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0014_));
 sky130_fd_sc_hd__inv_2 _2788_ (.A(_0596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0669_));
 sky130_fd_sc_hd__o221a_1 _2789_ (.A1(_0669_),
    .A2(_0637_),
    .B1(_0666_),
    .B2(net75),
    .C1(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0015_));
 sky130_fd_sc_hd__clkbuf_4 _2790_ (.A(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0670_));
 sky130_fd_sc_hd__nand4_1 _2791_ (.A(\genblk1[1].puf_buffer.cnt_2.ctr[15] ),
    .B(_0596_),
    .C(_0632_),
    .D(_0633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0671_));
 sky130_fd_sc_hd__a31o_1 _2792_ (.A1(_0596_),
    .A2(_0632_),
    .A3(_0633_),
    .B1(\genblk1[1].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0672_));
 sky130_fd_sc_hd__and3_1 _2793_ (.A(_0670_),
    .B(_0671_),
    .C(_0672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_1 _2794_ (.A(_0673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0016_));
 sky130_fd_sc_hd__and4_1 _2795_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[3] ),
    .B(\genblk1[1].puf_buffer.cnt_1.ctr[2] ),
    .C(\genblk1[1].puf_buffer.cnt_1.ctr[1] ),
    .D(\genblk1[1].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0674_));
 sky130_fd_sc_hd__and2_1 _2796_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[1].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0675_));
 sky130_fd_sc_hd__and4_1 _2797_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[1].puf_buffer.cnt_1.ctr[4] ),
    .C(_0674_),
    .D(_0675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0676_));
 sky130_fd_sc_hd__and3_1 _2798_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[9] ),
    .B(\genblk1[1].puf_buffer.cnt_1.ctr[8] ),
    .C(_0676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0677_));
 sky130_fd_sc_hd__and3_1 _2799_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[12] ),
    .B(\genblk1[1].puf_buffer.cnt_1.ctr[11] ),
    .C(\genblk1[1].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0678_));
 sky130_fd_sc_hd__and2_1 _2800_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[13] ),
    .B(_0678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0679_));
 sky130_fd_sc_hd__and3_1 _2801_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[14] ),
    .B(_0677_),
    .C(_0679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0680_));
 sky130_fd_sc_hd__a22o_1 _2802_ (.A1(_0589_),
    .A2(net165),
    .B1(_0680_),
    .B2(\genblk1[1].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0017_));
 sky130_fd_sc_hd__buf_2 _2803_ (.A(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0681_));
 sky130_fd_sc_hd__buf_2 _2804_ (.A(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0682_));
 sky130_fd_sc_hd__buf_2 _2805_ (.A(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0683_));
 sky130_fd_sc_hd__buf_2 _2806_ (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0684_));
 sky130_fd_sc_hd__or4_4 _2807_ (.A(_0681_),
    .B(_0682_),
    .C(_0683_),
    .D(_0684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0685_));
 sky130_fd_sc_hd__or2_2 _2808_ (.A(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0686_));
 sky130_fd_sc_hd__and4bb_4 _2809_ (.A_N(net4),
    .B_N(net2),
    .C(net3),
    .D(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0687_));
 sky130_fd_sc_hd__nor4b_4 _2810_ (.A(_0681_),
    .B(_0682_),
    .C(_0683_),
    .D_N(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0688_));
 sky130_fd_sc_hd__and4bb_4 _2811_ (.A_N(net5),
    .B_N(net2),
    .C(net3),
    .D(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0689_));
 sky130_fd_sc_hd__and4b_4 _2812_ (.A_N(net3),
    .B(_0684_),
    .C(net4),
    .D(_0682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0690_));
 sky130_fd_sc_hd__a22o_1 _2813_ (.A1(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .A2(_0689_),
    .B1(_0690_),
    .B2(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0691_));
 sky130_fd_sc_hd__a221o_1 _2814_ (.A1(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .A2(_0687_),
    .B1(net15),
    .B2(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .C1(_0691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0692_));
 sky130_fd_sc_hd__nor4b_2 _2815_ (.A(_0681_),
    .B(_0683_),
    .C(_0684_),
    .D_N(_0682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0693_));
 sky130_fd_sc_hd__and4bb_4 _2816_ (.A_N(net5),
    .B_N(net3),
    .C(net2),
    .D(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0694_));
 sky130_fd_sc_hd__and4_4 _2817_ (.A(_0681_),
    .B(_0682_),
    .C(_0683_),
    .D(_0684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0695_));
 sky130_fd_sc_hd__a22o_1 _2818_ (.A1(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .A2(_0694_),
    .B1(_0695_),
    .B2(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0696_));
 sky130_fd_sc_hd__nor4_1 _2819_ (.A(net4),
    .B(_0682_),
    .C(_0683_),
    .D(_0684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0697_));
 sky130_fd_sc_hd__a211o_1 _2820_ (.A1(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .A2(net13),
    .B1(_0696_),
    .C1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0698_));
 sky130_fd_sc_hd__and4b_4 _2821_ (.A_N(_0684_),
    .B(_0683_),
    .C(_0682_),
    .D(_0681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0699_));
 sky130_fd_sc_hd__and4b_4 _2822_ (.A_N(net5),
    .B(_0683_),
    .C(_0684_),
    .D(_0681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0700_));
 sky130_fd_sc_hd__a22o_1 _2823_ (.A1(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .A2(_0699_),
    .B1(_0700_),
    .B2(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0701_));
 sky130_fd_sc_hd__and4bb_4 _2824_ (.A_N(_0681_),
    .B_N(_0682_),
    .C(net3),
    .D(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0702_));
 sky130_fd_sc_hd__nor4b_1 _2825_ (.A(_0681_),
    .B(_0682_),
    .C(_0684_),
    .D_N(net3),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0703_));
 sky130_fd_sc_hd__a22o_1 _2826_ (.A1(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .A2(_0702_),
    .B1(net10),
    .B2(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0704_));
 sky130_fd_sc_hd__and4bb_4 _2827_ (.A_N(_0683_),
    .B_N(_0684_),
    .C(net4),
    .D(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0705_));
 sky130_fd_sc_hd__and4b_4 _2828_ (.A_N(_0681_),
    .B(_0682_),
    .C(_0683_),
    .D(_0684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0706_));
 sky130_fd_sc_hd__a22o_1 _2829_ (.A1(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .A2(_0705_),
    .B1(_0706_),
    .B2(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0707_));
 sky130_fd_sc_hd__nor4b_1 _2830_ (.A(net5),
    .B(net3),
    .C(net2),
    .D_N(net4),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0708_));
 sky130_fd_sc_hd__and4bb_4 _2831_ (.A_N(_0681_),
    .B_N(_0683_),
    .C(net2),
    .D(net5),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0709_));
 sky130_fd_sc_hd__a22o_1 _2832_ (.A1(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .A2(net23),
    .B1(_0709_),
    .B2(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0710_));
 sky130_fd_sc_hd__or4_1 _2833_ (.A(_0701_),
    .B(_0704_),
    .C(_0707_),
    .D(_0710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0711_));
 sky130_fd_sc_hd__or3_4 _2834_ (.A(_0692_),
    .B(_0698_),
    .C(_0711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0712_));
 sky130_fd_sc_hd__and3_1 _2835_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[0] ),
    .B(_0686_),
    .C(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0713_));
 sky130_fd_sc_hd__buf_2 _2836_ (.A(_0686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0714_));
 sky130_fd_sc_hd__buf_2 _2837_ (.A(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0715_));
 sky130_fd_sc_hd__a21o_1 _2838_ (.A1(_0714_),
    .A2(_0715_),
    .B1(\genblk1[1].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0716_));
 sky130_fd_sc_hd__and3b_1 _2839_ (.A_N(_0713_),
    .B(_0631_),
    .C(_0716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0717_));
 sky130_fd_sc_hd__clkbuf_1 _2840_ (.A(_0717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0018_));
 sky130_fd_sc_hd__nand2_1 _2841_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[1] ),
    .B(\genblk1[1].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0718_));
 sky130_fd_sc_hd__nand2_2 _2842_ (.A(_0714_),
    .B(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0719_));
 sky130_fd_sc_hd__o221a_1 _2843_ (.A1(_0718_),
    .A2(_0719_),
    .B1(_0713_),
    .B2(net223),
    .C1(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0019_));
 sky130_fd_sc_hd__inv_2 _2844_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0720_));
 sky130_fd_sc_hd__and4bb_1 _2845_ (.A_N(_0720_),
    .B_N(_0718_),
    .C(_0686_),
    .D(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0721_));
 sky130_fd_sc_hd__clkbuf_2 _2846_ (.A(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0722_));
 sky130_fd_sc_hd__a41o_1 _2847_ (.A1(\genblk1[1].puf_buffer.cnt_1.ctr[1] ),
    .A2(\genblk1[1].puf_buffer.cnt_1.ctr[0] ),
    .A3(_0686_),
    .A4(_0712_),
    .B1(\genblk1[1].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0723_));
 sky130_fd_sc_hd__and3b_1 _2848_ (.A_N(_0721_),
    .B(_0722_),
    .C(_0723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0724_));
 sky130_fd_sc_hd__clkbuf_1 _2849_ (.A(_0724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0020_));
 sky130_fd_sc_hd__inv_2 _2850_ (.A(_0674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0725_));
 sky130_fd_sc_hd__o221a_1 _2851_ (.A1(_0725_),
    .A2(_0719_),
    .B1(_0721_),
    .B2(net143),
    .C1(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0021_));
 sky130_fd_sc_hd__and4_1 _2852_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[4] ),
    .B(_0674_),
    .C(_0686_),
    .D(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0726_));
 sky130_fd_sc_hd__a31o_1 _2853_ (.A1(_0674_),
    .A2(_0714_),
    .A3(_0715_),
    .B1(\genblk1[1].puf_buffer.cnt_1.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0727_));
 sky130_fd_sc_hd__and3b_1 _2854_ (.A_N(_0726_),
    .B(_0722_),
    .C(_0727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0728_));
 sky130_fd_sc_hd__clkbuf_1 _2855_ (.A(_0728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0022_));
 sky130_fd_sc_hd__and3_1 _2856_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[1].puf_buffer.cnt_1.ctr[4] ),
    .C(_0674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0729_));
 sky130_fd_sc_hd__inv_2 _2857_ (.A(_0729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0730_));
 sky130_fd_sc_hd__o221a_1 _2858_ (.A1(_0730_),
    .A2(_0719_),
    .B1(_0726_),
    .B2(net177),
    .C1(_0639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0023_));
 sky130_fd_sc_hd__and4_1 _2859_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[6] ),
    .B(_0729_),
    .C(_0686_),
    .D(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0731_));
 sky130_fd_sc_hd__a31o_1 _2860_ (.A1(_0729_),
    .A2(_0714_),
    .A3(_0715_),
    .B1(\genblk1[1].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0732_));
 sky130_fd_sc_hd__and3b_1 _2861_ (.A_N(_0731_),
    .B(_0722_),
    .C(_0732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0733_));
 sky130_fd_sc_hd__clkbuf_1 _2862_ (.A(_0733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0024_));
 sky130_fd_sc_hd__inv_2 _2863_ (.A(_0676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0734_));
 sky130_fd_sc_hd__clkbuf_4 _2864_ (.A(_0638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0735_));
 sky130_fd_sc_hd__o221a_1 _2865_ (.A1(_0734_),
    .A2(_0719_),
    .B1(_0731_),
    .B2(net129),
    .C1(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0025_));
 sky130_fd_sc_hd__and4_1 _2866_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[8] ),
    .B(_0676_),
    .C(_0686_),
    .D(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0736_));
 sky130_fd_sc_hd__a31o_1 _2867_ (.A1(_0676_),
    .A2(_0714_),
    .A3(_0715_),
    .B1(\genblk1[1].puf_buffer.cnt_1.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0737_));
 sky130_fd_sc_hd__and3b_1 _2868_ (.A_N(_0736_),
    .B(_0722_),
    .C(_0737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0738_));
 sky130_fd_sc_hd__clkbuf_1 _2869_ (.A(_0738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0026_));
 sky130_fd_sc_hd__nand3_1 _2870_ (.A(_0677_),
    .B(_0714_),
    .C(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0739_));
 sky130_fd_sc_hd__o211a_1 _2871_ (.A1(net144),
    .A2(_0736_),
    .B1(_0739_),
    .C1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0027_));
 sky130_fd_sc_hd__and4_1 _2872_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[10] ),
    .B(_0677_),
    .C(_0686_),
    .D(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0740_));
 sky130_fd_sc_hd__a31o_1 _2873_ (.A1(_0677_),
    .A2(_0714_),
    .A3(_0715_),
    .B1(\genblk1[1].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0741_));
 sky130_fd_sc_hd__and3b_1 _2874_ (.A_N(_0740_),
    .B(_0722_),
    .C(_0741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0742_));
 sky130_fd_sc_hd__clkbuf_1 _2875_ (.A(_0742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0028_));
 sky130_fd_sc_hd__nand2_1 _2876_ (.A(net200),
    .B(\genblk1[1].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0743_));
 sky130_fd_sc_hd__o221a_1 _2877_ (.A1(_0743_),
    .A2(_0739_),
    .B1(_0740_),
    .B2(net200),
    .C1(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0029_));
 sky130_fd_sc_hd__inv_2 _2878_ (.A(_0678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0744_));
 sky130_fd_sc_hd__and2_1 _2879_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[11] ),
    .B(\genblk1[1].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0745_));
 sky130_fd_sc_hd__a41o_1 _2880_ (.A1(_0677_),
    .A2(_0745_),
    .A3(_0714_),
    .A4(_0715_),
    .B1(net221),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0746_));
 sky130_fd_sc_hd__o211a_1 _2881_ (.A1(_0744_),
    .A2(_0739_),
    .B1(_0746_),
    .C1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0030_));
 sky130_fd_sc_hd__and4_1 _2882_ (.A(_0677_),
    .B(_0679_),
    .C(_0686_),
    .D(_0712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0747_));
 sky130_fd_sc_hd__a41o_1 _2883_ (.A1(_0677_),
    .A2(_0678_),
    .A3(_0686_),
    .A4(_0712_),
    .B1(\genblk1[1].puf_buffer.cnt_1.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0748_));
 sky130_fd_sc_hd__and3b_1 _2884_ (.A_N(_0747_),
    .B(_0722_),
    .C(_0748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0749_));
 sky130_fd_sc_hd__clkbuf_1 _2885_ (.A(_0749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0031_));
 sky130_fd_sc_hd__inv_2 _2886_ (.A(_0680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0750_));
 sky130_fd_sc_hd__o221a_1 _2887_ (.A1(_0750_),
    .A2(_0719_),
    .B1(_0747_),
    .B2(net80),
    .C1(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0032_));
 sky130_fd_sc_hd__buf_2 _2888_ (.A(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0751_));
 sky130_fd_sc_hd__nand4_1 _2889_ (.A(\genblk1[1].puf_buffer.cnt_1.ctr[15] ),
    .B(_0680_),
    .C(_0714_),
    .D(_0715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0752_));
 sky130_fd_sc_hd__a31o_1 _2890_ (.A1(_0680_),
    .A2(_0714_),
    .A3(_0715_),
    .B1(\genblk1[1].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0753_));
 sky130_fd_sc_hd__and3_1 _2891_ (.A(_0751_),
    .B(_0752_),
    .C(_0753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0754_));
 sky130_fd_sc_hd__clkbuf_1 _2892_ (.A(_0754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0033_));
 sky130_fd_sc_hd__inv_2 _2893_ (.A(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0755_));
 sky130_fd_sc_hd__and3b_1 _2894_ (.A_N(\genblk1[2].puf_buffer.cnt_1.finish ),
    .B(\genblk1[2].puf_buffer.cnt_2.finish ),
    .C(_0325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0756_));
 sky130_fd_sc_hd__clkbuf_1 _2895_ (.A(_0756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0071_));
 sky130_fd_sc_hd__o21bai_1 _2896_ (.A1(_0755_),
    .A2(_0071_),
    .B1_N(\genblk1[2].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0034_));
 sky130_fd_sc_hd__and3b_1 _2897_ (.A_N(\genblk1[1].puf_buffer.cnt_1.finish ),
    .B(\genblk1[1].puf_buffer.cnt_2.finish ),
    .C(_0586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0757_));
 sky130_fd_sc_hd__clkbuf_1 _2898_ (.A(_0757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0035_));
 sky130_fd_sc_hd__and3_1 _2899_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[12] ),
    .B(\genblk1[2].puf_buffer.cnt_2.ctr[11] ),
    .C(\genblk1[2].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0758_));
 sky130_fd_sc_hd__and2_1 _2900_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[13] ),
    .B(_0758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0759_));
 sky130_fd_sc_hd__and2_1 _2901_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[9] ),
    .B(\genblk1[2].puf_buffer.cnt_2.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0760_));
 sky130_fd_sc_hd__and4_1 _2902_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[3] ),
    .B(\genblk1[2].puf_buffer.cnt_2.ctr[2] ),
    .C(\genblk1[2].puf_buffer.cnt_2.ctr[1] ),
    .D(\genblk1[2].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0761_));
 sky130_fd_sc_hd__and3_1 _2903_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[2].puf_buffer.cnt_2.ctr[4] ),
    .C(_0761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0762_));
 sky130_fd_sc_hd__and4_1 _2904_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[2].puf_buffer.cnt_2.ctr[6] ),
    .C(_0760_),
    .D(_0762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0763_));
 sky130_fd_sc_hd__and3_1 _2905_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[14] ),
    .B(_0759_),
    .C(_0763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0764_));
 sky130_fd_sc_hd__a22o_1 _2906_ (.A1(_0589_),
    .A2(\genblk1[2].puf_buffer.cnt_2.finish ),
    .B1(_0764_),
    .B2(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0036_));
 sky130_fd_sc_hd__or2_1 _2907_ (.A(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0765_));
 sky130_fd_sc_hd__buf_2 _2908_ (.A(_0765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0766_));
 sky130_fd_sc_hd__a22o_1 _2909_ (.A1(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .A2(_0621_),
    .B1(_0603_),
    .B2(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0767_));
 sky130_fd_sc_hd__a221o_1 _2910_ (.A1(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .A2(net18),
    .B1(_0625_),
    .B2(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .C1(_0767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0768_));
 sky130_fd_sc_hd__a22o_1 _2911_ (.A1(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .A2(_0611_),
    .B1(_0618_),
    .B2(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0769_));
 sky130_fd_sc_hd__a211o_1 _2912_ (.A1(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .A2(_0615_),
    .B1(_0769_),
    .C1(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0770_));
 sky130_fd_sc_hd__a22o_1 _2913_ (.A1(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .A2(_0624_),
    .B1(_0622_),
    .B2(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0771_));
 sky130_fd_sc_hd__a22o_1 _2914_ (.A1(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .A2(net25),
    .B1(_0604_),
    .B2(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0772_));
 sky130_fd_sc_hd__a22o_1 _2915_ (.A1(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .A2(_0610_),
    .B1(net16),
    .B2(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0773_));
 sky130_fd_sc_hd__a22o_1 _2916_ (.A1(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .A2(_0605_),
    .B1(net22),
    .B2(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0774_));
 sky130_fd_sc_hd__or4_1 _2917_ (.A(_0771_),
    .B(_0772_),
    .C(_0773_),
    .D(_0774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0775_));
 sky130_fd_sc_hd__or3_2 _2918_ (.A(_0768_),
    .B(_0770_),
    .C(_0775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0776_));
 sky130_fd_sc_hd__buf_2 _2919_ (.A(_0776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0777_));
 sky130_fd_sc_hd__and3_1 _2920_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[0] ),
    .B(_0766_),
    .C(_0777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0778_));
 sky130_fd_sc_hd__a21o_1 _2921_ (.A1(_0766_),
    .A2(_0777_),
    .B1(\genblk1[2].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0779_));
 sky130_fd_sc_hd__and3b_1 _2922_ (.A_N(_0778_),
    .B(_0722_),
    .C(_0779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0780_));
 sky130_fd_sc_hd__clkbuf_1 _2923_ (.A(_0780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0037_));
 sky130_fd_sc_hd__nand2_1 _2924_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[1] ),
    .B(\genblk1[2].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0781_));
 sky130_fd_sc_hd__buf_2 _2925_ (.A(_0765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0782_));
 sky130_fd_sc_hd__clkbuf_2 _2926_ (.A(_0776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0783_));
 sky130_fd_sc_hd__nand2_1 _2927_ (.A(_0782_),
    .B(_0783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0784_));
 sky130_fd_sc_hd__o221a_1 _2928_ (.A1(_0781_),
    .A2(_0784_),
    .B1(_0778_),
    .B2(net204),
    .C1(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0038_));
 sky130_fd_sc_hd__inv_2 _2929_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0785_));
 sky130_fd_sc_hd__and4bb_1 _2930_ (.A_N(_0785_),
    .B_N(_0781_),
    .C(_0765_),
    .D(_0776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0786_));
 sky130_fd_sc_hd__a41o_1 _2931_ (.A1(\genblk1[2].puf_buffer.cnt_2.ctr[1] ),
    .A2(\genblk1[2].puf_buffer.cnt_2.ctr[0] ),
    .A3(_0766_),
    .A4(_0777_),
    .B1(\genblk1[2].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0787_));
 sky130_fd_sc_hd__and3b_1 _2932_ (.A_N(_0786_),
    .B(_0722_),
    .C(_0787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0788_));
 sky130_fd_sc_hd__clkbuf_1 _2933_ (.A(_0788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0039_));
 sky130_fd_sc_hd__inv_2 _2934_ (.A(_0761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0789_));
 sky130_fd_sc_hd__o221a_1 _2935_ (.A1(_0789_),
    .A2(_0784_),
    .B1(_0786_),
    .B2(net133),
    .C1(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0040_));
 sky130_fd_sc_hd__and4_1 _2936_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[4] ),
    .B(_0761_),
    .C(_0765_),
    .D(_0776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0790_));
 sky130_fd_sc_hd__a31o_1 _2937_ (.A1(_0761_),
    .A2(_0766_),
    .A3(_0777_),
    .B1(\genblk1[2].puf_buffer.cnt_2.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0791_));
 sky130_fd_sc_hd__and3b_1 _2938_ (.A_N(_0790_),
    .B(_0722_),
    .C(_0791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0792_));
 sky130_fd_sc_hd__clkbuf_1 _2939_ (.A(_0792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0041_));
 sky130_fd_sc_hd__inv_2 _2940_ (.A(_0762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0793_));
 sky130_fd_sc_hd__o221a_1 _2941_ (.A1(_0793_),
    .A2(_0784_),
    .B1(_0790_),
    .B2(net110),
    .C1(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0042_));
 sky130_fd_sc_hd__and4_1 _2942_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[6] ),
    .B(_0762_),
    .C(_0766_),
    .D(_0777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0794_));
 sky130_fd_sc_hd__a31o_1 _2943_ (.A1(_0762_),
    .A2(_0766_),
    .A3(_0777_),
    .B1(\genblk1[2].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0795_));
 sky130_fd_sc_hd__and3b_1 _2944_ (.A_N(_0794_),
    .B(_0722_),
    .C(_0795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0796_));
 sky130_fd_sc_hd__clkbuf_1 _2945_ (.A(_0796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0043_));
 sky130_fd_sc_hd__and3_1 _2946_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[2].puf_buffer.cnt_2.ctr[6] ),
    .C(_0762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0797_));
 sky130_fd_sc_hd__nand3_1 _2947_ (.A(_0797_),
    .B(_0782_),
    .C(_0783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0798_));
 sky130_fd_sc_hd__o211a_1 _2948_ (.A1(net185),
    .A2(_0794_),
    .B1(_0798_),
    .C1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0044_));
 sky130_fd_sc_hd__and4_1 _2949_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[8] ),
    .B(_0797_),
    .C(_0766_),
    .D(_0777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0799_));
 sky130_fd_sc_hd__clkbuf_2 _2950_ (.A(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0800_));
 sky130_fd_sc_hd__a31o_1 _2951_ (.A1(_0797_),
    .A2(_0766_),
    .A3(_0777_),
    .B1(\genblk1[2].puf_buffer.cnt_2.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0801_));
 sky130_fd_sc_hd__and3b_1 _2952_ (.A_N(_0799_),
    .B(_0800_),
    .C(_0801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0802_));
 sky130_fd_sc_hd__clkbuf_1 _2953_ (.A(_0802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0045_));
 sky130_fd_sc_hd__and4_2 _2954_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[2].puf_buffer.cnt_2.ctr[6] ),
    .C(_0760_),
    .D(_0762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0803_));
 sky130_fd_sc_hd__inv_2 _2955_ (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0804_));
 sky130_fd_sc_hd__clkbuf_4 _2956_ (.A(_0804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0805_));
 sky130_fd_sc_hd__a31o_1 _2957_ (.A1(_0803_),
    .A2(_0782_),
    .A3(_0783_),
    .B1(_0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0806_));
 sky130_fd_sc_hd__o21ba_1 _2958_ (.A1(net48),
    .A2(_0799_),
    .B1_N(_0806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0046_));
 sky130_fd_sc_hd__a31o_1 _2959_ (.A1(_0803_),
    .A2(_0766_),
    .A3(_0777_),
    .B1(\genblk1[2].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0807_));
 sky130_fd_sc_hd__nand4_1 _2960_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[10] ),
    .B(_0803_),
    .C(_0782_),
    .D(_0783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0808_));
 sky130_fd_sc_hd__and3_1 _2961_ (.A(_0751_),
    .B(_0807_),
    .C(_0808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0809_));
 sky130_fd_sc_hd__clkbuf_1 _2962_ (.A(_0809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0047_));
 sky130_fd_sc_hd__inv_2 _2963_ (.A(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0810_));
 sky130_fd_sc_hd__and2_1 _2964_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[11] ),
    .B(\genblk1[2].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0811_));
 sky130_fd_sc_hd__and4_1 _2965_ (.A(_0811_),
    .B(_0803_),
    .C(_0782_),
    .D(_0783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0812_));
 sky130_fd_sc_hd__clkbuf_4 _2966_ (.A(_0804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0813_));
 sky130_fd_sc_hd__clkbuf_4 _2967_ (.A(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0814_));
 sky130_fd_sc_hd__a211oi_1 _2968_ (.A1(_0810_),
    .A2(_0808_),
    .B1(_0812_),
    .C1(_0814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0048_));
 sky130_fd_sc_hd__a41o_1 _2969_ (.A1(_0758_),
    .A2(_0803_),
    .A3(_0782_),
    .A4(_0783_),
    .B1(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0815_));
 sky130_fd_sc_hd__o21ba_1 _2970_ (.A1(net65),
    .A2(_0812_),
    .B1_N(_0815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0049_));
 sky130_fd_sc_hd__and4_1 _2971_ (.A(_0758_),
    .B(_0803_),
    .C(_0782_),
    .D(_0783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0816_));
 sky130_fd_sc_hd__nand4_1 _2972_ (.A(_0759_),
    .B(_0803_),
    .C(_0782_),
    .D(_0783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0817_));
 sky130_fd_sc_hd__o211a_1 _2973_ (.A1(net159),
    .A2(_0816_),
    .B1(_0817_),
    .C1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0050_));
 sky130_fd_sc_hd__inv_2 _2974_ (.A(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0818_));
 sky130_fd_sc_hd__and3_1 _2975_ (.A(_0764_),
    .B(_0782_),
    .C(_0783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0819_));
 sky130_fd_sc_hd__a211oi_1 _2976_ (.A1(_0818_),
    .A2(_0817_),
    .B1(_0819_),
    .C1(_0814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0051_));
 sky130_fd_sc_hd__a31o_1 _2977_ (.A1(_0764_),
    .A2(_0766_),
    .A3(_0777_),
    .B1(\genblk1[2].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0820_));
 sky130_fd_sc_hd__nand4_1 _2978_ (.A(\genblk1[2].puf_buffer.cnt_2.ctr[15] ),
    .B(_0764_),
    .C(_0782_),
    .D(_0783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0821_));
 sky130_fd_sc_hd__and3_1 _2979_ (.A(_0751_),
    .B(_0820_),
    .C(_0821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0822_));
 sky130_fd_sc_hd__clkbuf_1 _2980_ (.A(_0822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0052_));
 sky130_fd_sc_hd__and3_1 _2981_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[12] ),
    .B(\genblk1[2].puf_buffer.cnt_1.ctr[11] ),
    .C(\genblk1[2].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0823_));
 sky130_fd_sc_hd__and2_1 _2982_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[13] ),
    .B(_0823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0824_));
 sky130_fd_sc_hd__and2_1 _2983_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[9] ),
    .B(\genblk1[2].puf_buffer.cnt_1.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0825_));
 sky130_fd_sc_hd__and4_1 _2984_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[3] ),
    .B(\genblk1[2].puf_buffer.cnt_1.ctr[2] ),
    .C(\genblk1[2].puf_buffer.cnt_1.ctr[1] ),
    .D(\genblk1[2].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0826_));
 sky130_fd_sc_hd__and3_1 _2985_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[2].puf_buffer.cnt_1.ctr[4] ),
    .C(_0826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0827_));
 sky130_fd_sc_hd__and4_1 _2986_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[2].puf_buffer.cnt_1.ctr[6] ),
    .C(_0825_),
    .D(_0827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0828_));
 sky130_fd_sc_hd__and3_1 _2987_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[14] ),
    .B(_0824_),
    .C(_0828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0829_));
 sky130_fd_sc_hd__a22o_1 _2988_ (.A1(_0589_),
    .A2(\genblk1[2].puf_buffer.cnt_1.finish ),
    .B1(_0829_),
    .B2(net130),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0053_));
 sky130_fd_sc_hd__or2_1 _2989_ (.A(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0830_));
 sky130_fd_sc_hd__buf_2 _2990_ (.A(_0830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0831_));
 sky130_fd_sc_hd__a22o_1 _2991_ (.A1(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .A2(_0699_),
    .B1(_0695_),
    .B2(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0832_));
 sky130_fd_sc_hd__a22o_1 _2992_ (.A1(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .A2(_0705_),
    .B1(_0690_),
    .B2(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0833_));
 sky130_fd_sc_hd__a221o_1 _2993_ (.A1(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .A2(_0689_),
    .B1(net13),
    .B2(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .C1(_0833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0834_));
 sky130_fd_sc_hd__a22o_1 _2994_ (.A1(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .A2(net15),
    .B1(_0706_),
    .B2(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0835_));
 sky130_fd_sc_hd__a21o_1 _2995_ (.A1(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .A2(_0709_),
    .B1(_0835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0836_));
 sky130_fd_sc_hd__a221o_1 _2996_ (.A1(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .A2(net23),
    .B1(_0687_),
    .B2(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .C1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0837_));
 sky130_fd_sc_hd__a22o_1 _2997_ (.A1(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .A2(_0694_),
    .B1(_0702_),
    .B2(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0838_));
 sky130_fd_sc_hd__a22o_1 _2998_ (.A1(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .A2(_0700_),
    .B1(net10),
    .B2(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0839_));
 sky130_fd_sc_hd__or3_1 _2999_ (.A(_0837_),
    .B(_0838_),
    .C(_0839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0840_));
 sky130_fd_sc_hd__or4_2 _3000_ (.A(_0832_),
    .B(_0834_),
    .C(_0836_),
    .D(_0840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0841_));
 sky130_fd_sc_hd__buf_2 _3001_ (.A(_0841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0842_));
 sky130_fd_sc_hd__and3_1 _3002_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[0] ),
    .B(_0831_),
    .C(_0842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0843_));
 sky130_fd_sc_hd__a21o_1 _3003_ (.A1(_0831_),
    .A2(_0842_),
    .B1(\genblk1[2].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0844_));
 sky130_fd_sc_hd__and3b_1 _3004_ (.A_N(_0843_),
    .B(_0800_),
    .C(_0844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0845_));
 sky130_fd_sc_hd__clkbuf_1 _3005_ (.A(_0845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0054_));
 sky130_fd_sc_hd__nand2_1 _3006_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[1] ),
    .B(\genblk1[2].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0846_));
 sky130_fd_sc_hd__buf_2 _3007_ (.A(_0830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0847_));
 sky130_fd_sc_hd__buf_2 _3008_ (.A(_0841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0848_));
 sky130_fd_sc_hd__nand2_1 _3009_ (.A(_0847_),
    .B(_0848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0849_));
 sky130_fd_sc_hd__o221a_1 _3010_ (.A1(_0846_),
    .A2(_0849_),
    .B1(_0843_),
    .B2(net214),
    .C1(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0055_));
 sky130_fd_sc_hd__inv_2 _3011_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0850_));
 sky130_fd_sc_hd__and4bb_1 _3012_ (.A_N(_0850_),
    .B_N(_0846_),
    .C(_0830_),
    .D(_0841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0851_));
 sky130_fd_sc_hd__a41o_1 _3013_ (.A1(\genblk1[2].puf_buffer.cnt_1.ctr[1] ),
    .A2(\genblk1[2].puf_buffer.cnt_1.ctr[0] ),
    .A3(_0831_),
    .A4(_0842_),
    .B1(\genblk1[2].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0852_));
 sky130_fd_sc_hd__and3b_1 _3014_ (.A_N(_0851_),
    .B(_0800_),
    .C(_0852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0853_));
 sky130_fd_sc_hd__clkbuf_1 _3015_ (.A(_0853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0056_));
 sky130_fd_sc_hd__inv_2 _3016_ (.A(_0826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0854_));
 sky130_fd_sc_hd__o221a_1 _3017_ (.A1(_0854_),
    .A2(_0849_),
    .B1(_0851_),
    .B2(net109),
    .C1(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0057_));
 sky130_fd_sc_hd__and4_1 _3018_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[4] ),
    .B(_0826_),
    .C(_0830_),
    .D(_0841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0855_));
 sky130_fd_sc_hd__a31o_1 _3019_ (.A1(_0826_),
    .A2(_0831_),
    .A3(_0842_),
    .B1(\genblk1[2].puf_buffer.cnt_1.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0856_));
 sky130_fd_sc_hd__and3b_1 _3020_ (.A_N(_0855_),
    .B(_0800_),
    .C(_0856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0857_));
 sky130_fd_sc_hd__clkbuf_1 _3021_ (.A(_0857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0058_));
 sky130_fd_sc_hd__inv_2 _3022_ (.A(_0827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0858_));
 sky130_fd_sc_hd__o221a_1 _3023_ (.A1(_0858_),
    .A2(_0849_),
    .B1(_0855_),
    .B2(net120),
    .C1(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0059_));
 sky130_fd_sc_hd__and4_1 _3024_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[6] ),
    .B(_0827_),
    .C(_0831_),
    .D(_0842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0859_));
 sky130_fd_sc_hd__a31o_1 _3025_ (.A1(_0827_),
    .A2(_0831_),
    .A3(_0842_),
    .B1(\genblk1[2].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0860_));
 sky130_fd_sc_hd__and3b_1 _3026_ (.A_N(_0859_),
    .B(_0800_),
    .C(_0860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0861_));
 sky130_fd_sc_hd__clkbuf_1 _3027_ (.A(_0861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0060_));
 sky130_fd_sc_hd__and3_1 _3028_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[2].puf_buffer.cnt_1.ctr[6] ),
    .C(_0827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0862_));
 sky130_fd_sc_hd__nand3_1 _3029_ (.A(_0862_),
    .B(_0847_),
    .C(_0848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0863_));
 sky130_fd_sc_hd__o211a_1 _3030_ (.A1(net179),
    .A2(_0859_),
    .B1(_0863_),
    .C1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0061_));
 sky130_fd_sc_hd__and4_1 _3031_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[8] ),
    .B(_0862_),
    .C(_0831_),
    .D(_0842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0864_));
 sky130_fd_sc_hd__a31o_1 _3032_ (.A1(_0862_),
    .A2(_0831_),
    .A3(_0842_),
    .B1(\genblk1[2].puf_buffer.cnt_1.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0865_));
 sky130_fd_sc_hd__and3b_1 _3033_ (.A_N(_0864_),
    .B(_0800_),
    .C(_0865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0866_));
 sky130_fd_sc_hd__clkbuf_1 _3034_ (.A(_0866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0062_));
 sky130_fd_sc_hd__and4_2 _3035_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[2].puf_buffer.cnt_1.ctr[6] ),
    .C(_0825_),
    .D(_0827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0867_));
 sky130_fd_sc_hd__a31o_1 _3036_ (.A1(_0867_),
    .A2(_0847_),
    .A3(_0848_),
    .B1(_0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0868_));
 sky130_fd_sc_hd__o21ba_1 _3037_ (.A1(net49),
    .A2(_0864_),
    .B1_N(_0868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0063_));
 sky130_fd_sc_hd__a31o_1 _3038_ (.A1(_0867_),
    .A2(_0831_),
    .A3(_0842_),
    .B1(\genblk1[2].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0869_));
 sky130_fd_sc_hd__nand4_1 _3039_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[10] ),
    .B(_0867_),
    .C(_0847_),
    .D(_0848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0870_));
 sky130_fd_sc_hd__and3_1 _3040_ (.A(_0751_),
    .B(_0869_),
    .C(_0870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0871_));
 sky130_fd_sc_hd__clkbuf_1 _3041_ (.A(_0871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0064_));
 sky130_fd_sc_hd__inv_2 _3042_ (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0872_));
 sky130_fd_sc_hd__and2_1 _3043_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[11] ),
    .B(\genblk1[2].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0873_));
 sky130_fd_sc_hd__and4_1 _3044_ (.A(_0873_),
    .B(_0867_),
    .C(_0847_),
    .D(_0848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0874_));
 sky130_fd_sc_hd__a211oi_1 _3045_ (.A1(_0872_),
    .A2(_0870_),
    .B1(_0874_),
    .C1(_0814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0065_));
 sky130_fd_sc_hd__a41o_1 _3046_ (.A1(_0823_),
    .A2(_0867_),
    .A3(_0847_),
    .A4(_0848_),
    .B1(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0875_));
 sky130_fd_sc_hd__o21ba_1 _3047_ (.A1(net52),
    .A2(_0874_),
    .B1_N(_0875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0066_));
 sky130_fd_sc_hd__and4_1 _3048_ (.A(_0823_),
    .B(_0867_),
    .C(_0847_),
    .D(_0848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0876_));
 sky130_fd_sc_hd__nand4_1 _3049_ (.A(_0824_),
    .B(_0867_),
    .C(_0847_),
    .D(_0848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0877_));
 sky130_fd_sc_hd__o211a_1 _3050_ (.A1(net121),
    .A2(_0876_),
    .B1(_0877_),
    .C1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0067_));
 sky130_fd_sc_hd__inv_2 _3051_ (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0878_));
 sky130_fd_sc_hd__and3_1 _3052_ (.A(_0829_),
    .B(_0847_),
    .C(_0848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0879_));
 sky130_fd_sc_hd__a211oi_1 _3053_ (.A1(_0878_),
    .A2(_0877_),
    .B1(_0879_),
    .C1(_0814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0068_));
 sky130_fd_sc_hd__a31o_1 _3054_ (.A1(_0829_),
    .A2(_0831_),
    .A3(_0842_),
    .B1(\genblk1[2].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0880_));
 sky130_fd_sc_hd__nand4_1 _3055_ (.A(\genblk1[2].puf_buffer.cnt_1.ctr[15] ),
    .B(_0829_),
    .C(_0847_),
    .D(_0848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0881_));
 sky130_fd_sc_hd__and3_1 _3056_ (.A(_0751_),
    .B(_0880_),
    .C(_0881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0882_));
 sky130_fd_sc_hd__clkbuf_1 _3057_ (.A(_0882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0069_));
 sky130_fd_sc_hd__inv_2 _3058_ (.A(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0883_));
 sky130_fd_sc_hd__and3b_1 _3059_ (.A_N(\genblk1[3].puf_buffer.cnt_1.finish ),
    .B(\genblk1[3].puf_buffer.cnt_2.finish ),
    .C(_0363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0884_));
 sky130_fd_sc_hd__clkbuf_1 _3060_ (.A(_0884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0107_));
 sky130_fd_sc_hd__o21bai_1 _3061_ (.A1(_0883_),
    .A2(_0107_),
    .B1_N(\genblk1[3].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0070_));
 sky130_fd_sc_hd__and3_1 _3062_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[12] ),
    .B(\genblk1[3].puf_buffer.cnt_2.ctr[11] ),
    .C(\genblk1[3].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0885_));
 sky130_fd_sc_hd__and2_1 _3063_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[13] ),
    .B(_0885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0886_));
 sky130_fd_sc_hd__and4_1 _3064_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[3] ),
    .B(\genblk1[3].puf_buffer.cnt_2.ctr[2] ),
    .C(\genblk1[3].puf_buffer.cnt_2.ctr[1] ),
    .D(\genblk1[3].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0887_));
 sky130_fd_sc_hd__and4_1 _3065_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[3].puf_buffer.cnt_2.ctr[5] ),
    .C(\genblk1[3].puf_buffer.cnt_2.ctr[4] ),
    .D(_0887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0888_));
 sky130_fd_sc_hd__and4_1 _3066_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[9] ),
    .B(\genblk1[3].puf_buffer.cnt_2.ctr[8] ),
    .C(\genblk1[3].puf_buffer.cnt_2.ctr[6] ),
    .D(_0888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0889_));
 sky130_fd_sc_hd__clkbuf_2 _3067_ (.A(_0889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0890_));
 sky130_fd_sc_hd__and3_1 _3068_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[14] ),
    .B(_0886_),
    .C(_0890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0891_));
 sky130_fd_sc_hd__a22o_1 _3069_ (.A1(_0589_),
    .A2(net146),
    .B1(_0891_),
    .B2(\genblk1[3].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0072_));
 sky130_fd_sc_hd__or2_2 _3070_ (.A(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0892_));
 sky130_fd_sc_hd__buf_2 _3071_ (.A(_0892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0893_));
 sky130_fd_sc_hd__a22o_1 _3072_ (.A1(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .A2(net22),
    .B1(net16),
    .B2(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0894_));
 sky130_fd_sc_hd__a221o_1 _3073_ (.A1(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .A2(_0603_),
    .B1(_0604_),
    .B2(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .C1(_0894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0895_));
 sky130_fd_sc_hd__a22o_1 _3074_ (.A1(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .A2(_0610_),
    .B1(_0622_),
    .B2(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0896_));
 sky130_fd_sc_hd__a211o_1 _3075_ (.A1(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .A2(net25),
    .B1(_0896_),
    .C1(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0897_));
 sky130_fd_sc_hd__a22o_1 _3076_ (.A1(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .A2(_0611_),
    .B1(_0621_),
    .B2(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0898_));
 sky130_fd_sc_hd__a22o_1 _3077_ (.A1(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .A2(_0624_),
    .B1(_0625_),
    .B2(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0899_));
 sky130_fd_sc_hd__a22o_1 _3078_ (.A1(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .A2(_0615_),
    .B1(_0618_),
    .B2(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0900_));
 sky130_fd_sc_hd__a22o_1 _3079_ (.A1(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .A2(net18),
    .B1(_0605_),
    .B2(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0901_));
 sky130_fd_sc_hd__or4_1 _3080_ (.A(_0898_),
    .B(_0899_),
    .C(_0900_),
    .D(_0901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0902_));
 sky130_fd_sc_hd__or3_2 _3081_ (.A(_0895_),
    .B(_0897_),
    .C(_0902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0903_));
 sky130_fd_sc_hd__buf_2 _3082_ (.A(_0903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0904_));
 sky130_fd_sc_hd__and3_1 _3083_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[0] ),
    .B(_0893_),
    .C(_0904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0905_));
 sky130_fd_sc_hd__a21o_1 _3084_ (.A1(_0893_),
    .A2(_0904_),
    .B1(\genblk1[3].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0906_));
 sky130_fd_sc_hd__and3b_1 _3085_ (.A_N(_0905_),
    .B(_0800_),
    .C(_0906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0907_));
 sky130_fd_sc_hd__clkbuf_1 _3086_ (.A(_0907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0073_));
 sky130_fd_sc_hd__nand2_1 _3087_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[1] ),
    .B(\genblk1[3].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0908_));
 sky130_fd_sc_hd__buf_2 _3088_ (.A(_0892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0909_));
 sky130_fd_sc_hd__buf_2 _3089_ (.A(_0903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0910_));
 sky130_fd_sc_hd__nand2_1 _3090_ (.A(_0909_),
    .B(_0910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0911_));
 sky130_fd_sc_hd__o221a_1 _3091_ (.A1(_0908_),
    .A2(_0911_),
    .B1(_0905_),
    .B2(net219),
    .C1(_0735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0074_));
 sky130_fd_sc_hd__inv_2 _3092_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0912_));
 sky130_fd_sc_hd__and4bb_1 _3093_ (.A_N(_0912_),
    .B_N(_0908_),
    .C(_0892_),
    .D(_0903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0913_));
 sky130_fd_sc_hd__a41o_1 _3094_ (.A1(\genblk1[3].puf_buffer.cnt_2.ctr[1] ),
    .A2(\genblk1[3].puf_buffer.cnt_2.ctr[0] ),
    .A3(_0892_),
    .A4(_0903_),
    .B1(\genblk1[3].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0914_));
 sky130_fd_sc_hd__and3b_1 _3095_ (.A_N(_0913_),
    .B(_0800_),
    .C(_0914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0915_));
 sky130_fd_sc_hd__clkbuf_1 _3096_ (.A(_0915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0075_));
 sky130_fd_sc_hd__inv_2 _3097_ (.A(_0887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0916_));
 sky130_fd_sc_hd__clkbuf_4 _3098_ (.A(_0638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0917_));
 sky130_fd_sc_hd__o221a_1 _3099_ (.A1(_0916_),
    .A2(_0911_),
    .B1(_0913_),
    .B2(net111),
    .C1(_0917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0076_));
 sky130_fd_sc_hd__and4_1 _3100_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[4] ),
    .B(_0887_),
    .C(_0892_),
    .D(_0903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0918_));
 sky130_fd_sc_hd__a31o_1 _3101_ (.A1(_0887_),
    .A2(_0893_),
    .A3(_0904_),
    .B1(\genblk1[3].puf_buffer.cnt_2.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0919_));
 sky130_fd_sc_hd__and3b_1 _3102_ (.A_N(_0918_),
    .B(_0800_),
    .C(_0919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0920_));
 sky130_fd_sc_hd__clkbuf_1 _3103_ (.A(_0920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0077_));
 sky130_fd_sc_hd__and3_1 _3104_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[3].puf_buffer.cnt_2.ctr[4] ),
    .C(_0887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0921_));
 sky130_fd_sc_hd__a31o_1 _3105_ (.A1(_0921_),
    .A2(_0909_),
    .A3(_0910_),
    .B1(_0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0922_));
 sky130_fd_sc_hd__o21ba_1 _3106_ (.A1(net178),
    .A2(_0918_),
    .B1_N(_0922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0078_));
 sky130_fd_sc_hd__a41o_1 _3107_ (.A1(\genblk1[3].puf_buffer.cnt_2.ctr[6] ),
    .A2(_0921_),
    .A3(_0893_),
    .A4(_0904_),
    .B1(_0804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0923_));
 sky130_fd_sc_hd__and3_1 _3108_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[3].puf_buffer.cnt_2.ctr[4] ),
    .C(_0887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0924_));
 sky130_fd_sc_hd__a31o_1 _3109_ (.A1(_0924_),
    .A2(_0893_),
    .A3(_0904_),
    .B1(\genblk1[3].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0925_));
 sky130_fd_sc_hd__and2b_1 _3110_ (.A_N(_0923_),
    .B(_0925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0926_));
 sky130_fd_sc_hd__clkbuf_1 _3111_ (.A(_0926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0079_));
 sky130_fd_sc_hd__and3_1 _3112_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[3].puf_buffer.cnt_2.ctr[6] ),
    .C(_0921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0927_));
 sky130_fd_sc_hd__and3_1 _3113_ (.A(_0927_),
    .B(_0893_),
    .C(_0904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0928_));
 sky130_fd_sc_hd__a41o_1 _3114_ (.A1(\genblk1[3].puf_buffer.cnt_2.ctr[6] ),
    .A2(_0924_),
    .A3(_0892_),
    .A4(_0903_),
    .B1(\genblk1[3].puf_buffer.cnt_2.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0929_));
 sky130_fd_sc_hd__and3b_1 _3115_ (.A_N(_0928_),
    .B(_0800_),
    .C(_0929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0930_));
 sky130_fd_sc_hd__clkbuf_1 _3116_ (.A(_0930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0080_));
 sky130_fd_sc_hd__a41o_1 _3117_ (.A1(\genblk1[3].puf_buffer.cnt_2.ctr[8] ),
    .A2(_0927_),
    .A3(_0909_),
    .A4(_0910_),
    .B1(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0931_));
 sky130_fd_sc_hd__o21ba_1 _3118_ (.A1(net182),
    .A2(_0928_),
    .B1_N(_0931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0081_));
 sky130_fd_sc_hd__a31o_1 _3119_ (.A1(_0890_),
    .A2(_0893_),
    .A3(_0904_),
    .B1(_0804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0932_));
 sky130_fd_sc_hd__a41o_1 _3120_ (.A1(\genblk1[3].puf_buffer.cnt_2.ctr[8] ),
    .A2(_0927_),
    .A3(_0893_),
    .A4(_0904_),
    .B1(\genblk1[3].puf_buffer.cnt_2.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0933_));
 sky130_fd_sc_hd__and2b_1 _3121_ (.A_N(_0932_),
    .B(_0933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0934_));
 sky130_fd_sc_hd__clkbuf_1 _3122_ (.A(_0934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0082_));
 sky130_fd_sc_hd__a31o_1 _3123_ (.A1(_0890_),
    .A2(_0893_),
    .A3(_0904_),
    .B1(\genblk1[3].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0935_));
 sky130_fd_sc_hd__nand4_1 _3124_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[10] ),
    .B(_0890_),
    .C(_0909_),
    .D(_0910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0936_));
 sky130_fd_sc_hd__and3_1 _3125_ (.A(_0751_),
    .B(_0935_),
    .C(_0936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0937_));
 sky130_fd_sc_hd__clkbuf_1 _3126_ (.A(_0937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0083_));
 sky130_fd_sc_hd__inv_2 _3127_ (.A(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0938_));
 sky130_fd_sc_hd__and2_1 _3128_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[11] ),
    .B(\genblk1[3].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0939_));
 sky130_fd_sc_hd__and4_1 _3129_ (.A(_0939_),
    .B(_0890_),
    .C(_0909_),
    .D(_0910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0940_));
 sky130_fd_sc_hd__a211oi_1 _3130_ (.A1(_0938_),
    .A2(_0936_),
    .B1(_0940_),
    .C1(_0814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0084_));
 sky130_fd_sc_hd__a41o_1 _3131_ (.A1(_0885_),
    .A2(_0890_),
    .A3(_0909_),
    .A4(_0910_),
    .B1(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0941_));
 sky130_fd_sc_hd__o21ba_1 _3132_ (.A1(net57),
    .A2(_0940_),
    .B1_N(_0941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0085_));
 sky130_fd_sc_hd__and4_1 _3133_ (.A(_0885_),
    .B(_0890_),
    .C(_0909_),
    .D(_0910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0942_));
 sky130_fd_sc_hd__nand4_1 _3134_ (.A(_0886_),
    .B(_0890_),
    .C(_0909_),
    .D(_0910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0943_));
 sky130_fd_sc_hd__o211a_1 _3135_ (.A1(net117),
    .A2(_0942_),
    .B1(_0943_),
    .C1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0086_));
 sky130_fd_sc_hd__inv_2 _3136_ (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0944_));
 sky130_fd_sc_hd__a31o_1 _3137_ (.A1(_0891_),
    .A2(_0909_),
    .A3(_0910_),
    .B1(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0945_));
 sky130_fd_sc_hd__a21oi_1 _3138_ (.A1(_0944_),
    .A2(_0943_),
    .B1(_0945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0087_));
 sky130_fd_sc_hd__a31o_1 _3139_ (.A1(_0891_),
    .A2(_0893_),
    .A3(_0904_),
    .B1(\genblk1[3].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0946_));
 sky130_fd_sc_hd__nand4_1 _3140_ (.A(\genblk1[3].puf_buffer.cnt_2.ctr[15] ),
    .B(_0891_),
    .C(_0909_),
    .D(_0910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0947_));
 sky130_fd_sc_hd__and3_1 _3141_ (.A(_0751_),
    .B(_0946_),
    .C(_0947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0948_));
 sky130_fd_sc_hd__clkbuf_1 _3142_ (.A(_0948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0088_));
 sky130_fd_sc_hd__and4_1 _3143_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[3] ),
    .B(\genblk1[3].puf_buffer.cnt_1.ctr[2] ),
    .C(\genblk1[3].puf_buffer.cnt_1.ctr[1] ),
    .D(\genblk1[3].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0949_));
 sky130_fd_sc_hd__and2_1 _3144_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[3].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0950_));
 sky130_fd_sc_hd__and4_1 _3145_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[3].puf_buffer.cnt_1.ctr[4] ),
    .C(_0949_),
    .D(_0950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0951_));
 sky130_fd_sc_hd__and3_2 _3146_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[9] ),
    .B(\genblk1[3].puf_buffer.cnt_1.ctr[8] ),
    .C(_0951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0952_));
 sky130_fd_sc_hd__and3_1 _3147_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[12] ),
    .B(\genblk1[3].puf_buffer.cnt_1.ctr[11] ),
    .C(\genblk1[3].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0953_));
 sky130_fd_sc_hd__and2_1 _3148_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[13] ),
    .B(_0953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0954_));
 sky130_fd_sc_hd__and3_1 _3149_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[14] ),
    .B(_0952_),
    .C(_0954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0955_));
 sky130_fd_sc_hd__a22o_1 _3150_ (.A1(_0589_),
    .A2(\genblk1[3].puf_buffer.cnt_1.finish ),
    .B1(_0955_),
    .B2(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0089_));
 sky130_fd_sc_hd__or2_1 _3151_ (.A(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0956_));
 sky130_fd_sc_hd__clkbuf_2 _3152_ (.A(_0956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0957_));
 sky130_fd_sc_hd__a22o_1 _3153_ (.A1(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .A2(_0706_),
    .B1(_0709_),
    .B2(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0958_));
 sky130_fd_sc_hd__a22o_1 _3154_ (.A1(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .A2(_0699_),
    .B1(net10),
    .B2(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0959_));
 sky130_fd_sc_hd__a211o_1 _3155_ (.A1(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .A2(net15),
    .B1(_0958_),
    .C1(_0959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0960_));
 sky130_fd_sc_hd__a22o_1 _3156_ (.A1(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .A2(_0690_),
    .B1(_0702_),
    .B2(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0961_));
 sky130_fd_sc_hd__a221o_1 _3157_ (.A1(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .A2(_0695_),
    .B1(net13),
    .B2(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .C1(_0961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0962_));
 sky130_fd_sc_hd__a22o_1 _3158_ (.A1(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .A2(_0700_),
    .B1(_0705_),
    .B2(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0963_));
 sky130_fd_sc_hd__a221o_1 _3159_ (.A1(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .A2(_0694_),
    .B1(_0687_),
    .B2(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .C1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0964_));
 sky130_fd_sc_hd__a22o_1 _3160_ (.A1(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .A2(_0689_),
    .B1(net23),
    .B2(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0965_));
 sky130_fd_sc_hd__or3_1 _3161_ (.A(_0963_),
    .B(_0964_),
    .C(_0965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0966_));
 sky130_fd_sc_hd__or3_2 _3162_ (.A(_0960_),
    .B(_0962_),
    .C(_0966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0967_));
 sky130_fd_sc_hd__clkbuf_2 _3163_ (.A(_0967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0968_));
 sky130_fd_sc_hd__and3_1 _3164_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[0] ),
    .B(_0957_),
    .C(_0968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0969_));
 sky130_fd_sc_hd__clkbuf_2 _3165_ (.A(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0970_));
 sky130_fd_sc_hd__buf_2 _3166_ (.A(_0956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0971_));
 sky130_fd_sc_hd__buf_2 _3167_ (.A(_0967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0972_));
 sky130_fd_sc_hd__a21o_1 _3168_ (.A1(_0971_),
    .A2(_0972_),
    .B1(\genblk1[3].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0973_));
 sky130_fd_sc_hd__and3b_1 _3169_ (.A_N(_0969_),
    .B(_0970_),
    .C(_0973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0974_));
 sky130_fd_sc_hd__clkbuf_1 _3170_ (.A(_0974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0090_));
 sky130_fd_sc_hd__nand2_1 _3171_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[1] ),
    .B(\genblk1[3].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0975_));
 sky130_fd_sc_hd__nand2_1 _3172_ (.A(_0971_),
    .B(_0972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0976_));
 sky130_fd_sc_hd__o221a_1 _3173_ (.A1(_0975_),
    .A2(_0976_),
    .B1(_0969_),
    .B2(net225),
    .C1(_0917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0091_));
 sky130_fd_sc_hd__inv_2 _3174_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0977_));
 sky130_fd_sc_hd__and4bb_1 _3175_ (.A_N(_0977_),
    .B_N(_0975_),
    .C(_0956_),
    .D(_0967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0978_));
 sky130_fd_sc_hd__a41o_1 _3176_ (.A1(\genblk1[3].puf_buffer.cnt_1.ctr[1] ),
    .A2(\genblk1[3].puf_buffer.cnt_1.ctr[0] ),
    .A3(_0957_),
    .A4(_0968_),
    .B1(\genblk1[3].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0979_));
 sky130_fd_sc_hd__and3b_1 _3177_ (.A_N(_0978_),
    .B(_0970_),
    .C(_0979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_1 _3178_ (.A(_0980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0092_));
 sky130_fd_sc_hd__inv_2 _3179_ (.A(_0949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0981_));
 sky130_fd_sc_hd__o221a_1 _3180_ (.A1(_0981_),
    .A2(_0976_),
    .B1(_0978_),
    .B2(net89),
    .C1(_0917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0093_));
 sky130_fd_sc_hd__and4_1 _3181_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[4] ),
    .B(_0949_),
    .C(_0957_),
    .D(_0968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0982_));
 sky130_fd_sc_hd__a31o_1 _3182_ (.A1(_0949_),
    .A2(_0971_),
    .A3(_0972_),
    .B1(\genblk1[3].puf_buffer.cnt_1.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0983_));
 sky130_fd_sc_hd__and3b_1 _3183_ (.A_N(_0982_),
    .B(_0970_),
    .C(_0983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0984_));
 sky130_fd_sc_hd__clkbuf_1 _3184_ (.A(_0984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0094_));
 sky130_fd_sc_hd__and3_1 _3185_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[3].puf_buffer.cnt_1.ctr[4] ),
    .C(_0949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0985_));
 sky130_fd_sc_hd__inv_2 _3186_ (.A(_0985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0986_));
 sky130_fd_sc_hd__o221a_1 _3187_ (.A1(_0986_),
    .A2(_0976_),
    .B1(_0982_),
    .B2(net170),
    .C1(_0917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0095_));
 sky130_fd_sc_hd__and4_1 _3188_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[6] ),
    .B(_0985_),
    .C(_0957_),
    .D(_0968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0987_));
 sky130_fd_sc_hd__a31o_1 _3189_ (.A1(_0985_),
    .A2(_0971_),
    .A3(_0972_),
    .B1(\genblk1[3].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0988_));
 sky130_fd_sc_hd__and3b_1 _3190_ (.A_N(_0987_),
    .B(_0970_),
    .C(_0988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0989_));
 sky130_fd_sc_hd__clkbuf_1 _3191_ (.A(_0989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0096_));
 sky130_fd_sc_hd__inv_2 _3192_ (.A(_0951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0990_));
 sky130_fd_sc_hd__o221a_1 _3193_ (.A1(_0990_),
    .A2(_0976_),
    .B1(_0987_),
    .B2(net86),
    .C1(_0917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0097_));
 sky130_fd_sc_hd__and4_1 _3194_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[8] ),
    .B(_0951_),
    .C(_0957_),
    .D(_0968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0991_));
 sky130_fd_sc_hd__a31o_1 _3195_ (.A1(_0951_),
    .A2(_0971_),
    .A3(_0972_),
    .B1(\genblk1[3].puf_buffer.cnt_1.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0992_));
 sky130_fd_sc_hd__and3b_1 _3196_ (.A_N(_0991_),
    .B(_0970_),
    .C(_0992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0993_));
 sky130_fd_sc_hd__clkbuf_1 _3197_ (.A(_0993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0098_));
 sky130_fd_sc_hd__nand3_1 _3198_ (.A(_0952_),
    .B(_0971_),
    .C(_0972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0994_));
 sky130_fd_sc_hd__o211a_1 _3199_ (.A1(net95),
    .A2(_0991_),
    .B1(_0994_),
    .C1(_0658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0099_));
 sky130_fd_sc_hd__and4_1 _3200_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[10] ),
    .B(_0952_),
    .C(_0957_),
    .D(_0968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0995_));
 sky130_fd_sc_hd__a31o_1 _3201_ (.A1(_0952_),
    .A2(_0971_),
    .A3(_0968_),
    .B1(\genblk1[3].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0996_));
 sky130_fd_sc_hd__and3b_1 _3202_ (.A_N(_0995_),
    .B(_0970_),
    .C(_0996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0997_));
 sky130_fd_sc_hd__clkbuf_1 _3203_ (.A(_0997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_1 _3204_ (.A(net197),
    .B(\genblk1[3].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0998_));
 sky130_fd_sc_hd__o221a_1 _3205_ (.A1(_0998_),
    .A2(_0994_),
    .B1(_0995_),
    .B2(net197),
    .C1(_0917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0101_));
 sky130_fd_sc_hd__a41o_1 _3206_ (.A1(_0952_),
    .A2(_0953_),
    .A3(_0957_),
    .A4(_0972_),
    .B1(_0804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0999_));
 sky130_fd_sc_hd__and2_1 _3207_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[11] ),
    .B(\genblk1[3].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1000_));
 sky130_fd_sc_hd__a41o_1 _3208_ (.A1(_0952_),
    .A2(_1000_),
    .A3(_0957_),
    .A4(_0968_),
    .B1(\genblk1[3].puf_buffer.cnt_1.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1001_));
 sky130_fd_sc_hd__and2b_1 _3209_ (.A_N(_0999_),
    .B(_1001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1002_));
 sky130_fd_sc_hd__clkbuf_1 _3210_ (.A(_1002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0102_));
 sky130_fd_sc_hd__and4_1 _3211_ (.A(_0952_),
    .B(_0954_),
    .C(_0957_),
    .D(_0968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1003_));
 sky130_fd_sc_hd__a41o_1 _3212_ (.A1(_0952_),
    .A2(_0953_),
    .A3(_0957_),
    .A4(_0968_),
    .B1(\genblk1[3].puf_buffer.cnt_1.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1004_));
 sky130_fd_sc_hd__and3b_1 _3213_ (.A_N(_1003_),
    .B(_0970_),
    .C(_1004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1005_));
 sky130_fd_sc_hd__clkbuf_1 _3214_ (.A(_1005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0103_));
 sky130_fd_sc_hd__nand3_1 _3215_ (.A(_0955_),
    .B(_0971_),
    .C(_0972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1006_));
 sky130_fd_sc_hd__clkbuf_4 _3216_ (.A(_0631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1007_));
 sky130_fd_sc_hd__o211a_1 _3217_ (.A1(net124),
    .A2(_1003_),
    .B1(_1006_),
    .C1(_1007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0104_));
 sky130_fd_sc_hd__a31o_1 _3218_ (.A1(_0955_),
    .A2(_0971_),
    .A3(_0972_),
    .B1(\genblk1[3].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1008_));
 sky130_fd_sc_hd__nand4_1 _3219_ (.A(\genblk1[3].puf_buffer.cnt_1.ctr[15] ),
    .B(_0955_),
    .C(_0971_),
    .D(_0972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1009_));
 sky130_fd_sc_hd__and3_1 _3220_ (.A(_0751_),
    .B(_1008_),
    .C(_1009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1010_));
 sky130_fd_sc_hd__clkbuf_1 _3221_ (.A(_1010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0105_));
 sky130_fd_sc_hd__inv_2 _3222_ (.A(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1011_));
 sky130_fd_sc_hd__and3b_1 _3223_ (.A_N(\genblk1[4].puf_buffer.cnt_1.finish ),
    .B(\genblk1[4].puf_buffer.cnt_2.finish ),
    .C(_0400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1012_));
 sky130_fd_sc_hd__clkbuf_1 _3224_ (.A(_1012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0143_));
 sky130_fd_sc_hd__o21bai_1 _3225_ (.A1(_1011_),
    .A2(_0143_),
    .B1_N(\genblk1[4].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0106_));
 sky130_fd_sc_hd__and3_1 _3226_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[12] ),
    .B(\genblk1[4].puf_buffer.cnt_2.ctr[11] ),
    .C(\genblk1[4].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1013_));
 sky130_fd_sc_hd__and2_1 _3227_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[13] ),
    .B(_1013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1014_));
 sky130_fd_sc_hd__and2_1 _3228_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[9] ),
    .B(\genblk1[4].puf_buffer.cnt_2.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1015_));
 sky130_fd_sc_hd__and4_1 _3229_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[3] ),
    .B(\genblk1[4].puf_buffer.cnt_2.ctr[2] ),
    .C(\genblk1[4].puf_buffer.cnt_2.ctr[1] ),
    .D(\genblk1[4].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1016_));
 sky130_fd_sc_hd__and3_1 _3230_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[4].puf_buffer.cnt_2.ctr[4] ),
    .C(_1016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1017_));
 sky130_fd_sc_hd__and4_1 _3231_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[4].puf_buffer.cnt_2.ctr[6] ),
    .C(_1015_),
    .D(_1017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1018_));
 sky130_fd_sc_hd__and3_1 _3232_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[14] ),
    .B(_1014_),
    .C(_1018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1019_));
 sky130_fd_sc_hd__a22o_1 _3233_ (.A1(_0589_),
    .A2(\genblk1[4].puf_buffer.cnt_2.finish ),
    .B1(_1019_),
    .B2(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0108_));
 sky130_fd_sc_hd__or2_1 _3234_ (.A(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1020_));
 sky130_fd_sc_hd__buf_2 _3235_ (.A(_1020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1021_));
 sky130_fd_sc_hd__a22o_1 _3236_ (.A1(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .A2(_0605_),
    .B1(net25),
    .B2(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1022_));
 sky130_fd_sc_hd__a22o_1 _3237_ (.A1(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .A2(_0622_),
    .B1(_0603_),
    .B2(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1023_));
 sky130_fd_sc_hd__a211o_1 _3238_ (.A1(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .A2(_0625_),
    .B1(_1022_),
    .C1(_1023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1024_));
 sky130_fd_sc_hd__a22o_1 _3239_ (.A1(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .A2(_0610_),
    .B1(_0611_),
    .B2(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1025_));
 sky130_fd_sc_hd__a21o_1 _3240_ (.A1(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .A2(_0621_),
    .B1(_1025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1026_));
 sky130_fd_sc_hd__a22o_1 _3241_ (.A1(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .A2(_0615_),
    .B1(net18),
    .B2(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1027_));
 sky130_fd_sc_hd__a22o_1 _3242_ (.A1(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .A2(net22),
    .B1(net17),
    .B2(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1028_));
 sky130_fd_sc_hd__a221o_1 _3243_ (.A1(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .A2(_0618_),
    .B1(_0604_),
    .B2(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .C1(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1029_));
 sky130_fd_sc_hd__a2111o_1 _3244_ (.A1(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .A2(_0624_),
    .B1(_1027_),
    .C1(_1028_),
    .D1(_1029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1030_));
 sky130_fd_sc_hd__or3_2 _3245_ (.A(_1024_),
    .B(_1026_),
    .C(_1030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1031_));
 sky130_fd_sc_hd__buf_2 _3246_ (.A(_1031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1032_));
 sky130_fd_sc_hd__and3_1 _3247_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[0] ),
    .B(_1021_),
    .C(_1032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1033_));
 sky130_fd_sc_hd__a21o_1 _3248_ (.A1(_1021_),
    .A2(_1032_),
    .B1(\genblk1[4].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1034_));
 sky130_fd_sc_hd__and3b_1 _3249_ (.A_N(_1033_),
    .B(_0970_),
    .C(_1034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1035_));
 sky130_fd_sc_hd__clkbuf_1 _3250_ (.A(_1035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0109_));
 sky130_fd_sc_hd__nand2_1 _3251_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[1] ),
    .B(\genblk1[4].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1036_));
 sky130_fd_sc_hd__clkbuf_2 _3252_ (.A(_1020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1037_));
 sky130_fd_sc_hd__clkbuf_2 _3253_ (.A(_1031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1038_));
 sky130_fd_sc_hd__nand2_1 _3254_ (.A(_1037_),
    .B(_1038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1039_));
 sky130_fd_sc_hd__o221a_1 _3255_ (.A1(_1036_),
    .A2(_1039_),
    .B1(_1033_),
    .B2(net222),
    .C1(_0917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0110_));
 sky130_fd_sc_hd__inv_2 _3256_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1040_));
 sky130_fd_sc_hd__and4bb_1 _3257_ (.A_N(_1040_),
    .B_N(_1036_),
    .C(_1020_),
    .D(_1031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1041_));
 sky130_fd_sc_hd__a41o_1 _3258_ (.A1(\genblk1[4].puf_buffer.cnt_2.ctr[1] ),
    .A2(\genblk1[4].puf_buffer.cnt_2.ctr[0] ),
    .A3(_1021_),
    .A4(_1032_),
    .B1(\genblk1[4].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1042_));
 sky130_fd_sc_hd__and3b_1 _3259_ (.A_N(_1041_),
    .B(_0970_),
    .C(_1042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1043_));
 sky130_fd_sc_hd__clkbuf_1 _3260_ (.A(_1043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0111_));
 sky130_fd_sc_hd__inv_2 _3261_ (.A(_1016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1044_));
 sky130_fd_sc_hd__o221a_1 _3262_ (.A1(_1044_),
    .A2(_1039_),
    .B1(_1041_),
    .B2(net99),
    .C1(_0917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0112_));
 sky130_fd_sc_hd__and4_1 _3263_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[4] ),
    .B(_1016_),
    .C(_1020_),
    .D(_1031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1045_));
 sky130_fd_sc_hd__a31o_1 _3264_ (.A1(_1016_),
    .A2(_1021_),
    .A3(_1032_),
    .B1(\genblk1[4].puf_buffer.cnt_2.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1046_));
 sky130_fd_sc_hd__and3b_1 _3265_ (.A_N(_1045_),
    .B(_0970_),
    .C(_1046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1047_));
 sky130_fd_sc_hd__clkbuf_1 _3266_ (.A(_1047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0113_));
 sky130_fd_sc_hd__inv_2 _3267_ (.A(_1017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1048_));
 sky130_fd_sc_hd__o221a_1 _3268_ (.A1(_1048_),
    .A2(_1039_),
    .B1(_1045_),
    .B2(net87),
    .C1(_0917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0114_));
 sky130_fd_sc_hd__and4_1 _3269_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[6] ),
    .B(_1017_),
    .C(_1021_),
    .D(_1032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1049_));
 sky130_fd_sc_hd__clkbuf_2 _3270_ (.A(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1050_));
 sky130_fd_sc_hd__a31o_1 _3271_ (.A1(_1017_),
    .A2(_1021_),
    .A3(_1032_),
    .B1(\genblk1[4].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1051_));
 sky130_fd_sc_hd__and3b_1 _3272_ (.A_N(_1049_),
    .B(_1050_),
    .C(_1051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1052_));
 sky130_fd_sc_hd__clkbuf_1 _3273_ (.A(_1052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0115_));
 sky130_fd_sc_hd__and3_1 _3274_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[4].puf_buffer.cnt_2.ctr[6] ),
    .C(_1017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1053_));
 sky130_fd_sc_hd__nand3_1 _3275_ (.A(_1053_),
    .B(_1037_),
    .C(_1038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1054_));
 sky130_fd_sc_hd__o211a_1 _3276_ (.A1(net183),
    .A2(_1049_),
    .B1(_1054_),
    .C1(_1007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0116_));
 sky130_fd_sc_hd__and4_1 _3277_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[8] ),
    .B(_1053_),
    .C(_1021_),
    .D(_1032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1055_));
 sky130_fd_sc_hd__a31o_1 _3278_ (.A1(_1053_),
    .A2(_1021_),
    .A3(_1032_),
    .B1(\genblk1[4].puf_buffer.cnt_2.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1056_));
 sky130_fd_sc_hd__and3b_1 _3279_ (.A_N(_1055_),
    .B(_1050_),
    .C(_1056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1057_));
 sky130_fd_sc_hd__clkbuf_1 _3280_ (.A(_1057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0117_));
 sky130_fd_sc_hd__and4_2 _3281_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[4].puf_buffer.cnt_2.ctr[6] ),
    .C(_1015_),
    .D(_1017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1058_));
 sky130_fd_sc_hd__a31o_1 _3282_ (.A1(_1058_),
    .A2(_1037_),
    .A3(_1038_),
    .B1(_0805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1059_));
 sky130_fd_sc_hd__o21ba_1 _3283_ (.A1(net50),
    .A2(_1055_),
    .B1_N(_1059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0118_));
 sky130_fd_sc_hd__a31o_1 _3284_ (.A1(_1058_),
    .A2(_1021_),
    .A3(_1032_),
    .B1(\genblk1[4].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1060_));
 sky130_fd_sc_hd__nand4_1 _3285_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[10] ),
    .B(_1058_),
    .C(_1037_),
    .D(_1038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1061_));
 sky130_fd_sc_hd__and3_1 _3286_ (.A(_0751_),
    .B(_1060_),
    .C(_1061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1062_));
 sky130_fd_sc_hd__clkbuf_1 _3287_ (.A(_1062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0119_));
 sky130_fd_sc_hd__inv_2 _3288_ (.A(net112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1063_));
 sky130_fd_sc_hd__and2_1 _3289_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[11] ),
    .B(\genblk1[4].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1064_));
 sky130_fd_sc_hd__and4_1 _3290_ (.A(_1064_),
    .B(_1058_),
    .C(_1037_),
    .D(_1038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1065_));
 sky130_fd_sc_hd__a211oi_1 _3291_ (.A1(_1063_),
    .A2(_1061_),
    .B1(_1065_),
    .C1(_0814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0120_));
 sky130_fd_sc_hd__a41o_1 _3292_ (.A1(_1013_),
    .A2(_1058_),
    .A3(_1037_),
    .A4(_1038_),
    .B1(_0813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1066_));
 sky130_fd_sc_hd__o21ba_1 _3293_ (.A1(net59),
    .A2(_1065_),
    .B1_N(_1066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0121_));
 sky130_fd_sc_hd__and4_1 _3294_ (.A(_1013_),
    .B(_1058_),
    .C(_1037_),
    .D(_1038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1067_));
 sky130_fd_sc_hd__nand4_1 _3295_ (.A(_1014_),
    .B(_1058_),
    .C(_1037_),
    .D(_1038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1068_));
 sky130_fd_sc_hd__o211a_1 _3296_ (.A1(net125),
    .A2(_1067_),
    .B1(_1068_),
    .C1(_1007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0122_));
 sky130_fd_sc_hd__inv_2 _3297_ (.A(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1069_));
 sky130_fd_sc_hd__and3_1 _3298_ (.A(_1019_),
    .B(_1037_),
    .C(_1038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1070_));
 sky130_fd_sc_hd__a211oi_1 _3299_ (.A1(_1069_),
    .A2(_1068_),
    .B1(_1070_),
    .C1(_0814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0123_));
 sky130_fd_sc_hd__a31o_1 _3300_ (.A1(_1019_),
    .A2(_1021_),
    .A3(_1032_),
    .B1(\genblk1[4].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1071_));
 sky130_fd_sc_hd__nand4_1 _3301_ (.A(\genblk1[4].puf_buffer.cnt_2.ctr[15] ),
    .B(_1019_),
    .C(_1037_),
    .D(_1038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1072_));
 sky130_fd_sc_hd__and3_1 _3302_ (.A(_0751_),
    .B(_1071_),
    .C(_1072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1073_));
 sky130_fd_sc_hd__clkbuf_1 _3303_ (.A(_1073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0124_));
 sky130_fd_sc_hd__and4_1 _3304_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[3] ),
    .B(\genblk1[4].puf_buffer.cnt_1.ctr[2] ),
    .C(\genblk1[4].puf_buffer.cnt_1.ctr[1] ),
    .D(\genblk1[4].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1074_));
 sky130_fd_sc_hd__and2_1 _3305_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[4].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1075_));
 sky130_fd_sc_hd__and4_1 _3306_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[4].puf_buffer.cnt_1.ctr[4] ),
    .C(_1074_),
    .D(_1075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1076_));
 sky130_fd_sc_hd__and3_1 _3307_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[9] ),
    .B(\genblk1[4].puf_buffer.cnt_1.ctr[8] ),
    .C(_1076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1077_));
 sky130_fd_sc_hd__and3_1 _3308_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[12] ),
    .B(\genblk1[4].puf_buffer.cnt_1.ctr[11] ),
    .C(\genblk1[4].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1078_));
 sky130_fd_sc_hd__and2_1 _3309_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[13] ),
    .B(_1078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1079_));
 sky130_fd_sc_hd__and3_1 _3310_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[14] ),
    .B(_1077_),
    .C(_1079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1080_));
 sky130_fd_sc_hd__a22o_1 _3311_ (.A1(_0670_),
    .A2(net137),
    .B1(_1080_),
    .B2(\genblk1[4].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0125_));
 sky130_fd_sc_hd__or2_2 _3312_ (.A(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1081_));
 sky130_fd_sc_hd__a22o_1 _3313_ (.A1(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .A2(_0688_),
    .B1(_0709_),
    .B2(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1082_));
 sky130_fd_sc_hd__a221o_1 _3314_ (.A1(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .A2(_0687_),
    .B1(net14),
    .B2(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .C1(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1083_));
 sky130_fd_sc_hd__a211o_1 _3315_ (.A1(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .A2(_0706_),
    .B1(_1082_),
    .C1(_1083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1084_));
 sky130_fd_sc_hd__a22o_1 _3316_ (.A1(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .A2(_0700_),
    .B1(_0690_),
    .B2(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1085_));
 sky130_fd_sc_hd__a221o_1 _3317_ (.A1(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .A2(net24),
    .B1(_0702_),
    .B2(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .C1(_1085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1086_));
 sky130_fd_sc_hd__a22o_1 _3318_ (.A1(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .A2(_0699_),
    .B1(_0694_),
    .B2(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1087_));
 sky130_fd_sc_hd__a22o_1 _3319_ (.A1(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .A2(_0689_),
    .B1(net11),
    .B2(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1088_));
 sky130_fd_sc_hd__a22o_1 _3320_ (.A1(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .A2(_0705_),
    .B1(_0695_),
    .B2(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1089_));
 sky130_fd_sc_hd__or3_1 _3321_ (.A(_1087_),
    .B(_1088_),
    .C(_1089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1090_));
 sky130_fd_sc_hd__or3_4 _3322_ (.A(_1084_),
    .B(_1086_),
    .C(_1090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1091_));
 sky130_fd_sc_hd__and3_1 _3323_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[0] ),
    .B(_1081_),
    .C(_1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1092_));
 sky130_fd_sc_hd__buf_2 _3324_ (.A(_1081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1093_));
 sky130_fd_sc_hd__buf_2 _3325_ (.A(_1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1094_));
 sky130_fd_sc_hd__a21o_1 _3326_ (.A1(_1093_),
    .A2(_1094_),
    .B1(\genblk1[4].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1095_));
 sky130_fd_sc_hd__and3b_1 _3327_ (.A_N(_1092_),
    .B(_1050_),
    .C(_1095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1096_));
 sky130_fd_sc_hd__clkbuf_1 _3328_ (.A(_1096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0126_));
 sky130_fd_sc_hd__nand2_1 _3329_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[1] ),
    .B(\genblk1[4].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1097_));
 sky130_fd_sc_hd__nand2_2 _3330_ (.A(_1093_),
    .B(_1094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1098_));
 sky130_fd_sc_hd__o221a_1 _3331_ (.A1(_1097_),
    .A2(_1098_),
    .B1(_1092_),
    .B2(net212),
    .C1(_0917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0127_));
 sky130_fd_sc_hd__inv_2 _3332_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1099_));
 sky130_fd_sc_hd__and4bb_1 _3333_ (.A_N(_1099_),
    .B_N(_1097_),
    .C(_1081_),
    .D(_1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1100_));
 sky130_fd_sc_hd__a41o_1 _3334_ (.A1(\genblk1[4].puf_buffer.cnt_1.ctr[1] ),
    .A2(\genblk1[4].puf_buffer.cnt_1.ctr[0] ),
    .A3(_1081_),
    .A4(_1091_),
    .B1(\genblk1[4].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1101_));
 sky130_fd_sc_hd__and3b_1 _3335_ (.A_N(_1100_),
    .B(_1050_),
    .C(_1101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1102_));
 sky130_fd_sc_hd__clkbuf_1 _3336_ (.A(_1102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0128_));
 sky130_fd_sc_hd__inv_2 _3337_ (.A(_1074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1103_));
 sky130_fd_sc_hd__clkbuf_4 _3338_ (.A(_0638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1104_));
 sky130_fd_sc_hd__o221a_1 _3339_ (.A1(_1103_),
    .A2(_1098_),
    .B1(_1100_),
    .B2(net116),
    .C1(_1104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0129_));
 sky130_fd_sc_hd__and4_1 _3340_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[4] ),
    .B(_1074_),
    .C(_1081_),
    .D(_1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1105_));
 sky130_fd_sc_hd__a31o_1 _3341_ (.A1(_1074_),
    .A2(_1093_),
    .A3(_1094_),
    .B1(\genblk1[4].puf_buffer.cnt_1.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1106_));
 sky130_fd_sc_hd__and3b_1 _3342_ (.A_N(_1105_),
    .B(_1050_),
    .C(_1106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1107_));
 sky130_fd_sc_hd__clkbuf_1 _3343_ (.A(_1107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0130_));
 sky130_fd_sc_hd__and3_1 _3344_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[4].puf_buffer.cnt_1.ctr[4] ),
    .C(_1074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1108_));
 sky130_fd_sc_hd__inv_2 _3345_ (.A(_1108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1109_));
 sky130_fd_sc_hd__o221a_1 _3346_ (.A1(_1109_),
    .A2(_1098_),
    .B1(_1105_),
    .B2(net175),
    .C1(_1104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0131_));
 sky130_fd_sc_hd__and4_1 _3347_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[6] ),
    .B(_1108_),
    .C(_1081_),
    .D(_1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1110_));
 sky130_fd_sc_hd__a31o_1 _3348_ (.A1(_1108_),
    .A2(_1093_),
    .A3(_1094_),
    .B1(\genblk1[4].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1111_));
 sky130_fd_sc_hd__and3b_1 _3349_ (.A_N(_1110_),
    .B(_1050_),
    .C(_1111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1112_));
 sky130_fd_sc_hd__clkbuf_1 _3350_ (.A(_1112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0132_));
 sky130_fd_sc_hd__inv_2 _3351_ (.A(_1076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1113_));
 sky130_fd_sc_hd__o221a_1 _3352_ (.A1(_1113_),
    .A2(_1098_),
    .B1(_1110_),
    .B2(net102),
    .C1(_1104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0133_));
 sky130_fd_sc_hd__and4_1 _3353_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[8] ),
    .B(_1076_),
    .C(_1081_),
    .D(_1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1114_));
 sky130_fd_sc_hd__a31o_1 _3354_ (.A1(_1076_),
    .A2(_1093_),
    .A3(_1094_),
    .B1(\genblk1[4].puf_buffer.cnt_1.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1115_));
 sky130_fd_sc_hd__and3b_1 _3355_ (.A_N(_1114_),
    .B(_1050_),
    .C(_1115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1116_));
 sky130_fd_sc_hd__clkbuf_1 _3356_ (.A(_1116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0134_));
 sky130_fd_sc_hd__nand3_1 _3357_ (.A(_1077_),
    .B(_1093_),
    .C(_1094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1117_));
 sky130_fd_sc_hd__o211a_1 _3358_ (.A1(net141),
    .A2(_1114_),
    .B1(_1117_),
    .C1(_1007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0135_));
 sky130_fd_sc_hd__and4_1 _3359_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[10] ),
    .B(_1077_),
    .C(_1081_),
    .D(_1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1118_));
 sky130_fd_sc_hd__a31o_1 _3360_ (.A1(_1077_),
    .A2(_1093_),
    .A3(_1094_),
    .B1(\genblk1[4].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1119_));
 sky130_fd_sc_hd__and3b_1 _3361_ (.A_N(_1118_),
    .B(_1050_),
    .C(_1119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1120_));
 sky130_fd_sc_hd__clkbuf_1 _3362_ (.A(_1120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0136_));
 sky130_fd_sc_hd__nand2_1 _3363_ (.A(net195),
    .B(\genblk1[4].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1121_));
 sky130_fd_sc_hd__o221a_1 _3364_ (.A1(_1121_),
    .A2(_1117_),
    .B1(_1118_),
    .B2(net195),
    .C1(_1104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0137_));
 sky130_fd_sc_hd__inv_2 _3365_ (.A(_1078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1122_));
 sky130_fd_sc_hd__and2_1 _3366_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[11] ),
    .B(\genblk1[4].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1123_));
 sky130_fd_sc_hd__a41o_1 _3367_ (.A1(_1077_),
    .A2(_1123_),
    .A3(_1093_),
    .A4(_1094_),
    .B1(net211),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1124_));
 sky130_fd_sc_hd__o211a_1 _3368_ (.A1(_1122_),
    .A2(_1117_),
    .B1(_1124_),
    .C1(_1007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0138_));
 sky130_fd_sc_hd__and4_1 _3369_ (.A(_1077_),
    .B(_1079_),
    .C(_1081_),
    .D(_1091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1125_));
 sky130_fd_sc_hd__a41o_1 _3370_ (.A1(_1077_),
    .A2(_1078_),
    .A3(_1081_),
    .A4(_1091_),
    .B1(\genblk1[4].puf_buffer.cnt_1.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1126_));
 sky130_fd_sc_hd__and3b_1 _3371_ (.A_N(_1125_),
    .B(_1050_),
    .C(_1126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1127_));
 sky130_fd_sc_hd__clkbuf_1 _3372_ (.A(_1127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0139_));
 sky130_fd_sc_hd__inv_2 _3373_ (.A(_1080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1128_));
 sky130_fd_sc_hd__o221a_1 _3374_ (.A1(_1128_),
    .A2(_1098_),
    .B1(_1125_),
    .B2(net122),
    .C1(_1104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0140_));
 sky130_fd_sc_hd__buf_2 _3375_ (.A(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1129_));
 sky130_fd_sc_hd__nand4_1 _3376_ (.A(\genblk1[4].puf_buffer.cnt_1.ctr[15] ),
    .B(_1080_),
    .C(_1093_),
    .D(_1094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1130_));
 sky130_fd_sc_hd__a31o_1 _3377_ (.A1(_1080_),
    .A2(_1093_),
    .A3(_1094_),
    .B1(\genblk1[4].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1131_));
 sky130_fd_sc_hd__and3_1 _3378_ (.A(_1129_),
    .B(_1130_),
    .C(_1131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _3379_ (.A(_1132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0141_));
 sky130_fd_sc_hd__inv_2 _3380_ (.A(net169),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1133_));
 sky130_fd_sc_hd__and3b_1 _3381_ (.A_N(\genblk1[5].puf_buffer.cnt_1.finish ),
    .B(\genblk1[5].puf_buffer.cnt_2.finish ),
    .C(_0437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1134_));
 sky130_fd_sc_hd__clkbuf_1 _3382_ (.A(_1134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0179_));
 sky130_fd_sc_hd__o21bai_1 _3383_ (.A1(_1133_),
    .A2(_0179_),
    .B1_N(\genblk1[5].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_0142_));
 sky130_fd_sc_hd__and4_1 _3384_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[3] ),
    .B(\genblk1[5].puf_buffer.cnt_2.ctr[2] ),
    .C(\genblk1[5].puf_buffer.cnt_2.ctr[1] ),
    .D(\genblk1[5].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1135_));
 sky130_fd_sc_hd__and2_1 _3385_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[7] ),
    .B(\genblk1[5].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1136_));
 sky130_fd_sc_hd__and4_1 _3386_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[5].puf_buffer.cnt_2.ctr[4] ),
    .C(_1135_),
    .D(_1136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1137_));
 sky130_fd_sc_hd__and3_2 _3387_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[9] ),
    .B(\genblk1[5].puf_buffer.cnt_2.ctr[8] ),
    .C(_1137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1138_));
 sky130_fd_sc_hd__and3_1 _3388_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[12] ),
    .B(\genblk1[5].puf_buffer.cnt_2.ctr[11] ),
    .C(\genblk1[5].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1139_));
 sky130_fd_sc_hd__and2_1 _3389_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[13] ),
    .B(_1139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1140_));
 sky130_fd_sc_hd__and3_1 _3390_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[14] ),
    .B(_1138_),
    .C(_1140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1141_));
 sky130_fd_sc_hd__a22o_1 _3391_ (.A1(_0670_),
    .A2(\genblk1[5].puf_buffer.cnt_2.finish ),
    .B1(_1141_),
    .B2(net153),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0144_));
 sky130_fd_sc_hd__or2_1 _3392_ (.A(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[7] ),
    .B(_0601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1142_));
 sky130_fd_sc_hd__clkbuf_2 _3393_ (.A(_1142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1143_));
 sky130_fd_sc_hd__a22o_1 _3394_ (.A1(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[7] ),
    .A2(_0618_),
    .B1(_0624_),
    .B2(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1144_));
 sky130_fd_sc_hd__a221o_1 _3395_ (.A1(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[7] ),
    .A2(_0603_),
    .B1(_0604_),
    .B2(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[7] ),
    .C1(_1144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1145_));
 sky130_fd_sc_hd__a22o_1 _3396_ (.A1(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[7] ),
    .A2(_0615_),
    .B1(net19),
    .B2(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1146_));
 sky130_fd_sc_hd__a211o_1 _3397_ (.A1(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[7] ),
    .A2(_0610_),
    .B1(_1146_),
    .C1(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1147_));
 sky130_fd_sc_hd__a22o_1 _3398_ (.A1(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[7] ),
    .A2(_0611_),
    .B1(net17),
    .B2(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1148_));
 sky130_fd_sc_hd__a22o_1 _3399_ (.A1(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[7] ),
    .A2(_0622_),
    .B1(net26),
    .B2(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1149_));
 sky130_fd_sc_hd__a22o_1 _3400_ (.A1(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[7] ),
    .A2(_0605_),
    .B1(_0606_),
    .B2(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1150_));
 sky130_fd_sc_hd__a22o_1 _3401_ (.A1(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[7] ),
    .A2(_0621_),
    .B1(_0625_),
    .B2(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1151_));
 sky130_fd_sc_hd__or4_1 _3402_ (.A(_1148_),
    .B(_1149_),
    .C(_1150_),
    .D(_1151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1152_));
 sky130_fd_sc_hd__or3_2 _3403_ (.A(_1145_),
    .B(_1147_),
    .C(_1152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1153_));
 sky130_fd_sc_hd__clkbuf_2 _3404_ (.A(_1153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1154_));
 sky130_fd_sc_hd__and3_1 _3405_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[0] ),
    .B(_1143_),
    .C(_1154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1155_));
 sky130_fd_sc_hd__buf_2 _3406_ (.A(_1142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1156_));
 sky130_fd_sc_hd__buf_2 _3407_ (.A(_1153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1157_));
 sky130_fd_sc_hd__a21o_1 _3408_ (.A1(_1156_),
    .A2(_1157_),
    .B1(\genblk1[5].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1158_));
 sky130_fd_sc_hd__and3b_1 _3409_ (.A_N(_1155_),
    .B(_1050_),
    .C(_1158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1159_));
 sky130_fd_sc_hd__clkbuf_1 _3410_ (.A(_1159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0145_));
 sky130_fd_sc_hd__nand2_1 _3411_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[1] ),
    .B(\genblk1[5].puf_buffer.cnt_2.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1160_));
 sky130_fd_sc_hd__nand2_1 _3412_ (.A(_1156_),
    .B(_1157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1161_));
 sky130_fd_sc_hd__o221a_1 _3413_ (.A1(_1160_),
    .A2(_1161_),
    .B1(_1155_),
    .B2(net217),
    .C1(_1104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0146_));
 sky130_fd_sc_hd__inv_2 _3414_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1162_));
 sky130_fd_sc_hd__and4bb_1 _3415_ (.A_N(_1162_),
    .B_N(_1160_),
    .C(_1142_),
    .D(_1153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1163_));
 sky130_fd_sc_hd__clkbuf_2 _3416_ (.A(_0630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1164_));
 sky130_fd_sc_hd__a41o_1 _3417_ (.A1(\genblk1[5].puf_buffer.cnt_2.ctr[1] ),
    .A2(\genblk1[5].puf_buffer.cnt_2.ctr[0] ),
    .A3(_1143_),
    .A4(_1154_),
    .B1(\genblk1[5].puf_buffer.cnt_2.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1165_));
 sky130_fd_sc_hd__and3b_1 _3418_ (.A_N(_1163_),
    .B(_1164_),
    .C(_1165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1166_));
 sky130_fd_sc_hd__clkbuf_1 _3419_ (.A(_1166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0147_));
 sky130_fd_sc_hd__inv_2 _3420_ (.A(_1135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1167_));
 sky130_fd_sc_hd__o221a_1 _3421_ (.A1(_1167_),
    .A2(_1161_),
    .B1(_1163_),
    .B2(net134),
    .C1(_1104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0148_));
 sky130_fd_sc_hd__and4_1 _3422_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[4] ),
    .B(_1135_),
    .C(_1143_),
    .D(_1154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1168_));
 sky130_fd_sc_hd__a31o_1 _3423_ (.A1(_1135_),
    .A2(_1156_),
    .A3(_1157_),
    .B1(\genblk1[5].puf_buffer.cnt_2.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1169_));
 sky130_fd_sc_hd__and3b_1 _3424_ (.A_N(_1168_),
    .B(_1164_),
    .C(_1169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1170_));
 sky130_fd_sc_hd__clkbuf_1 _3425_ (.A(_1170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0149_));
 sky130_fd_sc_hd__and3_1 _3426_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[5] ),
    .B(\genblk1[5].puf_buffer.cnt_2.ctr[4] ),
    .C(_1135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1171_));
 sky130_fd_sc_hd__inv_2 _3427_ (.A(_1171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1172_));
 sky130_fd_sc_hd__o221a_1 _3428_ (.A1(_1172_),
    .A2(_1161_),
    .B1(_1168_),
    .B2(net173),
    .C1(_1104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0150_));
 sky130_fd_sc_hd__and4_1 _3429_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[6] ),
    .B(_1171_),
    .C(_1143_),
    .D(_1154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1173_));
 sky130_fd_sc_hd__a31o_1 _3430_ (.A1(_1171_),
    .A2(_1156_),
    .A3(_1157_),
    .B1(\genblk1[5].puf_buffer.cnt_2.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1174_));
 sky130_fd_sc_hd__and3b_1 _3431_ (.A_N(_1173_),
    .B(_1164_),
    .C(_1174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1175_));
 sky130_fd_sc_hd__clkbuf_1 _3432_ (.A(_1175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0151_));
 sky130_fd_sc_hd__inv_2 _3433_ (.A(_1137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1176_));
 sky130_fd_sc_hd__o221a_1 _3434_ (.A1(_1176_),
    .A2(_1161_),
    .B1(_1173_),
    .B2(net104),
    .C1(_1104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0152_));
 sky130_fd_sc_hd__and4_1 _3435_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[8] ),
    .B(_1137_),
    .C(_1143_),
    .D(_1154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1177_));
 sky130_fd_sc_hd__a31o_1 _3436_ (.A1(_1137_),
    .A2(_1156_),
    .A3(_1157_),
    .B1(\genblk1[5].puf_buffer.cnt_2.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1178_));
 sky130_fd_sc_hd__and3b_1 _3437_ (.A_N(_1177_),
    .B(_1164_),
    .C(_1178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1179_));
 sky130_fd_sc_hd__clkbuf_1 _3438_ (.A(_1179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0153_));
 sky130_fd_sc_hd__nand3_1 _3439_ (.A(_1138_),
    .B(_1156_),
    .C(_1157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1180_));
 sky130_fd_sc_hd__o211a_1 _3440_ (.A1(net156),
    .A2(_1177_),
    .B1(_1180_),
    .C1(_1007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0154_));
 sky130_fd_sc_hd__and4_1 _3441_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[10] ),
    .B(_1138_),
    .C(_1143_),
    .D(_1154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1181_));
 sky130_fd_sc_hd__a31o_1 _3442_ (.A1(_1138_),
    .A2(_1156_),
    .A3(_1154_),
    .B1(\genblk1[5].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1182_));
 sky130_fd_sc_hd__and3b_1 _3443_ (.A_N(_1181_),
    .B(_1164_),
    .C(_1182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1183_));
 sky130_fd_sc_hd__clkbuf_1 _3444_ (.A(_1183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0155_));
 sky130_fd_sc_hd__nand2_1 _3445_ (.A(net207),
    .B(\genblk1[5].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1184_));
 sky130_fd_sc_hd__o221a_1 _3446_ (.A1(_1184_),
    .A2(_1180_),
    .B1(_1181_),
    .B2(net207),
    .C1(_1104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0156_));
 sky130_fd_sc_hd__a41o_1 _3447_ (.A1(_1138_),
    .A2(_1139_),
    .A3(_1143_),
    .A4(_1157_),
    .B1(_0804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1185_));
 sky130_fd_sc_hd__and2_1 _3448_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[11] ),
    .B(\genblk1[5].puf_buffer.cnt_2.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1186_));
 sky130_fd_sc_hd__a41o_1 _3449_ (.A1(_1138_),
    .A2(_1186_),
    .A3(_1143_),
    .A4(_1154_),
    .B1(\genblk1[5].puf_buffer.cnt_2.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1187_));
 sky130_fd_sc_hd__and2b_1 _3450_ (.A_N(_1185_),
    .B(_1187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1188_));
 sky130_fd_sc_hd__clkbuf_1 _3451_ (.A(_1188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0157_));
 sky130_fd_sc_hd__and4_1 _3452_ (.A(_1138_),
    .B(_1140_),
    .C(_1143_),
    .D(_1154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1189_));
 sky130_fd_sc_hd__a41o_1 _3453_ (.A1(_1138_),
    .A2(_1139_),
    .A3(_1143_),
    .A4(_1154_),
    .B1(\genblk1[5].puf_buffer.cnt_2.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1190_));
 sky130_fd_sc_hd__and3b_1 _3454_ (.A_N(_1189_),
    .B(_1164_),
    .C(_1190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1191_));
 sky130_fd_sc_hd__clkbuf_1 _3455_ (.A(_1191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0158_));
 sky130_fd_sc_hd__nand3_1 _3456_ (.A(_1141_),
    .B(_1156_),
    .C(_1157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1192_));
 sky130_fd_sc_hd__o211a_1 _3457_ (.A1(net136),
    .A2(_1189_),
    .B1(_1192_),
    .C1(_1007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0159_));
 sky130_fd_sc_hd__a31o_1 _3458_ (.A1(_1141_),
    .A2(_1156_),
    .A3(_1157_),
    .B1(\genblk1[5].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1193_));
 sky130_fd_sc_hd__nand4_1 _3459_ (.A(\genblk1[5].puf_buffer.cnt_2.ctr[15] ),
    .B(_1141_),
    .C(_1156_),
    .D(_1157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1194_));
 sky130_fd_sc_hd__and3_1 _3460_ (.A(_1129_),
    .B(_1193_),
    .C(_1194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1195_));
 sky130_fd_sc_hd__clkbuf_1 _3461_ (.A(_1195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0160_));
 sky130_fd_sc_hd__and4_1 _3462_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[3] ),
    .B(\genblk1[5].puf_buffer.cnt_1.ctr[2] ),
    .C(\genblk1[5].puf_buffer.cnt_1.ctr[1] ),
    .D(\genblk1[5].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1196_));
 sky130_fd_sc_hd__and2_1 _3463_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[7] ),
    .B(\genblk1[5].puf_buffer.cnt_1.ctr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1197_));
 sky130_fd_sc_hd__and4_1 _3464_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[5] ),
    .B(\genblk1[5].puf_buffer.cnt_1.ctr[4] ),
    .C(_1196_),
    .D(_1197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1198_));
 sky130_fd_sc_hd__and3_2 _3465_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[9] ),
    .B(\genblk1[5].puf_buffer.cnt_1.ctr[8] ),
    .C(_1198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1199_));
 sky130_fd_sc_hd__and3_1 _3466_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[12] ),
    .B(\genblk1[5].puf_buffer.cnt_1.ctr[11] ),
    .C(\genblk1[5].puf_buffer.cnt_1.ctr[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1200_));
 sky130_fd_sc_hd__and2_1 _3467_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[13] ),
    .B(_1200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1201_));
 sky130_fd_sc_hd__and3_1 _3468_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[14] ),
    .B(_1199_),
    .C(_1201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1202_));
 sky130_fd_sc_hd__a22o_1 _3469_ (.A1(_0670_),
    .A2(net157),
    .B1(_1202_),
    .B2(\genblk1[5].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0161_));
 sky130_fd_sc_hd__or2_2 _3470_ (.A(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[7] ),
    .B(_0685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1203_));
 sky130_fd_sc_hd__a22o_1 _3471_ (.A1(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[7] ),
    .A2(_0706_),
    .B1(_0709_),
    .B2(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1204_));
 sky130_fd_sc_hd__a221o_1 _3472_ (.A1(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[7] ),
    .A2(_0688_),
    .B1(net11),
    .B2(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[7] ),
    .C1(_0697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1205_));
 sky130_fd_sc_hd__a211o_1 _3473_ (.A1(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[7] ),
    .A2(_0687_),
    .B1(_1204_),
    .C1(_1205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1206_));
 sky130_fd_sc_hd__a22o_1 _3474_ (.A1(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[7] ),
    .A2(_0695_),
    .B1(net231),
    .B2(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1207_));
 sky130_fd_sc_hd__a21o_1 _3475_ (.A1(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[7] ),
    .A2(_0699_),
    .B1(_1207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1208_));
 sky130_fd_sc_hd__a22o_1 _3476_ (.A1(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[7] ),
    .A2(_0694_),
    .B1(_0705_),
    .B2(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1209_));
 sky130_fd_sc_hd__a22o_1 _3477_ (.A1(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[7] ),
    .A2(_0700_),
    .B1(_0690_),
    .B2(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1210_));
 sky130_fd_sc_hd__a22o_1 _3478_ (.A1(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[7] ),
    .A2(_0702_),
    .B1(_0693_),
    .B2(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1211_));
 sky130_fd_sc_hd__a2111o_1 _3479_ (.A1(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[7] ),
    .A2(_0689_),
    .B1(_1209_),
    .C1(_1210_),
    .D1(_1211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1212_));
 sky130_fd_sc_hd__or3_4 _3480_ (.A(_1206_),
    .B(_1208_),
    .C(_1212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1213_));
 sky130_fd_sc_hd__and3_1 _3481_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[0] ),
    .B(_1203_),
    .C(_1213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1214_));
 sky130_fd_sc_hd__buf_2 _3482_ (.A(_1203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1215_));
 sky130_fd_sc_hd__buf_2 _3483_ (.A(_1213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1216_));
 sky130_fd_sc_hd__a21o_1 _3484_ (.A1(_1215_),
    .A2(_1216_),
    .B1(\genblk1[5].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1217_));
 sky130_fd_sc_hd__and3b_1 _3485_ (.A_N(_1214_),
    .B(_1164_),
    .C(_1217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1218_));
 sky130_fd_sc_hd__clkbuf_1 _3486_ (.A(_1218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0162_));
 sky130_fd_sc_hd__nand2_1 _3487_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[1] ),
    .B(\genblk1[5].puf_buffer.cnt_1.ctr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1219_));
 sky130_fd_sc_hd__nand2_2 _3488_ (.A(_1215_),
    .B(_1216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1220_));
 sky130_fd_sc_hd__buf_2 _3489_ (.A(_0638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1221_));
 sky130_fd_sc_hd__o221a_1 _3490_ (.A1(_1219_),
    .A2(_1220_),
    .B1(_1214_),
    .B2(net227),
    .C1(_1221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0163_));
 sky130_fd_sc_hd__inv_2 _3491_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1222_));
 sky130_fd_sc_hd__and4bb_1 _3492_ (.A_N(_1222_),
    .B_N(_1219_),
    .C(_1203_),
    .D(_1213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1223_));
 sky130_fd_sc_hd__a41o_1 _3493_ (.A1(\genblk1[5].puf_buffer.cnt_1.ctr[1] ),
    .A2(\genblk1[5].puf_buffer.cnt_1.ctr[0] ),
    .A3(_1203_),
    .A4(_1213_),
    .B1(\genblk1[5].puf_buffer.cnt_1.ctr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1224_));
 sky130_fd_sc_hd__and3b_1 _3494_ (.A_N(_1223_),
    .B(_1164_),
    .C(_1224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1225_));
 sky130_fd_sc_hd__clkbuf_1 _3495_ (.A(_1225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0164_));
 sky130_fd_sc_hd__inv_2 _3496_ (.A(_1196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_1226_));
 sky130_fd_sc_hd__o221a_1 _3497_ (.A1(_1226_),
    .A2(_1220_),
    .B1(_1223_),
    .B2(net114),
    .C1(_1221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_0165_));
 sky130_fd_sc_hd__and4_1 _3498_ (.A(\genblk1[5].puf_buffer.cnt_1.ctr[4] ),
    .B(_1196_),
    .C(_1203_),
    .D(_1213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1227_));
 sky130_fd_sc_hd__a31o_1 _3499_ (.A1(_1196_),
    .A2(_1215_),
    .A3(_1216_),
    .B1(\genblk1[5].puf_buffer.cnt_1.ctr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_1228_));
 sky130_fd_sc_hd__dfxtp_1 _3500_ (.CLK(clknet_leaf_11_clk),
    .D(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3501_ (.CLK(clknet_leaf_11_clk),
    .D(_0001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3502_ (.CLK(clknet_leaf_12_clk),
    .D(_0002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3503_ (.CLK(clknet_leaf_12_clk),
    .D(_0003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3504_ (.CLK(clknet_leaf_12_clk),
    .D(_0004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3505_ (.CLK(clknet_leaf_12_clk),
    .D(_0005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3506_ (.CLK(clknet_leaf_12_clk),
    .D(_0006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3507_ (.CLK(clknet_leaf_12_clk),
    .D(_0007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3508_ (.CLK(clknet_leaf_12_clk),
    .D(_0008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3509_ (.CLK(clknet_leaf_12_clk),
    .D(_0009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3510_ (.CLK(clknet_leaf_12_clk),
    .D(_0010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3511_ (.CLK(clknet_leaf_11_clk),
    .D(_0011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3512_ (.CLK(clknet_leaf_11_clk),
    .D(_0012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3513_ (.CLK(clknet_leaf_11_clk),
    .D(_0013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3514_ (.CLK(clknet_leaf_12_clk),
    .D(_0014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3515_ (.CLK(clknet_leaf_12_clk),
    .D(_0015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3516_ (.CLK(clknet_leaf_11_clk),
    .D(_0016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_2.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3517_ (.CLK(clknet_leaf_9_clk),
    .D(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3518_ (.CLK(clknet_leaf_10_clk),
    .D(_0018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3519_ (.CLK(clknet_leaf_9_clk),
    .D(net224),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3520_ (.CLK(clknet_leaf_10_clk),
    .D(_0020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3521_ (.CLK(clknet_leaf_9_clk),
    .D(_0021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3522_ (.CLK(clknet_leaf_9_clk),
    .D(_0022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3523_ (.CLK(clknet_leaf_9_clk),
    .D(_0023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3524_ (.CLK(clknet_leaf_9_clk),
    .D(_0024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3525_ (.CLK(clknet_leaf_9_clk),
    .D(_0025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3526_ (.CLK(clknet_leaf_9_clk),
    .D(_0026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3527_ (.CLK(clknet_leaf_9_clk),
    .D(_0027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3528_ (.CLK(clknet_leaf_9_clk),
    .D(_0028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3529_ (.CLK(clknet_leaf_9_clk),
    .D(_0029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3530_ (.CLK(clknet_leaf_9_clk),
    .D(_0030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3531_ (.CLK(clknet_leaf_9_clk),
    .D(_0031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3532_ (.CLK(clknet_leaf_10_clk),
    .D(_0032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3533_ (.CLK(clknet_leaf_9_clk),
    .D(_0033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.cnt_1.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3534_ (.CLK(clknet_leaf_8_clk),
    .D(_0034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.race_arb.resp ));
 sky130_fd_sc_hd__dfxtp_1 _3535_ (.CLK(clknet_leaf_9_clk),
    .D(_0035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.race_arb.marked_2 ));
 sky130_fd_sc_hd__dfxtp_1 _3536_ (.CLK(clknet_leaf_8_clk),
    .D(\genblk1[2].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.race_arb.marked_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3537_ (.CLK(clknet_leaf_10_clk),
    .D(net164),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3538_ (.CLK(clknet_leaf_11_clk),
    .D(_0037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3539_ (.CLK(clknet_leaf_10_clk),
    .D(_0038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3540_ (.CLK(clknet_leaf_10_clk),
    .D(_0039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3541_ (.CLK(clknet_leaf_9_clk),
    .D(_0040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3542_ (.CLK(clknet_leaf_10_clk),
    .D(_0041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3543_ (.CLK(clknet_leaf_9_clk),
    .D(_0042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3544_ (.CLK(clknet_leaf_11_clk),
    .D(_0043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3545_ (.CLK(clknet_leaf_11_clk),
    .D(_0044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3546_ (.CLK(clknet_leaf_11_clk),
    .D(_0045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3547_ (.CLK(clknet_leaf_11_clk),
    .D(_0046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3548_ (.CLK(clknet_leaf_10_clk),
    .D(_0047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3549_ (.CLK(clknet_leaf_11_clk),
    .D(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3550_ (.CLK(clknet_leaf_11_clk),
    .D(_0049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3551_ (.CLK(clknet_leaf_9_clk),
    .D(_0050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3552_ (.CLK(clknet_leaf_10_clk),
    .D(_0051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3553_ (.CLK(clknet_leaf_10_clk),
    .D(_0052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_2.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3554_ (.CLK(clknet_leaf_8_clk),
    .D(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3555_ (.CLK(clknet_leaf_10_clk),
    .D(_0054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3556_ (.CLK(clknet_leaf_9_clk),
    .D(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3557_ (.CLK(clknet_leaf_9_clk),
    .D(_0056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3558_ (.CLK(clknet_leaf_9_clk),
    .D(_0057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3559_ (.CLK(clknet_leaf_9_clk),
    .D(_0058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3560_ (.CLK(clknet_leaf_9_clk),
    .D(_0059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3561_ (.CLK(clknet_leaf_10_clk),
    .D(_0060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3562_ (.CLK(clknet_leaf_10_clk),
    .D(_0061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3563_ (.CLK(clknet_leaf_10_clk),
    .D(_0062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3564_ (.CLK(clknet_leaf_10_clk),
    .D(_0063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3565_ (.CLK(clknet_leaf_10_clk),
    .D(_0064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3566_ (.CLK(clknet_leaf_11_clk),
    .D(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3567_ (.CLK(clknet_leaf_11_clk),
    .D(_0066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3568_ (.CLK(clknet_leaf_10_clk),
    .D(_0067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3569_ (.CLK(clknet_leaf_10_clk),
    .D(_0068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3570_ (.CLK(clknet_leaf_8_clk),
    .D(_0069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.cnt_1.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3571_ (.CLK(clknet_leaf_1_clk),
    .D(_0070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.race_arb.resp ));
 sky130_fd_sc_hd__dfxtp_1 _3572_ (.CLK(clknet_leaf_8_clk),
    .D(_0071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[2].puf_buffer.race_arb.marked_2 ));
 sky130_fd_sc_hd__dfxtp_1 _3573_ (.CLK(clknet_leaf_1_clk),
    .D(\genblk1[3].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.race_arb.marked_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3574_ (.CLK(clknet_leaf_1_clk),
    .D(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3575_ (.CLK(clknet_leaf_10_clk),
    .D(_0073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3576_ (.CLK(clknet_leaf_11_clk),
    .D(net220),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3577_ (.CLK(clknet_leaf_11_clk),
    .D(_0075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3578_ (.CLK(clknet_leaf_11_clk),
    .D(_0076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3579_ (.CLK(clknet_leaf_11_clk),
    .D(_0077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3580_ (.CLK(clknet_leaf_11_clk),
    .D(_0078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3581_ (.CLK(clknet_leaf_11_clk),
    .D(_0079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3582_ (.CLK(clknet_leaf_11_clk),
    .D(_0080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3583_ (.CLK(clknet_leaf_1_clk),
    .D(_0081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3584_ (.CLK(clknet_leaf_1_clk),
    .D(_0082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3585_ (.CLK(clknet_leaf_11_clk),
    .D(_0083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3586_ (.CLK(clknet_leaf_0_clk),
    .D(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3587_ (.CLK(clknet_leaf_0_clk),
    .D(_0085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3588_ (.CLK(clknet_leaf_0_clk),
    .D(_0086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3589_ (.CLK(clknet_leaf_0_clk),
    .D(_0087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3590_ (.CLK(clknet_leaf_1_clk),
    .D(_0088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_2.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3591_ (.CLK(clknet_leaf_12_clk),
    .D(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3592_ (.CLK(clknet_leaf_12_clk),
    .D(_0090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3593_ (.CLK(clknet_leaf_12_clk),
    .D(_0091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3594_ (.CLK(clknet_leaf_12_clk),
    .D(_0092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3595_ (.CLK(clknet_leaf_12_clk),
    .D(_0093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3596_ (.CLK(clknet_leaf_12_clk),
    .D(_0094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3597_ (.CLK(clknet_leaf_12_clk),
    .D(_0095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3598_ (.CLK(clknet_leaf_12_clk),
    .D(_0096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3599_ (.CLK(clknet_leaf_12_clk),
    .D(_0097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3600_ (.CLK(clknet_leaf_12_clk),
    .D(_0098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3601_ (.CLK(clknet_leaf_12_clk),
    .D(_0099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3602_ (.CLK(clknet_leaf_0_clk),
    .D(_0100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3603_ (.CLK(clknet_leaf_0_clk),
    .D(_0101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3604_ (.CLK(clknet_leaf_0_clk),
    .D(_0102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3605_ (.CLK(clknet_leaf_0_clk),
    .D(_0103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3606_ (.CLK(clknet_leaf_0_clk),
    .D(_0104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3607_ (.CLK(clknet_leaf_0_clk),
    .D(_0105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.cnt_1.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3608_ (.CLK(clknet_leaf_1_clk),
    .D(_0106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.race_arb.resp ));
 sky130_fd_sc_hd__dfxtp_1 _3609_ (.CLK(clknet_leaf_1_clk),
    .D(_0107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[3].puf_buffer.race_arb.marked_2 ));
 sky130_fd_sc_hd__dfxtp_1 _3610_ (.CLK(clknet_leaf_1_clk),
    .D(\genblk1[4].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.race_arb.marked_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3611_ (.CLK(clknet_leaf_1_clk),
    .D(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3612_ (.CLK(clknet_leaf_0_clk),
    .D(_0109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3613_ (.CLK(clknet_leaf_0_clk),
    .D(_0110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3614_ (.CLK(clknet_leaf_0_clk),
    .D(_0111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3615_ (.CLK(clknet_leaf_0_clk),
    .D(_0112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3616_ (.CLK(clknet_leaf_0_clk),
    .D(_0113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3617_ (.CLK(clknet_leaf_0_clk),
    .D(_0114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3618_ (.CLK(clknet_leaf_0_clk),
    .D(_0115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3619_ (.CLK(clknet_leaf_0_clk),
    .D(_0116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3620_ (.CLK(clknet_leaf_0_clk),
    .D(_0117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3621_ (.CLK(clknet_leaf_0_clk),
    .D(_0118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3622_ (.CLK(clknet_leaf_0_clk),
    .D(_0119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3623_ (.CLK(clknet_leaf_1_clk),
    .D(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3624_ (.CLK(clknet_leaf_0_clk),
    .D(_0121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3625_ (.CLK(clknet_leaf_1_clk),
    .D(_0122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3626_ (.CLK(clknet_leaf_1_clk),
    .D(_0123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3627_ (.CLK(clknet_leaf_0_clk),
    .D(_0124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_2.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3628_ (.CLK(clknet_leaf_1_clk),
    .D(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3629_ (.CLK(clknet_leaf_2_clk),
    .D(_0126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3630_ (.CLK(clknet_leaf_1_clk),
    .D(net213),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3631_ (.CLK(clknet_leaf_0_clk),
    .D(_0128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3632_ (.CLK(clknet_leaf_2_clk),
    .D(_0129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3633_ (.CLK(clknet_leaf_2_clk),
    .D(_0130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3634_ (.CLK(clknet_leaf_2_clk),
    .D(_0131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3635_ (.CLK(clknet_leaf_2_clk),
    .D(_0132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3636_ (.CLK(clknet_leaf_2_clk),
    .D(_0133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3637_ (.CLK(clknet_leaf_2_clk),
    .D(_0134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3638_ (.CLK(clknet_leaf_2_clk),
    .D(_0135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3639_ (.CLK(clknet_leaf_2_clk),
    .D(_0136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3640_ (.CLK(clknet_leaf_2_clk),
    .D(_0137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3641_ (.CLK(clknet_leaf_2_clk),
    .D(_0138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3642_ (.CLK(clknet_leaf_2_clk),
    .D(_0139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3643_ (.CLK(clknet_leaf_1_clk),
    .D(_0140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3644_ (.CLK(clknet_leaf_1_clk),
    .D(_0141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.cnt_1.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3645_ (.CLK(clknet_leaf_4_clk),
    .D(_0142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.race_arb.resp ));
 sky130_fd_sc_hd__dfxtp_1 _3646_ (.CLK(clknet_leaf_1_clk),
    .D(_0143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[4].puf_buffer.race_arb.marked_2 ));
 sky130_fd_sc_hd__dfxtp_1 _3647_ (.CLK(clknet_leaf_4_clk),
    .D(\genblk1[5].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.race_arb.marked_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3648_ (.CLK(clknet_leaf_4_clk),
    .D(net154),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3649_ (.CLK(clknet_leaf_2_clk),
    .D(_0145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3650_ (.CLK(clknet_leaf_2_clk),
    .D(_0146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3651_ (.CLK(clknet_leaf_2_clk),
    .D(_0147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3652_ (.CLK(clknet_leaf_2_clk),
    .D(_0148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3653_ (.CLK(clknet_leaf_2_clk),
    .D(_0149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3654_ (.CLK(clknet_leaf_2_clk),
    .D(_0150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3655_ (.CLK(clknet_leaf_2_clk),
    .D(_0151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3656_ (.CLK(clknet_leaf_2_clk),
    .D(_0152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3657_ (.CLK(clknet_leaf_3_clk),
    .D(_0153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3658_ (.CLK(clknet_leaf_3_clk),
    .D(_0154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3659_ (.CLK(clknet_leaf_3_clk),
    .D(_0155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3660_ (.CLK(clknet_leaf_3_clk),
    .D(_0156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3661_ (.CLK(clknet_leaf_3_clk),
    .D(_0157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3662_ (.CLK(clknet_leaf_3_clk),
    .D(_0158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3663_ (.CLK(clknet_leaf_4_clk),
    .D(_0159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3664_ (.CLK(clknet_leaf_4_clk),
    .D(_0160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_2.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3665_ (.CLK(clknet_leaf_3_clk),
    .D(net158),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3666_ (.CLK(clknet_leaf_3_clk),
    .D(_0162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3667_ (.CLK(clknet_leaf_3_clk),
    .D(_0163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3668_ (.CLK(clknet_leaf_3_clk),
    .D(_0164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3669_ (.CLK(clknet_leaf_3_clk),
    .D(_0165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3670_ (.CLK(clknet_leaf_3_clk),
    .D(_0166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3671_ (.CLK(clknet_leaf_3_clk),
    .D(_0167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3672_ (.CLK(clknet_leaf_3_clk),
    .D(_0168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3673_ (.CLK(clknet_leaf_3_clk),
    .D(_0169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3674_ (.CLK(clknet_leaf_3_clk),
    .D(_0170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3675_ (.CLK(clknet_leaf_3_clk),
    .D(_0171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3676_ (.CLK(clknet_leaf_3_clk),
    .D(_0172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3677_ (.CLK(clknet_leaf_3_clk),
    .D(_0173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3678_ (.CLK(clknet_leaf_3_clk),
    .D(_0174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3679_ (.CLK(clknet_leaf_3_clk),
    .D(_0175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3680_ (.CLK(clknet_leaf_3_clk),
    .D(_0176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3681_ (.CLK(clknet_leaf_3_clk),
    .D(_0177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.cnt_1.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3682_ (.CLK(clknet_leaf_6_clk),
    .D(_0178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.race_arb.resp ));
 sky130_fd_sc_hd__dfxtp_1 _3683_ (.CLK(clknet_leaf_4_clk),
    .D(_0179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[5].puf_buffer.race_arb.marked_2 ));
 sky130_fd_sc_hd__dfxtp_1 _3684_ (.CLK(clknet_leaf_6_clk),
    .D(\genblk1[6].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.race_arb.marked_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3685_ (.CLK(clknet_leaf_4_clk),
    .D(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3686_ (.CLK(clknet_leaf_4_clk),
    .D(_0181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3687_ (.CLK(clknet_leaf_4_clk),
    .D(_0182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3688_ (.CLK(clknet_leaf_4_clk),
    .D(_0183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3689_ (.CLK(clknet_leaf_3_clk),
    .D(_0184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3690_ (.CLK(clknet_leaf_3_clk),
    .D(_0185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3691_ (.CLK(clknet_leaf_4_clk),
    .D(_0186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3692_ (.CLK(clknet_leaf_4_clk),
    .D(_0187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3693_ (.CLK(clknet_leaf_4_clk),
    .D(_0188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3694_ (.CLK(clknet_leaf_4_clk),
    .D(_0189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3695_ (.CLK(clknet_leaf_4_clk),
    .D(_0190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3696_ (.CLK(clknet_leaf_4_clk),
    .D(_0191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3697_ (.CLK(clknet_leaf_4_clk),
    .D(_0192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3698_ (.CLK(clknet_leaf_4_clk),
    .D(_0193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3699_ (.CLK(clknet_leaf_4_clk),
    .D(_0194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3700_ (.CLK(clknet_leaf_6_clk),
    .D(_0195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3701_ (.CLK(clknet_leaf_4_clk),
    .D(_0196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_2.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3702_ (.CLK(clknet_leaf_6_clk),
    .D(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3703_ (.CLK(clknet_leaf_6_clk),
    .D(_0198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3704_ (.CLK(clknet_leaf_6_clk),
    .D(_0199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3705_ (.CLK(clknet_leaf_6_clk),
    .D(_0200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3706_ (.CLK(clknet_leaf_6_clk),
    .D(_0201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3707_ (.CLK(clknet_leaf_6_clk),
    .D(_0202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3708_ (.CLK(clknet_leaf_6_clk),
    .D(_0203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3709_ (.CLK(clknet_leaf_6_clk),
    .D(_0204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3710_ (.CLK(clknet_leaf_6_clk),
    .D(_0205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3711_ (.CLK(clknet_leaf_6_clk),
    .D(_0206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3712_ (.CLK(clknet_leaf_6_clk),
    .D(_0207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3713_ (.CLK(clknet_leaf_6_clk),
    .D(_0208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3714_ (.CLK(clknet_leaf_6_clk),
    .D(_0209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3715_ (.CLK(clknet_leaf_5_clk),
    .D(_0210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3716_ (.CLK(clknet_leaf_6_clk),
    .D(_0211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3717_ (.CLK(clknet_leaf_6_clk),
    .D(_0212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3718_ (.CLK(clknet_leaf_5_clk),
    .D(_0213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.cnt_1.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3719_ (.CLK(clknet_leaf_6_clk),
    .D(_0214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.race_arb.resp ));
 sky130_fd_sc_hd__dfxtp_1 _3720_ (.CLK(clknet_leaf_6_clk),
    .D(_0215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[6].puf_buffer.race_arb.marked_2 ));
 sky130_fd_sc_hd__dfxtp_1 _3721_ (.CLK(clknet_leaf_5_clk),
    .D(\genblk1[7].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.race_arb.marked_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3722_ (.CLK(clknet_leaf_5_clk),
    .D(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3723_ (.CLK(clknet_leaf_7_clk),
    .D(_0217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3724_ (.CLK(clknet_leaf_7_clk),
    .D(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3725_ (.CLK(clknet_leaf_6_clk),
    .D(_0219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3726_ (.CLK(clknet_leaf_5_clk),
    .D(_0220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3727_ (.CLK(clknet_leaf_5_clk),
    .D(_0221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3728_ (.CLK(clknet_leaf_5_clk),
    .D(_0222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3729_ (.CLK(clknet_leaf_7_clk),
    .D(_0223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3730_ (.CLK(clknet_leaf_5_clk),
    .D(_0224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3731_ (.CLK(clknet_leaf_5_clk),
    .D(_0225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3732_ (.CLK(clknet_leaf_5_clk),
    .D(_0226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3733_ (.CLK(clknet_leaf_5_clk),
    .D(_0227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3734_ (.CLK(clknet_leaf_5_clk),
    .D(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3735_ (.CLK(clknet_leaf_4_clk),
    .D(_0229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3736_ (.CLK(clknet_leaf_4_clk),
    .D(_0230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3737_ (.CLK(clknet_leaf_5_clk),
    .D(_0231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3738_ (.CLK(clknet_leaf_5_clk),
    .D(_0232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_2.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3739_ (.CLK(clknet_leaf_5_clk),
    .D(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3740_ (.CLK(clknet_leaf_1_clk),
    .D(_0234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3741_ (.CLK(clknet_leaf_8_clk),
    .D(_0235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3742_ (.CLK(clknet_leaf_1_clk),
    .D(_0236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3743_ (.CLK(clknet_leaf_5_clk),
    .D(_0237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3744_ (.CLK(clknet_leaf_5_clk),
    .D(_0238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3745_ (.CLK(clknet_leaf_5_clk),
    .D(_0239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3746_ (.CLK(clknet_leaf_1_clk),
    .D(_0240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3747_ (.CLK(clknet_leaf_2_clk),
    .D(_0241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3748_ (.CLK(clknet_leaf_4_clk),
    .D(_0242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3749_ (.CLK(clknet_leaf_2_clk),
    .D(_0243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3750_ (.CLK(clknet_leaf_2_clk),
    .D(_0244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3751_ (.CLK(clknet_leaf_2_clk),
    .D(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3752_ (.CLK(clknet_leaf_2_clk),
    .D(_0246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3753_ (.CLK(clknet_leaf_5_clk),
    .D(_0247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3754_ (.CLK(clknet_leaf_4_clk),
    .D(_0248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3755_ (.CLK(clknet_leaf_4_clk),
    .D(_0249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.cnt_1.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3756_ (.CLK(clknet_leaf_5_clk),
    .D(_0250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[7].puf_buffer.race_arb.marked_2 ));
 sky130_fd_sc_hd__dfxtp_1 _3757_ (.CLK(clknet_leaf_7_clk),
    .D(_0251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.race_arb.resp ));
 sky130_fd_sc_hd__dfxtp_1 _3758_ (.CLK(clknet_leaf_7_clk),
    .D(\genblk1[0].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.race_arb.marked_1 ));
 sky130_fd_sc_hd__dfxtp_1 _3759_ (.CLK(clknet_leaf_5_clk),
    .D(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3760_ (.CLK(clknet_leaf_7_clk),
    .D(_0253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3761_ (.CLK(clknet_leaf_7_clk),
    .D(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3762_ (.CLK(clknet_leaf_7_clk),
    .D(_0255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3763_ (.CLK(clknet_leaf_7_clk),
    .D(_0256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3764_ (.CLK(clknet_leaf_7_clk),
    .D(_0257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3765_ (.CLK(clknet_leaf_7_clk),
    .D(_0258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3766_ (.CLK(clknet_leaf_7_clk),
    .D(_0259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3767_ (.CLK(clknet_leaf_7_clk),
    .D(_0260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3768_ (.CLK(clknet_leaf_8_clk),
    .D(_0261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3769_ (.CLK(clknet_leaf_8_clk),
    .D(_0262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3770_ (.CLK(clknet_leaf_8_clk),
    .D(_0263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3771_ (.CLK(clknet_leaf_5_clk),
    .D(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3772_ (.CLK(clknet_leaf_5_clk),
    .D(_0265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3773_ (.CLK(clknet_leaf_5_clk),
    .D(_0266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3774_ (.CLK(clknet_leaf_7_clk),
    .D(_0267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3775_ (.CLK(clknet_leaf_5_clk),
    .D(_0268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_2.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3776_ (.CLK(clknet_leaf_8_clk),
    .D(net168),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.finish ));
 sky130_fd_sc_hd__dfxtp_1 _3777_ (.CLK(clknet_leaf_8_clk),
    .D(_0270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3778_ (.CLK(clknet_leaf_8_clk),
    .D(_0271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3779_ (.CLK(clknet_leaf_8_clk),
    .D(_0272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3780_ (.CLK(clknet_leaf_8_clk),
    .D(_0273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3781_ (.CLK(clknet_leaf_8_clk),
    .D(_0274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3782_ (.CLK(clknet_leaf_8_clk),
    .D(_0275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3783_ (.CLK(clknet_leaf_8_clk),
    .D(_0276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3784_ (.CLK(clknet_leaf_8_clk),
    .D(_0277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3785_ (.CLK(clknet_leaf_8_clk),
    .D(_0278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3786_ (.CLK(clknet_leaf_8_clk),
    .D(_0279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3787_ (.CLK(clknet_leaf_1_clk),
    .D(_0280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3788_ (.CLK(clknet_leaf_1_clk),
    .D(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3789_ (.CLK(clknet_leaf_1_clk),
    .D(_0282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3790_ (.CLK(clknet_leaf_11_clk),
    .D(_0283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3791_ (.CLK(clknet_leaf_10_clk),
    .D(_0284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3792_ (.CLK(clknet_leaf_1_clk),
    .D(_0285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.cnt_1.ctr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3793_ (.CLK(clknet_leaf_9_clk),
    .D(_0286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.race_arb.resp ));
 sky130_fd_sc_hd__dfxtp_1 _3794_ (.CLK(clknet_leaf_7_clk),
    .D(_0287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[0].puf_buffer.race_arb.marked_2 ));
 sky130_fd_sc_hd__dfxtp_1 _3795_ (.CLK(clknet_leaf_9_clk),
    .D(\genblk1[1].puf_buffer.race_arb.win_1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\genblk1[1].puf_buffer.race_arb.marked_1 ));
 sky130_fd_sc_hd__buf_2 _3812_ (.A(\genblk1[0].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _3813_ (.A(\genblk1[1].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__buf_2 _3814_ (.A(\genblk1[2].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[2]));
 sky130_fd_sc_hd__clkbuf_4 _3815_ (.A(\genblk1[3].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[3]));
 sky130_fd_sc_hd__clkbuf_4 _3816_ (.A(\genblk1[4].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[4]));
 sky130_fd_sc_hd__clkbuf_4 _3817_ (.A(\genblk1[5].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__buf_2 _3818_ (.A(\genblk1[6].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__buf_2 _3819_ (.A(\genblk1[7].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_1_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_1_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[0].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[0].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[0].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[0].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[0].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[0].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[0].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[10].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[10].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[10].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[10].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[10].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[10].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[10].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[11].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[11].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[11].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[11].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[11].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[11].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[11].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[12].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[12].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[12].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[12].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[12].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[12].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[12].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[13].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[13].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[13].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[13].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[13].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[13].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[13].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[14].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[14].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[14].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[14].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[14].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[14].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[14].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[15].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[15].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[15].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[15].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[15].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[15].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[15].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[1].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[1].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[1].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[1].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[1].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[1].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[1].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[2].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[2].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[2].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[2].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[2].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[2].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[2].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[3].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[3].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[3].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[3].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[3].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[3].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[3].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[4].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[4].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[4].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[4].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[4].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[4].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[4].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[5].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[5].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[5].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[5].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[5].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[5].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[5].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[6].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[6].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[6].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[6].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[6].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[6].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[6].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[7].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[7].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[7].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[7].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[7].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[7].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[7].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[8].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[8].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[8].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[8].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[8].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[8].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[8].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[9].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[9].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[9].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[9].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[9].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[9].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_1[9].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_1[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[0].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[0].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[0].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[0].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[0].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[0].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[0].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[10].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[10].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[10].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[10].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[10].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[10].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[10].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[11].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[11].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[11].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[11].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[11].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[11].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[11].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[12].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[12].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[12].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[12].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[12].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[12].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[12].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[13].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[13].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[13].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[13].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[13].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[13].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[13].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[14].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[14].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[14].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[14].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[14].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[14].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[14].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[15].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[15].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[15].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[15].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[15].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[15].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[15].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[1].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[1].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[1].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[1].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[1].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[1].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[1].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[2].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[2].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[2].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[2].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[2].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[2].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[2].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[3].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[3].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[3].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[3].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[3].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[3].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[3].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[4].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[4].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[4].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[4].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[4].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[4].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[4].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[5].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[5].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[5].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[5].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[5].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[5].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[5].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[6].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[6].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[6].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[6].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[6].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[6].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[6].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[7].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[7].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[7].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[7].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[7].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[7].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[7].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[8].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[8].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[8].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[8].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[8].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[8].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[8].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[9].genblk1[0].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[9].genblk1[1].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[9].genblk1[2].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[9].genblk1[3].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[9].genblk1[4].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[9].genblk1[5].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[0].puf_buffer.ro_array_2[9].genblk1[6].inv  (.A(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[0].puf_buffer.ro_array_2[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[0].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[0].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[0].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[0].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[0].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[0].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[0].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[10].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[10].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[10].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[10].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[10].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[10].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[10].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[11].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[11].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[11].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[11].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[11].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[11].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[11].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[12].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[12].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[12].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[12].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[12].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[12].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[12].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[13].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[13].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[13].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[13].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[13].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[13].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[13].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[14].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[14].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[14].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[14].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[14].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[14].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[14].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[15].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[15].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[15].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[15].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[15].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[15].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[15].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[1].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[1].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[1].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[1].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[1].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[1].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[1].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[2].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[2].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[2].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[2].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[2].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[2].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[2].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[3].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[3].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[3].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[3].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[3].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[3].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[3].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[4].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[4].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[4].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[4].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[4].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[4].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[4].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[5].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[5].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[5].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[5].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[5].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[5].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[5].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[6].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[6].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[6].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[6].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[6].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[6].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[6].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[7].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[7].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[7].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[7].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[7].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[7].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[7].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[8].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[8].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[8].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[8].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[8].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[8].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[8].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[9].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[9].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[9].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[9].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[9].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[9].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_1[9].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_1[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[0].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[0].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[0].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[0].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[0].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[0].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[0].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[10].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[10].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[10].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[10].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[10].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[10].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[10].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[11].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[11].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[11].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[11].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[11].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[11].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[11].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[12].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[12].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[12].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[12].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[12].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[12].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[12].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[13].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[13].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[13].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[13].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[13].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[13].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[13].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[14].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[14].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[14].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[14].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[14].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[14].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[14].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[15].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[15].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[15].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[15].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[15].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[15].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[15].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[1].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[1].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[1].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[1].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[1].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[1].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[1].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[2].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[2].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[2].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[2].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[2].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[2].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[2].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[3].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[3].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[3].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[3].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[3].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[3].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[3].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[4].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[4].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[4].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[4].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[4].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[4].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[4].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[5].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[5].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[5].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[5].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[5].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[5].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[5].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[6].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[6].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[6].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[6].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[6].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[6].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[6].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[7].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[7].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[7].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[7].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[7].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[7].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[7].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[8].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[8].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[8].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[8].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[8].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[8].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[8].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[9].genblk1[0].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[9].genblk1[1].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[9].genblk1[2].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[9].genblk1[3].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[9].genblk1[4].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[9].genblk1[5].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[1].puf_buffer.ro_array_2[9].genblk1[6].inv  (.A(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[1].puf_buffer.ro_array_2[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[0].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[0].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[0].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[0].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[0].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[0].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[0].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[10].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[10].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[10].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[10].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[10].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[10].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[10].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[11].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[11].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[11].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[11].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[11].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[11].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[11].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[12].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[12].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[12].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[12].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[12].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[12].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[12].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[13].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[13].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[13].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[13].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[13].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[13].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[13].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[14].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[14].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[14].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[14].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[14].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[14].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[14].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[15].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[15].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[15].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[15].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[15].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[15].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[15].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[1].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[1].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[1].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[1].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[1].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[1].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[1].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[2].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[2].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[2].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[2].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[2].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[2].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[2].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[3].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[3].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[3].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[3].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[3].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[3].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[3].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[4].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[4].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[4].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[4].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[4].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[4].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[4].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[5].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[5].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[5].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[5].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[5].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[5].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[5].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[6].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[6].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[6].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[6].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[6].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[6].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[6].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[7].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[7].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[7].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[7].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[7].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[7].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[7].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[8].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[8].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[8].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[8].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[8].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[8].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[8].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[9].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[9].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[9].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[9].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[9].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[9].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_1[9].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_1[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[0].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[0].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[0].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[0].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[0].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[0].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[0].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[10].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[10].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[10].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[10].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[10].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[10].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[10].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[11].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[11].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[11].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[11].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[11].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[11].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[11].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[12].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[12].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[12].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[12].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[12].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[12].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[12].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[13].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[13].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[13].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[13].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[13].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[13].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[13].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[14].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[14].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[14].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[14].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[14].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[14].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[14].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[15].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[15].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[15].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[15].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[15].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[15].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[15].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[1].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[1].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[1].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[1].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[1].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[1].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[1].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[2].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[2].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[2].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[2].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[2].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[2].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[2].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[3].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[3].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[3].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[3].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[3].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[3].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[3].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[4].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[4].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[4].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[4].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[4].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[4].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[4].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[5].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[5].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[5].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[5].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[5].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[5].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[5].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[6].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[6].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[6].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[6].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[6].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[6].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[6].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[7].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[7].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[7].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[7].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[7].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[7].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[7].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[8].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[8].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[8].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[8].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[8].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[8].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[8].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[9].genblk1[0].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[9].genblk1[1].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[9].genblk1[2].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[9].genblk1[3].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[9].genblk1[4].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[9].genblk1[5].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[2].puf_buffer.ro_array_2[9].genblk1[6].inv  (.A(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[2].puf_buffer.ro_array_2[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[0].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[0].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[0].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[0].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[0].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[0].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[0].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[10].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[10].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[10].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[10].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[10].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[10].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[10].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[11].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[11].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[11].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[11].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[11].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[11].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[11].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[12].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[12].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[12].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[12].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[12].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[12].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[12].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[13].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[13].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[13].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[13].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[13].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[13].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[13].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[14].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[14].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[14].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[14].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[14].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[14].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[14].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[15].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[15].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[15].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[15].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[15].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[15].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[15].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[1].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[1].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[1].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[1].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[1].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[1].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[1].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[2].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[2].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[2].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[2].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[2].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[2].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[2].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[3].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[3].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[3].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[3].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[3].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[3].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[3].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[4].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[4].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[4].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[4].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[4].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[4].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[4].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[5].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[5].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[5].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[5].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[5].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[5].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[5].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[6].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[6].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[6].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[6].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[6].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[6].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[6].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[7].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[7].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[7].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[7].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[7].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[7].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[7].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[8].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[8].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[8].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[8].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[8].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[8].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[8].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[9].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[9].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[9].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[9].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[9].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[9].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_1[9].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_1[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[0].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[0].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[0].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[0].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[0].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[0].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[0].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[10].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[10].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[10].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[10].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[10].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[10].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[10].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[11].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[11].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[11].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[11].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[11].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[11].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[11].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[12].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[12].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[12].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[12].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[12].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[12].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[12].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[13].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[13].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[13].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[13].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[13].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[13].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[13].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[14].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[14].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[14].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[14].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[14].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[14].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[14].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[15].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[15].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[15].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[15].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[15].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[15].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[15].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[1].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[1].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[1].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[1].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[1].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[1].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[1].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[2].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[2].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[2].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[2].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[2].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[2].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[2].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[3].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[3].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[3].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[3].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[3].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[3].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[3].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[4].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[4].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[4].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[4].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[4].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[4].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[4].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[5].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[5].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[5].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[5].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[5].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[5].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[5].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[6].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[6].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[6].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[6].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[6].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[6].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[6].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[7].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[7].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[7].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[7].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[7].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[7].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[7].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[8].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[8].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[8].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[8].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[8].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[8].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[8].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[9].genblk1[0].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[9].genblk1[1].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[9].genblk1[2].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[9].genblk1[3].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[9].genblk1[4].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[9].genblk1[5].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[3].puf_buffer.ro_array_2[9].genblk1[6].inv  (.A(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[3].puf_buffer.ro_array_2[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[0].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[0].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[0].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[0].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[0].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[0].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[0].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[10].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[10].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[10].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[10].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[10].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[10].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[10].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[11].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[11].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[11].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[11].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[11].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[11].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[11].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[12].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[12].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[12].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[12].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[12].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[12].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[12].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[13].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[13].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[13].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[13].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[13].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[13].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[13].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[14].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[14].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[14].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[14].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[14].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[14].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[14].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[15].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[15].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[15].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[15].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[15].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[15].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[15].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[1].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[1].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[1].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[1].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[1].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[1].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[1].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[2].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[2].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[2].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[2].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[2].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[2].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[2].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[3].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[3].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[3].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[3].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[3].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[3].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[3].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[4].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[4].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[4].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[4].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[4].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[4].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[4].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[5].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[5].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[5].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[5].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[5].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[5].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[5].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[6].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[6].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[6].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[6].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[6].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[6].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[6].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[7].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[7].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[7].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[7].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[7].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[7].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[7].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[8].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[8].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[8].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[8].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[8].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[8].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[8].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[9].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[9].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[9].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[9].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[9].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[9].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_1[9].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_1[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[0].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[0].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[0].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[0].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[0].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[0].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[0].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[10].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[10].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[10].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[10].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[10].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[10].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[10].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[11].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[11].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[11].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[11].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[11].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[11].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[11].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[12].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[12].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[12].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[12].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[12].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[12].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[12].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[13].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[13].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[13].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[13].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[13].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[13].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[13].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[14].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[14].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[14].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[14].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[14].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[14].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[14].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[15].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[15].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[15].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[15].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[15].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[15].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[15].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[1].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[1].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[1].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[1].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[1].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[1].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[1].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[2].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[2].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[2].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[2].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[2].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[2].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[2].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[3].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[3].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[3].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[3].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[3].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[3].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[3].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[4].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[4].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[4].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[4].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[4].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[4].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[4].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[5].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[5].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[5].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[5].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[5].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[5].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[5].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[6].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[6].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[6].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[6].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[6].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[6].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[6].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[7].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[7].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[7].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[7].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[7].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[7].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[7].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[8].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[8].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[8].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[8].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[8].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[8].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[8].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[9].genblk1[0].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[9].genblk1[1].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[9].genblk1[2].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[9].genblk1[3].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[9].genblk1[4].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[9].genblk1[5].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[4].puf_buffer.ro_array_2[9].genblk1[6].inv  (.A(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[4].puf_buffer.ro_array_2[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[0].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[0].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[0].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[0].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[0].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[0].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[0].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[10].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[10].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[10].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[10].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[10].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[10].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[10].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[11].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[11].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[11].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[11].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[11].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[11].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[11].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[12].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[12].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[12].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[12].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[12].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[12].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[12].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[13].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[13].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[13].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[13].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[13].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[13].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[13].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[14].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[14].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[14].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[14].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[14].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[14].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[14].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[15].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[15].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[15].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[15].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[15].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[15].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[15].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[1].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[1].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[1].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[1].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[1].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[1].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[1].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[2].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[2].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[2].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[2].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[2].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[2].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[2].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[3].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[3].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[3].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[3].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[3].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[3].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[3].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[4].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[4].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[4].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[4].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[4].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[4].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[4].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[5].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[5].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[5].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[5].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[5].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[5].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[5].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[6].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[6].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[6].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[6].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[6].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[6].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[6].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[7].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[7].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[7].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[7].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[7].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[7].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[7].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[8].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[8].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[8].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[8].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[8].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[8].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[8].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[9].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[9].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[9].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[9].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[9].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[9].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_1[9].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_1[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[0].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[0].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[0].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[0].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[0].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[0].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[0].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[10].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[10].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[10].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[10].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[10].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[10].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[10].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[11].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[11].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[11].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[11].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[11].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[11].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[11].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[12].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[12].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[12].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[12].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[12].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[12].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[12].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[13].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[13].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[13].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[13].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[13].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[13].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[13].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[14].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[14].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[14].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[14].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[14].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[14].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[14].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[15].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[15].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[15].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[15].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[15].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[15].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[15].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[1].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[1].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[1].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[1].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[1].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[1].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[1].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[2].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[2].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[2].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[2].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[2].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[2].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[2].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[3].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[3].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[3].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[3].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[3].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[3].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[3].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[4].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[4].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[4].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[4].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[4].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[4].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[4].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[5].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[5].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[5].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[5].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[5].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[5].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[5].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[6].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[6].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[6].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[6].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[6].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[6].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[6].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[7].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[7].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[7].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[7].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[7].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[7].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[7].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[8].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[8].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[8].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[8].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[8].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[8].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[8].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[9].genblk1[0].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[9].genblk1[1].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[9].genblk1[2].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[9].genblk1[3].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[9].genblk1[4].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[9].genblk1[5].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[5].puf_buffer.ro_array_2[9].genblk1[6].inv  (.A(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[5].puf_buffer.ro_array_2[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[0].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[0].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[0].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[0].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[0].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[0].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[0].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[10].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[10].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[10].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[10].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[10].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[10].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[10].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[11].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[11].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[11].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[11].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[11].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[11].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[11].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[12].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[12].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[12].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[12].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[12].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[12].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[12].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[13].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[13].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[13].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[13].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[13].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[13].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[13].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[14].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[14].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[14].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[14].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[14].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[14].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[14].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[15].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[15].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[15].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[15].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[15].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[15].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[15].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[1].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[1].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[1].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[1].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[1].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[1].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[1].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[2].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[2].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[2].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[2].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[2].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[2].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[2].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[3].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[3].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[3].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[3].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[3].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[3].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[3].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[4].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[4].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[4].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[4].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[4].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[4].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[4].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[5].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[5].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[5].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[5].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[5].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[5].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[5].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[6].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[6].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[6].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[6].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[6].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[6].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[6].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[7].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[7].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[7].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[7].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[7].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[7].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[7].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[8].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[8].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[8].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[8].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[8].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[8].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[8].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[9].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[9].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[9].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[9].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[9].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[9].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_1[9].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_1[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[0].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[0].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[0].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[0].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[0].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[0].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[0].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[10].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[10].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[10].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[10].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[10].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[10].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[10].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[11].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[11].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[11].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[11].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[11].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[11].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[11].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[12].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[12].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[12].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[12].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[12].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[12].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[12].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[13].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[13].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[13].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[13].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[13].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[13].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[13].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[14].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[14].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[14].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[14].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[14].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[14].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[14].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[15].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[15].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[15].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[15].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[15].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[15].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[15].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[1].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[1].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[1].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[1].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[1].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[1].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[1].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[2].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[2].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[2].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[2].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[2].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[2].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[2].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[3].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[3].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[3].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[3].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[3].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[3].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[3].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[4].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[4].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[4].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[4].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[4].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[4].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[4].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[5].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[5].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[5].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[5].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[5].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[5].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[5].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[6].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[6].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[6].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[6].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[6].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[6].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[6].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[7].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[7].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[7].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[7].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[7].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[7].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[7].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[8].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[8].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[8].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[8].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[8].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[8].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[8].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[9].genblk1[0].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[9].genblk1[1].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[9].genblk1[2].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[9].genblk1[3].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[9].genblk1[4].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[9].genblk1[5].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[6].puf_buffer.ro_array_2[9].genblk1[6].inv  (.A(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[6].puf_buffer.ro_array_2[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[0].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[0].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[0].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[0].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[0].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[0].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[0].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[10].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[10].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[10].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[10].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[10].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[10].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[10].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[11].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[11].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[11].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[11].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[11].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[11].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[11].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[12].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[12].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[12].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[12].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[12].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[12].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[12].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[13].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[13].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[13].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[13].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[13].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[13].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[13].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[14].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[14].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[14].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[14].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[14].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[14].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[14].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[15].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[15].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[15].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[15].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[15].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[15].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[15].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[1].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[1].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[1].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[1].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[1].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[1].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[1].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[2].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[2].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[2].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[2].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[2].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[2].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[2].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[3].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[3].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[3].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[3].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[3].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[3].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[3].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[4].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[4].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[4].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[4].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[4].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[4].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[4].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[5].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[5].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[5].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[5].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[5].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[5].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[5].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[6].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[6].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[6].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[6].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[6].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[6].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[6].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[7].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[7].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[7].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[7].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[7].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[7].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[7].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[8].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[8].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[8].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[8].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[8].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[8].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[8].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[9].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[9].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[9].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[9].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[9].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[9].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_1[9].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_1[9].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[0].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[0].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[0].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[0].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[0].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[0].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[0].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[0].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[10].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[10].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[10].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[10].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[10].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[10].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[10].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[10].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[11].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[11].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[11].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[11].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[11].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[11].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[11].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[11].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[12].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[12].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[12].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[12].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[12].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[12].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[12].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[12].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[13].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[13].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[13].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[13].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[13].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[13].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[13].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[13].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[14].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[14].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[14].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[14].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[14].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[14].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[14].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[14].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[15].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[15].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[15].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[15].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[15].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[15].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[15].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[15].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[1].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[1].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[1].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[1].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[1].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[1].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[1].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[1].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[2].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[2].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[2].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[2].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[2].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[2].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[2].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[2].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[3].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[3].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[3].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[3].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[3].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[3].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[3].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[3].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[4].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[4].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[4].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[4].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[4].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[4].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[4].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[4].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[5].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[5].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[5].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[5].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[5].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[5].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[5].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[5].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[6].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[6].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[6].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[6].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[6].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[6].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[6].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[6].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[7].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[7].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[7].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[7].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[7].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[7].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[7].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[7].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[8].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[8].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[8].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[8].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[8].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[8].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[8].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[8].inter_wire[7] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[9].genblk1[0].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[1] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[9].genblk1[1].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[2] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[9].genblk1[2].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[3] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[9].genblk1[3].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[4] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[9].genblk1[4].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[5] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[9].genblk1[5].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[6] ));
 sky130_fd_sc_hd__inv_2 \genblk1[7].puf_buffer.ro_array_2[9].genblk1[6].inv  (.A(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\genblk1[7].puf_buffer.ro_array_2[9].inter_wire[7] ));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\genblk1[3].puf_buffer.cnt_2.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\genblk1[2].puf_buffer.cnt_1.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\genblk1[7].puf_buffer.cnt_2.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\genblk1[1].puf_buffer.cnt_1.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\genblk1[1].puf_buffer.cnt_1.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\genblk1[7].puf_buffer.cnt_2.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\genblk1[3].puf_buffer.cnt_2.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\genblk1[7].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\genblk1[6].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\genblk1[7].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\genblk1[5].puf_buffer.cnt_1.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\genblk1[5].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\genblk1[6].puf_buffer.cnt_2.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\genblk1[5].puf_buffer.cnt_2.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\genblk1[5].puf_buffer.cnt_1.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\genblk1[2].puf_buffer.cnt_2.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\genblk1[5].puf_buffer.cnt_1.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\genblk1[0].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\genblk1[0].puf_buffer.cnt_2.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\genblk1[2].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\genblk1[1].puf_buffer.cnt_1.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\genblk1[0].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\genblk1[5].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\genblk1[3].puf_buffer.cnt_1.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\genblk1[1].puf_buffer.cnt_2.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\genblk1[2].puf_buffer.cnt_1.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\genblk1[6].puf_buffer.cnt_1.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\genblk1[5].puf_buffer.cnt_2.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\genblk1[5].puf_buffer.cnt_1.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\genblk1[4].puf_buffer.cnt_1.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\genblk1[6].puf_buffer.cnt_2.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\genblk1[1].puf_buffer.cnt_1.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\genblk1[3].puf_buffer.cnt_2.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\genblk1[2].puf_buffer.cnt_1.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\genblk1[7].puf_buffer.cnt_1.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\genblk1[0].puf_buffer.cnt_1.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\genblk1[2].puf_buffer.cnt_2.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\genblk1[3].puf_buffer.cnt_2.ctr[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\genblk1[4].puf_buffer.cnt_2.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\genblk1[7].puf_buffer.cnt_2.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\genblk1[2].puf_buffer.cnt_2.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\genblk1[2].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\genblk1[0].puf_buffer.cnt_2.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\genblk1[5].puf_buffer.cnt_1.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\genblk1[0].puf_buffer.cnt_2.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_0264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\genblk1[3].puf_buffer.cnt_2.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\genblk1[6].puf_buffer.cnt_1.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\genblk1[7].puf_buffer.cnt_2.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\genblk1[4].puf_buffer.cnt_1.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\genblk1[4].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\genblk1[3].puf_buffer.cnt_1.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\genblk1[1].puf_buffer.cnt_2.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\genblk1[6].puf_buffer.cnt_2.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\genblk1[1].puf_buffer.cnt_1.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\genblk1[3].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\genblk1[6].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\genblk1[0].puf_buffer.cnt_1.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\genblk1[1].puf_buffer.cnt_2.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\genblk1[2].puf_buffer.cnt_2.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\genblk1[7].puf_buffer.cnt_1.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\genblk1[5].puf_buffer.cnt_1.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\genblk1[5].puf_buffer.cnt_2.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\genblk1[0].puf_buffer.cnt_2.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\genblk1[1].puf_buffer.cnt_2.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\genblk1[6].puf_buffer.cnt_1.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\genblk1[4].puf_buffer.cnt_1.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\genblk1[4].puf_buffer.cnt_2.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\genblk1[4].puf_buffer.cnt_1.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_0127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\genblk1[2].puf_buffer.cnt_1.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_0055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\genblk1[6].puf_buffer.cnt_2.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\genblk1[5].puf_buffer.cnt_2.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\genblk1[6].puf_buffer.cnt_2.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\genblk1[3].puf_buffer.cnt_2.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\genblk1[1].puf_buffer.cnt_1.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\genblk1[7].puf_buffer.cnt_2.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\genblk1[4].puf_buffer.cnt_2.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\genblk1[1].puf_buffer.cnt_1.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\genblk1[3].puf_buffer.cnt_1.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\genblk1[6].puf_buffer.cnt_1.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\genblk1[5].puf_buffer.cnt_1.ctr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\genblk1[1].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\genblk1[0].puf_buffer.cnt_1.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\genblk1[0].puf_buffer.cnt_1.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\genblk1[4].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\genblk1[0].puf_buffer.cnt_2.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\genblk1[2].puf_buffer.cnt_2.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\genblk1[7].puf_buffer.cnt_1.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\genblk1[7].puf_buffer.cnt_1.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\genblk1[0].puf_buffer.cnt_2.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\genblk1[7].puf_buffer.cnt_2.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\genblk1[3].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_0089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\genblk1[4].puf_buffer.cnt_2.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\genblk1[0].puf_buffer.cnt_2.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\genblk1[0].puf_buffer.cnt_1.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\genblk1[1].puf_buffer.cnt_2.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\genblk1[3].puf_buffer.cnt_2.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_0084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\genblk1[7].puf_buffer.cnt_1.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\genblk1[1].puf_buffer.cnt_1.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\genblk1[6].puf_buffer.cnt_1.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\genblk1[0].puf_buffer.cnt_1.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\genblk1[6].puf_buffer.cnt_2.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\genblk1[6].puf_buffer.cnt_1.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\genblk1[2].puf_buffer.cnt_1.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\genblk1[3].puf_buffer.cnt_1.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\genblk1[4].puf_buffer.cnt_2.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\genblk1[0].puf_buffer.cnt_2.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\genblk1[3].puf_buffer.cnt_1.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\genblk1[1].puf_buffer.cnt_2.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\genblk1[0].puf_buffer.cnt_1.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\genblk1[7].puf_buffer.cnt_2.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\genblk1[6].puf_buffer.cnt_1.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\genblk1[6].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\genblk1[3].puf_buffer.cnt_1.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\genblk1[2].puf_buffer.cnt_2.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\genblk1[7].puf_buffer.cnt_2.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\genblk1[4].puf_buffer.cnt_2.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\genblk1[6].puf_buffer.cnt_2.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\genblk1[1].puf_buffer.cnt_2.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\genblk1[2].puf_buffer.cnt_2.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\genblk1[4].puf_buffer.cnt_1.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\genblk1[5].puf_buffer.cnt_1.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\genblk1[5].puf_buffer.cnt_2.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\genblk1[7].puf_buffer.race_arb.resp ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\genblk1[6].puf_buffer.cnt_1.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\genblk1[7].puf_buffer.cnt_2.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\genblk1[2].puf_buffer.cnt_1.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\genblk1[2].puf_buffer.cnt_2.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\genblk1[3].puf_buffer.cnt_2.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\genblk1[2].puf_buffer.cnt_1.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\genblk1[4].puf_buffer.cnt_2.ctr[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\genblk1[5].puf_buffer.cnt_1.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\genblk1[7].puf_buffer.cnt_1.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\genblk1[4].puf_buffer.cnt_1.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\genblk1[3].puf_buffer.cnt_2.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\genblk1[6].puf_buffer.cnt_2.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\genblk1[7].puf_buffer.cnt_1.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\genblk1[2].puf_buffer.cnt_1.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\genblk1[2].puf_buffer.cnt_1.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\genblk1[4].puf_buffer.cnt_2.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\genblk1[4].puf_buffer.cnt_1.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\genblk1[1].puf_buffer.cnt_2.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\genblk1[3].puf_buffer.cnt_1.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\genblk1[4].puf_buffer.cnt_2.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\genblk1[7].puf_buffer.cnt_1.ctr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\genblk1[0].puf_buffer.cnt_2.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\genblk1[1].puf_buffer.cnt_1.ctr[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\genblk1[2].puf_buffer.cnt_1.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\genblk1[7].puf_buffer.cnt_1.ctr[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\genblk1[0].puf_buffer.cnt_1.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\genblk1[2].puf_buffer.cnt_2.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\genblk1[5].puf_buffer.cnt_2.ctr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\genblk1[0].puf_buffer.cnt_1.ctr[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\genblk1[5].puf_buffer.cnt_2.ctr[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\genblk1[4].puf_buffer.cnt_1.finish ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\genblk1[1].puf_buffer.cnt_2.ctr[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\genblk1[4].puf_buffer.cnt_1.ctr[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(ui_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(ui_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(ui_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(ui_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(ui_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(ui_in[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(ui_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(ui_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 max_cap10 (.A(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 max_cap11 (.A(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 max_cap14 (.A(_0693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 max_cap15 (.A(_0688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 max_cap16 (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 max_cap17 (.A(_0619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 max_cap18 (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 max_cap19 (.A(_0616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__buf_1 max_cap2 (.A(_0697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 max_cap20 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 max_cap21 (.A(_0613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 max_cap23 (.A(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 max_cap24 (.A(_0708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 max_cap25 (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 max_cap26 (.A(_0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 max_cap3 (.A(_0708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 max_cap4 (.A(_0609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net232));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net27));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net28));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net29));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net30));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net31));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net32));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net33));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net34));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net35));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net36));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net37));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net38));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net39));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net40));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net41));
 sky130_fd_sc_hd__conb_1 tt_um_litneet64_ro_puf_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net42));
 sky130_fd_sc_hd__clkbuf_1 wire1 (.A(_0703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 wire12 (.A(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 wire13 (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 wire22 (.A(_0606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 assign uio_oe[0] = net27;
 assign uio_oe[1] = net28;
 assign uio_oe[2] = net29;
 assign uio_oe[3] = net30;
 assign uio_oe[4] = net31;
 assign uio_oe[5] = net32;
 assign uio_oe[6] = net33;
 assign uio_oe[7] = net34;
 assign uio_out[0] = net35;
 assign uio_out[1] = net36;
 assign uio_out[2] = net37;
 assign uio_out[3] = net38;
 assign uio_out[4] = net39;
 assign uio_out[5] = net40;
 assign uio_out[6] = net41;
 assign uio_out[7] = net42;
endmodule
