VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_alfiero88_CurrentTrigger
  CLASS BLOCK ;
  FOREIGN tt_um_alfiero88_CurrentTrigger ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.350000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.530000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 10.312400 ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 41.144600 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 110.310 119.660 115.410 124.620 ;
        RECT 119.970 119.590 125.070 124.620 ;
      LAYER nwell ;
        RECT 129.100 118.470 134.290 124.620 ;
        RECT 137.490 119.550 142.680 124.510 ;
      LAYER pwell ;
        RECT 110.890 97.910 116.990 109.450 ;
        RECT 110.950 82.310 117.050 93.850 ;
      LAYER nwell ;
        RECT 121.720 86.310 125.410 105.800 ;
        RECT 129.550 86.310 133.240 105.800 ;
      LAYER pwell ;
        RECT 113.940 73.160 117.040 78.700 ;
      LAYER nwell ;
        RECT 127.080 73.060 131.410 79.210 ;
        RECT 137.390 71.150 141.580 102.430 ;
      LAYER pwell ;
        RECT 113.970 59.190 117.070 64.730 ;
        RECT 128.210 57.640 131.310 66.180 ;
      LAYER nwell ;
        RECT 137.040 61.760 140.900 65.350 ;
      LAYER pwell ;
        RECT 119.740 49.200 122.840 51.310 ;
      LAYER nwell ;
        RECT 125.070 49.050 129.260 51.360 ;
      LAYER pwell ;
        RECT 119.740 44.000 123.340 46.630 ;
      LAYER nwell ;
        RECT 125.070 43.630 129.260 47.220 ;
      LAYER pwell ;
        RECT 118.300 36.690 123.400 39.800 ;
      LAYER nwell ;
        RECT 125.070 35.490 130.260 41.000 ;
        RECT 136.840 35.380 141.030 56.790 ;
      LAYER li1 ;
        RECT 120.600 124.440 124.450 124.490 ;
        RECT 129.740 124.440 133.640 124.470 ;
        RECT 110.490 124.270 115.230 124.440 ;
        RECT 110.490 123.990 110.660 124.270 ;
        RECT 110.450 120.300 110.660 123.990 ;
        RECT 111.340 123.700 114.380 123.870 ;
        RECT 111.000 120.640 111.170 123.640 ;
        RECT 114.550 120.640 114.720 123.640 ;
        RECT 111.340 120.410 114.380 120.580 ;
        RECT 110.490 120.010 110.660 120.300 ;
        RECT 115.060 120.010 115.230 124.270 ;
        RECT 110.490 119.840 115.230 120.010 ;
        RECT 120.150 124.270 124.890 124.440 ;
        RECT 120.150 119.940 120.320 124.270 ;
        RECT 120.660 123.380 120.830 123.710 ;
        RECT 121.000 123.700 124.040 123.870 ;
        RECT 121.000 123.220 124.040 123.390 ;
        RECT 120.660 122.420 120.830 122.750 ;
        RECT 121.000 122.740 124.040 122.910 ;
        RECT 124.210 122.900 124.380 123.230 ;
        RECT 121.000 122.260 124.040 122.430 ;
        RECT 120.660 121.460 120.830 121.790 ;
        RECT 121.000 121.780 124.040 121.950 ;
        RECT 124.210 121.940 124.380 122.270 ;
        RECT 121.000 121.300 124.040 121.470 ;
        RECT 120.660 120.500 120.830 120.830 ;
        RECT 121.000 120.820 124.040 120.990 ;
        RECT 124.210 120.980 124.380 121.310 ;
        RECT 121.000 120.340 124.040 120.510 ;
        RECT 124.720 119.940 124.890 124.270 ;
        RECT 120.150 119.770 124.890 119.940 ;
        RECT 129.280 124.270 134.110 124.440 ;
        RECT 129.280 118.820 129.450 124.270 ;
        RECT 130.175 123.700 133.215 123.870 ;
        RECT 129.790 123.290 129.960 123.640 ;
        RECT 133.430 123.290 133.600 123.640 ;
        RECT 130.175 123.060 133.215 123.230 ;
        RECT 129.790 122.650 129.960 123.000 ;
        RECT 133.430 122.650 133.600 123.000 ;
        RECT 130.175 122.420 133.215 122.590 ;
        RECT 129.790 122.010 129.960 122.360 ;
        RECT 133.430 122.010 133.600 122.360 ;
        RECT 130.175 121.780 133.215 121.950 ;
        RECT 129.790 121.370 129.960 121.720 ;
        RECT 133.430 121.370 133.600 121.720 ;
        RECT 130.175 121.140 133.215 121.310 ;
        RECT 129.790 120.730 129.960 121.080 ;
        RECT 133.430 120.730 133.600 121.080 ;
        RECT 130.175 120.500 133.215 120.670 ;
        RECT 129.790 120.090 129.960 120.440 ;
        RECT 133.430 120.090 133.600 120.440 ;
        RECT 130.175 119.860 133.215 120.030 ;
        RECT 129.790 119.450 129.960 119.800 ;
        RECT 133.430 119.450 133.600 119.800 ;
        RECT 130.175 119.220 133.215 119.390 ;
        RECT 133.940 118.820 134.110 124.270 ;
        RECT 137.670 124.160 142.500 124.330 ;
        RECT 137.670 119.900 137.840 124.160 ;
        RECT 142.330 123.870 142.500 124.160 ;
        RECT 138.565 123.590 141.605 123.760 ;
        RECT 138.180 120.530 138.350 123.530 ;
        RECT 141.820 120.530 141.990 123.530 ;
        RECT 138.565 120.300 141.605 120.470 ;
        RECT 142.330 120.190 142.530 123.870 ;
        RECT 142.330 119.900 142.500 120.190 ;
        RECT 137.670 119.730 142.500 119.900 ;
        RECT 129.280 118.650 134.110 118.820 ;
        RECT 111.070 109.100 116.810 109.270 ;
        RECT 111.070 108.820 111.240 109.100 ;
        RECT 111.000 98.540 111.240 108.820 ;
        RECT 111.920 108.530 115.960 108.700 ;
        RECT 111.580 105.470 111.750 108.470 ;
        RECT 116.130 105.470 116.300 108.470 ;
        RECT 111.920 105.240 115.960 105.410 ;
        RECT 111.580 102.180 111.750 105.180 ;
        RECT 116.130 102.180 116.300 105.180 ;
        RECT 111.920 101.950 115.960 102.120 ;
        RECT 111.580 98.890 111.750 101.890 ;
        RECT 116.130 98.890 116.300 101.890 ;
        RECT 111.920 98.660 115.960 98.830 ;
        RECT 111.070 98.260 111.240 98.540 ;
        RECT 116.640 98.260 116.810 109.100 ;
        RECT 111.070 98.090 116.810 98.260 ;
        RECT 121.900 105.450 125.230 105.620 ;
        RECT 111.130 93.500 116.870 93.670 ;
        RECT 111.130 93.210 111.300 93.500 ;
        RECT 111.060 82.950 111.300 93.210 ;
        RECT 111.980 92.930 116.020 93.100 ;
        RECT 111.640 89.870 111.810 92.870 ;
        RECT 116.190 89.870 116.360 92.870 ;
        RECT 111.980 89.640 116.020 89.810 ;
        RECT 111.640 86.580 111.810 89.580 ;
        RECT 116.190 86.580 116.360 89.580 ;
        RECT 111.980 86.350 116.020 86.520 ;
        RECT 111.640 83.290 111.810 86.290 ;
        RECT 116.190 83.290 116.360 86.290 ;
        RECT 111.980 83.060 116.020 83.230 ;
        RECT 111.130 82.660 111.300 82.950 ;
        RECT 116.700 82.660 116.870 93.500 ;
        RECT 121.900 86.660 122.070 105.450 ;
        RECT 125.060 105.190 125.230 105.450 ;
        RECT 129.730 105.450 133.060 105.620 ;
        RECT 122.795 104.880 124.335 105.050 ;
        RECT 122.410 104.120 122.580 104.820 ;
        RECT 124.550 104.120 124.720 104.820 ;
        RECT 122.795 103.890 124.335 104.060 ;
        RECT 122.410 103.130 122.580 103.830 ;
        RECT 124.550 103.130 124.720 103.830 ;
        RECT 122.795 102.900 124.335 103.070 ;
        RECT 122.410 102.140 122.580 102.840 ;
        RECT 124.550 102.140 124.720 102.840 ;
        RECT 122.795 101.910 124.335 102.080 ;
        RECT 122.410 101.150 122.580 101.850 ;
        RECT 124.550 101.150 124.720 101.850 ;
        RECT 122.795 100.920 124.335 101.090 ;
        RECT 122.410 100.160 122.580 100.860 ;
        RECT 124.550 100.160 124.720 100.860 ;
        RECT 122.795 99.930 124.335 100.100 ;
        RECT 122.410 99.170 122.580 99.870 ;
        RECT 124.550 99.170 124.720 99.870 ;
        RECT 122.795 98.940 124.335 99.110 ;
        RECT 122.410 98.180 122.580 98.880 ;
        RECT 124.550 98.180 124.720 98.880 ;
        RECT 122.795 97.950 124.335 98.120 ;
        RECT 122.410 97.190 122.580 97.890 ;
        RECT 124.550 97.190 124.720 97.890 ;
        RECT 122.795 96.960 124.335 97.130 ;
        RECT 122.410 96.200 122.580 96.900 ;
        RECT 124.550 96.200 124.720 96.900 ;
        RECT 122.795 95.970 124.335 96.140 ;
        RECT 122.410 95.210 122.580 95.910 ;
        RECT 124.550 95.210 124.720 95.910 ;
        RECT 122.795 94.980 124.335 95.150 ;
        RECT 122.410 94.220 122.580 94.920 ;
        RECT 124.550 94.220 124.720 94.920 ;
        RECT 122.795 93.990 124.335 94.160 ;
        RECT 122.410 93.230 122.580 93.930 ;
        RECT 124.550 93.230 124.720 93.930 ;
        RECT 122.795 93.000 124.335 93.170 ;
        RECT 122.410 92.240 122.580 92.940 ;
        RECT 124.550 92.240 124.720 92.940 ;
        RECT 122.795 92.010 124.335 92.180 ;
        RECT 122.410 91.250 122.580 91.950 ;
        RECT 124.550 91.250 124.720 91.950 ;
        RECT 122.795 91.020 124.335 91.190 ;
        RECT 122.410 90.260 122.580 90.960 ;
        RECT 124.550 90.260 124.720 90.960 ;
        RECT 122.795 90.030 124.335 90.200 ;
        RECT 122.410 89.270 122.580 89.970 ;
        RECT 124.550 89.270 124.720 89.970 ;
        RECT 122.795 89.040 124.335 89.210 ;
        RECT 122.410 88.280 122.580 88.980 ;
        RECT 124.550 88.280 124.720 88.980 ;
        RECT 122.795 88.050 124.335 88.220 ;
        RECT 122.410 87.290 122.580 87.990 ;
        RECT 124.550 87.290 124.720 87.990 ;
        RECT 122.795 87.060 124.335 87.230 ;
        RECT 125.060 86.920 125.470 105.190 ;
        RECT 125.060 86.660 125.230 86.920 ;
        RECT 121.900 86.490 125.230 86.660 ;
        RECT 129.730 86.660 129.900 105.450 ;
        RECT 132.890 105.050 133.060 105.450 ;
        RECT 130.625 104.880 132.165 105.050 ;
        RECT 130.240 104.120 130.410 104.820 ;
        RECT 132.380 104.120 132.550 104.820 ;
        RECT 130.625 103.890 132.165 104.060 ;
        RECT 130.240 103.130 130.410 103.830 ;
        RECT 132.380 103.130 132.550 103.830 ;
        RECT 130.625 102.900 132.165 103.070 ;
        RECT 130.240 102.140 130.410 102.840 ;
        RECT 132.380 102.140 132.550 102.840 ;
        RECT 130.625 101.910 132.165 102.080 ;
        RECT 130.240 101.150 130.410 101.850 ;
        RECT 132.380 101.150 132.550 101.850 ;
        RECT 130.625 100.920 132.165 101.090 ;
        RECT 130.240 100.160 130.410 100.860 ;
        RECT 132.380 100.160 132.550 100.860 ;
        RECT 130.625 99.930 132.165 100.100 ;
        RECT 130.240 99.170 130.410 99.870 ;
        RECT 132.380 99.170 132.550 99.870 ;
        RECT 130.625 98.940 132.165 99.110 ;
        RECT 130.240 98.180 130.410 98.880 ;
        RECT 132.380 98.180 132.550 98.880 ;
        RECT 130.625 97.950 132.165 98.120 ;
        RECT 130.240 97.190 130.410 97.890 ;
        RECT 132.380 97.190 132.550 97.890 ;
        RECT 130.625 96.960 132.165 97.130 ;
        RECT 130.240 96.200 130.410 96.900 ;
        RECT 132.380 96.200 132.550 96.900 ;
        RECT 130.625 95.970 132.165 96.140 ;
        RECT 130.240 95.210 130.410 95.910 ;
        RECT 132.380 95.210 132.550 95.910 ;
        RECT 130.625 94.980 132.165 95.150 ;
        RECT 130.240 94.220 130.410 94.920 ;
        RECT 132.380 94.220 132.550 94.920 ;
        RECT 130.625 93.990 132.165 94.160 ;
        RECT 130.240 93.230 130.410 93.930 ;
        RECT 132.380 93.230 132.550 93.930 ;
        RECT 130.625 93.000 132.165 93.170 ;
        RECT 130.240 92.240 130.410 92.940 ;
        RECT 132.380 92.240 132.550 92.940 ;
        RECT 130.625 92.010 132.165 92.180 ;
        RECT 130.240 91.250 130.410 91.950 ;
        RECT 132.380 91.250 132.550 91.950 ;
        RECT 130.625 91.020 132.165 91.190 ;
        RECT 130.240 90.260 130.410 90.960 ;
        RECT 132.380 90.260 132.550 90.960 ;
        RECT 130.625 90.030 132.165 90.200 ;
        RECT 130.240 89.270 130.410 89.970 ;
        RECT 132.380 89.270 132.550 89.970 ;
        RECT 130.625 89.040 132.165 89.210 ;
        RECT 130.240 88.280 130.410 88.980 ;
        RECT 132.380 88.280 132.550 88.980 ;
        RECT 130.625 88.050 132.165 88.220 ;
        RECT 130.240 87.290 130.410 87.990 ;
        RECT 132.380 87.290 132.550 87.990 ;
        RECT 130.625 87.060 132.165 87.230 ;
        RECT 132.880 86.950 133.180 105.050 ;
        RECT 137.570 102.080 141.400 102.250 ;
        RECT 132.890 86.660 133.060 86.950 ;
        RECT 129.730 86.490 133.060 86.660 ;
        RECT 111.130 82.490 116.870 82.660 ;
        RECT 127.260 78.860 131.230 79.030 ;
        RECT 114.120 78.350 116.860 78.520 ;
        RECT 114.120 78.080 114.290 78.350 ;
        RECT 114.060 73.780 114.290 78.080 ;
        RECT 114.970 77.780 116.010 77.950 ;
        RECT 114.630 76.720 114.800 77.720 ;
        RECT 116.180 76.720 116.350 77.720 ;
        RECT 114.970 76.490 116.010 76.660 ;
        RECT 114.630 75.430 114.800 76.430 ;
        RECT 116.180 75.430 116.350 76.430 ;
        RECT 114.970 75.200 116.010 75.370 ;
        RECT 114.630 74.140 114.800 75.140 ;
        RECT 116.180 74.140 116.350 75.140 ;
        RECT 114.970 73.910 116.010 74.080 ;
        RECT 114.120 73.510 114.290 73.780 ;
        RECT 116.690 73.510 116.860 78.350 ;
        RECT 114.120 73.340 116.860 73.510 ;
        RECT 127.260 73.410 127.430 78.860 ;
        RECT 131.060 78.610 131.230 78.860 ;
        RECT 128.155 78.290 130.335 78.460 ;
        RECT 127.770 77.880 127.940 78.230 ;
        RECT 130.550 77.880 130.720 78.230 ;
        RECT 128.155 77.650 130.335 77.820 ;
        RECT 127.770 77.240 127.940 77.590 ;
        RECT 130.550 77.240 130.720 77.590 ;
        RECT 128.155 77.010 130.335 77.180 ;
        RECT 127.770 76.600 127.940 76.950 ;
        RECT 130.550 76.600 130.720 76.950 ;
        RECT 128.155 76.370 130.335 76.540 ;
        RECT 127.770 75.960 127.940 76.310 ;
        RECT 130.550 75.960 130.720 76.310 ;
        RECT 128.155 75.730 130.335 75.900 ;
        RECT 127.770 75.320 127.940 75.670 ;
        RECT 130.550 75.320 130.720 75.670 ;
        RECT 128.155 75.090 130.335 75.260 ;
        RECT 127.770 74.680 127.940 75.030 ;
        RECT 130.550 74.680 130.720 75.030 ;
        RECT 128.155 74.450 130.335 74.620 ;
        RECT 127.770 74.040 127.940 74.390 ;
        RECT 130.550 74.040 130.720 74.390 ;
        RECT 128.155 73.810 130.335 73.980 ;
        RECT 131.060 73.660 131.320 78.610 ;
        RECT 131.060 73.410 131.230 73.660 ;
        RECT 127.260 73.240 131.230 73.410 ;
        RECT 137.570 71.500 137.740 102.080 ;
        RECT 141.230 101.800 141.400 102.080 ;
        RECT 138.465 101.510 140.505 101.680 ;
        RECT 138.080 98.450 138.250 101.450 ;
        RECT 140.720 98.450 140.890 101.450 ;
        RECT 138.465 98.220 140.505 98.390 ;
        RECT 138.080 95.160 138.250 98.160 ;
        RECT 140.720 95.160 140.890 98.160 ;
        RECT 138.465 94.930 140.505 95.100 ;
        RECT 138.080 91.870 138.250 94.870 ;
        RECT 140.720 91.870 140.890 94.870 ;
        RECT 138.465 91.640 140.505 91.810 ;
        RECT 138.080 88.580 138.250 91.580 ;
        RECT 140.720 88.580 140.890 91.580 ;
        RECT 138.465 88.350 140.505 88.520 ;
        RECT 138.080 85.290 138.250 88.290 ;
        RECT 140.720 85.290 140.890 88.290 ;
        RECT 138.465 85.060 140.505 85.230 ;
        RECT 138.080 82.000 138.250 85.000 ;
        RECT 140.720 82.000 140.890 85.000 ;
        RECT 138.465 81.770 140.505 81.940 ;
        RECT 138.080 78.710 138.250 81.710 ;
        RECT 140.720 78.710 140.890 81.710 ;
        RECT 138.465 78.480 140.505 78.650 ;
        RECT 138.080 75.420 138.250 78.420 ;
        RECT 140.720 75.420 140.890 78.420 ;
        RECT 138.465 75.190 140.505 75.360 ;
        RECT 138.080 72.130 138.250 75.130 ;
        RECT 140.720 72.130 140.890 75.130 ;
        RECT 138.465 71.900 140.505 72.070 ;
        RECT 141.230 71.760 141.470 101.800 ;
        RECT 141.230 71.500 141.400 71.760 ;
        RECT 137.570 71.330 141.400 71.500 ;
        RECT 128.390 65.830 131.130 66.000 ;
        RECT 128.390 65.580 128.560 65.830 ;
        RECT 114.150 64.380 116.890 64.550 ;
        RECT 114.150 64.130 114.320 64.380 ;
        RECT 114.000 59.790 114.320 64.130 ;
        RECT 115.000 63.810 116.040 63.980 ;
        RECT 114.660 62.750 114.830 63.750 ;
        RECT 116.210 62.750 116.380 63.750 ;
        RECT 115.000 62.520 116.040 62.690 ;
        RECT 114.660 61.460 114.830 62.460 ;
        RECT 116.210 61.460 116.380 62.460 ;
        RECT 115.000 61.230 116.040 61.400 ;
        RECT 114.660 60.170 114.830 61.170 ;
        RECT 116.210 60.170 116.380 61.170 ;
        RECT 115.000 59.940 116.040 60.110 ;
        RECT 114.150 59.540 114.320 59.790 ;
        RECT 116.720 59.540 116.890 64.380 ;
        RECT 114.150 59.370 116.890 59.540 ;
        RECT 128.320 58.220 128.560 65.580 ;
        RECT 129.240 65.260 130.280 65.430 ;
        RECT 128.900 63.200 129.070 65.200 ;
        RECT 130.450 63.200 130.620 65.200 ;
        RECT 129.240 62.970 130.280 63.140 ;
        RECT 128.900 60.910 129.070 62.910 ;
        RECT 130.450 60.910 130.620 62.910 ;
        RECT 129.240 60.680 130.280 60.850 ;
        RECT 128.900 58.620 129.070 60.620 ;
        RECT 130.450 58.620 130.620 60.620 ;
        RECT 129.240 58.390 130.280 58.560 ;
        RECT 128.390 57.990 128.560 58.220 ;
        RECT 130.960 57.990 131.130 65.830 ;
        RECT 137.220 65.000 140.720 65.170 ;
        RECT 137.220 62.110 137.390 65.000 ;
        RECT 140.550 64.740 140.720 65.000 ;
        RECT 138.115 64.430 139.825 64.600 ;
        RECT 137.730 64.020 137.900 64.370 ;
        RECT 140.040 64.020 140.210 64.370 ;
        RECT 138.115 63.790 139.825 63.960 ;
        RECT 137.730 63.380 137.900 63.730 ;
        RECT 140.040 63.380 140.210 63.730 ;
        RECT 138.115 63.150 139.825 63.320 ;
        RECT 137.730 62.740 137.900 63.090 ;
        RECT 140.040 62.740 140.210 63.090 ;
        RECT 138.115 62.510 139.825 62.680 ;
        RECT 140.550 62.370 140.800 64.740 ;
        RECT 140.550 62.110 140.720 62.370 ;
        RECT 137.220 61.940 140.720 62.110 ;
        RECT 128.390 57.820 131.130 57.990 ;
        RECT 137.020 56.440 140.850 56.610 ;
        RECT 119.920 50.960 122.660 51.130 ;
        RECT 119.920 50.730 120.090 50.960 ;
        RECT 119.690 49.780 120.090 50.730 ;
        RECT 120.430 50.090 120.600 50.420 ;
        RECT 120.770 50.390 121.810 50.560 ;
        RECT 120.770 49.950 121.810 50.120 ;
        RECT 121.980 50.090 122.150 50.420 ;
        RECT 119.920 49.550 120.090 49.780 ;
        RECT 122.490 49.550 122.660 50.960 ;
        RECT 119.920 49.380 122.660 49.550 ;
        RECT 125.250 51.010 129.080 51.180 ;
        RECT 125.250 49.400 125.420 51.010 ;
        RECT 128.910 50.770 129.080 51.010 ;
        RECT 126.145 50.440 128.185 50.610 ;
        RECT 125.760 50.030 125.930 50.380 ;
        RECT 128.400 50.030 128.570 50.380 ;
        RECT 126.145 49.800 128.185 49.970 ;
        RECT 128.910 49.660 129.180 50.770 ;
        RECT 128.910 49.400 129.080 49.660 ;
        RECT 125.250 49.230 129.080 49.400 ;
        RECT 125.250 46.870 129.080 47.040 ;
        RECT 119.920 46.280 123.160 46.450 ;
        RECT 119.920 46.040 120.090 46.280 ;
        RECT 119.670 44.590 120.090 46.040 ;
        RECT 120.430 45.390 120.600 45.720 ;
        RECT 120.770 45.710 122.310 45.880 ;
        RECT 120.770 45.230 122.310 45.400 ;
        RECT 120.770 44.750 122.310 44.920 ;
        RECT 122.480 44.910 122.650 45.240 ;
        RECT 119.920 44.350 120.090 44.590 ;
        RECT 122.990 44.350 123.160 46.280 ;
        RECT 119.920 44.180 123.160 44.350 ;
        RECT 125.250 43.980 125.420 46.870 ;
        RECT 128.910 46.620 129.080 46.870 ;
        RECT 126.145 46.300 128.185 46.470 ;
        RECT 125.760 45.890 125.930 46.240 ;
        RECT 128.400 45.890 128.570 46.240 ;
        RECT 126.145 45.660 128.185 45.830 ;
        RECT 125.760 45.250 125.930 45.600 ;
        RECT 128.400 45.250 128.570 45.600 ;
        RECT 126.145 45.020 128.185 45.190 ;
        RECT 125.760 44.610 125.930 44.960 ;
        RECT 128.400 44.610 128.570 44.960 ;
        RECT 126.145 44.380 128.185 44.550 ;
        RECT 128.910 44.220 129.150 46.620 ;
        RECT 128.910 43.980 129.080 44.220 ;
        RECT 125.250 43.810 129.080 43.980 ;
        RECT 125.250 40.650 130.080 40.820 ;
        RECT 118.480 39.450 123.220 39.620 ;
        RECT 118.480 39.190 118.650 39.450 ;
        RECT 118.160 37.290 118.650 39.190 ;
        RECT 118.990 38.560 119.160 38.890 ;
        RECT 119.330 38.880 122.370 39.050 ;
        RECT 119.330 38.400 122.370 38.570 ;
        RECT 118.990 37.600 119.160 37.930 ;
        RECT 119.330 37.920 122.370 38.090 ;
        RECT 122.540 38.080 122.710 38.410 ;
        RECT 119.330 37.440 122.370 37.610 ;
        RECT 118.480 37.040 118.650 37.290 ;
        RECT 123.050 37.040 123.220 39.450 ;
        RECT 118.480 36.870 123.220 37.040 ;
        RECT 125.250 35.840 125.420 40.650 ;
        RECT 129.910 40.390 130.080 40.650 ;
        RECT 126.145 40.080 129.185 40.250 ;
        RECT 125.760 39.670 125.930 40.020 ;
        RECT 129.400 39.670 129.570 40.020 ;
        RECT 126.145 39.440 129.185 39.610 ;
        RECT 125.760 39.030 125.930 39.380 ;
        RECT 129.400 39.030 129.570 39.380 ;
        RECT 126.145 38.800 129.185 38.970 ;
        RECT 125.760 38.390 125.930 38.740 ;
        RECT 129.400 38.390 129.570 38.740 ;
        RECT 126.145 38.160 129.185 38.330 ;
        RECT 125.760 37.750 125.930 38.100 ;
        RECT 129.400 37.750 129.570 38.100 ;
        RECT 126.145 37.520 129.185 37.690 ;
        RECT 125.760 37.110 125.930 37.460 ;
        RECT 129.400 37.110 129.570 37.460 ;
        RECT 126.145 36.880 129.185 37.050 ;
        RECT 125.760 36.470 125.930 36.820 ;
        RECT 129.400 36.470 129.570 36.820 ;
        RECT 126.145 36.240 129.185 36.410 ;
        RECT 129.910 36.110 130.140 40.390 ;
        RECT 129.910 35.840 130.080 36.110 ;
        RECT 125.250 35.670 130.080 35.840 ;
        RECT 137.020 35.730 137.190 56.440 ;
        RECT 140.680 56.170 140.850 56.440 ;
        RECT 137.915 55.870 139.955 56.040 ;
        RECT 137.530 52.810 137.700 55.810 ;
        RECT 140.170 52.810 140.340 55.810 ;
        RECT 137.915 52.580 139.955 52.750 ;
        RECT 137.530 49.520 137.700 52.520 ;
        RECT 140.170 49.520 140.340 52.520 ;
        RECT 137.915 49.290 139.955 49.460 ;
        RECT 137.530 46.230 137.700 49.230 ;
        RECT 140.170 46.230 140.340 49.230 ;
        RECT 137.915 46.000 139.955 46.170 ;
        RECT 137.530 42.940 137.700 45.940 ;
        RECT 140.170 42.940 140.340 45.940 ;
        RECT 137.915 42.710 139.955 42.880 ;
        RECT 137.530 39.650 137.700 42.650 ;
        RECT 140.170 39.650 140.340 42.650 ;
        RECT 137.915 39.420 139.955 39.590 ;
        RECT 137.530 36.360 137.700 39.360 ;
        RECT 140.170 36.360 140.340 39.360 ;
        RECT 137.915 36.130 139.955 36.300 ;
        RECT 140.680 35.990 140.930 56.170 ;
        RECT 140.680 35.730 140.850 35.990 ;
        RECT 137.020 35.560 140.850 35.730 ;
      LAYER mcon ;
        RECT 111.420 123.700 114.300 123.870 ;
        RECT 111.000 120.720 111.170 123.560 ;
        RECT 114.550 120.720 114.720 123.560 ;
        RECT 111.420 120.410 114.300 120.580 ;
        RECT 120.600 124.270 124.450 124.490 ;
        RECT 121.080 123.700 123.960 123.870 ;
        RECT 120.660 123.460 120.830 123.630 ;
        RECT 121.080 123.220 123.960 123.390 ;
        RECT 124.210 122.980 124.380 123.150 ;
        RECT 121.080 122.740 123.960 122.910 ;
        RECT 120.660 122.500 120.830 122.670 ;
        RECT 121.080 122.260 123.960 122.430 ;
        RECT 124.210 122.020 124.380 122.190 ;
        RECT 121.080 121.780 123.960 121.950 ;
        RECT 120.660 121.540 120.830 121.710 ;
        RECT 121.080 121.300 123.960 121.470 ;
        RECT 124.210 121.060 124.380 121.230 ;
        RECT 121.080 120.820 123.960 120.990 ;
        RECT 120.660 120.580 120.830 120.750 ;
        RECT 121.080 120.340 123.960 120.510 ;
        RECT 129.740 124.270 133.640 124.470 ;
        RECT 130.255 123.700 133.135 123.870 ;
        RECT 129.790 123.370 129.960 123.560 ;
        RECT 133.430 123.370 133.600 123.560 ;
        RECT 130.255 123.060 133.135 123.230 ;
        RECT 129.790 122.730 129.960 122.920 ;
        RECT 133.430 122.730 133.600 122.920 ;
        RECT 130.255 122.420 133.135 122.590 ;
        RECT 129.790 122.090 129.960 122.280 ;
        RECT 133.430 122.090 133.600 122.280 ;
        RECT 130.255 121.780 133.135 121.950 ;
        RECT 129.790 121.450 129.960 121.640 ;
        RECT 133.430 121.450 133.600 121.640 ;
        RECT 130.255 121.140 133.135 121.310 ;
        RECT 129.790 120.810 129.960 121.000 ;
        RECT 133.430 120.810 133.600 121.000 ;
        RECT 130.255 120.500 133.135 120.670 ;
        RECT 129.790 120.170 129.960 120.360 ;
        RECT 133.430 120.170 133.600 120.360 ;
        RECT 130.255 119.860 133.135 120.030 ;
        RECT 129.790 119.530 129.960 119.720 ;
        RECT 133.430 119.530 133.600 119.720 ;
        RECT 130.255 119.220 133.135 119.390 ;
        RECT 138.645 123.590 141.525 123.760 ;
        RECT 138.180 120.610 138.350 123.450 ;
        RECT 141.820 120.610 141.990 123.450 ;
        RECT 138.645 120.300 141.525 120.470 ;
        RECT 112.000 108.530 115.880 108.700 ;
        RECT 111.580 105.550 111.750 108.390 ;
        RECT 116.130 105.550 116.300 108.390 ;
        RECT 112.000 105.240 115.880 105.410 ;
        RECT 111.580 102.260 111.750 105.100 ;
        RECT 116.130 102.260 116.300 105.100 ;
        RECT 112.000 101.950 115.880 102.120 ;
        RECT 111.580 98.970 111.750 101.810 ;
        RECT 116.130 98.970 116.300 101.810 ;
        RECT 112.000 98.660 115.880 98.830 ;
        RECT 112.060 92.930 115.940 93.100 ;
        RECT 111.640 89.950 111.810 92.790 ;
        RECT 116.190 89.950 116.360 92.790 ;
        RECT 112.060 89.640 115.940 89.810 ;
        RECT 111.640 86.660 111.810 89.500 ;
        RECT 116.190 86.660 116.360 89.500 ;
        RECT 112.060 86.350 115.940 86.520 ;
        RECT 111.640 83.370 111.810 86.210 ;
        RECT 116.190 83.370 116.360 86.210 ;
        RECT 112.060 83.060 115.940 83.230 ;
        RECT 122.875 104.880 124.255 105.050 ;
        RECT 122.410 104.200 122.580 104.740 ;
        RECT 124.550 104.200 124.720 104.740 ;
        RECT 122.875 103.890 124.255 104.060 ;
        RECT 122.410 103.210 122.580 103.750 ;
        RECT 124.550 103.210 124.720 103.750 ;
        RECT 122.875 102.900 124.255 103.070 ;
        RECT 122.410 102.220 122.580 102.760 ;
        RECT 124.550 102.220 124.720 102.760 ;
        RECT 122.875 101.910 124.255 102.080 ;
        RECT 122.410 101.230 122.580 101.770 ;
        RECT 124.550 101.230 124.720 101.770 ;
        RECT 122.875 100.920 124.255 101.090 ;
        RECT 122.410 100.240 122.580 100.780 ;
        RECT 124.550 100.240 124.720 100.780 ;
        RECT 122.875 99.930 124.255 100.100 ;
        RECT 122.410 99.250 122.580 99.790 ;
        RECT 124.550 99.250 124.720 99.790 ;
        RECT 122.875 98.940 124.255 99.110 ;
        RECT 122.410 98.260 122.580 98.800 ;
        RECT 124.550 98.260 124.720 98.800 ;
        RECT 122.875 97.950 124.255 98.120 ;
        RECT 122.410 97.270 122.580 97.810 ;
        RECT 124.550 97.270 124.720 97.810 ;
        RECT 122.875 96.960 124.255 97.130 ;
        RECT 122.410 96.280 122.580 96.820 ;
        RECT 124.550 96.280 124.720 96.820 ;
        RECT 122.875 95.970 124.255 96.140 ;
        RECT 122.410 95.290 122.580 95.830 ;
        RECT 124.550 95.290 124.720 95.830 ;
        RECT 122.875 94.980 124.255 95.150 ;
        RECT 122.410 94.300 122.580 94.840 ;
        RECT 124.550 94.300 124.720 94.840 ;
        RECT 122.875 93.990 124.255 94.160 ;
        RECT 122.410 93.310 122.580 93.850 ;
        RECT 124.550 93.310 124.720 93.850 ;
        RECT 122.875 93.000 124.255 93.170 ;
        RECT 122.410 92.320 122.580 92.860 ;
        RECT 124.550 92.320 124.720 92.860 ;
        RECT 122.875 92.010 124.255 92.180 ;
        RECT 122.410 91.330 122.580 91.870 ;
        RECT 124.550 91.330 124.720 91.870 ;
        RECT 122.875 91.020 124.255 91.190 ;
        RECT 122.410 90.340 122.580 90.880 ;
        RECT 124.550 90.340 124.720 90.880 ;
        RECT 122.875 90.030 124.255 90.200 ;
        RECT 122.410 89.350 122.580 89.890 ;
        RECT 124.550 89.350 124.720 89.890 ;
        RECT 122.875 89.040 124.255 89.210 ;
        RECT 122.410 88.360 122.580 88.900 ;
        RECT 124.550 88.360 124.720 88.900 ;
        RECT 122.875 88.050 124.255 88.220 ;
        RECT 122.410 87.370 122.580 87.910 ;
        RECT 124.550 87.370 124.720 87.910 ;
        RECT 122.875 87.060 124.255 87.230 ;
        RECT 130.705 104.880 132.085 105.050 ;
        RECT 130.240 104.200 130.410 104.740 ;
        RECT 132.380 104.200 132.550 104.740 ;
        RECT 130.705 103.890 132.085 104.060 ;
        RECT 130.240 103.210 130.410 103.750 ;
        RECT 132.380 103.210 132.550 103.750 ;
        RECT 130.705 102.900 132.085 103.070 ;
        RECT 130.240 102.220 130.410 102.760 ;
        RECT 132.380 102.220 132.550 102.760 ;
        RECT 130.705 101.910 132.085 102.080 ;
        RECT 130.240 101.230 130.410 101.770 ;
        RECT 132.380 101.230 132.550 101.770 ;
        RECT 130.705 100.920 132.085 101.090 ;
        RECT 130.240 100.240 130.410 100.780 ;
        RECT 132.380 100.240 132.550 100.780 ;
        RECT 130.705 99.930 132.085 100.100 ;
        RECT 130.240 99.250 130.410 99.790 ;
        RECT 132.380 99.250 132.550 99.790 ;
        RECT 130.705 98.940 132.085 99.110 ;
        RECT 130.240 98.260 130.410 98.800 ;
        RECT 132.380 98.260 132.550 98.800 ;
        RECT 130.705 97.950 132.085 98.120 ;
        RECT 130.240 97.270 130.410 97.810 ;
        RECT 132.380 97.270 132.550 97.810 ;
        RECT 130.705 96.960 132.085 97.130 ;
        RECT 130.240 96.280 130.410 96.820 ;
        RECT 132.380 96.280 132.550 96.820 ;
        RECT 130.705 95.970 132.085 96.140 ;
        RECT 130.240 95.290 130.410 95.830 ;
        RECT 132.380 95.290 132.550 95.830 ;
        RECT 130.705 94.980 132.085 95.150 ;
        RECT 130.240 94.300 130.410 94.840 ;
        RECT 132.380 94.300 132.550 94.840 ;
        RECT 130.705 93.990 132.085 94.160 ;
        RECT 130.240 93.310 130.410 93.850 ;
        RECT 132.380 93.310 132.550 93.850 ;
        RECT 130.705 93.000 132.085 93.170 ;
        RECT 130.240 92.320 130.410 92.860 ;
        RECT 132.380 92.320 132.550 92.860 ;
        RECT 130.705 92.010 132.085 92.180 ;
        RECT 130.240 91.330 130.410 91.870 ;
        RECT 132.380 91.330 132.550 91.870 ;
        RECT 130.705 91.020 132.085 91.190 ;
        RECT 130.240 90.340 130.410 90.880 ;
        RECT 132.380 90.340 132.550 90.880 ;
        RECT 130.705 90.030 132.085 90.200 ;
        RECT 130.240 89.350 130.410 89.890 ;
        RECT 132.380 89.350 132.550 89.890 ;
        RECT 130.705 89.040 132.085 89.210 ;
        RECT 130.240 88.360 130.410 88.900 ;
        RECT 132.380 88.360 132.550 88.900 ;
        RECT 130.705 88.050 132.085 88.220 ;
        RECT 130.240 87.370 130.410 87.910 ;
        RECT 132.380 87.370 132.550 87.910 ;
        RECT 130.705 87.060 132.085 87.230 ;
        RECT 115.050 77.780 115.930 77.950 ;
        RECT 114.630 76.800 114.800 77.640 ;
        RECT 116.180 76.800 116.350 77.640 ;
        RECT 115.050 76.490 115.930 76.660 ;
        RECT 114.630 75.510 114.800 76.350 ;
        RECT 116.180 75.510 116.350 76.350 ;
        RECT 115.050 75.200 115.930 75.370 ;
        RECT 114.630 74.220 114.800 75.060 ;
        RECT 116.180 74.220 116.350 75.060 ;
        RECT 115.050 73.910 115.930 74.080 ;
        RECT 128.235 78.290 130.255 78.460 ;
        RECT 127.770 77.960 127.940 78.150 ;
        RECT 130.550 77.960 130.720 78.150 ;
        RECT 128.235 77.650 130.255 77.820 ;
        RECT 127.770 77.320 127.940 77.510 ;
        RECT 130.550 77.320 130.720 77.510 ;
        RECT 128.235 77.010 130.255 77.180 ;
        RECT 127.770 76.680 127.940 76.870 ;
        RECT 130.550 76.680 130.720 76.870 ;
        RECT 128.235 76.370 130.255 76.540 ;
        RECT 127.770 76.040 127.940 76.230 ;
        RECT 130.550 76.040 130.720 76.230 ;
        RECT 128.235 75.730 130.255 75.900 ;
        RECT 127.770 75.400 127.940 75.590 ;
        RECT 130.550 75.400 130.720 75.590 ;
        RECT 128.235 75.090 130.255 75.260 ;
        RECT 127.770 74.760 127.940 74.950 ;
        RECT 130.550 74.760 130.720 74.950 ;
        RECT 128.235 74.450 130.255 74.620 ;
        RECT 127.770 74.120 127.940 74.310 ;
        RECT 130.550 74.120 130.720 74.310 ;
        RECT 128.235 73.810 130.255 73.980 ;
        RECT 138.545 101.510 140.425 101.680 ;
        RECT 138.080 98.530 138.250 101.370 ;
        RECT 140.720 98.530 140.890 101.370 ;
        RECT 138.545 98.220 140.425 98.390 ;
        RECT 138.080 95.240 138.250 98.080 ;
        RECT 140.720 95.240 140.890 98.080 ;
        RECT 138.545 94.930 140.425 95.100 ;
        RECT 138.080 91.950 138.250 94.790 ;
        RECT 140.720 91.950 140.890 94.790 ;
        RECT 138.545 91.640 140.425 91.810 ;
        RECT 138.080 88.660 138.250 91.500 ;
        RECT 140.720 88.660 140.890 91.500 ;
        RECT 138.545 88.350 140.425 88.520 ;
        RECT 138.080 85.370 138.250 88.210 ;
        RECT 140.720 85.370 140.890 88.210 ;
        RECT 138.545 85.060 140.425 85.230 ;
        RECT 138.080 82.080 138.250 84.920 ;
        RECT 140.720 82.080 140.890 84.920 ;
        RECT 138.545 81.770 140.425 81.940 ;
        RECT 138.080 78.790 138.250 81.630 ;
        RECT 140.720 78.790 140.890 81.630 ;
        RECT 138.545 78.480 140.425 78.650 ;
        RECT 138.080 75.500 138.250 78.340 ;
        RECT 140.720 75.500 140.890 78.340 ;
        RECT 138.545 75.190 140.425 75.360 ;
        RECT 138.080 72.210 138.250 75.050 ;
        RECT 140.720 72.210 140.890 75.050 ;
        RECT 138.545 71.900 140.425 72.070 ;
        RECT 115.080 63.810 115.960 63.980 ;
        RECT 114.660 62.830 114.830 63.670 ;
        RECT 116.210 62.830 116.380 63.670 ;
        RECT 115.080 62.520 115.960 62.690 ;
        RECT 114.660 61.540 114.830 62.380 ;
        RECT 116.210 61.540 116.380 62.380 ;
        RECT 115.080 61.230 115.960 61.400 ;
        RECT 114.660 60.250 114.830 61.090 ;
        RECT 116.210 60.250 116.380 61.090 ;
        RECT 115.080 59.940 115.960 60.110 ;
        RECT 129.320 65.260 130.200 65.430 ;
        RECT 128.900 63.280 129.070 65.120 ;
        RECT 130.450 63.280 130.620 65.120 ;
        RECT 129.320 62.970 130.200 63.140 ;
        RECT 128.900 60.990 129.070 62.830 ;
        RECT 130.450 60.990 130.620 62.830 ;
        RECT 129.320 60.680 130.200 60.850 ;
        RECT 128.900 58.700 129.070 60.540 ;
        RECT 130.450 58.700 130.620 60.540 ;
        RECT 129.320 58.390 130.200 58.560 ;
        RECT 138.195 64.430 139.745 64.600 ;
        RECT 137.730 64.100 137.900 64.290 ;
        RECT 140.040 64.100 140.210 64.290 ;
        RECT 138.195 63.790 139.745 63.960 ;
        RECT 137.730 63.460 137.900 63.650 ;
        RECT 140.040 63.460 140.210 63.650 ;
        RECT 138.195 63.150 139.745 63.320 ;
        RECT 137.730 62.820 137.900 63.010 ;
        RECT 140.040 62.820 140.210 63.010 ;
        RECT 138.195 62.510 139.745 62.680 ;
        RECT 120.850 50.390 121.730 50.560 ;
        RECT 120.430 50.170 120.600 50.340 ;
        RECT 121.980 50.170 122.150 50.340 ;
        RECT 120.850 49.950 121.730 50.120 ;
        RECT 126.225 50.440 128.105 50.610 ;
        RECT 125.760 50.110 125.930 50.300 ;
        RECT 128.400 50.110 128.570 50.300 ;
        RECT 126.225 49.800 128.105 49.970 ;
        RECT 120.850 45.710 122.230 45.880 ;
        RECT 120.430 45.470 120.600 45.640 ;
        RECT 120.850 45.230 122.230 45.400 ;
        RECT 122.480 44.990 122.650 45.160 ;
        RECT 120.850 44.750 122.230 44.920 ;
        RECT 126.225 46.300 128.105 46.470 ;
        RECT 125.760 45.970 125.930 46.160 ;
        RECT 128.400 45.970 128.570 46.160 ;
        RECT 126.225 45.660 128.105 45.830 ;
        RECT 125.760 45.330 125.930 45.520 ;
        RECT 128.400 45.330 128.570 45.520 ;
        RECT 126.225 45.020 128.105 45.190 ;
        RECT 125.760 44.690 125.930 44.880 ;
        RECT 128.400 44.690 128.570 44.880 ;
        RECT 126.225 44.380 128.105 44.550 ;
        RECT 119.410 38.880 122.290 39.050 ;
        RECT 118.990 38.640 119.160 38.810 ;
        RECT 119.410 38.400 122.290 38.570 ;
        RECT 122.540 38.160 122.710 38.330 ;
        RECT 119.410 37.920 122.290 38.090 ;
        RECT 118.990 37.680 119.160 37.850 ;
        RECT 119.410 37.440 122.290 37.610 ;
        RECT 126.225 40.080 129.105 40.250 ;
        RECT 125.760 39.750 125.930 39.940 ;
        RECT 129.400 39.750 129.570 39.940 ;
        RECT 126.225 39.440 129.105 39.610 ;
        RECT 125.760 39.110 125.930 39.300 ;
        RECT 129.400 39.110 129.570 39.300 ;
        RECT 126.225 38.800 129.105 38.970 ;
        RECT 125.760 38.470 125.930 38.660 ;
        RECT 129.400 38.470 129.570 38.660 ;
        RECT 126.225 38.160 129.105 38.330 ;
        RECT 125.760 37.830 125.930 38.020 ;
        RECT 129.400 37.830 129.570 38.020 ;
        RECT 126.225 37.520 129.105 37.690 ;
        RECT 125.760 37.190 125.930 37.380 ;
        RECT 129.400 37.190 129.570 37.380 ;
        RECT 126.225 36.880 129.105 37.050 ;
        RECT 125.760 36.550 125.930 36.740 ;
        RECT 129.400 36.550 129.570 36.740 ;
        RECT 126.225 36.240 129.105 36.410 ;
        RECT 137.995 55.870 139.875 56.040 ;
        RECT 137.530 52.890 137.700 55.730 ;
        RECT 140.170 52.890 140.340 55.730 ;
        RECT 137.995 52.580 139.875 52.750 ;
        RECT 137.530 49.600 137.700 52.440 ;
        RECT 140.170 49.600 140.340 52.440 ;
        RECT 137.995 49.290 139.875 49.460 ;
        RECT 137.530 46.310 137.700 49.150 ;
        RECT 140.170 46.310 140.340 49.150 ;
        RECT 137.995 46.000 139.875 46.170 ;
        RECT 137.530 43.020 137.700 45.860 ;
        RECT 140.170 43.020 140.340 45.860 ;
        RECT 137.995 42.710 139.875 42.880 ;
        RECT 137.530 39.730 137.700 42.570 ;
        RECT 140.170 39.730 140.340 42.570 ;
        RECT 137.995 39.420 139.875 39.590 ;
        RECT 137.530 36.440 137.700 39.280 ;
        RECT 140.170 36.440 140.340 39.280 ;
        RECT 137.995 36.130 139.875 36.300 ;
        RECT 140.690 35.990 140.930 56.170 ;
      LAYER met1 ;
        RECT 125.375 142.105 146.405 144.780 ;
        RECT 96.015 134.595 108.445 137.125 ;
        RECT 105.915 129.020 108.445 134.595 ;
        RECT 126.500 132.060 137.435 133.545 ;
        RECT 126.500 129.370 127.985 132.060 ;
        RECT 105.230 129.010 109.250 129.020 ;
        RECT 105.230 126.730 124.730 129.010 ;
        RECT 105.230 126.650 124.740 126.730 ;
        RECT 105.230 124.250 109.250 126.650 ;
        RECT 105.230 120.010 110.690 124.250 ;
        RECT 111.400 123.900 114.330 126.650 ;
        RECT 120.410 124.240 124.740 126.650 ;
        RECT 123.530 123.900 124.020 123.960 ;
        RECT 111.360 123.670 114.360 123.900 ;
        RECT 105.230 108.880 109.250 120.010 ;
        RECT 110.970 117.450 111.210 123.640 ;
        RECT 111.430 120.610 114.330 120.630 ;
        RECT 111.360 120.380 114.360 120.610 ;
        RECT 111.430 120.210 114.330 120.380 ;
        RECT 112.080 119.380 112.920 120.210 ;
        RECT 112.085 117.450 112.915 119.380 ;
        RECT 114.510 117.450 114.810 123.650 ;
        RECT 118.160 118.660 118.780 119.220 ;
        RECT 118.190 117.450 118.750 118.660 ;
        RECT 110.970 116.850 118.750 117.450 ;
        RECT 120.510 117.410 120.860 123.720 ;
        RECT 121.020 123.670 124.020 123.900 ;
        RECT 123.530 123.570 124.020 123.670 ;
        RECT 121.090 123.420 121.580 123.500 ;
        RECT 121.020 123.190 124.020 123.420 ;
        RECT 121.090 123.110 121.580 123.190 ;
        RECT 123.530 122.940 124.020 123.020 ;
        RECT 121.020 122.710 124.020 122.940 ;
        RECT 123.530 122.630 124.020 122.710 ;
        RECT 121.090 122.460 121.580 122.540 ;
        RECT 121.020 122.230 124.020 122.460 ;
        RECT 121.090 122.150 121.580 122.230 ;
        RECT 123.530 121.980 124.020 122.060 ;
        RECT 121.020 121.750 124.020 121.980 ;
        RECT 123.530 121.670 124.020 121.750 ;
        RECT 121.090 121.500 121.580 121.580 ;
        RECT 121.020 121.270 124.020 121.500 ;
        RECT 121.090 121.190 121.580 121.270 ;
        RECT 123.530 121.020 124.020 121.100 ;
        RECT 121.020 120.790 124.020 121.020 ;
        RECT 123.530 120.710 124.020 120.790 ;
        RECT 121.090 120.540 121.580 120.620 ;
        RECT 121.020 120.310 124.020 120.540 ;
        RECT 121.090 120.230 121.580 120.310 ;
        RECT 122.715 117.410 123.285 119.310 ;
        RECT 124.160 117.410 124.510 123.270 ;
        RECT 126.450 120.120 128.015 129.370 ;
        RECT 143.730 129.160 146.405 142.105 ;
        RECT 129.670 126.870 147.320 129.160 ;
        RECT 129.660 126.800 147.320 126.870 ;
        RECT 129.660 124.200 133.680 126.800 ;
        RECT 130.270 123.900 130.750 123.910 ;
        RECT 129.690 118.030 130.000 123.700 ;
        RECT 130.195 123.670 133.195 123.900 ;
        RECT 138.780 123.790 141.310 126.800 ;
        RECT 143.300 124.330 147.320 126.800 ;
        RECT 130.270 123.530 130.750 123.670 ;
        RECT 132.670 123.260 133.150 123.340 ;
        RECT 130.195 123.030 133.195 123.260 ;
        RECT 132.670 122.960 133.150 123.030 ;
        RECT 130.250 122.620 130.730 122.690 ;
        RECT 130.195 122.390 133.195 122.620 ;
        RECT 130.250 122.310 130.730 122.390 ;
        RECT 132.670 121.980 133.150 122.050 ;
        RECT 130.195 121.750 133.195 121.980 ;
        RECT 132.670 121.670 133.150 121.750 ;
        RECT 130.250 121.340 130.730 121.420 ;
        RECT 130.195 121.110 133.195 121.340 ;
        RECT 130.250 121.040 130.730 121.110 ;
        RECT 132.670 120.700 133.150 120.780 ;
        RECT 130.195 120.470 133.195 120.700 ;
        RECT 132.670 120.400 133.150 120.470 ;
        RECT 130.250 120.060 130.730 120.130 ;
        RECT 130.195 119.830 133.195 120.060 ;
        RECT 130.250 119.750 130.730 119.830 ;
        RECT 132.670 119.420 133.150 119.500 ;
        RECT 130.195 119.190 133.195 119.420 ;
        RECT 132.670 119.120 133.150 119.190 ;
        RECT 129.690 117.450 130.830 118.030 ;
        RECT 129.690 117.410 130.800 117.450 ;
        RECT 120.500 117.140 130.800 117.410 ;
        RECT 133.350 117.140 133.660 123.700 ;
        RECT 138.110 123.510 138.360 123.590 ;
        RECT 138.585 123.560 141.585 123.790 ;
        RECT 141.760 123.510 142.010 123.590 ;
        RECT 138.110 120.550 138.380 123.510 ;
        RECT 141.760 120.550 142.020 123.510 ;
        RECT 138.110 118.900 138.360 120.550 ;
        RECT 138.585 120.270 141.585 120.500 ;
        RECT 139.730 118.900 140.880 120.270 ;
        RECT 141.760 118.900 142.010 120.550 ;
        RECT 142.300 119.710 147.320 124.330 ;
        RECT 138.110 118.725 142.010 118.900 ;
        RECT 136.015 118.175 142.015 118.725 ;
        RECT 135.140 117.990 135.680 118.020 ;
        RECT 136.015 117.990 136.565 118.175 ;
        RECT 135.140 117.450 136.565 117.990 ;
        RECT 135.140 117.420 135.680 117.450 ;
        RECT 136.015 117.445 136.565 117.450 ;
        RECT 110.970 116.770 118.730 116.850 ;
        RECT 120.500 116.830 133.665 117.140 ;
        RECT 120.500 116.810 130.140 116.830 ;
        RECT 115.500 114.260 116.430 116.770 ;
        RECT 140.330 115.085 140.920 118.175 ;
        RECT 140.300 114.495 140.950 115.085 ;
        RECT 115.500 113.320 119.430 114.260 ;
        RECT 115.500 112.250 116.430 113.320 ;
        RECT 111.550 110.810 116.440 112.250 ;
        RECT 105.230 98.440 111.270 108.880 ;
        RECT 111.550 98.880 111.800 110.810 ;
        RECT 115.240 108.730 115.870 108.820 ;
        RECT 111.940 108.500 115.940 108.730 ;
        RECT 115.240 108.400 115.870 108.500 ;
        RECT 112.010 105.440 112.640 105.550 ;
        RECT 111.940 105.210 115.940 105.440 ;
        RECT 112.010 105.130 112.640 105.210 ;
        RECT 115.240 102.150 115.870 102.240 ;
        RECT 111.940 101.920 115.940 102.150 ;
        RECT 115.240 101.820 115.870 101.920 ;
        RECT 112.010 98.860 112.640 98.940 ;
        RECT 111.940 98.630 115.940 98.860 ;
        RECT 116.100 98.680 116.440 110.810 ;
        RECT 112.010 98.520 112.640 98.630 ;
        RECT 105.230 97.260 109.250 98.440 ;
        RECT 105.230 96.510 112.740 97.260 ;
        RECT 105.230 93.430 109.250 96.510 ;
        RECT 116.150 95.150 116.530 95.160 ;
        RECT 118.490 95.150 119.430 113.320 ;
        RECT 125.470 110.200 126.860 110.205 ;
        RECT 133.180 110.200 134.770 110.205 ;
        RECT 143.300 110.200 147.320 119.710 ;
        RECT 125.470 106.980 147.320 110.200 ;
        RECT 125.470 105.300 126.860 106.980 ;
        RECT 123.850 105.080 124.260 105.160 ;
        RECT 111.610 94.210 119.430 95.150 ;
        RECT 105.230 82.830 111.330 93.430 ;
        RECT 111.610 83.310 111.860 94.210 ;
        RECT 115.240 93.130 115.950 93.240 ;
        RECT 112.000 92.900 116.000 93.130 ;
        RECT 115.240 92.770 115.950 92.900 ;
        RECT 112.060 89.840 112.770 89.950 ;
        RECT 112.000 89.610 116.000 89.840 ;
        RECT 112.060 89.480 112.770 89.610 ;
        RECT 115.240 86.550 115.950 86.670 ;
        RECT 112.000 86.320 116.000 86.550 ;
        RECT 115.240 86.200 115.950 86.320 ;
        RECT 112.060 83.260 112.770 83.380 ;
        RECT 112.000 83.030 116.000 83.260 ;
        RECT 116.150 83.190 116.530 94.210 ;
        RECT 122.310 85.390 122.630 104.880 ;
        RECT 122.815 104.850 124.315 105.080 ;
        RECT 123.850 104.770 124.260 104.850 ;
        RECT 122.870 104.090 123.280 104.170 ;
        RECT 122.815 103.860 124.315 104.090 ;
        RECT 122.870 103.780 123.280 103.860 ;
        RECT 123.850 103.100 124.260 103.180 ;
        RECT 122.815 102.870 124.315 103.100 ;
        RECT 123.850 102.790 124.260 102.870 ;
        RECT 122.870 102.110 123.280 102.190 ;
        RECT 122.815 101.880 124.315 102.110 ;
        RECT 122.870 101.800 123.280 101.880 ;
        RECT 123.850 101.120 124.260 101.200 ;
        RECT 122.815 100.890 124.315 101.120 ;
        RECT 123.850 100.810 124.260 100.890 ;
        RECT 122.870 100.130 123.280 100.210 ;
        RECT 122.815 99.900 124.315 100.130 ;
        RECT 122.870 99.820 123.280 99.900 ;
        RECT 123.850 99.140 124.260 99.220 ;
        RECT 122.815 98.910 124.315 99.140 ;
        RECT 123.850 98.830 124.260 98.910 ;
        RECT 122.870 98.150 123.280 98.240 ;
        RECT 122.815 97.920 124.315 98.150 ;
        RECT 122.870 97.850 123.280 97.920 ;
        RECT 123.850 97.160 124.260 97.240 ;
        RECT 122.815 96.930 124.315 97.160 ;
        RECT 123.850 96.850 124.260 96.930 ;
        RECT 122.870 96.170 123.280 96.260 ;
        RECT 122.815 95.940 124.315 96.170 ;
        RECT 122.870 95.870 123.280 95.940 ;
        RECT 123.850 95.180 124.260 95.260 ;
        RECT 122.815 94.950 124.315 95.180 ;
        RECT 123.850 94.870 124.260 94.950 ;
        RECT 122.870 94.190 123.280 94.270 ;
        RECT 122.815 93.960 124.315 94.190 ;
        RECT 122.870 93.880 123.280 93.960 ;
        RECT 123.850 93.200 124.260 93.280 ;
        RECT 122.815 92.970 124.315 93.200 ;
        RECT 123.850 92.890 124.260 92.970 ;
        RECT 122.870 92.210 123.280 92.300 ;
        RECT 122.815 91.980 124.315 92.210 ;
        RECT 122.870 91.910 123.280 91.980 ;
        RECT 123.850 91.220 124.260 91.300 ;
        RECT 122.815 90.990 124.315 91.220 ;
        RECT 123.850 90.910 124.260 90.990 ;
        RECT 122.870 90.230 123.280 90.310 ;
        RECT 122.815 90.000 124.315 90.230 ;
        RECT 122.870 89.920 123.280 90.000 ;
        RECT 123.850 89.240 124.260 89.320 ;
        RECT 122.815 89.010 124.315 89.240 ;
        RECT 123.850 88.930 124.260 89.010 ;
        RECT 122.870 88.250 123.280 88.330 ;
        RECT 122.815 88.020 124.315 88.250 ;
        RECT 122.870 87.940 123.280 88.020 ;
        RECT 123.850 87.260 124.260 87.340 ;
        RECT 122.815 87.030 124.315 87.260 ;
        RECT 123.850 86.950 124.260 87.030 ;
        RECT 124.470 85.390 124.790 104.880 ;
        RECT 125.000 86.750 126.860 105.300 ;
        RECT 133.180 105.180 134.770 106.980 ;
        RECT 131.640 105.080 132.170 105.160 ;
        RECT 130.645 104.850 132.170 105.080 ;
        RECT 130.130 85.390 130.450 104.820 ;
        RECT 131.640 104.770 132.170 104.850 ;
        RECT 130.680 104.090 131.210 104.170 ;
        RECT 130.645 103.860 132.145 104.090 ;
        RECT 130.680 103.780 131.210 103.860 ;
        RECT 131.640 103.100 132.170 103.180 ;
        RECT 130.645 102.870 132.170 103.100 ;
        RECT 131.640 102.790 132.170 102.870 ;
        RECT 130.680 102.110 131.210 102.200 ;
        RECT 130.645 101.880 132.145 102.110 ;
        RECT 130.680 101.810 131.210 101.880 ;
        RECT 131.640 101.120 132.170 101.200 ;
        RECT 130.645 100.890 132.170 101.120 ;
        RECT 131.640 100.810 132.170 100.890 ;
        RECT 130.680 100.130 131.210 100.220 ;
        RECT 130.645 99.900 132.145 100.130 ;
        RECT 130.680 99.830 131.210 99.900 ;
        RECT 131.640 99.140 132.170 99.230 ;
        RECT 130.645 98.910 132.170 99.140 ;
        RECT 131.640 98.840 132.170 98.910 ;
        RECT 130.680 98.150 131.210 98.230 ;
        RECT 130.645 97.920 132.145 98.150 ;
        RECT 130.680 97.840 131.210 97.920 ;
        RECT 131.640 97.160 132.170 97.250 ;
        RECT 130.645 96.930 132.170 97.160 ;
        RECT 131.640 96.860 132.170 96.930 ;
        RECT 130.680 96.170 131.210 96.250 ;
        RECT 130.645 95.940 132.145 96.170 ;
        RECT 130.680 95.860 131.210 95.940 ;
        RECT 131.640 95.180 132.170 95.260 ;
        RECT 130.645 94.950 132.170 95.180 ;
        RECT 131.640 94.870 132.170 94.950 ;
        RECT 130.680 94.190 131.210 94.280 ;
        RECT 130.645 93.960 132.145 94.190 ;
        RECT 130.680 93.890 131.210 93.960 ;
        RECT 131.640 93.200 132.170 93.280 ;
        RECT 130.645 92.970 132.170 93.200 ;
        RECT 131.640 92.890 132.170 92.970 ;
        RECT 130.680 92.210 131.210 92.300 ;
        RECT 130.645 91.980 132.145 92.210 ;
        RECT 130.680 91.910 131.210 91.980 ;
        RECT 131.640 91.220 132.170 91.310 ;
        RECT 130.645 90.990 132.170 91.220 ;
        RECT 131.640 90.920 132.170 90.990 ;
        RECT 130.680 90.230 131.210 90.320 ;
        RECT 130.645 90.000 132.145 90.230 ;
        RECT 130.680 89.930 131.210 90.000 ;
        RECT 131.640 89.240 132.170 89.320 ;
        RECT 130.645 89.010 132.170 89.240 ;
        RECT 131.640 88.930 132.170 89.010 ;
        RECT 130.680 88.250 131.210 88.340 ;
        RECT 130.645 88.020 132.145 88.250 ;
        RECT 130.680 87.950 131.210 88.020 ;
        RECT 131.640 87.260 132.170 87.340 ;
        RECT 130.645 87.030 132.170 87.260 ;
        RECT 131.640 86.950 132.170 87.030 ;
        RECT 132.340 85.390 132.660 104.840 ;
        RECT 132.810 87.650 134.770 105.180 ;
        RECT 140.330 103.670 140.920 104.725 ;
        RECT 138.050 103.080 140.920 103.670 ;
        RECT 132.810 86.890 134.790 87.650 ;
        RECT 122.290 84.925 132.670 85.390 ;
        RECT 121.135 84.330 132.670 84.925 ;
        RECT 121.135 84.300 125.770 84.330 ;
        RECT 121.135 84.235 125.765 84.300 ;
        RECT 112.060 82.910 112.770 83.030 ;
        RECT 105.230 81.330 109.250 82.830 ;
        RECT 121.135 82.495 121.825 84.235 ;
        RECT 105.230 80.530 112.850 81.330 ;
        RECT 105.230 78.170 109.250 80.530 ;
        RECT 127.710 80.450 128.380 81.875 ;
        RECT 127.710 79.780 130.770 80.450 ;
        RECT 115.040 79.420 115.400 79.450 ;
        RECT 113.400 79.060 115.400 79.420 ;
        RECT 113.400 78.170 113.760 79.060 ;
        RECT 115.040 79.030 115.400 79.060 ;
        RECT 105.230 73.660 114.320 78.170 ;
        RECT 115.590 77.980 116.000 78.060 ;
        RECT 105.230 64.310 109.250 73.660 ;
        RECT 114.600 72.800 114.840 77.790 ;
        RECT 114.990 77.750 116.000 77.980 ;
        RECT 115.590 77.680 116.000 77.750 ;
        RECT 115.000 76.690 115.410 76.760 ;
        RECT 114.990 76.460 115.990 76.690 ;
        RECT 115.000 76.380 115.410 76.460 ;
        RECT 115.590 75.400 116.000 75.470 ;
        RECT 114.990 75.170 116.000 75.400 ;
        RECT 115.590 75.090 116.000 75.170 ;
        RECT 114.990 74.110 115.400 74.190 ;
        RECT 114.990 73.880 115.990 74.110 ;
        RECT 114.990 73.810 115.400 73.880 ;
        RECT 116.140 72.800 116.380 77.790 ;
        RECT 127.710 73.960 127.980 79.780 ;
        RECT 129.670 78.490 130.330 78.580 ;
        RECT 128.175 78.260 130.330 78.490 ;
        RECT 129.670 78.180 130.330 78.260 ;
        RECT 128.180 77.850 128.840 77.940 ;
        RECT 128.175 77.620 130.315 77.850 ;
        RECT 128.180 77.540 128.840 77.620 ;
        RECT 129.670 77.210 130.330 77.300 ;
        RECT 128.175 76.980 130.330 77.210 ;
        RECT 129.670 76.900 130.330 76.980 ;
        RECT 128.180 76.570 128.840 76.650 ;
        RECT 128.175 76.340 130.315 76.570 ;
        RECT 128.180 76.250 128.840 76.340 ;
        RECT 129.670 75.930 130.330 76.020 ;
        RECT 128.175 75.700 130.330 75.930 ;
        RECT 129.670 75.620 130.330 75.700 ;
        RECT 128.170 75.290 128.830 75.380 ;
        RECT 128.170 75.060 130.315 75.290 ;
        RECT 128.170 74.980 128.830 75.060 ;
        RECT 129.670 74.650 130.330 74.740 ;
        RECT 128.175 74.420 130.330 74.650 ;
        RECT 129.670 74.340 130.330 74.420 ;
        RECT 128.180 74.010 128.840 74.100 ;
        RECT 128.175 73.780 130.315 74.010 ;
        RECT 130.500 73.960 130.770 79.780 ;
        RECT 133.630 78.700 134.790 86.890 ;
        RECT 131.030 77.540 134.790 78.700 ;
        RECT 128.180 73.700 128.840 73.780 ;
        RECT 131.030 73.540 132.480 77.540 ;
        RECT 114.600 72.710 116.380 72.800 ;
        RECT 118.525 72.710 119.255 72.740 ;
        RECT 114.600 71.980 119.255 72.710 ;
        RECT 138.050 72.090 138.280 103.080 ;
        RECT 139.890 101.710 140.490 101.790 ;
        RECT 138.485 101.480 140.490 101.710 ;
        RECT 139.890 101.400 140.490 101.480 ;
        RECT 138.490 98.420 139.090 98.500 ;
        RECT 138.485 98.190 140.485 98.420 ;
        RECT 138.490 98.110 139.090 98.190 ;
        RECT 139.890 95.130 140.490 95.210 ;
        RECT 138.485 94.900 140.490 95.130 ;
        RECT 139.890 94.820 140.490 94.900 ;
        RECT 138.490 91.840 139.090 91.930 ;
        RECT 138.485 91.610 140.485 91.840 ;
        RECT 138.490 91.540 139.090 91.610 ;
        RECT 139.890 88.550 140.490 88.640 ;
        RECT 138.485 88.320 140.490 88.550 ;
        RECT 139.890 88.250 140.490 88.320 ;
        RECT 138.490 85.260 139.090 85.340 ;
        RECT 138.485 85.030 140.485 85.260 ;
        RECT 138.490 84.950 139.090 85.030 ;
        RECT 139.890 81.970 140.490 82.050 ;
        RECT 138.485 81.740 140.490 81.970 ;
        RECT 139.890 81.660 140.490 81.740 ;
        RECT 138.490 78.680 139.090 78.760 ;
        RECT 138.485 78.450 140.485 78.680 ;
        RECT 138.490 78.370 139.090 78.450 ;
        RECT 139.890 75.390 140.490 75.480 ;
        RECT 138.485 75.160 140.490 75.390 ;
        RECT 139.890 75.090 140.490 75.160 ;
        RECT 138.490 72.100 139.090 72.180 ;
        RECT 114.600 71.940 116.380 71.980 ;
        RECT 118.525 71.950 119.255 71.980 ;
        RECT 138.485 71.870 140.485 72.100 ;
        RECT 140.690 72.090 140.920 103.080 ;
        RECT 143.300 101.930 147.320 106.980 ;
        RECT 138.490 71.790 139.090 71.870 ;
        RECT 141.200 71.640 147.320 101.930 ;
        RECT 115.130 69.530 124.830 69.680 ;
        RECT 111.090 68.140 124.830 69.530 ;
        RECT 143.300 68.900 147.320 71.640 ;
        RECT 139.820 68.200 147.320 68.900 ;
        RECT 111.090 68.070 116.770 68.140 ;
        RECT 112.675 64.310 113.405 66.535 ;
        RECT 143.300 66.435 147.320 68.200 ;
        RECT 140.725 65.745 147.320 66.435 ;
        RECT 114.630 65.110 120.895 65.620 ;
        RECT 105.230 59.610 114.340 64.310 ;
        RECT 114.630 60.130 114.870 65.110 ;
        RECT 115.020 64.010 115.390 64.090 ;
        RECT 115.020 63.780 116.020 64.010 ;
        RECT 115.020 63.710 115.390 63.780 ;
        RECT 115.650 62.720 116.020 62.800 ;
        RECT 115.020 62.490 116.020 62.720 ;
        RECT 115.650 62.420 116.020 62.490 ;
        RECT 115.010 61.430 115.380 61.510 ;
        RECT 115.010 61.200 116.020 61.430 ;
        RECT 115.010 61.130 115.380 61.200 ;
        RECT 115.650 60.140 116.020 60.220 ;
        RECT 115.020 59.910 116.020 60.140 ;
        RECT 116.160 60.130 116.430 65.110 ;
        RECT 115.650 59.840 116.020 59.910 ;
        RECT 105.230 56.325 109.250 59.610 ;
        RECT 127.420 58.050 128.590 65.720 ;
        RECT 129.860 65.460 130.260 65.550 ;
        RECT 129.260 65.230 130.260 65.460 ;
        RECT 105.230 56.070 125.505 56.325 ;
        RECT 127.420 56.070 128.320 58.050 ;
        RECT 128.860 57.380 129.110 65.220 ;
        RECT 129.860 65.150 130.260 65.230 ;
        RECT 129.250 63.170 129.650 63.260 ;
        RECT 129.250 62.940 130.260 63.170 ;
        RECT 129.250 62.860 129.650 62.940 ;
        RECT 129.870 60.880 130.270 60.970 ;
        RECT 129.260 60.650 130.270 60.880 ;
        RECT 129.870 60.570 130.270 60.650 ;
        RECT 129.250 58.590 129.650 58.680 ;
        RECT 129.250 58.360 130.260 58.590 ;
        RECT 129.250 58.280 129.650 58.360 ;
        RECT 130.410 57.380 130.660 65.220 ;
        RECT 143.300 64.880 147.320 65.745 ;
        RECT 139.300 64.630 139.810 64.710 ;
        RECT 138.135 64.400 139.810 64.630 ;
        RECT 135.595 62.155 136.645 63.145 ;
        RECT 135.625 58.375 136.615 62.155 ;
        RECT 137.680 61.200 137.960 64.400 ;
        RECT 139.300 64.320 139.810 64.400 ;
        RECT 138.150 63.990 138.660 64.070 ;
        RECT 138.135 63.760 139.805 63.990 ;
        RECT 138.150 63.680 138.660 63.760 ;
        RECT 139.300 63.350 139.810 63.430 ;
        RECT 138.135 63.120 139.810 63.350 ;
        RECT 139.300 63.040 139.810 63.120 ;
        RECT 138.150 62.710 138.660 62.790 ;
        RECT 138.135 62.480 139.805 62.710 ;
        RECT 138.150 62.400 138.660 62.480 ;
        RECT 139.990 61.200 140.270 64.400 ;
        RECT 140.500 62.200 147.320 64.880 ;
        RECT 137.680 60.920 140.270 61.200 ;
        RECT 137.730 59.540 138.010 60.920 ;
        RECT 135.625 57.385 140.385 58.375 ;
        RECT 128.860 56.790 130.660 57.380 ;
        RECT 105.230 55.170 128.320 56.070 ;
        RECT 129.860 56.690 130.660 56.790 ;
        RECT 137.480 57.330 140.380 57.385 ;
        RECT 129.860 55.670 134.190 56.690 ;
        RECT 105.230 54.915 125.505 55.170 ;
        RECT 105.230 32.190 109.250 54.915 ;
        RECT 126.270 52.860 127.010 53.540 ;
        RECT 116.500 50.860 117.710 50.870 ;
        RECT 118.740 50.860 119.425 52.790 ;
        RECT 120.600 52.020 125.965 52.030 ;
        RECT 126.300 52.020 126.980 52.860 ;
        RECT 120.340 51.600 128.630 52.020 ;
        RECT 116.500 49.630 120.150 50.860 ;
        RECT 120.340 50.030 120.630 51.600 ;
        RECT 120.790 50.590 121.200 50.680 ;
        RECT 120.790 50.360 121.790 50.590 ;
        RECT 120.790 50.310 121.200 50.360 ;
        RECT 121.380 50.150 121.790 50.210 ;
        RECT 120.790 49.920 121.790 50.150 ;
        RECT 121.940 50.030 122.230 51.600 ;
        RECT 125.680 49.980 125.970 51.600 ;
        RECT 127.550 50.640 128.170 50.720 ;
        RECT 126.165 50.410 128.170 50.640 ;
        RECT 127.550 50.340 128.170 50.410 ;
        RECT 126.180 50.000 126.800 50.080 ;
        RECT 121.380 49.840 121.790 49.920 ;
        RECT 126.165 49.770 128.165 50.000 ;
        RECT 128.340 49.980 128.630 51.600 ;
        RECT 129.525 50.920 130.420 52.905 ;
        RECT 126.180 49.700 126.800 49.770 ;
        RECT 116.500 46.180 119.280 49.630 ;
        RECT 128.850 49.510 131.950 50.920 ;
        RECT 123.700 47.980 124.385 49.155 ;
        RECT 120.600 47.970 128.640 47.980 ;
        RECT 120.370 47.540 128.640 47.970 ;
        RECT 120.370 47.520 125.970 47.540 ;
        RECT 116.500 44.470 120.130 46.180 ;
        RECT 120.370 45.360 120.650 47.520 ;
        RECT 121.820 45.910 122.250 45.990 ;
        RECT 120.790 45.680 122.290 45.910 ;
        RECT 121.820 45.590 122.250 45.680 ;
        RECT 120.840 45.430 121.270 45.510 ;
        RECT 120.790 45.200 122.290 45.430 ;
        RECT 120.840 45.110 121.270 45.200 ;
        RECT 121.820 44.950 122.250 45.040 ;
        RECT 120.790 44.720 122.290 44.950 ;
        RECT 122.430 44.880 122.720 47.520 ;
        RECT 121.820 44.640 122.250 44.720 ;
        RECT 125.680 44.590 125.960 47.520 ;
        RECT 127.600 46.500 128.160 46.590 ;
        RECT 126.165 46.270 128.165 46.500 ;
        RECT 127.600 46.190 128.160 46.270 ;
        RECT 126.180 45.860 126.740 45.940 ;
        RECT 126.165 45.630 128.165 45.860 ;
        RECT 126.180 45.540 126.740 45.630 ;
        RECT 127.600 45.220 128.160 45.310 ;
        RECT 126.165 44.990 128.165 45.220 ;
        RECT 127.600 44.910 128.160 44.990 ;
        RECT 126.180 44.580 126.740 44.660 ;
        RECT 128.350 44.590 128.630 47.540 ;
        RECT 130.030 46.770 131.950 49.510 ;
        RECT 116.500 39.340 117.710 44.470 ;
        RECT 126.165 44.350 128.165 44.580 ;
        RECT 126.180 44.260 126.740 44.350 ;
        RECT 128.840 44.080 131.950 46.770 ;
        RECT 118.730 42.280 121.120 42.960 ;
        RECT 123.625 42.280 124.500 43.780 ;
        RECT 118.730 42.260 126.085 42.280 ;
        RECT 118.730 41.590 129.620 42.260 ;
        RECT 118.730 41.570 126.085 41.590 ;
        RECT 118.730 41.415 121.120 41.570 ;
        RECT 116.500 37.150 118.690 39.340 ;
        RECT 118.930 37.580 119.200 41.415 ;
        RECT 119.410 39.080 119.920 39.180 ;
        RECT 119.350 38.850 122.350 39.080 ;
        RECT 119.410 38.750 119.920 38.850 ;
        RECT 121.790 38.600 122.300 38.700 ;
        RECT 119.350 38.370 122.350 38.600 ;
        RECT 121.790 38.270 122.300 38.370 ;
        RECT 119.420 38.120 119.930 38.220 ;
        RECT 119.350 37.890 122.350 38.120 ;
        RECT 122.500 38.060 122.770 41.570 ;
        RECT 119.420 37.790 119.930 37.890 ;
        RECT 121.790 37.640 122.300 37.740 ;
        RECT 119.350 37.410 122.350 37.640 ;
        RECT 121.790 37.310 122.300 37.410 ;
        RECT 116.500 32.190 118.160 37.150 ;
        RECT 125.680 36.420 125.960 41.570 ;
        RECT 128.560 40.280 129.160 40.360 ;
        RECT 126.165 40.050 129.165 40.280 ;
        RECT 128.560 39.960 129.160 40.050 ;
        RECT 126.200 39.640 126.800 39.720 ;
        RECT 126.165 39.410 129.165 39.640 ;
        RECT 126.200 39.320 126.800 39.410 ;
        RECT 128.560 39.000 129.160 39.090 ;
        RECT 126.165 38.770 129.165 39.000 ;
        RECT 128.560 38.690 129.160 38.770 ;
        RECT 126.200 38.360 126.800 38.450 ;
        RECT 126.165 38.130 129.165 38.360 ;
        RECT 126.200 38.050 126.800 38.130 ;
        RECT 128.560 37.720 129.160 37.800 ;
        RECT 126.165 37.490 129.165 37.720 ;
        RECT 128.560 37.400 129.160 37.490 ;
        RECT 126.200 37.080 126.800 37.170 ;
        RECT 126.165 36.850 129.165 37.080 ;
        RECT 126.200 36.770 126.800 36.850 ;
        RECT 128.560 36.440 129.160 36.530 ;
        RECT 126.165 36.210 129.165 36.440 ;
        RECT 129.340 36.420 129.620 41.590 ;
        RECT 130.800 40.480 131.950 44.080 ;
        RECT 128.560 36.130 129.160 36.210 ;
        RECT 129.870 35.960 131.950 40.480 ;
        RECT 133.170 39.295 134.190 55.670 ;
        RECT 105.230 30.530 118.160 32.190 ;
        RECT 123.180 31.985 124.260 34.260 ;
        RECT 130.140 32.015 131.950 35.960 ;
        RECT 133.035 34.305 134.245 39.295 ;
        RECT 137.480 36.320 137.740 57.330 ;
        RECT 137.950 56.070 138.520 56.170 ;
        RECT 137.935 55.840 139.935 56.070 ;
        RECT 137.950 55.750 138.520 55.840 ;
        RECT 139.370 52.780 139.940 52.880 ;
        RECT 137.935 52.550 139.940 52.780 ;
        RECT 139.370 52.460 139.940 52.550 ;
        RECT 137.950 49.490 138.520 49.600 ;
        RECT 137.935 49.260 139.935 49.490 ;
        RECT 137.950 49.180 138.520 49.260 ;
        RECT 139.380 46.200 139.950 46.300 ;
        RECT 137.935 45.970 139.950 46.200 ;
        RECT 139.380 45.880 139.950 45.970 ;
        RECT 137.950 42.910 138.520 43.010 ;
        RECT 137.935 42.680 139.935 42.910 ;
        RECT 137.950 42.590 138.520 42.680 ;
        RECT 139.380 39.620 139.950 39.720 ;
        RECT 137.935 39.390 139.950 39.620 ;
        RECT 139.380 39.300 139.950 39.390 ;
        RECT 137.950 36.330 138.520 36.420 ;
        RECT 137.935 36.100 139.935 36.330 ;
        RECT 140.120 36.320 140.380 57.330 ;
        RECT 143.300 56.330 147.320 62.200 ;
        RECT 137.950 36.000 138.520 36.100 ;
        RECT 140.660 35.800 147.320 56.330 ;
        RECT 143.300 34.295 147.320 35.800 ;
        RECT 139.255 33.480 147.320 34.295 ;
        RECT 143.300 32.015 147.320 33.480 ;
        RECT 105.230 29.730 109.250 30.530 ;
        RECT 122.895 25.485 124.305 31.985 ;
        RECT 130.140 30.205 147.320 32.015 ;
        RECT 143.300 29.730 147.320 30.205 ;
      LAYER via ;
        RECT 125.960 142.690 127.460 144.190 ;
        RECT 96.530 135.110 98.030 136.610 ;
        RECT 136.240 132.350 137.140 133.250 ;
        RECT 118.190 118.660 118.750 119.220 ;
        RECT 123.530 123.620 124.020 123.910 ;
        RECT 121.090 123.160 121.580 123.450 ;
        RECT 123.530 122.680 124.020 122.970 ;
        RECT 121.090 122.200 121.580 122.490 ;
        RECT 123.530 121.720 124.020 122.010 ;
        RECT 121.090 121.240 121.580 121.530 ;
        RECT 123.530 120.760 124.020 121.050 ;
        RECT 121.090 120.280 121.580 120.570 ;
        RECT 122.715 118.710 123.285 119.280 ;
        RECT 126.450 120.150 128.015 121.715 ;
        RECT 130.270 123.580 130.750 123.860 ;
        RECT 132.670 123.010 133.150 123.290 ;
        RECT 130.250 122.360 130.730 122.640 ;
        RECT 132.670 121.720 133.150 122.000 ;
        RECT 130.250 121.090 130.730 121.370 ;
        RECT 132.670 120.450 133.150 120.730 ;
        RECT 130.250 119.800 130.730 120.080 ;
        RECT 132.670 119.170 133.150 119.450 ;
        RECT 130.220 117.450 130.800 118.030 ;
        RECT 140.330 114.495 140.920 115.085 ;
        RECT 115.240 108.450 115.870 108.770 ;
        RECT 112.010 105.180 112.640 105.500 ;
        RECT 115.240 101.870 115.870 102.190 ;
        RECT 112.010 98.570 112.640 98.890 ;
        RECT 111.960 96.510 112.710 97.260 ;
        RECT 115.240 92.820 115.950 93.190 ;
        RECT 112.060 89.530 112.770 89.900 ;
        RECT 115.240 86.250 115.950 86.620 ;
        RECT 112.060 82.960 112.770 83.330 ;
        RECT 123.850 104.820 124.260 105.110 ;
        RECT 122.870 103.830 123.280 104.120 ;
        RECT 123.850 102.840 124.260 103.130 ;
        RECT 122.870 101.850 123.280 102.140 ;
        RECT 123.850 100.860 124.260 101.150 ;
        RECT 122.870 99.870 123.280 100.160 ;
        RECT 123.850 98.880 124.260 99.170 ;
        RECT 122.870 97.900 123.280 98.190 ;
        RECT 123.850 96.900 124.260 97.190 ;
        RECT 122.870 95.920 123.280 96.210 ;
        RECT 123.850 94.920 124.260 95.210 ;
        RECT 122.870 93.930 123.280 94.220 ;
        RECT 123.850 92.940 124.260 93.230 ;
        RECT 122.870 91.960 123.280 92.250 ;
        RECT 123.850 90.960 124.260 91.250 ;
        RECT 122.870 89.970 123.280 90.260 ;
        RECT 123.850 88.980 124.260 89.270 ;
        RECT 122.870 87.990 123.280 88.280 ;
        RECT 123.850 87.000 124.260 87.290 ;
        RECT 131.640 104.820 132.170 105.110 ;
        RECT 130.680 103.830 131.210 104.120 ;
        RECT 131.640 102.840 132.170 103.130 ;
        RECT 130.680 101.860 131.210 102.150 ;
        RECT 131.640 100.860 132.170 101.150 ;
        RECT 130.680 99.880 131.210 100.170 ;
        RECT 131.640 98.890 132.170 99.180 ;
        RECT 130.680 97.890 131.210 98.180 ;
        RECT 131.640 96.910 132.170 97.200 ;
        RECT 130.680 95.910 131.210 96.200 ;
        RECT 131.640 94.920 132.170 95.210 ;
        RECT 130.680 93.940 131.210 94.230 ;
        RECT 131.640 92.940 132.170 93.230 ;
        RECT 130.680 91.960 131.210 92.250 ;
        RECT 131.640 90.970 132.170 91.260 ;
        RECT 130.680 89.980 131.210 90.270 ;
        RECT 131.640 88.980 132.170 89.270 ;
        RECT 130.680 88.000 131.210 88.290 ;
        RECT 131.640 87.000 132.170 87.290 ;
        RECT 140.330 104.105 140.920 104.695 ;
        RECT 121.135 82.525 121.825 83.215 ;
        RECT 112.020 80.530 112.820 81.330 ;
        RECT 127.710 81.175 128.380 81.845 ;
        RECT 115.040 79.060 115.400 79.420 ;
        RECT 115.590 77.730 116.000 78.010 ;
        RECT 115.000 76.430 115.410 76.710 ;
        RECT 115.590 75.140 116.000 75.420 ;
        RECT 114.990 73.860 115.400 74.140 ;
        RECT 129.670 78.230 130.330 78.530 ;
        RECT 128.180 77.590 128.840 77.890 ;
        RECT 129.670 76.950 130.330 77.250 ;
        RECT 128.180 76.300 128.840 76.600 ;
        RECT 129.670 75.670 130.330 75.970 ;
        RECT 128.170 75.030 128.830 75.330 ;
        RECT 129.670 74.390 130.330 74.690 ;
        RECT 128.180 73.750 128.840 74.050 ;
        RECT 115.650 72.255 116.040 72.645 ;
        RECT 118.525 71.980 119.255 72.710 ;
        RECT 139.890 101.450 140.490 101.740 ;
        RECT 138.490 98.160 139.090 98.450 ;
        RECT 139.890 94.870 140.490 95.160 ;
        RECT 138.490 91.590 139.090 91.880 ;
        RECT 139.890 88.300 140.490 88.590 ;
        RECT 138.490 85.000 139.090 85.290 ;
        RECT 139.890 81.710 140.490 82.000 ;
        RECT 138.490 78.420 139.090 78.710 ;
        RECT 139.890 75.140 140.490 75.430 ;
        RECT 138.490 71.840 139.090 72.130 ;
        RECT 111.370 68.350 112.270 69.250 ;
        RECT 123.260 68.140 124.800 69.680 ;
        RECT 139.850 68.200 140.550 68.900 ;
        RECT 112.675 65.775 113.405 66.505 ;
        RECT 140.780 65.800 141.360 66.380 ;
        RECT 120.355 65.110 120.865 65.620 ;
        RECT 115.020 63.760 115.390 64.040 ;
        RECT 115.650 62.470 116.020 62.750 ;
        RECT 115.010 61.180 115.380 61.460 ;
        RECT 115.650 59.890 116.020 60.170 ;
        RECT 129.860 65.200 130.260 65.500 ;
        RECT 129.250 62.910 129.650 63.210 ;
        RECT 129.870 60.620 130.270 60.920 ;
        RECT 129.250 58.330 129.650 58.630 ;
        RECT 135.625 62.155 136.615 63.145 ;
        RECT 139.300 64.370 139.810 64.660 ;
        RECT 138.150 63.730 138.660 64.020 ;
        RECT 139.300 63.090 139.810 63.380 ;
        RECT 138.150 62.450 138.660 62.740 ;
        RECT 137.730 59.570 138.010 59.850 ;
        RECT 126.300 52.860 126.980 53.540 ;
        RECT 118.825 52.195 119.335 52.705 ;
        RECT 129.605 52.095 130.335 52.825 ;
        RECT 121.380 49.890 121.790 50.160 ;
        RECT 127.550 50.390 128.170 50.670 ;
        RECT 126.180 49.750 126.800 50.030 ;
        RECT 123.775 48.550 124.305 49.080 ;
        RECT 118.130 46.720 118.650 47.240 ;
        RECT 130.435 47.665 131.085 48.315 ;
        RECT 121.820 45.640 122.250 45.940 ;
        RECT 120.840 45.160 121.270 45.460 ;
        RECT 121.820 44.690 122.250 44.990 ;
        RECT 127.600 46.240 128.160 46.540 ;
        RECT 126.180 45.590 126.740 45.890 ;
        RECT 127.600 44.960 128.160 45.260 ;
        RECT 126.180 44.310 126.740 44.610 ;
        RECT 123.735 43.020 124.385 43.670 ;
        RECT 118.935 41.625 120.065 42.755 ;
        RECT 119.410 38.800 119.920 39.130 ;
        RECT 121.790 38.320 122.300 38.650 ;
        RECT 119.420 37.840 119.930 38.170 ;
        RECT 121.790 37.360 122.300 37.690 ;
        RECT 128.560 40.010 129.160 40.310 ;
        RECT 126.200 39.370 126.800 39.670 ;
        RECT 128.560 38.740 129.160 39.040 ;
        RECT 126.200 38.100 126.800 38.400 ;
        RECT 128.560 37.450 129.160 37.750 ;
        RECT 126.200 36.820 126.800 37.120 ;
        RECT 128.560 36.180 129.160 36.480 ;
        RECT 117.145 35.320 117.775 35.950 ;
        RECT 130.555 34.340 131.325 35.110 ;
        RECT 123.405 33.405 124.035 34.035 ;
        RECT 137.950 55.800 138.520 56.120 ;
        RECT 139.370 52.510 139.940 52.830 ;
        RECT 137.950 49.230 138.520 49.550 ;
        RECT 139.380 45.930 139.950 46.250 ;
        RECT 137.950 42.640 138.520 42.960 ;
        RECT 139.380 39.350 139.950 39.670 ;
        RECT 137.950 36.050 138.520 36.370 ;
        RECT 133.190 34.460 134.090 35.360 ;
        RECT 139.340 33.570 139.980 34.210 ;
        RECT 123.150 25.740 124.050 26.640 ;
      LAYER met2 ;
        RECT 87.225 144.190 88.675 144.210 ;
        RECT 87.200 142.690 127.490 144.190 ;
        RECT 87.225 142.670 88.675 142.690 ;
        RECT 86.935 136.610 88.385 136.630 ;
        RECT 86.910 135.110 98.060 136.610 ;
        RECT 86.935 135.090 88.385 135.110 ;
        RECT 136.210 132.350 157.310 133.250 ;
        RECT 123.480 123.620 124.070 123.910 ;
        RECT 121.040 123.160 121.630 123.450 ;
        RECT 121.070 122.490 121.630 123.160 ;
        RECT 123.500 122.970 124.070 123.620 ;
        RECT 123.480 122.680 124.070 122.970 ;
        RECT 121.040 122.200 121.630 122.490 ;
        RECT 121.070 121.530 121.630 122.200 ;
        RECT 123.500 122.010 124.070 122.680 ;
        RECT 130.220 122.640 130.800 123.870 ;
        RECT 132.640 123.290 133.180 123.350 ;
        RECT 132.620 123.010 133.200 123.290 ;
        RECT 130.200 122.360 130.800 122.640 ;
        RECT 123.480 121.720 124.070 122.010 ;
        RECT 121.040 121.240 121.630 121.530 ;
        RECT 121.070 120.570 121.630 121.240 ;
        RECT 123.500 121.050 124.070 121.720 ;
        RECT 123.480 120.760 124.070 121.050 ;
        RECT 121.040 120.280 121.630 120.570 ;
        RECT 118.190 119.220 118.750 119.250 ;
        RECT 121.070 119.220 121.630 120.280 ;
        RECT 123.500 119.280 124.070 120.760 ;
        RECT 126.420 120.150 128.045 121.715 ;
        RECT 130.220 121.370 130.800 122.360 ;
        RECT 132.640 122.000 133.180 123.010 ;
        RECT 132.620 121.720 133.200 122.000 ;
        RECT 130.200 121.090 130.800 121.370 ;
        RECT 118.190 118.660 121.630 119.220 ;
        RECT 122.685 118.710 124.070 119.280 ;
        RECT 118.190 118.630 118.750 118.660 ;
        RECT 126.450 112.505 128.015 120.150 ;
        RECT 130.220 120.080 130.800 121.090 ;
        RECT 132.640 120.730 133.180 121.720 ;
        RECT 132.620 120.450 133.200 120.730 ;
        RECT 130.200 119.800 130.800 120.080 ;
        RECT 130.220 117.420 130.800 119.800 ;
        RECT 132.640 119.450 133.180 120.450 ;
        RECT 132.620 119.170 133.200 119.450 ;
        RECT 132.640 117.990 133.180 119.170 ;
        RECT 132.640 117.450 135.710 117.990 ;
        RECT 156.410 116.055 157.310 132.350 ;
        RECT 156.390 115.205 157.330 116.055 ;
        RECT 156.410 115.180 157.310 115.205 ;
        RECT 115.190 110.300 124.405 111.010 ;
        RECT 126.450 110.940 132.660 112.505 ;
        RECT 115.190 108.770 115.900 110.300 ;
        RECT 115.190 108.450 115.920 108.770 ;
        RECT 111.960 96.480 112.710 105.570 ;
        RECT 115.190 102.190 115.900 108.450 ;
        RECT 123.695 107.925 124.405 110.300 ;
        RECT 131.095 108.790 132.660 110.940 ;
        RECT 130.640 107.925 131.230 107.950 ;
        RECT 123.695 107.215 131.230 107.925 ;
        RECT 123.810 105.110 124.320 105.160 ;
        RECT 123.800 104.820 124.320 105.110 ;
        RECT 115.190 101.870 115.920 102.190 ;
        RECT 115.190 101.470 115.900 101.870 ;
        RECT 115.170 93.190 115.970 93.300 ;
        RECT 115.170 92.820 116.000 93.190 ;
        RECT 112.020 89.900 112.820 90.010 ;
        RECT 112.010 89.530 112.820 89.900 ;
        RECT 112.020 83.330 112.820 89.530 ;
        RECT 112.010 82.960 112.820 83.330 ;
        RECT 112.020 80.500 112.820 82.960 ;
        RECT 115.170 86.620 115.970 92.820 ;
        RECT 115.170 86.250 116.000 86.620 ;
        RECT 115.170 81.520 115.970 86.250 ;
        RECT 122.760 83.380 123.420 104.320 ;
        RECT 123.810 103.130 124.320 104.820 ;
        RECT 123.800 102.840 124.320 103.130 ;
        RECT 123.810 101.150 124.320 102.840 ;
        RECT 123.800 100.860 124.320 101.150 ;
        RECT 123.810 99.170 124.320 100.860 ;
        RECT 123.800 98.880 124.320 99.170 ;
        RECT 123.810 97.190 124.320 98.880 ;
        RECT 123.800 96.900 124.320 97.190 ;
        RECT 123.810 95.210 124.320 96.900 ;
        RECT 123.800 94.920 124.320 95.210 ;
        RECT 123.810 93.230 124.320 94.920 ;
        RECT 123.800 92.940 124.320 93.230 ;
        RECT 123.810 91.250 124.320 92.940 ;
        RECT 123.800 90.960 124.320 91.250 ;
        RECT 123.810 89.270 124.320 90.960 ;
        RECT 123.800 88.980 124.320 89.270 ;
        RECT 123.810 87.290 124.320 88.980 ;
        RECT 123.800 87.000 124.320 87.290 ;
        RECT 122.760 83.215 123.450 83.380 ;
        RECT 121.105 82.525 123.450 83.215 ;
        RECT 122.760 82.320 123.450 82.525 ;
        RECT 122.760 81.520 123.420 82.320 ;
        RECT 115.170 80.720 123.490 81.520 ;
        RECT 123.810 80.315 124.320 87.000 ;
        RECT 127.710 81.845 128.380 107.215 ;
        RECT 130.640 104.120 131.230 107.215 ;
        RECT 131.540 105.110 132.210 108.790 ;
        RECT 135.625 105.735 136.615 105.935 ;
        RECT 140.330 105.735 140.920 115.115 ;
        RECT 135.625 105.145 140.920 105.735 ;
        RECT 131.540 104.820 132.220 105.110 ;
        RECT 130.630 103.830 131.260 104.120 ;
        RECT 130.640 102.150 131.230 103.830 ;
        RECT 131.540 103.130 132.210 104.820 ;
        RECT 131.540 102.840 132.220 103.130 ;
        RECT 130.630 101.860 131.260 102.150 ;
        RECT 130.640 100.170 131.230 101.860 ;
        RECT 131.540 101.150 132.210 102.840 ;
        RECT 131.540 100.860 132.220 101.150 ;
        RECT 130.630 99.880 131.260 100.170 ;
        RECT 130.640 98.180 131.230 99.880 ;
        RECT 131.540 99.180 132.210 100.860 ;
        RECT 131.540 98.890 132.220 99.180 ;
        RECT 130.630 97.890 131.260 98.180 ;
        RECT 130.640 96.200 131.230 97.890 ;
        RECT 131.540 97.200 132.210 98.890 ;
        RECT 131.540 96.910 132.220 97.200 ;
        RECT 130.630 95.910 131.260 96.200 ;
        RECT 130.640 94.230 131.230 95.910 ;
        RECT 131.540 95.210 132.210 96.910 ;
        RECT 131.540 94.920 132.220 95.210 ;
        RECT 130.630 93.940 131.260 94.230 ;
        RECT 130.640 92.250 131.230 93.940 ;
        RECT 131.540 93.230 132.210 94.920 ;
        RECT 131.540 92.940 132.220 93.230 ;
        RECT 130.630 91.960 131.260 92.250 ;
        RECT 130.640 90.270 131.230 91.960 ;
        RECT 131.540 91.260 132.210 92.940 ;
        RECT 131.540 90.970 132.220 91.260 ;
        RECT 130.630 89.980 131.260 90.270 ;
        RECT 130.640 88.290 131.230 89.980 ;
        RECT 131.540 89.270 132.210 90.970 ;
        RECT 131.540 88.980 132.220 89.270 ;
        RECT 130.630 88.000 131.260 88.290 ;
        RECT 130.640 87.880 131.230 88.000 ;
        RECT 131.540 87.290 132.210 88.980 ;
        RECT 131.540 87.000 132.220 87.290 ;
        RECT 131.540 86.965 132.210 87.000 ;
        RECT 127.680 81.175 128.410 81.845 ;
        RECT 123.810 79.805 134.105 80.315 ;
        RECT 115.010 79.060 115.430 79.420 ;
        RECT 115.040 76.710 115.400 79.060 ;
        RECT 115.540 77.730 116.050 78.010 ;
        RECT 128.190 77.890 128.920 77.940 ;
        RECT 114.950 76.430 115.460 76.710 ;
        RECT 115.040 74.140 115.400 76.430 ;
        RECT 115.650 75.420 116.040 77.730 ;
        RECT 128.130 77.590 128.920 77.890 ;
        RECT 128.190 76.600 128.920 77.590 ;
        RECT 128.130 76.300 128.920 76.600 ;
        RECT 115.540 75.140 116.050 75.420 ;
        RECT 128.190 75.330 128.920 76.300 ;
        RECT 114.940 73.860 115.450 74.140 ;
        RECT 115.040 73.850 115.400 73.860 ;
        RECT 115.650 72.225 116.040 75.140 ;
        RECT 128.120 75.030 128.920 75.330 ;
        RECT 128.190 74.050 128.920 75.030 ;
        RECT 129.610 74.240 130.380 79.805 ;
        RECT 128.130 73.750 128.920 74.050 ;
        RECT 128.190 72.710 128.920 73.750 ;
        RECT 118.495 71.980 128.920 72.710 ;
        RECT 90.170 68.350 112.300 69.250 ;
        RECT 90.170 64.285 91.070 68.350 ;
        RECT 112.645 66.370 114.115 66.505 ;
        RECT 112.645 65.910 115.430 66.370 ;
        RECT 112.645 65.775 114.115 65.910 ;
        RECT 90.150 63.435 91.090 64.285 ;
        RECT 114.970 64.040 115.430 65.910 ;
        RECT 120.210 64.960 121.015 71.980 ;
        RECT 133.595 71.545 134.105 79.805 ;
        RECT 135.625 73.460 136.615 105.145 ;
        RECT 140.330 104.695 140.920 105.145 ;
        RECT 140.300 104.105 140.950 104.695 ;
        RECT 139.850 101.740 140.550 101.800 ;
        RECT 139.840 101.450 140.550 101.740 ;
        RECT 138.450 98.450 139.150 98.550 ;
        RECT 138.440 98.160 139.150 98.450 ;
        RECT 138.450 91.880 139.150 98.160 ;
        RECT 139.850 95.160 140.550 101.450 ;
        RECT 139.840 94.870 140.550 95.160 ;
        RECT 138.440 91.590 139.150 91.880 ;
        RECT 138.450 85.290 139.150 91.590 ;
        RECT 139.850 88.590 140.550 94.870 ;
        RECT 139.840 88.300 140.550 88.590 ;
        RECT 138.440 85.000 139.150 85.290 ;
        RECT 138.450 78.710 139.150 85.000 ;
        RECT 139.850 82.000 140.550 88.300 ;
        RECT 139.840 81.710 140.550 82.000 ;
        RECT 138.440 78.420 139.150 78.710 ;
        RECT 138.450 72.130 139.150 78.420 ;
        RECT 139.850 75.430 140.550 81.710 ;
        RECT 139.840 75.140 140.550 75.430 ;
        RECT 138.440 71.840 139.150 72.130 ;
        RECT 133.585 70.975 134.105 71.545 ;
        RECT 133.585 70.040 134.095 70.975 ;
        RECT 138.450 70.040 139.150 71.840 ;
        RECT 123.260 69.680 124.800 69.710 ;
        RECT 123.260 69.650 129.670 69.680 ;
        RECT 133.580 69.650 139.150 70.040 ;
        RECT 123.260 68.205 139.150 69.650 ;
        RECT 123.260 68.140 129.670 68.205 ;
        RECT 133.580 68.200 139.150 68.205 ;
        RECT 139.850 68.170 140.550 75.140 ;
        RECT 123.260 68.110 124.800 68.140 ;
        RECT 114.970 63.760 115.440 64.040 ;
        RECT 90.170 63.410 91.070 63.435 ;
        RECT 114.970 61.460 115.430 63.760 ;
        RECT 129.190 63.210 129.650 68.140 ;
        RECT 129.860 66.410 138.700 66.860 ;
        RECT 129.860 65.500 130.310 66.410 ;
        RECT 129.810 65.200 130.310 65.500 ;
        RECT 129.190 62.910 129.700 63.210 ;
        RECT 115.620 62.750 116.070 62.780 ;
        RECT 115.600 62.470 116.070 62.750 ;
        RECT 114.960 61.180 115.430 61.460 ;
        RECT 114.970 61.150 115.430 61.180 ;
        RECT 115.620 60.170 116.070 62.470 ;
        RECT 115.600 59.890 116.070 60.170 ;
        RECT 115.620 58.110 116.070 59.890 ;
        RECT 129.190 58.630 129.650 62.910 ;
        RECT 129.860 60.920 130.310 65.200 ;
        RECT 135.625 64.590 136.615 64.615 ;
        RECT 129.820 60.620 130.320 60.920 ;
        RECT 133.045 60.695 134.175 64.580 ;
        RECT 135.605 63.650 136.635 64.590 ;
        RECT 138.090 64.020 138.700 66.410 ;
        RECT 139.280 65.800 141.390 66.380 ;
        RECT 139.280 64.660 139.860 65.800 ;
        RECT 139.250 64.370 139.860 64.660 ;
        RECT 138.090 63.730 138.710 64.020 ;
        RECT 135.625 62.125 136.615 63.650 ;
        RECT 138.090 62.740 138.700 63.730 ;
        RECT 139.280 63.380 139.860 64.370 ;
        RECT 139.250 63.090 139.860 63.380 ;
        RECT 139.280 63.050 139.860 63.090 ;
        RECT 138.090 62.450 138.710 62.740 ;
        RECT 138.090 62.430 138.700 62.450 ;
        RECT 129.860 60.520 130.310 60.620 ;
        RECT 133.300 60.020 133.925 60.695 ;
        RECT 133.300 59.395 138.185 60.020 ;
        RECT 129.190 58.330 129.700 58.630 ;
        RECT 129.190 58.290 129.650 58.330 ;
        RECT 115.620 56.845 126.980 58.110 ;
        RECT 116.000 56.820 126.980 56.845 ;
        RECT 126.290 54.760 126.970 56.820 ;
        RECT 126.290 54.170 131.830 54.760 ;
        RECT 126.290 54.155 134.430 54.170 ;
        RECT 126.290 54.080 136.425 54.155 ;
        RECT 126.300 52.830 126.980 54.080 ;
        RECT 131.150 53.490 136.425 54.080 ;
        RECT 133.885 53.465 136.425 53.490 ;
        RECT 118.795 52.195 121.250 52.705 ;
        RECT 120.740 50.360 121.250 52.195 ;
        RECT 127.500 52.095 130.365 52.825 ;
        RECT 127.500 50.390 128.230 52.095 ;
        RECT 121.330 49.080 121.860 50.160 ;
        RECT 126.120 49.080 126.850 50.040 ;
        RECT 121.330 48.550 126.850 49.080 ;
        RECT 127.560 47.665 131.115 48.315 ;
        RECT 118.100 46.720 121.310 47.240 ;
        RECT 120.790 45.460 121.310 46.720 ;
        RECT 127.560 46.540 128.210 47.665 ;
        RECT 127.550 46.240 128.210 46.540 ;
        RECT 121.800 45.940 122.300 45.960 ;
        RECT 121.770 45.640 122.300 45.940 ;
        RECT 120.790 45.160 121.320 45.460 ;
        RECT 120.790 45.130 121.310 45.160 ;
        RECT 121.800 44.990 122.300 45.640 ;
        RECT 121.770 44.690 122.300 44.990 ;
        RECT 121.800 43.670 122.300 44.690 ;
        RECT 126.130 45.890 126.780 45.930 ;
        RECT 126.130 45.590 126.790 45.890 ;
        RECT 126.130 44.610 126.780 45.590 ;
        RECT 127.560 45.260 128.210 46.240 ;
        RECT 127.550 44.960 128.210 45.260 ;
        RECT 127.560 44.940 128.210 44.960 ;
        RECT 126.130 44.310 126.790 44.610 ;
        RECT 123.735 43.670 124.385 43.700 ;
        RECT 126.130 43.670 126.780 44.310 ;
        RECT 121.795 43.020 126.780 43.670 ;
        RECT 121.800 43.000 122.300 43.020 ;
        RECT 123.735 42.990 124.385 43.020 ;
        RECT 113.275 42.730 120.095 42.755 ;
        RECT 113.255 41.650 120.095 42.730 ;
        RECT 113.275 41.625 120.095 41.650 ;
        RECT 119.350 35.950 119.980 39.180 ;
        RECT 117.115 35.320 119.980 35.950 ;
        RECT 121.720 34.960 122.350 38.660 ;
        RECT 126.150 34.960 126.860 39.680 ;
        RECT 121.720 34.330 126.860 34.960 ;
        RECT 128.450 35.110 129.220 40.370 ;
        RECT 128.450 34.340 131.355 35.110 ;
        RECT 123.405 33.375 124.035 34.330 ;
        RECT 123.150 21.225 124.050 26.670 ;
        RECT 133.190 21.955 134.090 35.390 ;
        RECT 135.735 34.940 136.425 53.465 ;
        RECT 137.880 34.940 138.570 56.180 ;
        RECT 139.340 52.830 139.980 52.920 ;
        RECT 139.320 52.510 139.990 52.830 ;
        RECT 139.340 46.250 139.980 52.510 ;
        RECT 139.330 45.930 140.000 46.250 ;
        RECT 139.340 39.670 139.980 45.930 ;
        RECT 139.330 39.350 140.000 39.670 ;
        RECT 135.735 34.250 138.570 34.940 ;
        RECT 139.340 34.210 139.980 39.350 ;
        RECT 139.310 33.570 140.010 34.210 ;
        RECT 123.130 20.375 124.070 21.225 ;
        RECT 133.170 21.105 134.110 21.955 ;
        RECT 133.190 21.080 134.090 21.105 ;
        RECT 123.150 20.350 124.050 20.375 ;
      LAYER via2 ;
        RECT 87.225 142.715 88.675 144.165 ;
        RECT 86.935 135.135 88.385 136.585 ;
        RECT 156.435 115.205 157.285 116.055 ;
        RECT 90.195 63.435 91.045 64.285 ;
        RECT 135.625 73.505 136.615 74.495 ;
        RECT 133.045 63.405 134.175 64.535 ;
        RECT 135.650 63.650 136.590 64.590 ;
        RECT 113.300 41.650 114.380 42.730 ;
        RECT 123.175 20.375 124.025 21.225 ;
        RECT 133.215 21.105 134.065 21.955 ;
      LAYER met3 ;
        RECT 28.925 144.190 30.415 144.215 ;
        RECT 28.920 142.690 88.700 144.190 ;
        RECT 28.925 142.665 30.415 142.690 ;
        RECT 78.465 136.610 79.955 136.635 ;
        RECT 78.460 135.110 88.410 136.610 ;
        RECT 78.465 135.085 79.955 135.110 ;
        RECT 135.600 73.480 136.640 74.520 ;
        RECT 125.525 67.285 134.175 68.415 ;
        RECT 90.170 37.245 91.070 64.310 ;
        RECT 125.525 61.675 126.655 67.285 ;
        RECT 133.045 64.560 134.175 67.285 ;
        RECT 133.020 63.380 134.200 64.560 ;
        RECT 135.625 63.625 136.615 73.480 ;
        RECT 156.410 69.220 157.310 116.080 ;
        RECT 156.415 69.195 157.305 69.220 ;
        RECT 119.555 60.545 126.655 61.675 ;
        RECT 119.555 55.775 120.685 60.545 ;
        RECT 113.275 54.645 120.685 55.775 ;
        RECT 113.275 41.625 114.405 54.645 ;
        RECT 90.145 36.355 91.095 37.245 ;
        RECT 90.170 36.350 91.070 36.355 ;
        RECT 123.150 13.975 124.050 21.250 ;
        RECT 133.190 15.435 134.090 21.980 ;
        RECT 133.165 14.545 134.115 15.435 ;
        RECT 133.190 14.540 134.090 14.545 ;
        RECT 123.125 13.085 124.075 13.975 ;
        RECT 123.150 13.080 124.050 13.085 ;
      LAYER via3 ;
        RECT 28.925 142.695 30.415 144.185 ;
        RECT 78.465 135.115 79.955 136.605 ;
        RECT 156.415 69.225 157.305 70.115 ;
        RECT 90.175 36.355 91.065 37.245 ;
        RECT 133.195 14.545 134.085 15.435 ;
        RECT 123.155 13.085 124.045 13.975 ;
      LAYER met4 ;
        RECT 3.990 224.110 4.290 224.760 ;
        RECT 7.670 224.110 7.970 224.760 ;
        RECT 11.350 224.110 11.650 224.760 ;
        RECT 15.030 224.110 15.330 224.760 ;
        RECT 18.710 224.110 19.010 224.760 ;
        RECT 22.390 224.110 22.690 224.760 ;
        RECT 26.070 224.110 26.370 224.760 ;
        RECT 29.750 224.110 30.050 224.760 ;
        RECT 33.430 224.110 33.730 224.760 ;
        RECT 37.110 224.110 37.410 224.760 ;
        RECT 40.790 224.110 41.090 224.760 ;
        RECT 44.470 224.110 44.770 224.760 ;
        RECT 48.150 224.110 48.450 224.760 ;
        RECT 51.830 224.110 52.130 224.760 ;
        RECT 55.510 224.110 55.810 224.760 ;
        RECT 59.190 224.110 59.490 224.760 ;
        RECT 62.870 224.110 63.170 224.760 ;
        RECT 66.550 224.110 66.850 224.760 ;
        RECT 70.230 224.110 70.530 224.760 ;
        RECT 73.910 224.110 74.210 224.760 ;
        RECT 77.590 224.110 77.890 224.760 ;
        RECT 81.270 224.110 81.570 224.760 ;
        RECT 84.950 224.110 85.250 224.760 ;
        RECT 88.630 224.110 88.930 224.760 ;
        RECT 3.100 222.640 89.260 224.110 ;
        RECT 49.000 220.760 50.500 222.640 ;
        RECT 2.500 142.690 30.420 144.190 ;
        RECT 50.500 135.110 79.960 136.610 ;
        RECT 90.170 1.000 91.070 37.250 ;
        RECT 123.150 6.860 124.050 13.980 ;
        RECT 133.190 10.200 134.090 15.440 ;
        RECT 133.190 9.300 135.230 10.200 ;
        RECT 112.250 5.960 124.050 6.860 ;
        RECT 112.250 1.000 113.150 5.960 ;
        RECT 134.330 1.000 135.230 9.300 ;
        RECT 156.410 1.000 157.310 70.120 ;
  END
END tt_um_alfiero88_CurrentTrigger
END LIBRARY

