VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_htfab_fprn
  CLASS BLOCK ;
  FOREIGN tt_um_htfab_fprn ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.785000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.785000 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 28.709999 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.785000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 43.064999 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 43.064999 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 43.064999 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 43.064999 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 43.064999 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 43.064999 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.785000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.785000 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.475000 ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.785000 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 129.700 1.535 131.300 216.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.275 1.535 105.875 216.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.850 1.535 80.450 216.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.425 1.535 55.025 216.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.000 1.535 29.600 216.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.575 1.535 4.175 216.550 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 140.400 1.535 142.000 216.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.975 1.535 116.575 216.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.550 1.535 91.150 216.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.125 1.535 65.725 216.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.700 1.535 40.300 216.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.275 1.535 14.875 216.550 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 8.500 203.995 11.580 212.995 ;
        RECT 16.600 209.025 30.975 212.995 ;
        RECT 16.600 203.995 22.380 209.025 ;
      LAYER pwell ;
        RECT 22.645 205.525 30.825 208.755 ;
      LAYER nwell ;
        RECT 33.925 203.995 37.005 212.995 ;
        RECT 42.025 203.995 47.805 212.995 ;
        RECT 59.350 203.995 62.430 212.995 ;
        RECT 67.450 209.025 81.825 212.995 ;
        RECT 67.450 203.995 73.230 209.025 ;
      LAYER pwell ;
        RECT 73.495 205.525 81.675 208.755 ;
      LAYER nwell ;
        RECT 84.775 203.995 87.855 212.995 ;
        RECT 92.875 203.995 98.655 212.995 ;
        RECT 110.200 203.995 113.280 212.995 ;
        RECT 118.300 209.025 132.675 212.995 ;
        RECT 118.300 203.995 124.080 209.025 ;
      LAYER pwell ;
        RECT 124.345 205.525 132.525 208.755 ;
      LAYER nwell ;
        RECT 135.625 203.995 138.705 212.995 ;
        RECT 143.725 203.995 149.505 212.995 ;
        RECT 5.800 200.025 22.380 203.995 ;
        RECT 31.225 200.025 47.805 203.995 ;
        RECT 56.650 200.025 73.230 203.995 ;
        RECT 82.075 200.025 98.655 203.995 ;
        RECT 107.500 200.025 124.080 203.995 ;
        RECT 132.925 200.025 149.505 203.995 ;
      LAYER pwell ;
        RECT 5.950 196.525 22.230 199.755 ;
        RECT 31.375 196.525 47.655 199.755 ;
        RECT 56.800 196.525 73.080 199.755 ;
        RECT 82.225 196.525 98.505 199.755 ;
        RECT 107.650 196.525 123.930 199.755 ;
        RECT 133.075 196.525 149.355 199.755 ;
        RECT 8.650 190.675 11.430 196.525 ;
        RECT 16.750 190.675 22.230 196.525 ;
        RECT 34.075 190.675 36.855 196.525 ;
        RECT 42.175 190.675 47.655 196.525 ;
        RECT 59.500 190.675 62.280 196.525 ;
        RECT 67.600 190.675 73.080 196.525 ;
        RECT 84.925 190.675 87.705 196.525 ;
        RECT 93.025 190.675 98.505 196.525 ;
        RECT 110.350 190.675 113.130 196.525 ;
        RECT 118.450 190.675 123.930 196.525 ;
        RECT 135.775 190.675 138.555 196.525 ;
        RECT 143.875 190.675 149.355 196.525 ;
      LAYER nwell ;
        RECT 8.500 181.420 11.580 190.420 ;
        RECT 16.600 181.420 22.380 190.420 ;
        RECT 33.925 181.420 37.005 190.420 ;
        RECT 42.025 181.420 47.805 190.420 ;
        RECT 59.350 181.420 62.430 190.420 ;
        RECT 67.450 181.420 73.230 190.420 ;
        RECT 84.775 181.420 87.855 190.420 ;
        RECT 92.875 181.420 98.655 190.420 ;
        RECT 110.200 181.420 113.280 190.420 ;
        RECT 118.300 181.420 124.080 190.420 ;
        RECT 135.625 181.420 138.705 190.420 ;
        RECT 143.725 181.420 149.505 190.420 ;
        RECT 5.800 177.450 22.380 181.420 ;
        RECT 31.225 177.450 47.805 181.420 ;
        RECT 56.650 177.450 73.230 181.420 ;
        RECT 82.075 177.450 98.655 181.420 ;
        RECT 107.500 177.450 124.080 181.420 ;
        RECT 132.925 177.450 149.505 181.420 ;
      LAYER pwell ;
        RECT 5.950 173.950 22.230 177.180 ;
        RECT 31.375 173.950 47.655 177.180 ;
        RECT 56.800 173.950 73.080 177.180 ;
        RECT 82.225 173.950 98.505 177.180 ;
        RECT 107.650 173.950 123.930 177.180 ;
        RECT 133.075 173.950 149.355 177.180 ;
        RECT 8.650 168.100 11.430 173.950 ;
        RECT 16.750 168.100 22.230 173.950 ;
      LAYER nwell ;
        RECT 8.500 158.845 11.580 167.845 ;
        RECT 16.600 158.845 22.380 167.845 ;
        RECT 5.800 154.875 22.380 158.845 ;
      LAYER pwell ;
        RECT 5.950 151.375 22.230 154.605 ;
        RECT 22.650 153.450 24.660 168.180 ;
        RECT 34.075 168.100 36.855 173.950 ;
        RECT 42.175 168.100 47.655 173.950 ;
      LAYER nwell ;
        RECT 33.925 158.845 37.005 167.845 ;
        RECT 42.025 158.845 47.805 167.845 ;
        RECT 31.225 154.875 47.805 158.845 ;
      LAYER pwell ;
        RECT 31.375 151.375 47.655 154.605 ;
        RECT 48.075 153.450 50.085 168.180 ;
        RECT 59.500 168.100 62.280 173.950 ;
        RECT 67.600 168.100 73.080 173.950 ;
      LAYER nwell ;
        RECT 59.350 158.845 62.430 167.845 ;
        RECT 67.450 158.845 73.230 167.845 ;
        RECT 56.650 154.875 73.230 158.845 ;
      LAYER pwell ;
        RECT 56.800 151.375 73.080 154.605 ;
        RECT 73.500 153.450 75.510 168.180 ;
        RECT 84.925 168.100 87.705 173.950 ;
        RECT 93.025 168.100 98.505 173.950 ;
      LAYER nwell ;
        RECT 84.775 158.845 87.855 167.845 ;
        RECT 92.875 158.845 98.655 167.845 ;
        RECT 82.075 154.875 98.655 158.845 ;
      LAYER pwell ;
        RECT 82.225 151.375 98.505 154.605 ;
        RECT 98.925 153.450 100.935 168.180 ;
        RECT 110.350 168.100 113.130 173.950 ;
        RECT 118.450 168.100 123.930 173.950 ;
      LAYER nwell ;
        RECT 110.200 158.845 113.280 167.845 ;
        RECT 118.300 158.845 124.080 167.845 ;
        RECT 107.500 154.875 124.080 158.845 ;
      LAYER pwell ;
        RECT 107.650 151.375 123.930 154.605 ;
        RECT 124.350 153.450 126.360 168.180 ;
        RECT 135.775 168.100 138.555 173.950 ;
        RECT 143.875 168.100 149.355 173.950 ;
      LAYER nwell ;
        RECT 135.625 158.845 138.705 167.845 ;
        RECT 143.725 158.845 149.505 167.845 ;
        RECT 132.925 154.875 149.505 158.845 ;
      LAYER pwell ;
        RECT 133.075 151.375 149.355 154.605 ;
        RECT 149.775 153.450 151.785 168.180 ;
        RECT 8.650 145.525 11.430 151.375 ;
        RECT 16.750 145.525 22.230 151.375 ;
        RECT 34.075 145.525 36.855 151.375 ;
        RECT 42.175 145.525 47.655 151.375 ;
        RECT 59.500 145.525 62.280 151.375 ;
        RECT 67.600 145.525 73.080 151.375 ;
        RECT 84.925 145.525 87.705 151.375 ;
        RECT 93.025 145.525 98.505 151.375 ;
        RECT 110.350 145.525 113.130 151.375 ;
        RECT 118.450 145.525 123.930 151.375 ;
        RECT 135.775 145.525 138.555 151.375 ;
        RECT 143.875 145.525 149.355 151.375 ;
      LAYER nwell ;
        RECT 8.500 131.995 11.580 140.995 ;
        RECT 16.600 137.025 30.975 140.995 ;
        RECT 16.600 131.995 22.380 137.025 ;
      LAYER pwell ;
        RECT 22.645 133.525 30.825 136.755 ;
      LAYER nwell ;
        RECT 33.925 131.995 37.005 140.995 ;
        RECT 42.025 131.995 47.805 140.995 ;
        RECT 59.350 131.995 62.430 140.995 ;
        RECT 67.450 137.025 81.825 140.995 ;
        RECT 67.450 131.995 73.230 137.025 ;
      LAYER pwell ;
        RECT 73.495 133.525 81.675 136.755 ;
      LAYER nwell ;
        RECT 84.775 131.995 87.855 140.995 ;
        RECT 92.875 131.995 98.655 140.995 ;
        RECT 110.200 131.995 113.280 140.995 ;
        RECT 118.300 137.025 132.675 140.995 ;
        RECT 118.300 131.995 124.080 137.025 ;
      LAYER pwell ;
        RECT 124.345 133.525 132.525 136.755 ;
      LAYER nwell ;
        RECT 135.625 131.995 138.705 140.995 ;
        RECT 143.725 131.995 149.505 140.995 ;
        RECT 5.800 128.025 22.380 131.995 ;
        RECT 31.225 128.025 47.805 131.995 ;
        RECT 56.650 128.025 73.230 131.995 ;
        RECT 82.075 128.025 98.655 131.995 ;
        RECT 107.500 128.025 124.080 131.995 ;
        RECT 132.925 128.025 149.505 131.995 ;
      LAYER pwell ;
        RECT 5.950 124.525 22.230 127.755 ;
        RECT 31.375 124.525 47.655 127.755 ;
        RECT 56.800 124.525 73.080 127.755 ;
        RECT 82.225 124.525 98.505 127.755 ;
        RECT 107.650 124.525 123.930 127.755 ;
        RECT 133.075 124.525 149.355 127.755 ;
        RECT 8.650 118.675 11.430 124.525 ;
        RECT 16.750 118.675 22.230 124.525 ;
        RECT 34.075 118.675 36.855 124.525 ;
        RECT 42.175 118.675 47.655 124.525 ;
        RECT 59.500 118.675 62.280 124.525 ;
        RECT 67.600 118.675 73.080 124.525 ;
        RECT 84.925 118.675 87.705 124.525 ;
        RECT 93.025 118.675 98.505 124.525 ;
        RECT 110.350 118.675 113.130 124.525 ;
        RECT 118.450 118.675 123.930 124.525 ;
        RECT 135.775 118.675 138.555 124.525 ;
        RECT 143.875 118.675 149.355 124.525 ;
      LAYER nwell ;
        RECT 8.500 109.420 11.580 118.420 ;
        RECT 16.600 109.420 22.380 118.420 ;
        RECT 33.925 109.420 37.005 118.420 ;
        RECT 42.025 109.420 47.805 118.420 ;
        RECT 59.350 109.420 62.430 118.420 ;
        RECT 67.450 109.420 73.230 118.420 ;
        RECT 84.775 109.420 87.855 118.420 ;
        RECT 92.875 109.420 98.655 118.420 ;
        RECT 110.200 109.420 113.280 118.420 ;
        RECT 118.300 109.420 124.080 118.420 ;
        RECT 135.625 109.420 138.705 118.420 ;
        RECT 143.725 109.420 149.505 118.420 ;
        RECT 5.800 105.450 22.380 109.420 ;
        RECT 31.225 105.450 47.805 109.420 ;
        RECT 56.650 105.450 73.230 109.420 ;
        RECT 82.075 105.450 98.655 109.420 ;
        RECT 107.500 105.450 124.080 109.420 ;
        RECT 132.925 105.450 149.505 109.420 ;
      LAYER pwell ;
        RECT 5.950 101.950 22.230 105.180 ;
        RECT 31.375 101.950 47.655 105.180 ;
        RECT 56.800 101.950 73.080 105.180 ;
        RECT 82.225 101.950 98.505 105.180 ;
        RECT 107.650 101.950 123.930 105.180 ;
        RECT 133.075 101.950 149.355 105.180 ;
        RECT 8.650 96.100 11.430 101.950 ;
        RECT 16.750 96.100 22.230 101.950 ;
      LAYER nwell ;
        RECT 8.500 86.845 11.580 95.845 ;
        RECT 16.600 86.845 22.380 95.845 ;
        RECT 5.800 82.875 22.380 86.845 ;
      LAYER pwell ;
        RECT 5.950 79.375 22.230 82.605 ;
        RECT 22.650 81.450 24.660 96.180 ;
        RECT 34.075 96.100 36.855 101.950 ;
        RECT 42.175 96.100 47.655 101.950 ;
      LAYER nwell ;
        RECT 33.925 86.845 37.005 95.845 ;
        RECT 42.025 86.845 47.805 95.845 ;
        RECT 31.225 82.875 47.805 86.845 ;
      LAYER pwell ;
        RECT 31.375 79.375 47.655 82.605 ;
        RECT 48.075 81.450 50.085 96.180 ;
        RECT 59.500 96.100 62.280 101.950 ;
        RECT 67.600 96.100 73.080 101.950 ;
      LAYER nwell ;
        RECT 59.350 86.845 62.430 95.845 ;
        RECT 67.450 86.845 73.230 95.845 ;
        RECT 56.650 82.875 73.230 86.845 ;
      LAYER pwell ;
        RECT 56.800 79.375 73.080 82.605 ;
        RECT 73.500 81.450 75.510 96.180 ;
        RECT 84.925 96.100 87.705 101.950 ;
        RECT 93.025 96.100 98.505 101.950 ;
      LAYER nwell ;
        RECT 84.775 86.845 87.855 95.845 ;
        RECT 92.875 86.845 98.655 95.845 ;
        RECT 82.075 82.875 98.655 86.845 ;
      LAYER pwell ;
        RECT 82.225 79.375 98.505 82.605 ;
        RECT 98.925 81.450 100.935 96.180 ;
        RECT 110.350 96.100 113.130 101.950 ;
        RECT 118.450 96.100 123.930 101.950 ;
      LAYER nwell ;
        RECT 110.200 86.845 113.280 95.845 ;
        RECT 118.300 86.845 124.080 95.845 ;
        RECT 107.500 82.875 124.080 86.845 ;
      LAYER pwell ;
        RECT 107.650 79.375 123.930 82.605 ;
        RECT 124.350 81.450 126.360 96.180 ;
        RECT 135.775 96.100 138.555 101.950 ;
        RECT 143.875 96.100 149.355 101.950 ;
      LAYER nwell ;
        RECT 135.625 86.845 138.705 95.845 ;
        RECT 143.725 86.845 149.505 95.845 ;
        RECT 132.925 82.875 149.505 86.845 ;
      LAYER pwell ;
        RECT 133.075 79.375 149.355 82.605 ;
        RECT 149.775 81.450 151.785 96.180 ;
        RECT 8.650 73.525 11.430 79.375 ;
        RECT 16.750 73.525 22.230 79.375 ;
        RECT 34.075 73.525 36.855 79.375 ;
        RECT 42.175 73.525 47.655 79.375 ;
        RECT 59.500 73.525 62.280 79.375 ;
        RECT 67.600 73.525 73.080 79.375 ;
        RECT 84.925 73.525 87.705 79.375 ;
        RECT 93.025 73.525 98.505 79.375 ;
        RECT 110.350 73.525 113.130 79.375 ;
        RECT 118.450 73.525 123.930 79.375 ;
        RECT 135.775 73.525 138.555 79.375 ;
        RECT 143.875 73.525 149.355 79.375 ;
      LAYER nwell ;
        RECT 8.500 59.995 11.580 68.995 ;
        RECT 16.600 65.025 30.975 68.995 ;
        RECT 16.600 59.995 22.380 65.025 ;
      LAYER pwell ;
        RECT 22.645 61.525 30.825 64.755 ;
      LAYER nwell ;
        RECT 33.925 59.995 37.005 68.995 ;
        RECT 42.025 59.995 47.805 68.995 ;
        RECT 59.350 59.995 62.430 68.995 ;
        RECT 67.450 65.025 81.825 68.995 ;
        RECT 67.450 59.995 73.230 65.025 ;
      LAYER pwell ;
        RECT 73.495 61.525 81.675 64.755 ;
      LAYER nwell ;
        RECT 84.775 59.995 87.855 68.995 ;
        RECT 92.875 59.995 98.655 68.995 ;
        RECT 110.200 59.995 113.280 68.995 ;
        RECT 118.300 65.025 132.675 68.995 ;
        RECT 118.300 59.995 124.080 65.025 ;
      LAYER pwell ;
        RECT 124.345 61.525 132.525 64.755 ;
      LAYER nwell ;
        RECT 135.625 59.995 138.705 68.995 ;
        RECT 143.725 59.995 149.505 68.995 ;
        RECT 5.800 56.025 22.380 59.995 ;
        RECT 31.225 56.025 47.805 59.995 ;
        RECT 56.650 56.025 73.230 59.995 ;
        RECT 82.075 56.025 98.655 59.995 ;
        RECT 107.500 56.025 124.080 59.995 ;
        RECT 132.925 56.025 149.505 59.995 ;
      LAYER pwell ;
        RECT 5.950 52.525 22.230 55.755 ;
        RECT 31.375 52.525 47.655 55.755 ;
        RECT 56.800 52.525 73.080 55.755 ;
        RECT 82.225 52.525 98.505 55.755 ;
        RECT 107.650 52.525 123.930 55.755 ;
        RECT 133.075 52.525 149.355 55.755 ;
        RECT 8.650 46.675 11.430 52.525 ;
        RECT 16.750 46.675 22.230 52.525 ;
        RECT 34.075 46.675 36.855 52.525 ;
        RECT 42.175 46.675 47.655 52.525 ;
        RECT 59.500 46.675 62.280 52.525 ;
        RECT 67.600 46.675 73.080 52.525 ;
        RECT 84.925 46.675 87.705 52.525 ;
        RECT 93.025 46.675 98.505 52.525 ;
        RECT 110.350 46.675 113.130 52.525 ;
        RECT 118.450 46.675 123.930 52.525 ;
        RECT 135.775 46.675 138.555 52.525 ;
        RECT 143.875 46.675 149.355 52.525 ;
      LAYER nwell ;
        RECT 8.500 37.420 11.580 46.420 ;
        RECT 16.600 37.420 22.380 46.420 ;
        RECT 33.925 37.420 37.005 46.420 ;
        RECT 42.025 37.420 47.805 46.420 ;
        RECT 59.350 37.420 62.430 46.420 ;
        RECT 67.450 37.420 73.230 46.420 ;
        RECT 84.775 37.420 87.855 46.420 ;
        RECT 92.875 37.420 98.655 46.420 ;
        RECT 110.200 37.420 113.280 46.420 ;
        RECT 118.300 37.420 124.080 46.420 ;
        RECT 135.625 37.420 138.705 46.420 ;
        RECT 143.725 37.420 149.505 46.420 ;
        RECT 5.800 33.450 22.380 37.420 ;
        RECT 31.225 33.450 47.805 37.420 ;
        RECT 56.650 33.450 73.230 37.420 ;
        RECT 82.075 33.450 98.655 37.420 ;
        RECT 107.500 33.450 124.080 37.420 ;
        RECT 132.925 33.450 149.505 37.420 ;
      LAYER pwell ;
        RECT 5.950 29.950 22.230 33.180 ;
        RECT 31.375 29.950 47.655 33.180 ;
        RECT 56.800 29.950 73.080 33.180 ;
        RECT 82.225 29.950 98.505 33.180 ;
        RECT 107.650 29.950 123.930 33.180 ;
        RECT 133.075 29.950 149.355 33.180 ;
        RECT 8.650 24.100 11.430 29.950 ;
        RECT 16.750 24.100 22.230 29.950 ;
      LAYER nwell ;
        RECT 8.500 14.845 11.580 23.845 ;
        RECT 16.600 14.845 22.380 23.845 ;
        RECT 5.800 10.875 22.380 14.845 ;
      LAYER pwell ;
        RECT 5.950 7.375 22.230 10.605 ;
        RECT 22.650 9.450 24.660 24.180 ;
        RECT 34.075 24.100 36.855 29.950 ;
        RECT 42.175 24.100 47.655 29.950 ;
      LAYER nwell ;
        RECT 33.925 14.845 37.005 23.845 ;
        RECT 42.025 14.845 47.805 23.845 ;
        RECT 31.225 10.875 47.805 14.845 ;
      LAYER pwell ;
        RECT 31.375 7.375 47.655 10.605 ;
        RECT 48.075 9.450 50.085 24.180 ;
        RECT 59.500 24.100 62.280 29.950 ;
        RECT 67.600 24.100 73.080 29.950 ;
      LAYER nwell ;
        RECT 59.350 14.845 62.430 23.845 ;
        RECT 67.450 14.845 73.230 23.845 ;
        RECT 56.650 10.875 73.230 14.845 ;
      LAYER pwell ;
        RECT 56.800 7.375 73.080 10.605 ;
        RECT 73.500 9.450 75.510 24.180 ;
        RECT 84.925 24.100 87.705 29.950 ;
        RECT 93.025 24.100 98.505 29.950 ;
      LAYER nwell ;
        RECT 84.775 14.845 87.855 23.845 ;
        RECT 92.875 14.845 98.655 23.845 ;
        RECT 82.075 10.875 98.655 14.845 ;
      LAYER pwell ;
        RECT 82.225 7.375 98.505 10.605 ;
        RECT 98.925 9.450 100.935 24.180 ;
        RECT 110.350 24.100 113.130 29.950 ;
        RECT 118.450 24.100 123.930 29.950 ;
      LAYER nwell ;
        RECT 110.200 14.845 113.280 23.845 ;
        RECT 118.300 14.845 124.080 23.845 ;
        RECT 107.500 10.875 124.080 14.845 ;
      LAYER pwell ;
        RECT 107.650 7.375 123.930 10.605 ;
        RECT 124.350 9.450 126.360 24.180 ;
        RECT 135.775 24.100 138.555 29.950 ;
        RECT 143.875 24.100 149.355 29.950 ;
      LAYER nwell ;
        RECT 135.625 14.845 138.705 23.845 ;
        RECT 143.725 14.845 149.505 23.845 ;
        RECT 132.925 10.875 149.505 14.845 ;
      LAYER pwell ;
        RECT 133.075 7.375 149.355 10.605 ;
        RECT 149.775 9.450 151.785 24.180 ;
        RECT 8.650 1.525 11.430 7.375 ;
        RECT 16.750 1.525 22.230 7.375 ;
        RECT 34.075 1.525 36.855 7.375 ;
        RECT 42.175 1.525 47.655 7.375 ;
        RECT 59.500 1.525 62.280 7.375 ;
        RECT 67.600 1.525 73.080 7.375 ;
        RECT 84.925 1.525 87.705 7.375 ;
        RECT 93.025 1.525 98.505 7.375 ;
        RECT 110.350 1.525 113.130 7.375 ;
        RECT 118.450 1.525 123.930 7.375 ;
        RECT 135.775 1.525 138.555 7.375 ;
        RECT 143.875 1.525 149.355 7.375 ;
      LAYER li1 ;
        RECT 8.890 212.435 11.190 212.605 ;
        RECT 6.190 203.435 8.490 203.605 ;
        RECT 6.190 202.500 6.360 203.435 ;
        RECT 7.090 202.745 7.590 202.915 ;
        RECT 6.860 202.500 7.030 202.530 ;
        RECT 6.135 201.520 7.030 202.500 ;
        RECT 6.190 200.585 6.360 201.520 ;
        RECT 6.860 201.490 7.030 201.520 ;
        RECT 7.650 201.490 7.820 202.530 ;
        RECT 6.675 201.105 7.590 201.275 ;
        RECT 6.675 200.900 7.510 201.105 ;
        RECT 8.320 200.585 8.490 203.435 ;
        RECT 6.190 200.415 8.490 200.585 ;
        RECT 8.890 200.585 9.060 212.435 ;
        RECT 9.550 211.725 10.550 212.175 ;
        RECT 9.560 201.490 9.730 211.530 ;
        RECT 10.350 201.490 10.520 211.530 ;
        RECT 9.790 201.105 10.290 201.275 ;
        RECT 11.020 200.585 11.190 212.435 ;
        RECT 16.990 212.435 19.290 212.605 ;
        RECT 11.590 203.435 13.890 203.605 ;
        RECT 11.590 202.500 11.760 203.435 ;
        RECT 12.490 202.745 12.990 202.915 ;
        RECT 12.260 202.500 12.430 202.530 ;
        RECT 11.535 201.520 12.430 202.500 ;
        RECT 8.890 200.415 11.190 200.585 ;
        RECT 11.590 200.585 11.760 201.520 ;
        RECT 12.260 201.490 12.430 201.520 ;
        RECT 13.050 201.490 13.220 202.530 ;
        RECT 12.075 201.105 12.990 201.275 ;
        RECT 12.075 200.900 12.910 201.105 ;
        RECT 13.720 200.585 13.890 203.435 ;
        RECT 14.290 203.435 16.590 203.605 ;
        RECT 14.290 202.500 14.460 203.435 ;
        RECT 15.190 202.745 15.690 202.915 ;
        RECT 14.960 202.500 15.130 202.530 ;
        RECT 14.235 201.520 15.130 202.500 ;
        RECT 11.590 200.415 13.890 200.585 ;
        RECT 14.290 200.585 14.460 201.520 ;
        RECT 14.960 201.490 15.130 201.520 ;
        RECT 15.750 201.490 15.920 202.530 ;
        RECT 14.775 201.105 15.690 201.275 ;
        RECT 14.775 200.900 15.610 201.105 ;
        RECT 16.420 200.585 16.590 203.435 ;
        RECT 14.290 200.415 16.590 200.585 ;
        RECT 16.990 200.585 17.160 212.435 ;
        RECT 17.650 211.725 18.650 212.175 ;
        RECT 17.660 201.490 17.830 211.530 ;
        RECT 18.450 201.490 18.620 211.530 ;
        RECT 17.890 201.105 18.390 201.275 ;
        RECT 19.120 200.585 19.290 212.435 ;
        RECT 16.990 200.415 19.290 200.585 ;
        RECT 19.690 212.435 21.990 212.605 ;
        RECT 19.690 200.585 19.860 212.435 ;
        RECT 20.350 211.725 21.350 212.175 ;
        RECT 20.360 201.490 20.530 211.530 ;
        RECT 21.150 201.490 21.320 211.530 ;
        RECT 20.590 201.105 21.090 201.275 ;
        RECT 21.820 200.585 21.990 212.435 ;
        RECT 22.885 212.435 25.185 212.605 ;
        RECT 22.885 211.450 23.055 212.435 ;
        RECT 23.785 211.745 24.285 211.915 ;
        RECT 23.555 211.450 23.725 211.530 ;
        RECT 24.345 211.525 24.515 211.530 ;
        RECT 22.885 210.575 23.725 211.450 ;
        RECT 22.885 209.585 23.055 210.575 ;
        RECT 23.555 210.490 23.725 210.575 ;
        RECT 24.295 210.495 24.770 211.525 ;
        RECT 24.345 210.490 24.515 210.495 ;
        RECT 23.545 209.850 24.520 210.300 ;
        RECT 25.015 209.585 25.185 212.435 ;
        RECT 22.885 209.415 25.185 209.585 ;
        RECT 25.585 212.435 27.885 212.605 ;
        RECT 25.585 209.585 25.755 212.435 ;
        RECT 26.485 211.745 26.985 211.915 ;
        RECT 26.255 211.525 26.425 211.530 ;
        RECT 25.980 210.495 26.475 211.525 ;
        RECT 27.045 211.500 27.215 211.530 ;
        RECT 27.715 211.500 27.885 212.435 ;
        RECT 28.285 212.435 30.585 212.605 ;
        RECT 28.285 211.500 28.455 212.435 ;
        RECT 29.185 211.745 29.685 211.915 ;
        RECT 28.955 211.500 29.125 211.530 ;
        RECT 26.970 210.570 27.890 211.500 ;
        RECT 26.255 210.490 26.425 210.495 ;
        RECT 27.045 210.490 27.215 210.570 ;
        RECT 26.245 209.850 27.220 210.300 ;
        RECT 27.715 209.585 27.885 210.570 ;
        RECT 28.230 210.520 29.125 211.500 ;
        RECT 25.585 209.415 27.885 209.585 ;
        RECT 28.285 209.585 28.455 210.520 ;
        RECT 28.955 210.490 29.125 210.520 ;
        RECT 29.745 210.490 29.915 211.530 ;
        RECT 28.770 210.105 29.685 210.275 ;
        RECT 28.770 209.900 29.605 210.105 ;
        RECT 30.415 209.585 30.585 212.435 ;
        RECT 28.285 209.415 30.585 209.585 ;
        RECT 34.315 212.435 36.615 212.605 ;
        RECT 22.885 208.345 25.185 208.515 ;
        RECT 22.885 205.935 23.055 208.345 ;
        RECT 23.545 207.675 24.520 208.100 ;
        RECT 25.015 208.035 25.185 208.345 ;
        RECT 25.585 208.345 27.885 208.515 ;
        RECT 25.585 208.035 25.755 208.345 ;
        RECT 23.785 207.655 24.285 207.675 ;
        RECT 23.555 207.480 23.725 207.485 ;
        RECT 24.345 207.480 24.515 207.485 ;
        RECT 23.455 206.800 23.825 207.480 ;
        RECT 24.245 206.800 24.615 207.480 ;
        RECT 23.555 206.795 23.725 206.800 ;
        RECT 24.345 206.795 24.515 206.800 ;
        RECT 23.785 206.455 24.285 206.625 ;
        RECT 25.015 206.245 25.755 208.035 ;
        RECT 26.245 207.675 27.220 208.100 ;
        RECT 26.485 207.655 26.985 207.675 ;
        RECT 26.255 207.480 26.425 207.485 ;
        RECT 26.155 206.800 26.525 207.480 ;
        RECT 27.045 207.405 27.215 207.485 ;
        RECT 27.715 207.405 27.885 208.345 ;
        RECT 28.285 208.345 30.585 208.515 ;
        RECT 28.285 207.405 28.455 208.345 ;
        RECT 28.665 207.655 29.705 208.100 ;
        RECT 28.955 207.405 29.125 207.485 ;
        RECT 26.970 206.825 27.890 207.405 ;
        RECT 28.280 206.875 29.125 207.405 ;
        RECT 26.255 206.795 26.425 206.800 ;
        RECT 27.045 206.795 27.215 206.825 ;
        RECT 26.485 206.455 26.985 206.625 ;
        RECT 25.015 205.935 25.185 206.245 ;
        RECT 22.885 205.765 25.185 205.935 ;
        RECT 25.585 205.935 25.755 206.245 ;
        RECT 27.715 205.935 27.885 206.825 ;
        RECT 25.585 205.765 27.885 205.935 ;
        RECT 28.285 205.935 28.455 206.875 ;
        RECT 28.955 206.795 29.125 206.875 ;
        RECT 29.745 206.795 29.915 207.485 ;
        RECT 29.185 206.455 29.685 206.625 ;
        RECT 30.415 205.935 30.585 208.345 ;
        RECT 28.285 205.765 30.585 205.935 ;
        RECT 31.615 203.435 33.915 203.605 ;
        RECT 31.615 202.500 31.785 203.435 ;
        RECT 32.515 202.745 33.015 202.915 ;
        RECT 32.285 202.500 32.455 202.530 ;
        RECT 31.560 201.520 32.455 202.500 ;
        RECT 19.690 200.415 21.990 200.585 ;
        RECT 31.615 200.585 31.785 201.520 ;
        RECT 32.285 201.490 32.455 201.520 ;
        RECT 33.075 201.490 33.245 202.530 ;
        RECT 32.100 201.105 33.015 201.275 ;
        RECT 32.100 200.900 32.935 201.105 ;
        RECT 33.745 200.585 33.915 203.435 ;
        RECT 31.615 200.415 33.915 200.585 ;
        RECT 34.315 200.585 34.485 212.435 ;
        RECT 34.975 211.725 35.975 212.175 ;
        RECT 34.985 201.490 35.155 211.530 ;
        RECT 35.775 201.490 35.945 211.530 ;
        RECT 35.215 201.105 35.715 201.275 ;
        RECT 36.445 200.585 36.615 212.435 ;
        RECT 42.415 212.435 44.715 212.605 ;
        RECT 37.015 203.435 39.315 203.605 ;
        RECT 37.015 202.500 37.185 203.435 ;
        RECT 37.915 202.745 38.415 202.915 ;
        RECT 37.685 202.500 37.855 202.530 ;
        RECT 36.960 201.520 37.855 202.500 ;
        RECT 34.315 200.415 36.615 200.585 ;
        RECT 37.015 200.585 37.185 201.520 ;
        RECT 37.685 201.490 37.855 201.520 ;
        RECT 38.475 201.490 38.645 202.530 ;
        RECT 37.500 201.105 38.415 201.275 ;
        RECT 37.500 200.900 38.335 201.105 ;
        RECT 39.145 200.585 39.315 203.435 ;
        RECT 39.715 203.435 42.015 203.605 ;
        RECT 39.715 202.500 39.885 203.435 ;
        RECT 40.615 202.745 41.115 202.915 ;
        RECT 40.385 202.500 40.555 202.530 ;
        RECT 39.660 201.520 40.555 202.500 ;
        RECT 37.015 200.415 39.315 200.585 ;
        RECT 39.715 200.585 39.885 201.520 ;
        RECT 40.385 201.490 40.555 201.520 ;
        RECT 41.175 201.490 41.345 202.530 ;
        RECT 40.200 201.105 41.115 201.275 ;
        RECT 40.200 200.900 41.035 201.105 ;
        RECT 41.845 200.585 42.015 203.435 ;
        RECT 39.715 200.415 42.015 200.585 ;
        RECT 42.415 200.585 42.585 212.435 ;
        RECT 43.075 211.725 44.075 212.175 ;
        RECT 43.085 201.490 43.255 211.530 ;
        RECT 43.875 201.490 44.045 211.530 ;
        RECT 43.315 201.105 43.815 201.275 ;
        RECT 44.545 200.585 44.715 212.435 ;
        RECT 42.415 200.415 44.715 200.585 ;
        RECT 45.115 212.435 47.415 212.605 ;
        RECT 45.115 200.585 45.285 212.435 ;
        RECT 45.775 211.725 46.775 212.175 ;
        RECT 45.785 201.490 45.955 211.530 ;
        RECT 46.575 201.490 46.745 211.530 ;
        RECT 46.015 201.105 46.515 201.275 ;
        RECT 47.245 200.585 47.415 212.435 ;
        RECT 59.740 212.435 62.040 212.605 ;
        RECT 57.040 203.435 59.340 203.605 ;
        RECT 57.040 202.500 57.210 203.435 ;
        RECT 57.940 202.745 58.440 202.915 ;
        RECT 57.710 202.500 57.880 202.530 ;
        RECT 56.985 201.520 57.880 202.500 ;
        RECT 45.115 200.415 47.415 200.585 ;
        RECT 57.040 200.585 57.210 201.520 ;
        RECT 57.710 201.490 57.880 201.520 ;
        RECT 58.500 201.490 58.670 202.530 ;
        RECT 57.525 201.105 58.440 201.275 ;
        RECT 57.525 200.900 58.360 201.105 ;
        RECT 59.170 200.585 59.340 203.435 ;
        RECT 57.040 200.415 59.340 200.585 ;
        RECT 59.740 200.585 59.910 212.435 ;
        RECT 60.400 211.725 61.400 212.175 ;
        RECT 60.410 201.490 60.580 211.530 ;
        RECT 61.200 201.490 61.370 211.530 ;
        RECT 60.640 201.105 61.140 201.275 ;
        RECT 61.870 200.585 62.040 212.435 ;
        RECT 67.840 212.435 70.140 212.605 ;
        RECT 62.440 203.435 64.740 203.605 ;
        RECT 62.440 202.500 62.610 203.435 ;
        RECT 63.340 202.745 63.840 202.915 ;
        RECT 63.110 202.500 63.280 202.530 ;
        RECT 62.385 201.520 63.280 202.500 ;
        RECT 59.740 200.415 62.040 200.585 ;
        RECT 62.440 200.585 62.610 201.520 ;
        RECT 63.110 201.490 63.280 201.520 ;
        RECT 63.900 201.490 64.070 202.530 ;
        RECT 62.925 201.105 63.840 201.275 ;
        RECT 62.925 200.900 63.760 201.105 ;
        RECT 64.570 200.585 64.740 203.435 ;
        RECT 65.140 203.435 67.440 203.605 ;
        RECT 65.140 202.500 65.310 203.435 ;
        RECT 66.040 202.745 66.540 202.915 ;
        RECT 65.810 202.500 65.980 202.530 ;
        RECT 65.085 201.520 65.980 202.500 ;
        RECT 62.440 200.415 64.740 200.585 ;
        RECT 65.140 200.585 65.310 201.520 ;
        RECT 65.810 201.490 65.980 201.520 ;
        RECT 66.600 201.490 66.770 202.530 ;
        RECT 65.625 201.105 66.540 201.275 ;
        RECT 65.625 200.900 66.460 201.105 ;
        RECT 67.270 200.585 67.440 203.435 ;
        RECT 65.140 200.415 67.440 200.585 ;
        RECT 67.840 200.585 68.010 212.435 ;
        RECT 68.500 211.725 69.500 212.175 ;
        RECT 68.510 201.490 68.680 211.530 ;
        RECT 69.300 201.490 69.470 211.530 ;
        RECT 68.740 201.105 69.240 201.275 ;
        RECT 69.970 200.585 70.140 212.435 ;
        RECT 67.840 200.415 70.140 200.585 ;
        RECT 70.540 212.435 72.840 212.605 ;
        RECT 70.540 200.585 70.710 212.435 ;
        RECT 71.200 211.725 72.200 212.175 ;
        RECT 71.210 201.490 71.380 211.530 ;
        RECT 72.000 201.490 72.170 211.530 ;
        RECT 71.440 201.105 71.940 201.275 ;
        RECT 72.670 200.585 72.840 212.435 ;
        RECT 73.735 212.435 76.035 212.605 ;
        RECT 73.735 211.450 73.905 212.435 ;
        RECT 74.635 211.745 75.135 211.915 ;
        RECT 74.405 211.450 74.575 211.530 ;
        RECT 75.195 211.525 75.365 211.530 ;
        RECT 73.735 210.575 74.575 211.450 ;
        RECT 73.735 209.585 73.905 210.575 ;
        RECT 74.405 210.490 74.575 210.575 ;
        RECT 75.145 210.495 75.620 211.525 ;
        RECT 75.195 210.490 75.365 210.495 ;
        RECT 74.395 209.850 75.370 210.300 ;
        RECT 75.865 209.585 76.035 212.435 ;
        RECT 73.735 209.415 76.035 209.585 ;
        RECT 76.435 212.435 78.735 212.605 ;
        RECT 76.435 209.585 76.605 212.435 ;
        RECT 77.335 211.745 77.835 211.915 ;
        RECT 77.105 211.525 77.275 211.530 ;
        RECT 76.830 210.495 77.325 211.525 ;
        RECT 77.895 211.500 78.065 211.530 ;
        RECT 78.565 211.500 78.735 212.435 ;
        RECT 79.135 212.435 81.435 212.605 ;
        RECT 79.135 211.500 79.305 212.435 ;
        RECT 80.035 211.745 80.535 211.915 ;
        RECT 79.805 211.500 79.975 211.530 ;
        RECT 77.820 210.570 78.740 211.500 ;
        RECT 77.105 210.490 77.275 210.495 ;
        RECT 77.895 210.490 78.065 210.570 ;
        RECT 77.095 209.850 78.070 210.300 ;
        RECT 78.565 209.585 78.735 210.570 ;
        RECT 79.080 210.520 79.975 211.500 ;
        RECT 76.435 209.415 78.735 209.585 ;
        RECT 79.135 209.585 79.305 210.520 ;
        RECT 79.805 210.490 79.975 210.520 ;
        RECT 80.595 210.490 80.765 211.530 ;
        RECT 79.620 210.105 80.535 210.275 ;
        RECT 79.620 209.900 80.455 210.105 ;
        RECT 81.265 209.585 81.435 212.435 ;
        RECT 79.135 209.415 81.435 209.585 ;
        RECT 85.165 212.435 87.465 212.605 ;
        RECT 73.735 208.345 76.035 208.515 ;
        RECT 73.735 205.935 73.905 208.345 ;
        RECT 74.395 207.675 75.370 208.100 ;
        RECT 75.865 208.035 76.035 208.345 ;
        RECT 76.435 208.345 78.735 208.515 ;
        RECT 76.435 208.035 76.605 208.345 ;
        RECT 74.635 207.655 75.135 207.675 ;
        RECT 74.405 207.480 74.575 207.485 ;
        RECT 75.195 207.480 75.365 207.485 ;
        RECT 74.305 206.800 74.675 207.480 ;
        RECT 75.095 206.800 75.465 207.480 ;
        RECT 74.405 206.795 74.575 206.800 ;
        RECT 75.195 206.795 75.365 206.800 ;
        RECT 74.635 206.455 75.135 206.625 ;
        RECT 75.865 206.245 76.605 208.035 ;
        RECT 77.095 207.675 78.070 208.100 ;
        RECT 77.335 207.655 77.835 207.675 ;
        RECT 77.105 207.480 77.275 207.485 ;
        RECT 77.005 206.800 77.375 207.480 ;
        RECT 77.895 207.405 78.065 207.485 ;
        RECT 78.565 207.405 78.735 208.345 ;
        RECT 79.135 208.345 81.435 208.515 ;
        RECT 79.135 207.405 79.305 208.345 ;
        RECT 79.515 207.655 80.555 208.100 ;
        RECT 79.805 207.405 79.975 207.485 ;
        RECT 77.820 206.825 78.740 207.405 ;
        RECT 79.130 206.875 79.975 207.405 ;
        RECT 77.105 206.795 77.275 206.800 ;
        RECT 77.895 206.795 78.065 206.825 ;
        RECT 77.335 206.455 77.835 206.625 ;
        RECT 75.865 205.935 76.035 206.245 ;
        RECT 73.735 205.765 76.035 205.935 ;
        RECT 76.435 205.935 76.605 206.245 ;
        RECT 78.565 205.935 78.735 206.825 ;
        RECT 76.435 205.765 78.735 205.935 ;
        RECT 79.135 205.935 79.305 206.875 ;
        RECT 79.805 206.795 79.975 206.875 ;
        RECT 80.595 206.795 80.765 207.485 ;
        RECT 80.035 206.455 80.535 206.625 ;
        RECT 81.265 205.935 81.435 208.345 ;
        RECT 79.135 205.765 81.435 205.935 ;
        RECT 82.465 203.435 84.765 203.605 ;
        RECT 82.465 202.500 82.635 203.435 ;
        RECT 83.365 202.745 83.865 202.915 ;
        RECT 83.135 202.500 83.305 202.530 ;
        RECT 82.410 201.520 83.305 202.500 ;
        RECT 70.540 200.415 72.840 200.585 ;
        RECT 82.465 200.585 82.635 201.520 ;
        RECT 83.135 201.490 83.305 201.520 ;
        RECT 83.925 201.490 84.095 202.530 ;
        RECT 82.950 201.105 83.865 201.275 ;
        RECT 82.950 200.900 83.785 201.105 ;
        RECT 84.595 200.585 84.765 203.435 ;
        RECT 82.465 200.415 84.765 200.585 ;
        RECT 85.165 200.585 85.335 212.435 ;
        RECT 85.825 211.725 86.825 212.175 ;
        RECT 85.835 201.490 86.005 211.530 ;
        RECT 86.625 201.490 86.795 211.530 ;
        RECT 86.065 201.105 86.565 201.275 ;
        RECT 87.295 200.585 87.465 212.435 ;
        RECT 93.265 212.435 95.565 212.605 ;
        RECT 87.865 203.435 90.165 203.605 ;
        RECT 87.865 202.500 88.035 203.435 ;
        RECT 88.765 202.745 89.265 202.915 ;
        RECT 88.535 202.500 88.705 202.530 ;
        RECT 87.810 201.520 88.705 202.500 ;
        RECT 85.165 200.415 87.465 200.585 ;
        RECT 87.865 200.585 88.035 201.520 ;
        RECT 88.535 201.490 88.705 201.520 ;
        RECT 89.325 201.490 89.495 202.530 ;
        RECT 88.350 201.105 89.265 201.275 ;
        RECT 88.350 200.900 89.185 201.105 ;
        RECT 89.995 200.585 90.165 203.435 ;
        RECT 90.565 203.435 92.865 203.605 ;
        RECT 90.565 202.500 90.735 203.435 ;
        RECT 91.465 202.745 91.965 202.915 ;
        RECT 91.235 202.500 91.405 202.530 ;
        RECT 90.510 201.520 91.405 202.500 ;
        RECT 87.865 200.415 90.165 200.585 ;
        RECT 90.565 200.585 90.735 201.520 ;
        RECT 91.235 201.490 91.405 201.520 ;
        RECT 92.025 201.490 92.195 202.530 ;
        RECT 91.050 201.105 91.965 201.275 ;
        RECT 91.050 200.900 91.885 201.105 ;
        RECT 92.695 200.585 92.865 203.435 ;
        RECT 90.565 200.415 92.865 200.585 ;
        RECT 93.265 200.585 93.435 212.435 ;
        RECT 93.925 211.725 94.925 212.175 ;
        RECT 93.935 201.490 94.105 211.530 ;
        RECT 94.725 201.490 94.895 211.530 ;
        RECT 94.165 201.105 94.665 201.275 ;
        RECT 95.395 200.585 95.565 212.435 ;
        RECT 93.265 200.415 95.565 200.585 ;
        RECT 95.965 212.435 98.265 212.605 ;
        RECT 95.965 200.585 96.135 212.435 ;
        RECT 96.625 211.725 97.625 212.175 ;
        RECT 96.635 201.490 96.805 211.530 ;
        RECT 97.425 201.490 97.595 211.530 ;
        RECT 96.865 201.105 97.365 201.275 ;
        RECT 98.095 200.585 98.265 212.435 ;
        RECT 110.590 212.435 112.890 212.605 ;
        RECT 107.890 203.435 110.190 203.605 ;
        RECT 107.890 202.500 108.060 203.435 ;
        RECT 108.790 202.745 109.290 202.915 ;
        RECT 108.560 202.500 108.730 202.530 ;
        RECT 107.835 201.520 108.730 202.500 ;
        RECT 95.965 200.415 98.265 200.585 ;
        RECT 107.890 200.585 108.060 201.520 ;
        RECT 108.560 201.490 108.730 201.520 ;
        RECT 109.350 201.490 109.520 202.530 ;
        RECT 108.375 201.105 109.290 201.275 ;
        RECT 108.375 200.900 109.210 201.105 ;
        RECT 110.020 200.585 110.190 203.435 ;
        RECT 107.890 200.415 110.190 200.585 ;
        RECT 110.590 200.585 110.760 212.435 ;
        RECT 111.250 211.725 112.250 212.175 ;
        RECT 111.260 201.490 111.430 211.530 ;
        RECT 112.050 201.490 112.220 211.530 ;
        RECT 111.490 201.105 111.990 201.275 ;
        RECT 112.720 200.585 112.890 212.435 ;
        RECT 118.690 212.435 120.990 212.605 ;
        RECT 113.290 203.435 115.590 203.605 ;
        RECT 113.290 202.500 113.460 203.435 ;
        RECT 114.190 202.745 114.690 202.915 ;
        RECT 113.960 202.500 114.130 202.530 ;
        RECT 113.235 201.520 114.130 202.500 ;
        RECT 110.590 200.415 112.890 200.585 ;
        RECT 113.290 200.585 113.460 201.520 ;
        RECT 113.960 201.490 114.130 201.520 ;
        RECT 114.750 201.490 114.920 202.530 ;
        RECT 113.775 201.105 114.690 201.275 ;
        RECT 113.775 200.900 114.610 201.105 ;
        RECT 115.420 200.585 115.590 203.435 ;
        RECT 115.990 203.435 118.290 203.605 ;
        RECT 115.990 202.500 116.160 203.435 ;
        RECT 116.890 202.745 117.390 202.915 ;
        RECT 116.660 202.500 116.830 202.530 ;
        RECT 115.935 201.520 116.830 202.500 ;
        RECT 113.290 200.415 115.590 200.585 ;
        RECT 115.990 200.585 116.160 201.520 ;
        RECT 116.660 201.490 116.830 201.520 ;
        RECT 117.450 201.490 117.620 202.530 ;
        RECT 116.475 201.105 117.390 201.275 ;
        RECT 116.475 200.900 117.310 201.105 ;
        RECT 118.120 200.585 118.290 203.435 ;
        RECT 115.990 200.415 118.290 200.585 ;
        RECT 118.690 200.585 118.860 212.435 ;
        RECT 119.350 211.725 120.350 212.175 ;
        RECT 119.360 201.490 119.530 211.530 ;
        RECT 120.150 201.490 120.320 211.530 ;
        RECT 119.590 201.105 120.090 201.275 ;
        RECT 120.820 200.585 120.990 212.435 ;
        RECT 118.690 200.415 120.990 200.585 ;
        RECT 121.390 212.435 123.690 212.605 ;
        RECT 121.390 200.585 121.560 212.435 ;
        RECT 122.050 211.725 123.050 212.175 ;
        RECT 122.060 201.490 122.230 211.530 ;
        RECT 122.850 201.490 123.020 211.530 ;
        RECT 122.290 201.105 122.790 201.275 ;
        RECT 123.520 200.585 123.690 212.435 ;
        RECT 124.585 212.435 126.885 212.605 ;
        RECT 124.585 211.450 124.755 212.435 ;
        RECT 125.485 211.745 125.985 211.915 ;
        RECT 125.255 211.450 125.425 211.530 ;
        RECT 126.045 211.525 126.215 211.530 ;
        RECT 124.585 210.575 125.425 211.450 ;
        RECT 124.585 209.585 124.755 210.575 ;
        RECT 125.255 210.490 125.425 210.575 ;
        RECT 125.995 210.495 126.470 211.525 ;
        RECT 126.045 210.490 126.215 210.495 ;
        RECT 125.245 209.850 126.220 210.300 ;
        RECT 126.715 209.585 126.885 212.435 ;
        RECT 124.585 209.415 126.885 209.585 ;
        RECT 127.285 212.435 129.585 212.605 ;
        RECT 127.285 209.585 127.455 212.435 ;
        RECT 128.185 211.745 128.685 211.915 ;
        RECT 127.955 211.525 128.125 211.530 ;
        RECT 127.680 210.495 128.175 211.525 ;
        RECT 128.745 211.500 128.915 211.530 ;
        RECT 129.415 211.500 129.585 212.435 ;
        RECT 129.985 212.435 132.285 212.605 ;
        RECT 129.985 211.500 130.155 212.435 ;
        RECT 130.885 211.745 131.385 211.915 ;
        RECT 130.655 211.500 130.825 211.530 ;
        RECT 128.670 210.570 129.590 211.500 ;
        RECT 127.955 210.490 128.125 210.495 ;
        RECT 128.745 210.490 128.915 210.570 ;
        RECT 127.945 209.850 128.920 210.300 ;
        RECT 129.415 209.585 129.585 210.570 ;
        RECT 129.930 210.520 130.825 211.500 ;
        RECT 127.285 209.415 129.585 209.585 ;
        RECT 129.985 209.585 130.155 210.520 ;
        RECT 130.655 210.490 130.825 210.520 ;
        RECT 131.445 210.490 131.615 211.530 ;
        RECT 130.470 210.105 131.385 210.275 ;
        RECT 130.470 209.900 131.305 210.105 ;
        RECT 132.115 209.585 132.285 212.435 ;
        RECT 129.985 209.415 132.285 209.585 ;
        RECT 136.015 212.435 138.315 212.605 ;
        RECT 124.585 208.345 126.885 208.515 ;
        RECT 124.585 205.935 124.755 208.345 ;
        RECT 125.245 207.675 126.220 208.100 ;
        RECT 126.715 208.035 126.885 208.345 ;
        RECT 127.285 208.345 129.585 208.515 ;
        RECT 127.285 208.035 127.455 208.345 ;
        RECT 125.485 207.655 125.985 207.675 ;
        RECT 125.255 207.480 125.425 207.485 ;
        RECT 126.045 207.480 126.215 207.485 ;
        RECT 125.155 206.800 125.525 207.480 ;
        RECT 125.945 206.800 126.315 207.480 ;
        RECT 125.255 206.795 125.425 206.800 ;
        RECT 126.045 206.795 126.215 206.800 ;
        RECT 125.485 206.455 125.985 206.625 ;
        RECT 126.715 206.245 127.455 208.035 ;
        RECT 127.945 207.675 128.920 208.100 ;
        RECT 128.185 207.655 128.685 207.675 ;
        RECT 127.955 207.480 128.125 207.485 ;
        RECT 127.855 206.800 128.225 207.480 ;
        RECT 128.745 207.405 128.915 207.485 ;
        RECT 129.415 207.405 129.585 208.345 ;
        RECT 129.985 208.345 132.285 208.515 ;
        RECT 129.985 207.405 130.155 208.345 ;
        RECT 130.365 207.655 131.405 208.100 ;
        RECT 130.655 207.405 130.825 207.485 ;
        RECT 128.670 206.825 129.590 207.405 ;
        RECT 129.980 206.875 130.825 207.405 ;
        RECT 127.955 206.795 128.125 206.800 ;
        RECT 128.745 206.795 128.915 206.825 ;
        RECT 128.185 206.455 128.685 206.625 ;
        RECT 126.715 205.935 126.885 206.245 ;
        RECT 124.585 205.765 126.885 205.935 ;
        RECT 127.285 205.935 127.455 206.245 ;
        RECT 129.415 205.935 129.585 206.825 ;
        RECT 127.285 205.765 129.585 205.935 ;
        RECT 129.985 205.935 130.155 206.875 ;
        RECT 130.655 206.795 130.825 206.875 ;
        RECT 131.445 206.795 131.615 207.485 ;
        RECT 130.885 206.455 131.385 206.625 ;
        RECT 132.115 205.935 132.285 208.345 ;
        RECT 129.985 205.765 132.285 205.935 ;
        RECT 133.315 203.435 135.615 203.605 ;
        RECT 133.315 202.500 133.485 203.435 ;
        RECT 134.215 202.745 134.715 202.915 ;
        RECT 133.985 202.500 134.155 202.530 ;
        RECT 133.260 201.520 134.155 202.500 ;
        RECT 121.390 200.415 123.690 200.585 ;
        RECT 133.315 200.585 133.485 201.520 ;
        RECT 133.985 201.490 134.155 201.520 ;
        RECT 134.775 201.490 134.945 202.530 ;
        RECT 133.800 201.105 134.715 201.275 ;
        RECT 133.800 200.900 134.635 201.105 ;
        RECT 135.445 200.585 135.615 203.435 ;
        RECT 133.315 200.415 135.615 200.585 ;
        RECT 136.015 200.585 136.185 212.435 ;
        RECT 136.675 211.725 137.675 212.175 ;
        RECT 136.685 201.490 136.855 211.530 ;
        RECT 137.475 201.490 137.645 211.530 ;
        RECT 136.915 201.105 137.415 201.275 ;
        RECT 138.145 200.585 138.315 212.435 ;
        RECT 144.115 212.435 146.415 212.605 ;
        RECT 138.715 203.435 141.015 203.605 ;
        RECT 138.715 202.500 138.885 203.435 ;
        RECT 139.615 202.745 140.115 202.915 ;
        RECT 139.385 202.500 139.555 202.530 ;
        RECT 138.660 201.520 139.555 202.500 ;
        RECT 136.015 200.415 138.315 200.585 ;
        RECT 138.715 200.585 138.885 201.520 ;
        RECT 139.385 201.490 139.555 201.520 ;
        RECT 140.175 201.490 140.345 202.530 ;
        RECT 139.200 201.105 140.115 201.275 ;
        RECT 139.200 200.900 140.035 201.105 ;
        RECT 140.845 200.585 141.015 203.435 ;
        RECT 141.415 203.435 143.715 203.605 ;
        RECT 141.415 202.500 141.585 203.435 ;
        RECT 142.315 202.745 142.815 202.915 ;
        RECT 142.085 202.500 142.255 202.530 ;
        RECT 141.360 201.520 142.255 202.500 ;
        RECT 138.715 200.415 141.015 200.585 ;
        RECT 141.415 200.585 141.585 201.520 ;
        RECT 142.085 201.490 142.255 201.520 ;
        RECT 142.875 201.490 143.045 202.530 ;
        RECT 141.900 201.105 142.815 201.275 ;
        RECT 141.900 200.900 142.735 201.105 ;
        RECT 143.545 200.585 143.715 203.435 ;
        RECT 141.415 200.415 143.715 200.585 ;
        RECT 144.115 200.585 144.285 212.435 ;
        RECT 144.775 211.725 145.775 212.175 ;
        RECT 144.785 201.490 144.955 211.530 ;
        RECT 145.575 201.490 145.745 211.530 ;
        RECT 145.015 201.105 145.515 201.275 ;
        RECT 146.245 200.585 146.415 212.435 ;
        RECT 144.115 200.415 146.415 200.585 ;
        RECT 146.815 212.435 149.115 212.605 ;
        RECT 146.815 200.585 146.985 212.435 ;
        RECT 147.475 211.725 148.475 212.175 ;
        RECT 147.485 201.490 147.655 211.530 ;
        RECT 148.275 201.490 148.445 211.530 ;
        RECT 147.715 201.105 148.215 201.275 ;
        RECT 148.945 200.585 149.115 212.435 ;
        RECT 146.815 200.415 149.115 200.585 ;
        RECT 6.190 199.345 8.490 199.515 ;
        RECT 6.190 198.405 6.360 199.345 ;
        RECT 6.570 198.655 7.610 199.100 ;
        RECT 6.860 198.405 7.030 198.485 ;
        RECT 6.185 197.875 7.030 198.405 ;
        RECT 6.190 196.935 6.360 197.875 ;
        RECT 6.860 197.795 7.030 197.875 ;
        RECT 7.650 197.795 7.820 198.485 ;
        RECT 7.090 197.455 7.590 197.625 ;
        RECT 8.320 196.935 8.490 199.345 ;
        RECT 6.190 196.765 8.490 196.935 ;
        RECT 8.890 199.345 11.190 199.515 ;
        RECT 8.890 191.085 9.060 199.345 ;
        RECT 9.790 198.655 10.290 198.825 ;
        RECT 9.560 191.945 9.730 198.485 ;
        RECT 10.350 191.945 10.520 198.485 ;
        RECT 9.550 191.375 10.550 191.775 ;
        RECT 11.020 191.085 11.190 199.345 ;
        RECT 11.590 199.345 13.890 199.515 ;
        RECT 11.590 198.405 11.760 199.345 ;
        RECT 11.970 198.655 13.010 199.100 ;
        RECT 12.260 198.405 12.430 198.485 ;
        RECT 11.585 197.875 12.430 198.405 ;
        RECT 11.590 196.935 11.760 197.875 ;
        RECT 12.260 197.795 12.430 197.875 ;
        RECT 13.050 197.795 13.220 198.485 ;
        RECT 12.490 197.455 12.990 197.625 ;
        RECT 13.720 196.935 13.890 199.345 ;
        RECT 14.290 199.345 16.590 199.515 ;
        RECT 14.290 198.405 14.460 199.345 ;
        RECT 14.670 198.655 15.710 199.100 ;
        RECT 14.960 198.405 15.130 198.485 ;
        RECT 14.285 197.875 15.130 198.405 ;
        RECT 11.590 196.765 13.890 196.935 ;
        RECT 14.290 196.935 14.460 197.875 ;
        RECT 14.960 197.795 15.130 197.875 ;
        RECT 15.750 197.795 15.920 198.485 ;
        RECT 15.190 197.455 15.690 197.625 ;
        RECT 16.420 196.935 16.590 199.345 ;
        RECT 14.290 196.765 16.590 196.935 ;
        RECT 16.990 199.345 19.290 199.515 ;
        RECT 8.890 190.915 11.190 191.085 ;
        RECT 16.990 191.085 17.160 199.345 ;
        RECT 17.890 198.655 18.390 198.825 ;
        RECT 17.660 191.945 17.830 198.485 ;
        RECT 18.450 191.945 18.620 198.485 ;
        RECT 17.650 191.375 18.650 191.775 ;
        RECT 19.120 191.085 19.290 199.345 ;
        RECT 16.990 190.915 19.290 191.085 ;
        RECT 19.690 199.345 21.990 199.515 ;
        RECT 19.690 191.085 19.860 199.345 ;
        RECT 20.590 198.655 21.090 198.825 ;
        RECT 20.360 191.945 20.530 198.485 ;
        RECT 21.150 191.945 21.320 198.485 ;
        RECT 20.350 191.375 21.350 191.775 ;
        RECT 21.820 191.085 21.990 199.345 ;
        RECT 31.615 199.345 33.915 199.515 ;
        RECT 31.615 198.405 31.785 199.345 ;
        RECT 31.995 198.655 33.035 199.100 ;
        RECT 32.285 198.405 32.455 198.485 ;
        RECT 31.610 197.875 32.455 198.405 ;
        RECT 31.615 196.935 31.785 197.875 ;
        RECT 32.285 197.795 32.455 197.875 ;
        RECT 33.075 197.795 33.245 198.485 ;
        RECT 32.515 197.455 33.015 197.625 ;
        RECT 33.745 196.935 33.915 199.345 ;
        RECT 31.615 196.765 33.915 196.935 ;
        RECT 34.315 199.345 36.615 199.515 ;
        RECT 19.690 190.915 21.990 191.085 ;
        RECT 34.315 191.085 34.485 199.345 ;
        RECT 35.215 198.655 35.715 198.825 ;
        RECT 34.985 191.945 35.155 198.485 ;
        RECT 35.775 191.945 35.945 198.485 ;
        RECT 34.975 191.375 35.975 191.775 ;
        RECT 36.445 191.085 36.615 199.345 ;
        RECT 37.015 199.345 39.315 199.515 ;
        RECT 37.015 198.405 37.185 199.345 ;
        RECT 37.395 198.655 38.435 199.100 ;
        RECT 37.685 198.405 37.855 198.485 ;
        RECT 37.010 197.875 37.855 198.405 ;
        RECT 37.015 196.935 37.185 197.875 ;
        RECT 37.685 197.795 37.855 197.875 ;
        RECT 38.475 197.795 38.645 198.485 ;
        RECT 37.915 197.455 38.415 197.625 ;
        RECT 39.145 196.935 39.315 199.345 ;
        RECT 39.715 199.345 42.015 199.515 ;
        RECT 39.715 198.405 39.885 199.345 ;
        RECT 40.095 198.655 41.135 199.100 ;
        RECT 40.385 198.405 40.555 198.485 ;
        RECT 39.710 197.875 40.555 198.405 ;
        RECT 37.015 196.765 39.315 196.935 ;
        RECT 39.715 196.935 39.885 197.875 ;
        RECT 40.385 197.795 40.555 197.875 ;
        RECT 41.175 197.795 41.345 198.485 ;
        RECT 40.615 197.455 41.115 197.625 ;
        RECT 41.845 196.935 42.015 199.345 ;
        RECT 39.715 196.765 42.015 196.935 ;
        RECT 42.415 199.345 44.715 199.515 ;
        RECT 34.315 190.915 36.615 191.085 ;
        RECT 42.415 191.085 42.585 199.345 ;
        RECT 43.315 198.655 43.815 198.825 ;
        RECT 43.085 191.945 43.255 198.485 ;
        RECT 43.875 191.945 44.045 198.485 ;
        RECT 43.075 191.375 44.075 191.775 ;
        RECT 44.545 191.085 44.715 199.345 ;
        RECT 42.415 190.915 44.715 191.085 ;
        RECT 45.115 199.345 47.415 199.515 ;
        RECT 45.115 191.085 45.285 199.345 ;
        RECT 46.015 198.655 46.515 198.825 ;
        RECT 45.785 191.945 45.955 198.485 ;
        RECT 46.575 191.945 46.745 198.485 ;
        RECT 45.775 191.375 46.775 191.775 ;
        RECT 47.245 191.085 47.415 199.345 ;
        RECT 57.040 199.345 59.340 199.515 ;
        RECT 57.040 198.405 57.210 199.345 ;
        RECT 57.420 198.655 58.460 199.100 ;
        RECT 57.710 198.405 57.880 198.485 ;
        RECT 57.035 197.875 57.880 198.405 ;
        RECT 57.040 196.935 57.210 197.875 ;
        RECT 57.710 197.795 57.880 197.875 ;
        RECT 58.500 197.795 58.670 198.485 ;
        RECT 57.940 197.455 58.440 197.625 ;
        RECT 59.170 196.935 59.340 199.345 ;
        RECT 57.040 196.765 59.340 196.935 ;
        RECT 59.740 199.345 62.040 199.515 ;
        RECT 45.115 190.915 47.415 191.085 ;
        RECT 59.740 191.085 59.910 199.345 ;
        RECT 60.640 198.655 61.140 198.825 ;
        RECT 60.410 191.945 60.580 198.485 ;
        RECT 61.200 191.945 61.370 198.485 ;
        RECT 60.400 191.375 61.400 191.775 ;
        RECT 61.870 191.085 62.040 199.345 ;
        RECT 62.440 199.345 64.740 199.515 ;
        RECT 62.440 198.405 62.610 199.345 ;
        RECT 62.820 198.655 63.860 199.100 ;
        RECT 63.110 198.405 63.280 198.485 ;
        RECT 62.435 197.875 63.280 198.405 ;
        RECT 62.440 196.935 62.610 197.875 ;
        RECT 63.110 197.795 63.280 197.875 ;
        RECT 63.900 197.795 64.070 198.485 ;
        RECT 63.340 197.455 63.840 197.625 ;
        RECT 64.570 196.935 64.740 199.345 ;
        RECT 65.140 199.345 67.440 199.515 ;
        RECT 65.140 198.405 65.310 199.345 ;
        RECT 65.520 198.655 66.560 199.100 ;
        RECT 65.810 198.405 65.980 198.485 ;
        RECT 65.135 197.875 65.980 198.405 ;
        RECT 62.440 196.765 64.740 196.935 ;
        RECT 65.140 196.935 65.310 197.875 ;
        RECT 65.810 197.795 65.980 197.875 ;
        RECT 66.600 197.795 66.770 198.485 ;
        RECT 66.040 197.455 66.540 197.625 ;
        RECT 67.270 196.935 67.440 199.345 ;
        RECT 65.140 196.765 67.440 196.935 ;
        RECT 67.840 199.345 70.140 199.515 ;
        RECT 59.740 190.915 62.040 191.085 ;
        RECT 67.840 191.085 68.010 199.345 ;
        RECT 68.740 198.655 69.240 198.825 ;
        RECT 68.510 191.945 68.680 198.485 ;
        RECT 69.300 191.945 69.470 198.485 ;
        RECT 68.500 191.375 69.500 191.775 ;
        RECT 69.970 191.085 70.140 199.345 ;
        RECT 67.840 190.915 70.140 191.085 ;
        RECT 70.540 199.345 72.840 199.515 ;
        RECT 70.540 191.085 70.710 199.345 ;
        RECT 71.440 198.655 71.940 198.825 ;
        RECT 71.210 191.945 71.380 198.485 ;
        RECT 72.000 191.945 72.170 198.485 ;
        RECT 71.200 191.375 72.200 191.775 ;
        RECT 72.670 191.085 72.840 199.345 ;
        RECT 82.465 199.345 84.765 199.515 ;
        RECT 82.465 198.405 82.635 199.345 ;
        RECT 82.845 198.655 83.885 199.100 ;
        RECT 83.135 198.405 83.305 198.485 ;
        RECT 82.460 197.875 83.305 198.405 ;
        RECT 82.465 196.935 82.635 197.875 ;
        RECT 83.135 197.795 83.305 197.875 ;
        RECT 83.925 197.795 84.095 198.485 ;
        RECT 83.365 197.455 83.865 197.625 ;
        RECT 84.595 196.935 84.765 199.345 ;
        RECT 82.465 196.765 84.765 196.935 ;
        RECT 85.165 199.345 87.465 199.515 ;
        RECT 70.540 190.915 72.840 191.085 ;
        RECT 85.165 191.085 85.335 199.345 ;
        RECT 86.065 198.655 86.565 198.825 ;
        RECT 85.835 191.945 86.005 198.485 ;
        RECT 86.625 191.945 86.795 198.485 ;
        RECT 85.825 191.375 86.825 191.775 ;
        RECT 87.295 191.085 87.465 199.345 ;
        RECT 87.865 199.345 90.165 199.515 ;
        RECT 87.865 198.405 88.035 199.345 ;
        RECT 88.245 198.655 89.285 199.100 ;
        RECT 88.535 198.405 88.705 198.485 ;
        RECT 87.860 197.875 88.705 198.405 ;
        RECT 87.865 196.935 88.035 197.875 ;
        RECT 88.535 197.795 88.705 197.875 ;
        RECT 89.325 197.795 89.495 198.485 ;
        RECT 88.765 197.455 89.265 197.625 ;
        RECT 89.995 196.935 90.165 199.345 ;
        RECT 90.565 199.345 92.865 199.515 ;
        RECT 90.565 198.405 90.735 199.345 ;
        RECT 90.945 198.655 91.985 199.100 ;
        RECT 91.235 198.405 91.405 198.485 ;
        RECT 90.560 197.875 91.405 198.405 ;
        RECT 87.865 196.765 90.165 196.935 ;
        RECT 90.565 196.935 90.735 197.875 ;
        RECT 91.235 197.795 91.405 197.875 ;
        RECT 92.025 197.795 92.195 198.485 ;
        RECT 91.465 197.455 91.965 197.625 ;
        RECT 92.695 196.935 92.865 199.345 ;
        RECT 90.565 196.765 92.865 196.935 ;
        RECT 93.265 199.345 95.565 199.515 ;
        RECT 85.165 190.915 87.465 191.085 ;
        RECT 93.265 191.085 93.435 199.345 ;
        RECT 94.165 198.655 94.665 198.825 ;
        RECT 93.935 191.945 94.105 198.485 ;
        RECT 94.725 191.945 94.895 198.485 ;
        RECT 93.925 191.375 94.925 191.775 ;
        RECT 95.395 191.085 95.565 199.345 ;
        RECT 93.265 190.915 95.565 191.085 ;
        RECT 95.965 199.345 98.265 199.515 ;
        RECT 95.965 191.085 96.135 199.345 ;
        RECT 96.865 198.655 97.365 198.825 ;
        RECT 96.635 191.945 96.805 198.485 ;
        RECT 97.425 191.945 97.595 198.485 ;
        RECT 96.625 191.375 97.625 191.775 ;
        RECT 98.095 191.085 98.265 199.345 ;
        RECT 107.890 199.345 110.190 199.515 ;
        RECT 107.890 198.405 108.060 199.345 ;
        RECT 108.270 198.655 109.310 199.100 ;
        RECT 108.560 198.405 108.730 198.485 ;
        RECT 107.885 197.875 108.730 198.405 ;
        RECT 107.890 196.935 108.060 197.875 ;
        RECT 108.560 197.795 108.730 197.875 ;
        RECT 109.350 197.795 109.520 198.485 ;
        RECT 108.790 197.455 109.290 197.625 ;
        RECT 110.020 196.935 110.190 199.345 ;
        RECT 107.890 196.765 110.190 196.935 ;
        RECT 110.590 199.345 112.890 199.515 ;
        RECT 95.965 190.915 98.265 191.085 ;
        RECT 110.590 191.085 110.760 199.345 ;
        RECT 111.490 198.655 111.990 198.825 ;
        RECT 111.260 191.945 111.430 198.485 ;
        RECT 112.050 191.945 112.220 198.485 ;
        RECT 111.250 191.375 112.250 191.775 ;
        RECT 112.720 191.085 112.890 199.345 ;
        RECT 113.290 199.345 115.590 199.515 ;
        RECT 113.290 198.405 113.460 199.345 ;
        RECT 113.670 198.655 114.710 199.100 ;
        RECT 113.960 198.405 114.130 198.485 ;
        RECT 113.285 197.875 114.130 198.405 ;
        RECT 113.290 196.935 113.460 197.875 ;
        RECT 113.960 197.795 114.130 197.875 ;
        RECT 114.750 197.795 114.920 198.485 ;
        RECT 114.190 197.455 114.690 197.625 ;
        RECT 115.420 196.935 115.590 199.345 ;
        RECT 115.990 199.345 118.290 199.515 ;
        RECT 115.990 198.405 116.160 199.345 ;
        RECT 116.370 198.655 117.410 199.100 ;
        RECT 116.660 198.405 116.830 198.485 ;
        RECT 115.985 197.875 116.830 198.405 ;
        RECT 113.290 196.765 115.590 196.935 ;
        RECT 115.990 196.935 116.160 197.875 ;
        RECT 116.660 197.795 116.830 197.875 ;
        RECT 117.450 197.795 117.620 198.485 ;
        RECT 116.890 197.455 117.390 197.625 ;
        RECT 118.120 196.935 118.290 199.345 ;
        RECT 115.990 196.765 118.290 196.935 ;
        RECT 118.690 199.345 120.990 199.515 ;
        RECT 110.590 190.915 112.890 191.085 ;
        RECT 118.690 191.085 118.860 199.345 ;
        RECT 119.590 198.655 120.090 198.825 ;
        RECT 119.360 191.945 119.530 198.485 ;
        RECT 120.150 191.945 120.320 198.485 ;
        RECT 119.350 191.375 120.350 191.775 ;
        RECT 120.820 191.085 120.990 199.345 ;
        RECT 118.690 190.915 120.990 191.085 ;
        RECT 121.390 199.345 123.690 199.515 ;
        RECT 121.390 191.085 121.560 199.345 ;
        RECT 122.290 198.655 122.790 198.825 ;
        RECT 122.060 191.945 122.230 198.485 ;
        RECT 122.850 191.945 123.020 198.485 ;
        RECT 122.050 191.375 123.050 191.775 ;
        RECT 123.520 191.085 123.690 199.345 ;
        RECT 133.315 199.345 135.615 199.515 ;
        RECT 133.315 198.405 133.485 199.345 ;
        RECT 133.695 198.655 134.735 199.100 ;
        RECT 133.985 198.405 134.155 198.485 ;
        RECT 133.310 197.875 134.155 198.405 ;
        RECT 133.315 196.935 133.485 197.875 ;
        RECT 133.985 197.795 134.155 197.875 ;
        RECT 134.775 197.795 134.945 198.485 ;
        RECT 134.215 197.455 134.715 197.625 ;
        RECT 135.445 196.935 135.615 199.345 ;
        RECT 133.315 196.765 135.615 196.935 ;
        RECT 136.015 199.345 138.315 199.515 ;
        RECT 121.390 190.915 123.690 191.085 ;
        RECT 136.015 191.085 136.185 199.345 ;
        RECT 136.915 198.655 137.415 198.825 ;
        RECT 136.685 191.945 136.855 198.485 ;
        RECT 137.475 191.945 137.645 198.485 ;
        RECT 136.675 191.375 137.675 191.775 ;
        RECT 138.145 191.085 138.315 199.345 ;
        RECT 138.715 199.345 141.015 199.515 ;
        RECT 138.715 198.405 138.885 199.345 ;
        RECT 139.095 198.655 140.135 199.100 ;
        RECT 139.385 198.405 139.555 198.485 ;
        RECT 138.710 197.875 139.555 198.405 ;
        RECT 138.715 196.935 138.885 197.875 ;
        RECT 139.385 197.795 139.555 197.875 ;
        RECT 140.175 197.795 140.345 198.485 ;
        RECT 139.615 197.455 140.115 197.625 ;
        RECT 140.845 196.935 141.015 199.345 ;
        RECT 141.415 199.345 143.715 199.515 ;
        RECT 141.415 198.405 141.585 199.345 ;
        RECT 141.795 198.655 142.835 199.100 ;
        RECT 142.085 198.405 142.255 198.485 ;
        RECT 141.410 197.875 142.255 198.405 ;
        RECT 138.715 196.765 141.015 196.935 ;
        RECT 141.415 196.935 141.585 197.875 ;
        RECT 142.085 197.795 142.255 197.875 ;
        RECT 142.875 197.795 143.045 198.485 ;
        RECT 142.315 197.455 142.815 197.625 ;
        RECT 143.545 196.935 143.715 199.345 ;
        RECT 141.415 196.765 143.715 196.935 ;
        RECT 144.115 199.345 146.415 199.515 ;
        RECT 136.015 190.915 138.315 191.085 ;
        RECT 144.115 191.085 144.285 199.345 ;
        RECT 145.015 198.655 145.515 198.825 ;
        RECT 144.785 191.945 144.955 198.485 ;
        RECT 145.575 191.945 145.745 198.485 ;
        RECT 144.775 191.375 145.775 191.775 ;
        RECT 146.245 191.085 146.415 199.345 ;
        RECT 144.115 190.915 146.415 191.085 ;
        RECT 146.815 199.345 149.115 199.515 ;
        RECT 146.815 191.085 146.985 199.345 ;
        RECT 147.715 198.655 148.215 198.825 ;
        RECT 147.485 191.945 147.655 198.485 ;
        RECT 148.275 191.945 148.445 198.485 ;
        RECT 147.475 191.375 148.475 191.775 ;
        RECT 148.945 191.085 149.115 199.345 ;
        RECT 146.815 190.915 149.115 191.085 ;
        RECT 8.890 189.860 11.190 190.030 ;
        RECT 6.190 180.860 8.490 181.030 ;
        RECT 6.190 179.925 6.360 180.860 ;
        RECT 7.090 180.170 7.590 180.340 ;
        RECT 6.860 179.925 7.030 179.955 ;
        RECT 6.135 178.945 7.030 179.925 ;
        RECT 6.190 178.010 6.360 178.945 ;
        RECT 6.860 178.915 7.030 178.945 ;
        RECT 7.650 178.915 7.820 179.955 ;
        RECT 6.675 178.530 7.590 178.700 ;
        RECT 6.675 178.325 7.510 178.530 ;
        RECT 8.320 178.010 8.490 180.860 ;
        RECT 6.190 177.840 8.490 178.010 ;
        RECT 8.890 178.010 9.060 189.860 ;
        RECT 9.550 189.150 10.550 189.600 ;
        RECT 9.560 178.915 9.730 188.955 ;
        RECT 10.350 178.915 10.520 188.955 ;
        RECT 9.790 178.530 10.290 178.700 ;
        RECT 11.020 178.010 11.190 189.860 ;
        RECT 16.990 189.860 19.290 190.030 ;
        RECT 11.590 180.860 13.890 181.030 ;
        RECT 11.590 179.925 11.760 180.860 ;
        RECT 12.490 180.170 12.990 180.340 ;
        RECT 12.260 179.925 12.430 179.955 ;
        RECT 11.535 178.945 12.430 179.925 ;
        RECT 8.890 177.840 11.190 178.010 ;
        RECT 11.590 178.010 11.760 178.945 ;
        RECT 12.260 178.915 12.430 178.945 ;
        RECT 13.050 178.915 13.220 179.955 ;
        RECT 12.075 178.530 12.990 178.700 ;
        RECT 12.075 178.325 12.910 178.530 ;
        RECT 13.720 178.010 13.890 180.860 ;
        RECT 14.290 180.860 16.590 181.030 ;
        RECT 14.290 179.925 14.460 180.860 ;
        RECT 15.190 180.170 15.690 180.340 ;
        RECT 14.960 179.925 15.130 179.955 ;
        RECT 14.235 178.945 15.130 179.925 ;
        RECT 11.590 177.840 13.890 178.010 ;
        RECT 14.290 178.010 14.460 178.945 ;
        RECT 14.960 178.915 15.130 178.945 ;
        RECT 15.750 178.915 15.920 179.955 ;
        RECT 14.775 178.530 15.690 178.700 ;
        RECT 14.775 178.325 15.610 178.530 ;
        RECT 16.420 178.010 16.590 180.860 ;
        RECT 14.290 177.840 16.590 178.010 ;
        RECT 16.990 178.010 17.160 189.860 ;
        RECT 17.650 189.150 18.650 189.600 ;
        RECT 17.660 178.915 17.830 188.955 ;
        RECT 18.450 178.915 18.620 188.955 ;
        RECT 17.890 178.530 18.390 178.700 ;
        RECT 19.120 178.010 19.290 189.860 ;
        RECT 16.990 177.840 19.290 178.010 ;
        RECT 19.690 189.860 21.990 190.030 ;
        RECT 19.690 178.010 19.860 189.860 ;
        RECT 20.350 189.150 21.350 189.600 ;
        RECT 20.360 178.915 20.530 188.955 ;
        RECT 21.150 178.915 21.320 188.955 ;
        RECT 20.590 178.530 21.090 178.700 ;
        RECT 21.820 178.010 21.990 189.860 ;
        RECT 34.315 189.860 36.615 190.030 ;
        RECT 31.615 180.860 33.915 181.030 ;
        RECT 31.615 179.925 31.785 180.860 ;
        RECT 32.515 180.170 33.015 180.340 ;
        RECT 32.285 179.925 32.455 179.955 ;
        RECT 31.560 178.945 32.455 179.925 ;
        RECT 19.690 177.840 21.990 178.010 ;
        RECT 31.615 178.010 31.785 178.945 ;
        RECT 32.285 178.915 32.455 178.945 ;
        RECT 33.075 178.915 33.245 179.955 ;
        RECT 32.100 178.530 33.015 178.700 ;
        RECT 32.100 178.325 32.935 178.530 ;
        RECT 33.745 178.010 33.915 180.860 ;
        RECT 31.615 177.840 33.915 178.010 ;
        RECT 34.315 178.010 34.485 189.860 ;
        RECT 34.975 189.150 35.975 189.600 ;
        RECT 34.985 178.915 35.155 188.955 ;
        RECT 35.775 178.915 35.945 188.955 ;
        RECT 35.215 178.530 35.715 178.700 ;
        RECT 36.445 178.010 36.615 189.860 ;
        RECT 42.415 189.860 44.715 190.030 ;
        RECT 37.015 180.860 39.315 181.030 ;
        RECT 37.015 179.925 37.185 180.860 ;
        RECT 37.915 180.170 38.415 180.340 ;
        RECT 37.685 179.925 37.855 179.955 ;
        RECT 36.960 178.945 37.855 179.925 ;
        RECT 34.315 177.840 36.615 178.010 ;
        RECT 37.015 178.010 37.185 178.945 ;
        RECT 37.685 178.915 37.855 178.945 ;
        RECT 38.475 178.915 38.645 179.955 ;
        RECT 37.500 178.530 38.415 178.700 ;
        RECT 37.500 178.325 38.335 178.530 ;
        RECT 39.145 178.010 39.315 180.860 ;
        RECT 39.715 180.860 42.015 181.030 ;
        RECT 39.715 179.925 39.885 180.860 ;
        RECT 40.615 180.170 41.115 180.340 ;
        RECT 40.385 179.925 40.555 179.955 ;
        RECT 39.660 178.945 40.555 179.925 ;
        RECT 37.015 177.840 39.315 178.010 ;
        RECT 39.715 178.010 39.885 178.945 ;
        RECT 40.385 178.915 40.555 178.945 ;
        RECT 41.175 178.915 41.345 179.955 ;
        RECT 40.200 178.530 41.115 178.700 ;
        RECT 40.200 178.325 41.035 178.530 ;
        RECT 41.845 178.010 42.015 180.860 ;
        RECT 39.715 177.840 42.015 178.010 ;
        RECT 42.415 178.010 42.585 189.860 ;
        RECT 43.075 189.150 44.075 189.600 ;
        RECT 43.085 178.915 43.255 188.955 ;
        RECT 43.875 178.915 44.045 188.955 ;
        RECT 43.315 178.530 43.815 178.700 ;
        RECT 44.545 178.010 44.715 189.860 ;
        RECT 42.415 177.840 44.715 178.010 ;
        RECT 45.115 189.860 47.415 190.030 ;
        RECT 45.115 178.010 45.285 189.860 ;
        RECT 45.775 189.150 46.775 189.600 ;
        RECT 45.785 178.915 45.955 188.955 ;
        RECT 46.575 178.915 46.745 188.955 ;
        RECT 46.015 178.530 46.515 178.700 ;
        RECT 47.245 178.010 47.415 189.860 ;
        RECT 59.740 189.860 62.040 190.030 ;
        RECT 57.040 180.860 59.340 181.030 ;
        RECT 57.040 179.925 57.210 180.860 ;
        RECT 57.940 180.170 58.440 180.340 ;
        RECT 57.710 179.925 57.880 179.955 ;
        RECT 56.985 178.945 57.880 179.925 ;
        RECT 45.115 177.840 47.415 178.010 ;
        RECT 57.040 178.010 57.210 178.945 ;
        RECT 57.710 178.915 57.880 178.945 ;
        RECT 58.500 178.915 58.670 179.955 ;
        RECT 57.525 178.530 58.440 178.700 ;
        RECT 57.525 178.325 58.360 178.530 ;
        RECT 59.170 178.010 59.340 180.860 ;
        RECT 57.040 177.840 59.340 178.010 ;
        RECT 59.740 178.010 59.910 189.860 ;
        RECT 60.400 189.150 61.400 189.600 ;
        RECT 60.410 178.915 60.580 188.955 ;
        RECT 61.200 178.915 61.370 188.955 ;
        RECT 60.640 178.530 61.140 178.700 ;
        RECT 61.870 178.010 62.040 189.860 ;
        RECT 67.840 189.860 70.140 190.030 ;
        RECT 62.440 180.860 64.740 181.030 ;
        RECT 62.440 179.925 62.610 180.860 ;
        RECT 63.340 180.170 63.840 180.340 ;
        RECT 63.110 179.925 63.280 179.955 ;
        RECT 62.385 178.945 63.280 179.925 ;
        RECT 59.740 177.840 62.040 178.010 ;
        RECT 62.440 178.010 62.610 178.945 ;
        RECT 63.110 178.915 63.280 178.945 ;
        RECT 63.900 178.915 64.070 179.955 ;
        RECT 62.925 178.530 63.840 178.700 ;
        RECT 62.925 178.325 63.760 178.530 ;
        RECT 64.570 178.010 64.740 180.860 ;
        RECT 65.140 180.860 67.440 181.030 ;
        RECT 65.140 179.925 65.310 180.860 ;
        RECT 66.040 180.170 66.540 180.340 ;
        RECT 65.810 179.925 65.980 179.955 ;
        RECT 65.085 178.945 65.980 179.925 ;
        RECT 62.440 177.840 64.740 178.010 ;
        RECT 65.140 178.010 65.310 178.945 ;
        RECT 65.810 178.915 65.980 178.945 ;
        RECT 66.600 178.915 66.770 179.955 ;
        RECT 65.625 178.530 66.540 178.700 ;
        RECT 65.625 178.325 66.460 178.530 ;
        RECT 67.270 178.010 67.440 180.860 ;
        RECT 65.140 177.840 67.440 178.010 ;
        RECT 67.840 178.010 68.010 189.860 ;
        RECT 68.500 189.150 69.500 189.600 ;
        RECT 68.510 178.915 68.680 188.955 ;
        RECT 69.300 178.915 69.470 188.955 ;
        RECT 68.740 178.530 69.240 178.700 ;
        RECT 69.970 178.010 70.140 189.860 ;
        RECT 67.840 177.840 70.140 178.010 ;
        RECT 70.540 189.860 72.840 190.030 ;
        RECT 70.540 178.010 70.710 189.860 ;
        RECT 71.200 189.150 72.200 189.600 ;
        RECT 71.210 178.915 71.380 188.955 ;
        RECT 72.000 178.915 72.170 188.955 ;
        RECT 71.440 178.530 71.940 178.700 ;
        RECT 72.670 178.010 72.840 189.860 ;
        RECT 85.165 189.860 87.465 190.030 ;
        RECT 82.465 180.860 84.765 181.030 ;
        RECT 82.465 179.925 82.635 180.860 ;
        RECT 83.365 180.170 83.865 180.340 ;
        RECT 83.135 179.925 83.305 179.955 ;
        RECT 82.410 178.945 83.305 179.925 ;
        RECT 70.540 177.840 72.840 178.010 ;
        RECT 82.465 178.010 82.635 178.945 ;
        RECT 83.135 178.915 83.305 178.945 ;
        RECT 83.925 178.915 84.095 179.955 ;
        RECT 82.950 178.530 83.865 178.700 ;
        RECT 82.950 178.325 83.785 178.530 ;
        RECT 84.595 178.010 84.765 180.860 ;
        RECT 82.465 177.840 84.765 178.010 ;
        RECT 85.165 178.010 85.335 189.860 ;
        RECT 85.825 189.150 86.825 189.600 ;
        RECT 85.835 178.915 86.005 188.955 ;
        RECT 86.625 178.915 86.795 188.955 ;
        RECT 86.065 178.530 86.565 178.700 ;
        RECT 87.295 178.010 87.465 189.860 ;
        RECT 93.265 189.860 95.565 190.030 ;
        RECT 87.865 180.860 90.165 181.030 ;
        RECT 87.865 179.925 88.035 180.860 ;
        RECT 88.765 180.170 89.265 180.340 ;
        RECT 88.535 179.925 88.705 179.955 ;
        RECT 87.810 178.945 88.705 179.925 ;
        RECT 85.165 177.840 87.465 178.010 ;
        RECT 87.865 178.010 88.035 178.945 ;
        RECT 88.535 178.915 88.705 178.945 ;
        RECT 89.325 178.915 89.495 179.955 ;
        RECT 88.350 178.530 89.265 178.700 ;
        RECT 88.350 178.325 89.185 178.530 ;
        RECT 89.995 178.010 90.165 180.860 ;
        RECT 90.565 180.860 92.865 181.030 ;
        RECT 90.565 179.925 90.735 180.860 ;
        RECT 91.465 180.170 91.965 180.340 ;
        RECT 91.235 179.925 91.405 179.955 ;
        RECT 90.510 178.945 91.405 179.925 ;
        RECT 87.865 177.840 90.165 178.010 ;
        RECT 90.565 178.010 90.735 178.945 ;
        RECT 91.235 178.915 91.405 178.945 ;
        RECT 92.025 178.915 92.195 179.955 ;
        RECT 91.050 178.530 91.965 178.700 ;
        RECT 91.050 178.325 91.885 178.530 ;
        RECT 92.695 178.010 92.865 180.860 ;
        RECT 90.565 177.840 92.865 178.010 ;
        RECT 93.265 178.010 93.435 189.860 ;
        RECT 93.925 189.150 94.925 189.600 ;
        RECT 93.935 178.915 94.105 188.955 ;
        RECT 94.725 178.915 94.895 188.955 ;
        RECT 94.165 178.530 94.665 178.700 ;
        RECT 95.395 178.010 95.565 189.860 ;
        RECT 93.265 177.840 95.565 178.010 ;
        RECT 95.965 189.860 98.265 190.030 ;
        RECT 95.965 178.010 96.135 189.860 ;
        RECT 96.625 189.150 97.625 189.600 ;
        RECT 96.635 178.915 96.805 188.955 ;
        RECT 97.425 178.915 97.595 188.955 ;
        RECT 96.865 178.530 97.365 178.700 ;
        RECT 98.095 178.010 98.265 189.860 ;
        RECT 110.590 189.860 112.890 190.030 ;
        RECT 107.890 180.860 110.190 181.030 ;
        RECT 107.890 179.925 108.060 180.860 ;
        RECT 108.790 180.170 109.290 180.340 ;
        RECT 108.560 179.925 108.730 179.955 ;
        RECT 107.835 178.945 108.730 179.925 ;
        RECT 95.965 177.840 98.265 178.010 ;
        RECT 107.890 178.010 108.060 178.945 ;
        RECT 108.560 178.915 108.730 178.945 ;
        RECT 109.350 178.915 109.520 179.955 ;
        RECT 108.375 178.530 109.290 178.700 ;
        RECT 108.375 178.325 109.210 178.530 ;
        RECT 110.020 178.010 110.190 180.860 ;
        RECT 107.890 177.840 110.190 178.010 ;
        RECT 110.590 178.010 110.760 189.860 ;
        RECT 111.250 189.150 112.250 189.600 ;
        RECT 111.260 178.915 111.430 188.955 ;
        RECT 112.050 178.915 112.220 188.955 ;
        RECT 111.490 178.530 111.990 178.700 ;
        RECT 112.720 178.010 112.890 189.860 ;
        RECT 118.690 189.860 120.990 190.030 ;
        RECT 113.290 180.860 115.590 181.030 ;
        RECT 113.290 179.925 113.460 180.860 ;
        RECT 114.190 180.170 114.690 180.340 ;
        RECT 113.960 179.925 114.130 179.955 ;
        RECT 113.235 178.945 114.130 179.925 ;
        RECT 110.590 177.840 112.890 178.010 ;
        RECT 113.290 178.010 113.460 178.945 ;
        RECT 113.960 178.915 114.130 178.945 ;
        RECT 114.750 178.915 114.920 179.955 ;
        RECT 113.775 178.530 114.690 178.700 ;
        RECT 113.775 178.325 114.610 178.530 ;
        RECT 115.420 178.010 115.590 180.860 ;
        RECT 115.990 180.860 118.290 181.030 ;
        RECT 115.990 179.925 116.160 180.860 ;
        RECT 116.890 180.170 117.390 180.340 ;
        RECT 116.660 179.925 116.830 179.955 ;
        RECT 115.935 178.945 116.830 179.925 ;
        RECT 113.290 177.840 115.590 178.010 ;
        RECT 115.990 178.010 116.160 178.945 ;
        RECT 116.660 178.915 116.830 178.945 ;
        RECT 117.450 178.915 117.620 179.955 ;
        RECT 116.475 178.530 117.390 178.700 ;
        RECT 116.475 178.325 117.310 178.530 ;
        RECT 118.120 178.010 118.290 180.860 ;
        RECT 115.990 177.840 118.290 178.010 ;
        RECT 118.690 178.010 118.860 189.860 ;
        RECT 119.350 189.150 120.350 189.600 ;
        RECT 119.360 178.915 119.530 188.955 ;
        RECT 120.150 178.915 120.320 188.955 ;
        RECT 119.590 178.530 120.090 178.700 ;
        RECT 120.820 178.010 120.990 189.860 ;
        RECT 118.690 177.840 120.990 178.010 ;
        RECT 121.390 189.860 123.690 190.030 ;
        RECT 121.390 178.010 121.560 189.860 ;
        RECT 122.050 189.150 123.050 189.600 ;
        RECT 122.060 178.915 122.230 188.955 ;
        RECT 122.850 178.915 123.020 188.955 ;
        RECT 122.290 178.530 122.790 178.700 ;
        RECT 123.520 178.010 123.690 189.860 ;
        RECT 136.015 189.860 138.315 190.030 ;
        RECT 133.315 180.860 135.615 181.030 ;
        RECT 133.315 179.925 133.485 180.860 ;
        RECT 134.215 180.170 134.715 180.340 ;
        RECT 133.985 179.925 134.155 179.955 ;
        RECT 133.260 178.945 134.155 179.925 ;
        RECT 121.390 177.840 123.690 178.010 ;
        RECT 133.315 178.010 133.485 178.945 ;
        RECT 133.985 178.915 134.155 178.945 ;
        RECT 134.775 178.915 134.945 179.955 ;
        RECT 133.800 178.530 134.715 178.700 ;
        RECT 133.800 178.325 134.635 178.530 ;
        RECT 135.445 178.010 135.615 180.860 ;
        RECT 133.315 177.840 135.615 178.010 ;
        RECT 136.015 178.010 136.185 189.860 ;
        RECT 136.675 189.150 137.675 189.600 ;
        RECT 136.685 178.915 136.855 188.955 ;
        RECT 137.475 178.915 137.645 188.955 ;
        RECT 136.915 178.530 137.415 178.700 ;
        RECT 138.145 178.010 138.315 189.860 ;
        RECT 144.115 189.860 146.415 190.030 ;
        RECT 138.715 180.860 141.015 181.030 ;
        RECT 138.715 179.925 138.885 180.860 ;
        RECT 139.615 180.170 140.115 180.340 ;
        RECT 139.385 179.925 139.555 179.955 ;
        RECT 138.660 178.945 139.555 179.925 ;
        RECT 136.015 177.840 138.315 178.010 ;
        RECT 138.715 178.010 138.885 178.945 ;
        RECT 139.385 178.915 139.555 178.945 ;
        RECT 140.175 178.915 140.345 179.955 ;
        RECT 139.200 178.530 140.115 178.700 ;
        RECT 139.200 178.325 140.035 178.530 ;
        RECT 140.845 178.010 141.015 180.860 ;
        RECT 141.415 180.860 143.715 181.030 ;
        RECT 141.415 179.925 141.585 180.860 ;
        RECT 142.315 180.170 142.815 180.340 ;
        RECT 142.085 179.925 142.255 179.955 ;
        RECT 141.360 178.945 142.255 179.925 ;
        RECT 138.715 177.840 141.015 178.010 ;
        RECT 141.415 178.010 141.585 178.945 ;
        RECT 142.085 178.915 142.255 178.945 ;
        RECT 142.875 178.915 143.045 179.955 ;
        RECT 141.900 178.530 142.815 178.700 ;
        RECT 141.900 178.325 142.735 178.530 ;
        RECT 143.545 178.010 143.715 180.860 ;
        RECT 141.415 177.840 143.715 178.010 ;
        RECT 144.115 178.010 144.285 189.860 ;
        RECT 144.775 189.150 145.775 189.600 ;
        RECT 144.785 178.915 144.955 188.955 ;
        RECT 145.575 178.915 145.745 188.955 ;
        RECT 145.015 178.530 145.515 178.700 ;
        RECT 146.245 178.010 146.415 189.860 ;
        RECT 144.115 177.840 146.415 178.010 ;
        RECT 146.815 189.860 149.115 190.030 ;
        RECT 146.815 178.010 146.985 189.860 ;
        RECT 147.475 189.150 148.475 189.600 ;
        RECT 147.485 178.915 147.655 188.955 ;
        RECT 148.275 178.915 148.445 188.955 ;
        RECT 147.715 178.530 148.215 178.700 ;
        RECT 148.945 178.010 149.115 189.860 ;
        RECT 146.815 177.840 149.115 178.010 ;
        RECT 6.190 176.770 8.490 176.940 ;
        RECT 6.190 175.830 6.360 176.770 ;
        RECT 6.570 176.080 7.610 176.525 ;
        RECT 6.860 175.830 7.030 175.910 ;
        RECT 6.185 175.300 7.030 175.830 ;
        RECT 6.190 174.360 6.360 175.300 ;
        RECT 6.860 175.220 7.030 175.300 ;
        RECT 7.650 175.220 7.820 175.910 ;
        RECT 7.090 174.880 7.590 175.050 ;
        RECT 8.320 174.360 8.490 176.770 ;
        RECT 6.190 174.190 8.490 174.360 ;
        RECT 8.890 176.770 11.190 176.940 ;
        RECT 8.890 168.510 9.060 176.770 ;
        RECT 9.790 176.080 10.290 176.250 ;
        RECT 9.560 169.370 9.730 175.910 ;
        RECT 10.350 169.370 10.520 175.910 ;
        RECT 9.550 168.800 10.550 169.200 ;
        RECT 11.020 168.510 11.190 176.770 ;
        RECT 11.590 176.770 13.890 176.940 ;
        RECT 11.590 175.830 11.760 176.770 ;
        RECT 11.970 176.080 13.010 176.525 ;
        RECT 12.260 175.830 12.430 175.910 ;
        RECT 11.585 175.300 12.430 175.830 ;
        RECT 11.590 174.360 11.760 175.300 ;
        RECT 12.260 175.220 12.430 175.300 ;
        RECT 13.050 175.220 13.220 175.910 ;
        RECT 12.490 174.880 12.990 175.050 ;
        RECT 13.720 174.360 13.890 176.770 ;
        RECT 14.290 176.770 16.590 176.940 ;
        RECT 14.290 175.830 14.460 176.770 ;
        RECT 14.670 176.080 15.710 176.525 ;
        RECT 14.960 175.830 15.130 175.910 ;
        RECT 14.285 175.300 15.130 175.830 ;
        RECT 11.590 174.190 13.890 174.360 ;
        RECT 14.290 174.360 14.460 175.300 ;
        RECT 14.960 175.220 15.130 175.300 ;
        RECT 15.750 175.220 15.920 175.910 ;
        RECT 15.190 174.880 15.690 175.050 ;
        RECT 16.420 174.360 16.590 176.770 ;
        RECT 14.290 174.190 16.590 174.360 ;
        RECT 16.990 176.770 19.290 176.940 ;
        RECT 8.890 168.340 11.190 168.510 ;
        RECT 16.990 168.510 17.160 176.770 ;
        RECT 17.890 176.080 18.390 176.250 ;
        RECT 17.660 169.370 17.830 175.910 ;
        RECT 18.450 169.370 18.620 175.910 ;
        RECT 17.650 168.800 18.650 169.200 ;
        RECT 19.120 168.510 19.290 176.770 ;
        RECT 16.990 168.340 19.290 168.510 ;
        RECT 19.690 176.770 21.990 176.940 ;
        RECT 19.690 168.510 19.860 176.770 ;
        RECT 20.590 176.080 21.090 176.250 ;
        RECT 20.360 169.370 20.530 175.910 ;
        RECT 21.150 169.370 21.320 175.910 ;
        RECT 20.350 168.800 21.350 169.200 ;
        RECT 21.820 168.510 21.990 176.770 ;
        RECT 31.615 176.770 33.915 176.940 ;
        RECT 31.615 175.830 31.785 176.770 ;
        RECT 31.995 176.080 33.035 176.525 ;
        RECT 32.285 175.830 32.455 175.910 ;
        RECT 31.610 175.300 32.455 175.830 ;
        RECT 31.615 174.360 31.785 175.300 ;
        RECT 32.285 175.220 32.455 175.300 ;
        RECT 33.075 175.220 33.245 175.910 ;
        RECT 32.515 174.880 33.015 175.050 ;
        RECT 33.745 174.360 33.915 176.770 ;
        RECT 31.615 174.190 33.915 174.360 ;
        RECT 34.315 176.770 36.615 176.940 ;
        RECT 19.690 168.340 21.990 168.510 ;
        RECT 34.315 168.510 34.485 176.770 ;
        RECT 35.215 176.080 35.715 176.250 ;
        RECT 34.985 169.370 35.155 175.910 ;
        RECT 35.775 169.370 35.945 175.910 ;
        RECT 34.975 168.800 35.975 169.200 ;
        RECT 36.445 168.510 36.615 176.770 ;
        RECT 37.015 176.770 39.315 176.940 ;
        RECT 37.015 175.830 37.185 176.770 ;
        RECT 37.395 176.080 38.435 176.525 ;
        RECT 37.685 175.830 37.855 175.910 ;
        RECT 37.010 175.300 37.855 175.830 ;
        RECT 37.015 174.360 37.185 175.300 ;
        RECT 37.685 175.220 37.855 175.300 ;
        RECT 38.475 175.220 38.645 175.910 ;
        RECT 37.915 174.880 38.415 175.050 ;
        RECT 39.145 174.360 39.315 176.770 ;
        RECT 39.715 176.770 42.015 176.940 ;
        RECT 39.715 175.830 39.885 176.770 ;
        RECT 40.095 176.080 41.135 176.525 ;
        RECT 40.385 175.830 40.555 175.910 ;
        RECT 39.710 175.300 40.555 175.830 ;
        RECT 37.015 174.190 39.315 174.360 ;
        RECT 39.715 174.360 39.885 175.300 ;
        RECT 40.385 175.220 40.555 175.300 ;
        RECT 41.175 175.220 41.345 175.910 ;
        RECT 40.615 174.880 41.115 175.050 ;
        RECT 41.845 174.360 42.015 176.770 ;
        RECT 39.715 174.190 42.015 174.360 ;
        RECT 42.415 176.770 44.715 176.940 ;
        RECT 34.315 168.340 36.615 168.510 ;
        RECT 42.415 168.510 42.585 176.770 ;
        RECT 43.315 176.080 43.815 176.250 ;
        RECT 43.085 169.370 43.255 175.910 ;
        RECT 43.875 169.370 44.045 175.910 ;
        RECT 43.075 168.800 44.075 169.200 ;
        RECT 44.545 168.510 44.715 176.770 ;
        RECT 42.415 168.340 44.715 168.510 ;
        RECT 45.115 176.770 47.415 176.940 ;
        RECT 45.115 168.510 45.285 176.770 ;
        RECT 46.015 176.080 46.515 176.250 ;
        RECT 45.785 169.370 45.955 175.910 ;
        RECT 46.575 169.370 46.745 175.910 ;
        RECT 45.775 168.800 46.775 169.200 ;
        RECT 47.245 168.510 47.415 176.770 ;
        RECT 57.040 176.770 59.340 176.940 ;
        RECT 57.040 175.830 57.210 176.770 ;
        RECT 57.420 176.080 58.460 176.525 ;
        RECT 57.710 175.830 57.880 175.910 ;
        RECT 57.035 175.300 57.880 175.830 ;
        RECT 57.040 174.360 57.210 175.300 ;
        RECT 57.710 175.220 57.880 175.300 ;
        RECT 58.500 175.220 58.670 175.910 ;
        RECT 57.940 174.880 58.440 175.050 ;
        RECT 59.170 174.360 59.340 176.770 ;
        RECT 57.040 174.190 59.340 174.360 ;
        RECT 59.740 176.770 62.040 176.940 ;
        RECT 45.115 168.340 47.415 168.510 ;
        RECT 59.740 168.510 59.910 176.770 ;
        RECT 60.640 176.080 61.140 176.250 ;
        RECT 60.410 169.370 60.580 175.910 ;
        RECT 61.200 169.370 61.370 175.910 ;
        RECT 60.400 168.800 61.400 169.200 ;
        RECT 61.870 168.510 62.040 176.770 ;
        RECT 62.440 176.770 64.740 176.940 ;
        RECT 62.440 175.830 62.610 176.770 ;
        RECT 62.820 176.080 63.860 176.525 ;
        RECT 63.110 175.830 63.280 175.910 ;
        RECT 62.435 175.300 63.280 175.830 ;
        RECT 62.440 174.360 62.610 175.300 ;
        RECT 63.110 175.220 63.280 175.300 ;
        RECT 63.900 175.220 64.070 175.910 ;
        RECT 63.340 174.880 63.840 175.050 ;
        RECT 64.570 174.360 64.740 176.770 ;
        RECT 65.140 176.770 67.440 176.940 ;
        RECT 65.140 175.830 65.310 176.770 ;
        RECT 65.520 176.080 66.560 176.525 ;
        RECT 65.810 175.830 65.980 175.910 ;
        RECT 65.135 175.300 65.980 175.830 ;
        RECT 62.440 174.190 64.740 174.360 ;
        RECT 65.140 174.360 65.310 175.300 ;
        RECT 65.810 175.220 65.980 175.300 ;
        RECT 66.600 175.220 66.770 175.910 ;
        RECT 66.040 174.880 66.540 175.050 ;
        RECT 67.270 174.360 67.440 176.770 ;
        RECT 65.140 174.190 67.440 174.360 ;
        RECT 67.840 176.770 70.140 176.940 ;
        RECT 59.740 168.340 62.040 168.510 ;
        RECT 67.840 168.510 68.010 176.770 ;
        RECT 68.740 176.080 69.240 176.250 ;
        RECT 68.510 169.370 68.680 175.910 ;
        RECT 69.300 169.370 69.470 175.910 ;
        RECT 68.500 168.800 69.500 169.200 ;
        RECT 69.970 168.510 70.140 176.770 ;
        RECT 67.840 168.340 70.140 168.510 ;
        RECT 70.540 176.770 72.840 176.940 ;
        RECT 70.540 168.510 70.710 176.770 ;
        RECT 71.440 176.080 71.940 176.250 ;
        RECT 71.210 169.370 71.380 175.910 ;
        RECT 72.000 169.370 72.170 175.910 ;
        RECT 71.200 168.800 72.200 169.200 ;
        RECT 72.670 168.510 72.840 176.770 ;
        RECT 82.465 176.770 84.765 176.940 ;
        RECT 82.465 175.830 82.635 176.770 ;
        RECT 82.845 176.080 83.885 176.525 ;
        RECT 83.135 175.830 83.305 175.910 ;
        RECT 82.460 175.300 83.305 175.830 ;
        RECT 82.465 174.360 82.635 175.300 ;
        RECT 83.135 175.220 83.305 175.300 ;
        RECT 83.925 175.220 84.095 175.910 ;
        RECT 83.365 174.880 83.865 175.050 ;
        RECT 84.595 174.360 84.765 176.770 ;
        RECT 82.465 174.190 84.765 174.360 ;
        RECT 85.165 176.770 87.465 176.940 ;
        RECT 70.540 168.340 72.840 168.510 ;
        RECT 85.165 168.510 85.335 176.770 ;
        RECT 86.065 176.080 86.565 176.250 ;
        RECT 85.835 169.370 86.005 175.910 ;
        RECT 86.625 169.370 86.795 175.910 ;
        RECT 85.825 168.800 86.825 169.200 ;
        RECT 87.295 168.510 87.465 176.770 ;
        RECT 87.865 176.770 90.165 176.940 ;
        RECT 87.865 175.830 88.035 176.770 ;
        RECT 88.245 176.080 89.285 176.525 ;
        RECT 88.535 175.830 88.705 175.910 ;
        RECT 87.860 175.300 88.705 175.830 ;
        RECT 87.865 174.360 88.035 175.300 ;
        RECT 88.535 175.220 88.705 175.300 ;
        RECT 89.325 175.220 89.495 175.910 ;
        RECT 88.765 174.880 89.265 175.050 ;
        RECT 89.995 174.360 90.165 176.770 ;
        RECT 90.565 176.770 92.865 176.940 ;
        RECT 90.565 175.830 90.735 176.770 ;
        RECT 90.945 176.080 91.985 176.525 ;
        RECT 91.235 175.830 91.405 175.910 ;
        RECT 90.560 175.300 91.405 175.830 ;
        RECT 87.865 174.190 90.165 174.360 ;
        RECT 90.565 174.360 90.735 175.300 ;
        RECT 91.235 175.220 91.405 175.300 ;
        RECT 92.025 175.220 92.195 175.910 ;
        RECT 91.465 174.880 91.965 175.050 ;
        RECT 92.695 174.360 92.865 176.770 ;
        RECT 90.565 174.190 92.865 174.360 ;
        RECT 93.265 176.770 95.565 176.940 ;
        RECT 85.165 168.340 87.465 168.510 ;
        RECT 93.265 168.510 93.435 176.770 ;
        RECT 94.165 176.080 94.665 176.250 ;
        RECT 93.935 169.370 94.105 175.910 ;
        RECT 94.725 169.370 94.895 175.910 ;
        RECT 93.925 168.800 94.925 169.200 ;
        RECT 95.395 168.510 95.565 176.770 ;
        RECT 93.265 168.340 95.565 168.510 ;
        RECT 95.965 176.770 98.265 176.940 ;
        RECT 95.965 168.510 96.135 176.770 ;
        RECT 96.865 176.080 97.365 176.250 ;
        RECT 96.635 169.370 96.805 175.910 ;
        RECT 97.425 169.370 97.595 175.910 ;
        RECT 96.625 168.800 97.625 169.200 ;
        RECT 98.095 168.510 98.265 176.770 ;
        RECT 107.890 176.770 110.190 176.940 ;
        RECT 107.890 175.830 108.060 176.770 ;
        RECT 108.270 176.080 109.310 176.525 ;
        RECT 108.560 175.830 108.730 175.910 ;
        RECT 107.885 175.300 108.730 175.830 ;
        RECT 107.890 174.360 108.060 175.300 ;
        RECT 108.560 175.220 108.730 175.300 ;
        RECT 109.350 175.220 109.520 175.910 ;
        RECT 108.790 174.880 109.290 175.050 ;
        RECT 110.020 174.360 110.190 176.770 ;
        RECT 107.890 174.190 110.190 174.360 ;
        RECT 110.590 176.770 112.890 176.940 ;
        RECT 95.965 168.340 98.265 168.510 ;
        RECT 110.590 168.510 110.760 176.770 ;
        RECT 111.490 176.080 111.990 176.250 ;
        RECT 111.260 169.370 111.430 175.910 ;
        RECT 112.050 169.370 112.220 175.910 ;
        RECT 111.250 168.800 112.250 169.200 ;
        RECT 112.720 168.510 112.890 176.770 ;
        RECT 113.290 176.770 115.590 176.940 ;
        RECT 113.290 175.830 113.460 176.770 ;
        RECT 113.670 176.080 114.710 176.525 ;
        RECT 113.960 175.830 114.130 175.910 ;
        RECT 113.285 175.300 114.130 175.830 ;
        RECT 113.290 174.360 113.460 175.300 ;
        RECT 113.960 175.220 114.130 175.300 ;
        RECT 114.750 175.220 114.920 175.910 ;
        RECT 114.190 174.880 114.690 175.050 ;
        RECT 115.420 174.360 115.590 176.770 ;
        RECT 115.990 176.770 118.290 176.940 ;
        RECT 115.990 175.830 116.160 176.770 ;
        RECT 116.370 176.080 117.410 176.525 ;
        RECT 116.660 175.830 116.830 175.910 ;
        RECT 115.985 175.300 116.830 175.830 ;
        RECT 113.290 174.190 115.590 174.360 ;
        RECT 115.990 174.360 116.160 175.300 ;
        RECT 116.660 175.220 116.830 175.300 ;
        RECT 117.450 175.220 117.620 175.910 ;
        RECT 116.890 174.880 117.390 175.050 ;
        RECT 118.120 174.360 118.290 176.770 ;
        RECT 115.990 174.190 118.290 174.360 ;
        RECT 118.690 176.770 120.990 176.940 ;
        RECT 110.590 168.340 112.890 168.510 ;
        RECT 118.690 168.510 118.860 176.770 ;
        RECT 119.590 176.080 120.090 176.250 ;
        RECT 119.360 169.370 119.530 175.910 ;
        RECT 120.150 169.370 120.320 175.910 ;
        RECT 119.350 168.800 120.350 169.200 ;
        RECT 120.820 168.510 120.990 176.770 ;
        RECT 118.690 168.340 120.990 168.510 ;
        RECT 121.390 176.770 123.690 176.940 ;
        RECT 121.390 168.510 121.560 176.770 ;
        RECT 122.290 176.080 122.790 176.250 ;
        RECT 122.060 169.370 122.230 175.910 ;
        RECT 122.850 169.370 123.020 175.910 ;
        RECT 122.050 168.800 123.050 169.200 ;
        RECT 123.520 168.510 123.690 176.770 ;
        RECT 133.315 176.770 135.615 176.940 ;
        RECT 133.315 175.830 133.485 176.770 ;
        RECT 133.695 176.080 134.735 176.525 ;
        RECT 133.985 175.830 134.155 175.910 ;
        RECT 133.310 175.300 134.155 175.830 ;
        RECT 133.315 174.360 133.485 175.300 ;
        RECT 133.985 175.220 134.155 175.300 ;
        RECT 134.775 175.220 134.945 175.910 ;
        RECT 134.215 174.880 134.715 175.050 ;
        RECT 135.445 174.360 135.615 176.770 ;
        RECT 133.315 174.190 135.615 174.360 ;
        RECT 136.015 176.770 138.315 176.940 ;
        RECT 121.390 168.340 123.690 168.510 ;
        RECT 136.015 168.510 136.185 176.770 ;
        RECT 136.915 176.080 137.415 176.250 ;
        RECT 136.685 169.370 136.855 175.910 ;
        RECT 137.475 169.370 137.645 175.910 ;
        RECT 136.675 168.800 137.675 169.200 ;
        RECT 138.145 168.510 138.315 176.770 ;
        RECT 138.715 176.770 141.015 176.940 ;
        RECT 138.715 175.830 138.885 176.770 ;
        RECT 139.095 176.080 140.135 176.525 ;
        RECT 139.385 175.830 139.555 175.910 ;
        RECT 138.710 175.300 139.555 175.830 ;
        RECT 138.715 174.360 138.885 175.300 ;
        RECT 139.385 175.220 139.555 175.300 ;
        RECT 140.175 175.220 140.345 175.910 ;
        RECT 139.615 174.880 140.115 175.050 ;
        RECT 140.845 174.360 141.015 176.770 ;
        RECT 141.415 176.770 143.715 176.940 ;
        RECT 141.415 175.830 141.585 176.770 ;
        RECT 141.795 176.080 142.835 176.525 ;
        RECT 142.085 175.830 142.255 175.910 ;
        RECT 141.410 175.300 142.255 175.830 ;
        RECT 138.715 174.190 141.015 174.360 ;
        RECT 141.415 174.360 141.585 175.300 ;
        RECT 142.085 175.220 142.255 175.300 ;
        RECT 142.875 175.220 143.045 175.910 ;
        RECT 142.315 174.880 142.815 175.050 ;
        RECT 143.545 174.360 143.715 176.770 ;
        RECT 141.415 174.190 143.715 174.360 ;
        RECT 144.115 176.770 146.415 176.940 ;
        RECT 136.015 168.340 138.315 168.510 ;
        RECT 144.115 168.510 144.285 176.770 ;
        RECT 145.015 176.080 145.515 176.250 ;
        RECT 144.785 169.370 144.955 175.910 ;
        RECT 145.575 169.370 145.745 175.910 ;
        RECT 144.775 168.800 145.775 169.200 ;
        RECT 146.245 168.510 146.415 176.770 ;
        RECT 144.115 168.340 146.415 168.510 ;
        RECT 146.815 176.770 149.115 176.940 ;
        RECT 146.815 168.510 146.985 176.770 ;
        RECT 147.715 176.080 148.215 176.250 ;
        RECT 147.485 169.370 147.655 175.910 ;
        RECT 148.275 169.370 148.445 175.910 ;
        RECT 147.475 168.800 148.475 169.200 ;
        RECT 148.945 168.510 149.115 176.770 ;
        RECT 146.815 168.340 149.115 168.510 ;
        RECT 23.235 168.000 24.075 168.050 ;
        RECT 48.660 168.000 49.500 168.050 ;
        RECT 74.085 168.000 74.925 168.050 ;
        RECT 99.510 168.000 100.350 168.050 ;
        RECT 124.935 168.000 125.775 168.050 ;
        RECT 150.360 168.000 151.200 168.050 ;
        RECT 22.830 167.830 24.480 168.000 ;
        RECT 8.890 167.285 11.190 167.455 ;
        RECT 6.190 158.285 8.490 158.455 ;
        RECT 6.190 157.350 6.360 158.285 ;
        RECT 7.090 157.595 7.590 157.765 ;
        RECT 6.860 157.350 7.030 157.380 ;
        RECT 6.135 156.370 7.030 157.350 ;
        RECT 6.190 155.435 6.360 156.370 ;
        RECT 6.860 156.340 7.030 156.370 ;
        RECT 7.650 156.340 7.820 157.380 ;
        RECT 6.675 155.955 7.590 156.125 ;
        RECT 6.675 155.750 7.510 155.955 ;
        RECT 8.320 155.435 8.490 158.285 ;
        RECT 6.190 155.265 8.490 155.435 ;
        RECT 8.890 155.435 9.060 167.285 ;
        RECT 9.550 166.575 10.550 167.025 ;
        RECT 9.560 156.340 9.730 166.380 ;
        RECT 10.350 156.340 10.520 166.380 ;
        RECT 9.790 155.955 10.290 156.125 ;
        RECT 11.020 155.435 11.190 167.285 ;
        RECT 16.990 167.285 19.290 167.455 ;
        RECT 11.590 158.285 13.890 158.455 ;
        RECT 11.590 157.350 11.760 158.285 ;
        RECT 12.490 157.595 12.990 157.765 ;
        RECT 12.260 157.350 12.430 157.380 ;
        RECT 11.535 156.370 12.430 157.350 ;
        RECT 8.890 155.265 11.190 155.435 ;
        RECT 11.590 155.435 11.760 156.370 ;
        RECT 12.260 156.340 12.430 156.370 ;
        RECT 13.050 156.340 13.220 157.380 ;
        RECT 12.075 155.955 12.990 156.125 ;
        RECT 12.075 155.750 12.910 155.955 ;
        RECT 13.720 155.435 13.890 158.285 ;
        RECT 14.290 158.285 16.590 158.455 ;
        RECT 14.290 157.350 14.460 158.285 ;
        RECT 15.190 157.595 15.690 157.765 ;
        RECT 14.960 157.350 15.130 157.380 ;
        RECT 14.235 156.370 15.130 157.350 ;
        RECT 11.590 155.265 13.890 155.435 ;
        RECT 14.290 155.435 14.460 156.370 ;
        RECT 14.960 156.340 15.130 156.370 ;
        RECT 15.750 156.340 15.920 157.380 ;
        RECT 14.775 155.955 15.690 156.125 ;
        RECT 14.775 155.750 15.610 155.955 ;
        RECT 16.420 155.435 16.590 158.285 ;
        RECT 14.290 155.265 16.590 155.435 ;
        RECT 16.990 155.435 17.160 167.285 ;
        RECT 17.650 166.575 18.650 167.025 ;
        RECT 17.660 156.340 17.830 166.380 ;
        RECT 18.450 156.340 18.620 166.380 ;
        RECT 17.890 155.955 18.390 156.125 ;
        RECT 19.120 155.435 19.290 167.285 ;
        RECT 16.990 155.265 19.290 155.435 ;
        RECT 19.690 167.285 21.990 167.455 ;
        RECT 19.690 155.435 19.860 167.285 ;
        RECT 20.350 166.575 21.350 167.025 ;
        RECT 20.360 156.340 20.530 166.380 ;
        RECT 21.150 156.340 21.320 166.380 ;
        RECT 20.590 155.955 21.090 156.125 ;
        RECT 21.820 155.435 21.990 167.285 ;
        RECT 19.690 155.265 21.990 155.435 ;
        RECT 6.190 154.195 8.490 154.365 ;
        RECT 6.190 153.255 6.360 154.195 ;
        RECT 6.570 153.505 7.610 153.950 ;
        RECT 6.860 153.255 7.030 153.335 ;
        RECT 6.185 152.725 7.030 153.255 ;
        RECT 6.190 151.785 6.360 152.725 ;
        RECT 6.860 152.645 7.030 152.725 ;
        RECT 7.650 152.645 7.820 153.335 ;
        RECT 7.090 152.305 7.590 152.475 ;
        RECT 8.320 151.785 8.490 154.195 ;
        RECT 6.190 151.615 8.490 151.785 ;
        RECT 8.890 154.195 11.190 154.365 ;
        RECT 8.890 145.935 9.060 154.195 ;
        RECT 9.790 153.505 10.290 153.675 ;
        RECT 9.560 146.795 9.730 153.335 ;
        RECT 10.350 146.795 10.520 153.335 ;
        RECT 9.550 146.225 10.550 146.625 ;
        RECT 11.020 145.935 11.190 154.195 ;
        RECT 11.590 154.195 13.890 154.365 ;
        RECT 11.590 153.255 11.760 154.195 ;
        RECT 11.970 153.505 13.010 153.950 ;
        RECT 12.260 153.255 12.430 153.335 ;
        RECT 11.585 152.725 12.430 153.255 ;
        RECT 11.590 151.785 11.760 152.725 ;
        RECT 12.260 152.645 12.430 152.725 ;
        RECT 13.050 152.645 13.220 153.335 ;
        RECT 12.490 152.305 12.990 152.475 ;
        RECT 13.720 151.785 13.890 154.195 ;
        RECT 14.290 154.195 16.590 154.365 ;
        RECT 14.290 153.255 14.460 154.195 ;
        RECT 14.670 153.505 15.710 153.950 ;
        RECT 14.960 153.255 15.130 153.335 ;
        RECT 14.285 152.725 15.130 153.255 ;
        RECT 11.590 151.615 13.890 151.785 ;
        RECT 14.290 151.785 14.460 152.725 ;
        RECT 14.960 152.645 15.130 152.725 ;
        RECT 15.750 152.645 15.920 153.335 ;
        RECT 15.190 152.305 15.690 152.475 ;
        RECT 16.420 151.785 16.590 154.195 ;
        RECT 14.290 151.615 16.590 151.785 ;
        RECT 16.990 154.195 19.290 154.365 ;
        RECT 8.890 145.765 11.190 145.935 ;
        RECT 16.990 145.935 17.160 154.195 ;
        RECT 17.890 153.505 18.390 153.675 ;
        RECT 17.660 146.795 17.830 153.335 ;
        RECT 18.450 146.795 18.620 153.335 ;
        RECT 17.650 146.225 18.650 146.625 ;
        RECT 19.120 145.935 19.290 154.195 ;
        RECT 16.990 145.765 19.290 145.935 ;
        RECT 19.690 154.195 21.990 154.365 ;
        RECT 19.690 145.935 19.860 154.195 ;
        RECT 20.590 153.505 21.090 153.675 ;
        RECT 20.360 146.795 20.530 153.335 ;
        RECT 21.150 146.795 21.320 153.335 ;
        RECT 20.350 146.225 21.350 146.625 ;
        RECT 21.820 145.935 21.990 154.195 ;
        RECT 22.830 153.800 23.000 167.830 ;
        RECT 23.235 167.780 24.075 167.830 ;
        RECT 23.430 165.115 23.880 167.425 ;
        RECT 23.430 154.205 23.880 156.515 ;
        RECT 23.260 153.800 24.050 153.850 ;
        RECT 24.310 153.800 24.480 167.830 ;
        RECT 48.255 167.830 49.905 168.000 ;
        RECT 34.315 167.285 36.615 167.455 ;
        RECT 31.615 158.285 33.915 158.455 ;
        RECT 31.615 157.350 31.785 158.285 ;
        RECT 32.515 157.595 33.015 157.765 ;
        RECT 32.285 157.350 32.455 157.380 ;
        RECT 31.560 156.370 32.455 157.350 ;
        RECT 31.615 155.435 31.785 156.370 ;
        RECT 32.285 156.340 32.455 156.370 ;
        RECT 33.075 156.340 33.245 157.380 ;
        RECT 32.100 155.955 33.015 156.125 ;
        RECT 32.100 155.750 32.935 155.955 ;
        RECT 33.745 155.435 33.915 158.285 ;
        RECT 31.615 155.265 33.915 155.435 ;
        RECT 34.315 155.435 34.485 167.285 ;
        RECT 34.975 166.575 35.975 167.025 ;
        RECT 34.985 156.340 35.155 166.380 ;
        RECT 35.775 156.340 35.945 166.380 ;
        RECT 35.215 155.955 35.715 156.125 ;
        RECT 36.445 155.435 36.615 167.285 ;
        RECT 42.415 167.285 44.715 167.455 ;
        RECT 37.015 158.285 39.315 158.455 ;
        RECT 37.015 157.350 37.185 158.285 ;
        RECT 37.915 157.595 38.415 157.765 ;
        RECT 37.685 157.350 37.855 157.380 ;
        RECT 36.960 156.370 37.855 157.350 ;
        RECT 34.315 155.265 36.615 155.435 ;
        RECT 37.015 155.435 37.185 156.370 ;
        RECT 37.685 156.340 37.855 156.370 ;
        RECT 38.475 156.340 38.645 157.380 ;
        RECT 37.500 155.955 38.415 156.125 ;
        RECT 37.500 155.750 38.335 155.955 ;
        RECT 39.145 155.435 39.315 158.285 ;
        RECT 39.715 158.285 42.015 158.455 ;
        RECT 39.715 157.350 39.885 158.285 ;
        RECT 40.615 157.595 41.115 157.765 ;
        RECT 40.385 157.350 40.555 157.380 ;
        RECT 39.660 156.370 40.555 157.350 ;
        RECT 37.015 155.265 39.315 155.435 ;
        RECT 39.715 155.435 39.885 156.370 ;
        RECT 40.385 156.340 40.555 156.370 ;
        RECT 41.175 156.340 41.345 157.380 ;
        RECT 40.200 155.955 41.115 156.125 ;
        RECT 40.200 155.750 41.035 155.955 ;
        RECT 41.845 155.435 42.015 158.285 ;
        RECT 39.715 155.265 42.015 155.435 ;
        RECT 42.415 155.435 42.585 167.285 ;
        RECT 43.075 166.575 44.075 167.025 ;
        RECT 43.085 156.340 43.255 166.380 ;
        RECT 43.875 156.340 44.045 166.380 ;
        RECT 43.315 155.955 43.815 156.125 ;
        RECT 44.545 155.435 44.715 167.285 ;
        RECT 42.415 155.265 44.715 155.435 ;
        RECT 45.115 167.285 47.415 167.455 ;
        RECT 45.115 155.435 45.285 167.285 ;
        RECT 45.775 166.575 46.775 167.025 ;
        RECT 45.785 156.340 45.955 166.380 ;
        RECT 46.575 156.340 46.745 166.380 ;
        RECT 46.015 155.955 46.515 156.125 ;
        RECT 47.245 155.435 47.415 167.285 ;
        RECT 45.115 155.265 47.415 155.435 ;
        RECT 22.830 153.630 24.480 153.800 ;
        RECT 31.615 154.195 33.915 154.365 ;
        RECT 23.260 153.580 24.050 153.630 ;
        RECT 31.615 153.255 31.785 154.195 ;
        RECT 31.995 153.505 33.035 153.950 ;
        RECT 32.285 153.255 32.455 153.335 ;
        RECT 31.610 152.725 32.455 153.255 ;
        RECT 31.615 151.785 31.785 152.725 ;
        RECT 32.285 152.645 32.455 152.725 ;
        RECT 33.075 152.645 33.245 153.335 ;
        RECT 32.515 152.305 33.015 152.475 ;
        RECT 33.745 151.785 33.915 154.195 ;
        RECT 31.615 151.615 33.915 151.785 ;
        RECT 34.315 154.195 36.615 154.365 ;
        RECT 19.690 145.765 21.990 145.935 ;
        RECT 34.315 145.935 34.485 154.195 ;
        RECT 35.215 153.505 35.715 153.675 ;
        RECT 34.985 146.795 35.155 153.335 ;
        RECT 35.775 146.795 35.945 153.335 ;
        RECT 34.975 146.225 35.975 146.625 ;
        RECT 36.445 145.935 36.615 154.195 ;
        RECT 37.015 154.195 39.315 154.365 ;
        RECT 37.015 153.255 37.185 154.195 ;
        RECT 37.395 153.505 38.435 153.950 ;
        RECT 37.685 153.255 37.855 153.335 ;
        RECT 37.010 152.725 37.855 153.255 ;
        RECT 37.015 151.785 37.185 152.725 ;
        RECT 37.685 152.645 37.855 152.725 ;
        RECT 38.475 152.645 38.645 153.335 ;
        RECT 37.915 152.305 38.415 152.475 ;
        RECT 39.145 151.785 39.315 154.195 ;
        RECT 39.715 154.195 42.015 154.365 ;
        RECT 39.715 153.255 39.885 154.195 ;
        RECT 40.095 153.505 41.135 153.950 ;
        RECT 40.385 153.255 40.555 153.335 ;
        RECT 39.710 152.725 40.555 153.255 ;
        RECT 37.015 151.615 39.315 151.785 ;
        RECT 39.715 151.785 39.885 152.725 ;
        RECT 40.385 152.645 40.555 152.725 ;
        RECT 41.175 152.645 41.345 153.335 ;
        RECT 40.615 152.305 41.115 152.475 ;
        RECT 41.845 151.785 42.015 154.195 ;
        RECT 39.715 151.615 42.015 151.785 ;
        RECT 42.415 154.195 44.715 154.365 ;
        RECT 34.315 145.765 36.615 145.935 ;
        RECT 42.415 145.935 42.585 154.195 ;
        RECT 43.315 153.505 43.815 153.675 ;
        RECT 43.085 146.795 43.255 153.335 ;
        RECT 43.875 146.795 44.045 153.335 ;
        RECT 43.075 146.225 44.075 146.625 ;
        RECT 44.545 145.935 44.715 154.195 ;
        RECT 42.415 145.765 44.715 145.935 ;
        RECT 45.115 154.195 47.415 154.365 ;
        RECT 45.115 145.935 45.285 154.195 ;
        RECT 46.015 153.505 46.515 153.675 ;
        RECT 45.785 146.795 45.955 153.335 ;
        RECT 46.575 146.795 46.745 153.335 ;
        RECT 45.775 146.225 46.775 146.625 ;
        RECT 47.245 145.935 47.415 154.195 ;
        RECT 48.255 153.800 48.425 167.830 ;
        RECT 48.660 167.780 49.500 167.830 ;
        RECT 48.855 165.115 49.305 167.425 ;
        RECT 48.855 154.205 49.305 156.515 ;
        RECT 48.685 153.800 49.475 153.850 ;
        RECT 49.735 153.800 49.905 167.830 ;
        RECT 73.680 167.830 75.330 168.000 ;
        RECT 59.740 167.285 62.040 167.455 ;
        RECT 57.040 158.285 59.340 158.455 ;
        RECT 57.040 157.350 57.210 158.285 ;
        RECT 57.940 157.595 58.440 157.765 ;
        RECT 57.710 157.350 57.880 157.380 ;
        RECT 56.985 156.370 57.880 157.350 ;
        RECT 57.040 155.435 57.210 156.370 ;
        RECT 57.710 156.340 57.880 156.370 ;
        RECT 58.500 156.340 58.670 157.380 ;
        RECT 57.525 155.955 58.440 156.125 ;
        RECT 57.525 155.750 58.360 155.955 ;
        RECT 59.170 155.435 59.340 158.285 ;
        RECT 57.040 155.265 59.340 155.435 ;
        RECT 59.740 155.435 59.910 167.285 ;
        RECT 60.400 166.575 61.400 167.025 ;
        RECT 60.410 156.340 60.580 166.380 ;
        RECT 61.200 156.340 61.370 166.380 ;
        RECT 60.640 155.955 61.140 156.125 ;
        RECT 61.870 155.435 62.040 167.285 ;
        RECT 67.840 167.285 70.140 167.455 ;
        RECT 62.440 158.285 64.740 158.455 ;
        RECT 62.440 157.350 62.610 158.285 ;
        RECT 63.340 157.595 63.840 157.765 ;
        RECT 63.110 157.350 63.280 157.380 ;
        RECT 62.385 156.370 63.280 157.350 ;
        RECT 59.740 155.265 62.040 155.435 ;
        RECT 62.440 155.435 62.610 156.370 ;
        RECT 63.110 156.340 63.280 156.370 ;
        RECT 63.900 156.340 64.070 157.380 ;
        RECT 62.925 155.955 63.840 156.125 ;
        RECT 62.925 155.750 63.760 155.955 ;
        RECT 64.570 155.435 64.740 158.285 ;
        RECT 65.140 158.285 67.440 158.455 ;
        RECT 65.140 157.350 65.310 158.285 ;
        RECT 66.040 157.595 66.540 157.765 ;
        RECT 65.810 157.350 65.980 157.380 ;
        RECT 65.085 156.370 65.980 157.350 ;
        RECT 62.440 155.265 64.740 155.435 ;
        RECT 65.140 155.435 65.310 156.370 ;
        RECT 65.810 156.340 65.980 156.370 ;
        RECT 66.600 156.340 66.770 157.380 ;
        RECT 65.625 155.955 66.540 156.125 ;
        RECT 65.625 155.750 66.460 155.955 ;
        RECT 67.270 155.435 67.440 158.285 ;
        RECT 65.140 155.265 67.440 155.435 ;
        RECT 67.840 155.435 68.010 167.285 ;
        RECT 68.500 166.575 69.500 167.025 ;
        RECT 68.510 156.340 68.680 166.380 ;
        RECT 69.300 156.340 69.470 166.380 ;
        RECT 68.740 155.955 69.240 156.125 ;
        RECT 69.970 155.435 70.140 167.285 ;
        RECT 67.840 155.265 70.140 155.435 ;
        RECT 70.540 167.285 72.840 167.455 ;
        RECT 70.540 155.435 70.710 167.285 ;
        RECT 71.200 166.575 72.200 167.025 ;
        RECT 71.210 156.340 71.380 166.380 ;
        RECT 72.000 156.340 72.170 166.380 ;
        RECT 71.440 155.955 71.940 156.125 ;
        RECT 72.670 155.435 72.840 167.285 ;
        RECT 70.540 155.265 72.840 155.435 ;
        RECT 48.255 153.630 49.905 153.800 ;
        RECT 57.040 154.195 59.340 154.365 ;
        RECT 48.685 153.580 49.475 153.630 ;
        RECT 57.040 153.255 57.210 154.195 ;
        RECT 57.420 153.505 58.460 153.950 ;
        RECT 57.710 153.255 57.880 153.335 ;
        RECT 57.035 152.725 57.880 153.255 ;
        RECT 57.040 151.785 57.210 152.725 ;
        RECT 57.710 152.645 57.880 152.725 ;
        RECT 58.500 152.645 58.670 153.335 ;
        RECT 57.940 152.305 58.440 152.475 ;
        RECT 59.170 151.785 59.340 154.195 ;
        RECT 57.040 151.615 59.340 151.785 ;
        RECT 59.740 154.195 62.040 154.365 ;
        RECT 45.115 145.765 47.415 145.935 ;
        RECT 59.740 145.935 59.910 154.195 ;
        RECT 60.640 153.505 61.140 153.675 ;
        RECT 60.410 146.795 60.580 153.335 ;
        RECT 61.200 146.795 61.370 153.335 ;
        RECT 60.400 146.225 61.400 146.625 ;
        RECT 61.870 145.935 62.040 154.195 ;
        RECT 62.440 154.195 64.740 154.365 ;
        RECT 62.440 153.255 62.610 154.195 ;
        RECT 62.820 153.505 63.860 153.950 ;
        RECT 63.110 153.255 63.280 153.335 ;
        RECT 62.435 152.725 63.280 153.255 ;
        RECT 62.440 151.785 62.610 152.725 ;
        RECT 63.110 152.645 63.280 152.725 ;
        RECT 63.900 152.645 64.070 153.335 ;
        RECT 63.340 152.305 63.840 152.475 ;
        RECT 64.570 151.785 64.740 154.195 ;
        RECT 65.140 154.195 67.440 154.365 ;
        RECT 65.140 153.255 65.310 154.195 ;
        RECT 65.520 153.505 66.560 153.950 ;
        RECT 65.810 153.255 65.980 153.335 ;
        RECT 65.135 152.725 65.980 153.255 ;
        RECT 62.440 151.615 64.740 151.785 ;
        RECT 65.140 151.785 65.310 152.725 ;
        RECT 65.810 152.645 65.980 152.725 ;
        RECT 66.600 152.645 66.770 153.335 ;
        RECT 66.040 152.305 66.540 152.475 ;
        RECT 67.270 151.785 67.440 154.195 ;
        RECT 65.140 151.615 67.440 151.785 ;
        RECT 67.840 154.195 70.140 154.365 ;
        RECT 59.740 145.765 62.040 145.935 ;
        RECT 67.840 145.935 68.010 154.195 ;
        RECT 68.740 153.505 69.240 153.675 ;
        RECT 68.510 146.795 68.680 153.335 ;
        RECT 69.300 146.795 69.470 153.335 ;
        RECT 68.500 146.225 69.500 146.625 ;
        RECT 69.970 145.935 70.140 154.195 ;
        RECT 67.840 145.765 70.140 145.935 ;
        RECT 70.540 154.195 72.840 154.365 ;
        RECT 70.540 145.935 70.710 154.195 ;
        RECT 71.440 153.505 71.940 153.675 ;
        RECT 71.210 146.795 71.380 153.335 ;
        RECT 72.000 146.795 72.170 153.335 ;
        RECT 71.200 146.225 72.200 146.625 ;
        RECT 72.670 145.935 72.840 154.195 ;
        RECT 73.680 153.800 73.850 167.830 ;
        RECT 74.085 167.780 74.925 167.830 ;
        RECT 74.280 165.115 74.730 167.425 ;
        RECT 74.280 154.205 74.730 156.515 ;
        RECT 74.110 153.800 74.900 153.850 ;
        RECT 75.160 153.800 75.330 167.830 ;
        RECT 99.105 167.830 100.755 168.000 ;
        RECT 85.165 167.285 87.465 167.455 ;
        RECT 82.465 158.285 84.765 158.455 ;
        RECT 82.465 157.350 82.635 158.285 ;
        RECT 83.365 157.595 83.865 157.765 ;
        RECT 83.135 157.350 83.305 157.380 ;
        RECT 82.410 156.370 83.305 157.350 ;
        RECT 82.465 155.435 82.635 156.370 ;
        RECT 83.135 156.340 83.305 156.370 ;
        RECT 83.925 156.340 84.095 157.380 ;
        RECT 82.950 155.955 83.865 156.125 ;
        RECT 82.950 155.750 83.785 155.955 ;
        RECT 84.595 155.435 84.765 158.285 ;
        RECT 82.465 155.265 84.765 155.435 ;
        RECT 85.165 155.435 85.335 167.285 ;
        RECT 85.825 166.575 86.825 167.025 ;
        RECT 85.835 156.340 86.005 166.380 ;
        RECT 86.625 156.340 86.795 166.380 ;
        RECT 86.065 155.955 86.565 156.125 ;
        RECT 87.295 155.435 87.465 167.285 ;
        RECT 93.265 167.285 95.565 167.455 ;
        RECT 87.865 158.285 90.165 158.455 ;
        RECT 87.865 157.350 88.035 158.285 ;
        RECT 88.765 157.595 89.265 157.765 ;
        RECT 88.535 157.350 88.705 157.380 ;
        RECT 87.810 156.370 88.705 157.350 ;
        RECT 85.165 155.265 87.465 155.435 ;
        RECT 87.865 155.435 88.035 156.370 ;
        RECT 88.535 156.340 88.705 156.370 ;
        RECT 89.325 156.340 89.495 157.380 ;
        RECT 88.350 155.955 89.265 156.125 ;
        RECT 88.350 155.750 89.185 155.955 ;
        RECT 89.995 155.435 90.165 158.285 ;
        RECT 90.565 158.285 92.865 158.455 ;
        RECT 90.565 157.350 90.735 158.285 ;
        RECT 91.465 157.595 91.965 157.765 ;
        RECT 91.235 157.350 91.405 157.380 ;
        RECT 90.510 156.370 91.405 157.350 ;
        RECT 87.865 155.265 90.165 155.435 ;
        RECT 90.565 155.435 90.735 156.370 ;
        RECT 91.235 156.340 91.405 156.370 ;
        RECT 92.025 156.340 92.195 157.380 ;
        RECT 91.050 155.955 91.965 156.125 ;
        RECT 91.050 155.750 91.885 155.955 ;
        RECT 92.695 155.435 92.865 158.285 ;
        RECT 90.565 155.265 92.865 155.435 ;
        RECT 93.265 155.435 93.435 167.285 ;
        RECT 93.925 166.575 94.925 167.025 ;
        RECT 93.935 156.340 94.105 166.380 ;
        RECT 94.725 156.340 94.895 166.380 ;
        RECT 94.165 155.955 94.665 156.125 ;
        RECT 95.395 155.435 95.565 167.285 ;
        RECT 93.265 155.265 95.565 155.435 ;
        RECT 95.965 167.285 98.265 167.455 ;
        RECT 95.965 155.435 96.135 167.285 ;
        RECT 96.625 166.575 97.625 167.025 ;
        RECT 96.635 156.340 96.805 166.380 ;
        RECT 97.425 156.340 97.595 166.380 ;
        RECT 96.865 155.955 97.365 156.125 ;
        RECT 98.095 155.435 98.265 167.285 ;
        RECT 95.965 155.265 98.265 155.435 ;
        RECT 73.680 153.630 75.330 153.800 ;
        RECT 82.465 154.195 84.765 154.365 ;
        RECT 74.110 153.580 74.900 153.630 ;
        RECT 82.465 153.255 82.635 154.195 ;
        RECT 82.845 153.505 83.885 153.950 ;
        RECT 83.135 153.255 83.305 153.335 ;
        RECT 82.460 152.725 83.305 153.255 ;
        RECT 82.465 151.785 82.635 152.725 ;
        RECT 83.135 152.645 83.305 152.725 ;
        RECT 83.925 152.645 84.095 153.335 ;
        RECT 83.365 152.305 83.865 152.475 ;
        RECT 84.595 151.785 84.765 154.195 ;
        RECT 82.465 151.615 84.765 151.785 ;
        RECT 85.165 154.195 87.465 154.365 ;
        RECT 70.540 145.765 72.840 145.935 ;
        RECT 85.165 145.935 85.335 154.195 ;
        RECT 86.065 153.505 86.565 153.675 ;
        RECT 85.835 146.795 86.005 153.335 ;
        RECT 86.625 146.795 86.795 153.335 ;
        RECT 85.825 146.225 86.825 146.625 ;
        RECT 87.295 145.935 87.465 154.195 ;
        RECT 87.865 154.195 90.165 154.365 ;
        RECT 87.865 153.255 88.035 154.195 ;
        RECT 88.245 153.505 89.285 153.950 ;
        RECT 88.535 153.255 88.705 153.335 ;
        RECT 87.860 152.725 88.705 153.255 ;
        RECT 87.865 151.785 88.035 152.725 ;
        RECT 88.535 152.645 88.705 152.725 ;
        RECT 89.325 152.645 89.495 153.335 ;
        RECT 88.765 152.305 89.265 152.475 ;
        RECT 89.995 151.785 90.165 154.195 ;
        RECT 90.565 154.195 92.865 154.365 ;
        RECT 90.565 153.255 90.735 154.195 ;
        RECT 90.945 153.505 91.985 153.950 ;
        RECT 91.235 153.255 91.405 153.335 ;
        RECT 90.560 152.725 91.405 153.255 ;
        RECT 87.865 151.615 90.165 151.785 ;
        RECT 90.565 151.785 90.735 152.725 ;
        RECT 91.235 152.645 91.405 152.725 ;
        RECT 92.025 152.645 92.195 153.335 ;
        RECT 91.465 152.305 91.965 152.475 ;
        RECT 92.695 151.785 92.865 154.195 ;
        RECT 90.565 151.615 92.865 151.785 ;
        RECT 93.265 154.195 95.565 154.365 ;
        RECT 85.165 145.765 87.465 145.935 ;
        RECT 93.265 145.935 93.435 154.195 ;
        RECT 94.165 153.505 94.665 153.675 ;
        RECT 93.935 146.795 94.105 153.335 ;
        RECT 94.725 146.795 94.895 153.335 ;
        RECT 93.925 146.225 94.925 146.625 ;
        RECT 95.395 145.935 95.565 154.195 ;
        RECT 93.265 145.765 95.565 145.935 ;
        RECT 95.965 154.195 98.265 154.365 ;
        RECT 95.965 145.935 96.135 154.195 ;
        RECT 96.865 153.505 97.365 153.675 ;
        RECT 96.635 146.795 96.805 153.335 ;
        RECT 97.425 146.795 97.595 153.335 ;
        RECT 96.625 146.225 97.625 146.625 ;
        RECT 98.095 145.935 98.265 154.195 ;
        RECT 99.105 153.800 99.275 167.830 ;
        RECT 99.510 167.780 100.350 167.830 ;
        RECT 99.705 165.115 100.155 167.425 ;
        RECT 99.705 154.205 100.155 156.515 ;
        RECT 99.535 153.800 100.325 153.850 ;
        RECT 100.585 153.800 100.755 167.830 ;
        RECT 124.530 167.830 126.180 168.000 ;
        RECT 110.590 167.285 112.890 167.455 ;
        RECT 107.890 158.285 110.190 158.455 ;
        RECT 107.890 157.350 108.060 158.285 ;
        RECT 108.790 157.595 109.290 157.765 ;
        RECT 108.560 157.350 108.730 157.380 ;
        RECT 107.835 156.370 108.730 157.350 ;
        RECT 107.890 155.435 108.060 156.370 ;
        RECT 108.560 156.340 108.730 156.370 ;
        RECT 109.350 156.340 109.520 157.380 ;
        RECT 108.375 155.955 109.290 156.125 ;
        RECT 108.375 155.750 109.210 155.955 ;
        RECT 110.020 155.435 110.190 158.285 ;
        RECT 107.890 155.265 110.190 155.435 ;
        RECT 110.590 155.435 110.760 167.285 ;
        RECT 111.250 166.575 112.250 167.025 ;
        RECT 111.260 156.340 111.430 166.380 ;
        RECT 112.050 156.340 112.220 166.380 ;
        RECT 111.490 155.955 111.990 156.125 ;
        RECT 112.720 155.435 112.890 167.285 ;
        RECT 118.690 167.285 120.990 167.455 ;
        RECT 113.290 158.285 115.590 158.455 ;
        RECT 113.290 157.350 113.460 158.285 ;
        RECT 114.190 157.595 114.690 157.765 ;
        RECT 113.960 157.350 114.130 157.380 ;
        RECT 113.235 156.370 114.130 157.350 ;
        RECT 110.590 155.265 112.890 155.435 ;
        RECT 113.290 155.435 113.460 156.370 ;
        RECT 113.960 156.340 114.130 156.370 ;
        RECT 114.750 156.340 114.920 157.380 ;
        RECT 113.775 155.955 114.690 156.125 ;
        RECT 113.775 155.750 114.610 155.955 ;
        RECT 115.420 155.435 115.590 158.285 ;
        RECT 115.990 158.285 118.290 158.455 ;
        RECT 115.990 157.350 116.160 158.285 ;
        RECT 116.890 157.595 117.390 157.765 ;
        RECT 116.660 157.350 116.830 157.380 ;
        RECT 115.935 156.370 116.830 157.350 ;
        RECT 113.290 155.265 115.590 155.435 ;
        RECT 115.990 155.435 116.160 156.370 ;
        RECT 116.660 156.340 116.830 156.370 ;
        RECT 117.450 156.340 117.620 157.380 ;
        RECT 116.475 155.955 117.390 156.125 ;
        RECT 116.475 155.750 117.310 155.955 ;
        RECT 118.120 155.435 118.290 158.285 ;
        RECT 115.990 155.265 118.290 155.435 ;
        RECT 118.690 155.435 118.860 167.285 ;
        RECT 119.350 166.575 120.350 167.025 ;
        RECT 119.360 156.340 119.530 166.380 ;
        RECT 120.150 156.340 120.320 166.380 ;
        RECT 119.590 155.955 120.090 156.125 ;
        RECT 120.820 155.435 120.990 167.285 ;
        RECT 118.690 155.265 120.990 155.435 ;
        RECT 121.390 167.285 123.690 167.455 ;
        RECT 121.390 155.435 121.560 167.285 ;
        RECT 122.050 166.575 123.050 167.025 ;
        RECT 122.060 156.340 122.230 166.380 ;
        RECT 122.850 156.340 123.020 166.380 ;
        RECT 122.290 155.955 122.790 156.125 ;
        RECT 123.520 155.435 123.690 167.285 ;
        RECT 121.390 155.265 123.690 155.435 ;
        RECT 99.105 153.630 100.755 153.800 ;
        RECT 107.890 154.195 110.190 154.365 ;
        RECT 99.535 153.580 100.325 153.630 ;
        RECT 107.890 153.255 108.060 154.195 ;
        RECT 108.270 153.505 109.310 153.950 ;
        RECT 108.560 153.255 108.730 153.335 ;
        RECT 107.885 152.725 108.730 153.255 ;
        RECT 107.890 151.785 108.060 152.725 ;
        RECT 108.560 152.645 108.730 152.725 ;
        RECT 109.350 152.645 109.520 153.335 ;
        RECT 108.790 152.305 109.290 152.475 ;
        RECT 110.020 151.785 110.190 154.195 ;
        RECT 107.890 151.615 110.190 151.785 ;
        RECT 110.590 154.195 112.890 154.365 ;
        RECT 95.965 145.765 98.265 145.935 ;
        RECT 110.590 145.935 110.760 154.195 ;
        RECT 111.490 153.505 111.990 153.675 ;
        RECT 111.260 146.795 111.430 153.335 ;
        RECT 112.050 146.795 112.220 153.335 ;
        RECT 111.250 146.225 112.250 146.625 ;
        RECT 112.720 145.935 112.890 154.195 ;
        RECT 113.290 154.195 115.590 154.365 ;
        RECT 113.290 153.255 113.460 154.195 ;
        RECT 113.670 153.505 114.710 153.950 ;
        RECT 113.960 153.255 114.130 153.335 ;
        RECT 113.285 152.725 114.130 153.255 ;
        RECT 113.290 151.785 113.460 152.725 ;
        RECT 113.960 152.645 114.130 152.725 ;
        RECT 114.750 152.645 114.920 153.335 ;
        RECT 114.190 152.305 114.690 152.475 ;
        RECT 115.420 151.785 115.590 154.195 ;
        RECT 115.990 154.195 118.290 154.365 ;
        RECT 115.990 153.255 116.160 154.195 ;
        RECT 116.370 153.505 117.410 153.950 ;
        RECT 116.660 153.255 116.830 153.335 ;
        RECT 115.985 152.725 116.830 153.255 ;
        RECT 113.290 151.615 115.590 151.785 ;
        RECT 115.990 151.785 116.160 152.725 ;
        RECT 116.660 152.645 116.830 152.725 ;
        RECT 117.450 152.645 117.620 153.335 ;
        RECT 116.890 152.305 117.390 152.475 ;
        RECT 118.120 151.785 118.290 154.195 ;
        RECT 115.990 151.615 118.290 151.785 ;
        RECT 118.690 154.195 120.990 154.365 ;
        RECT 110.590 145.765 112.890 145.935 ;
        RECT 118.690 145.935 118.860 154.195 ;
        RECT 119.590 153.505 120.090 153.675 ;
        RECT 119.360 146.795 119.530 153.335 ;
        RECT 120.150 146.795 120.320 153.335 ;
        RECT 119.350 146.225 120.350 146.625 ;
        RECT 120.820 145.935 120.990 154.195 ;
        RECT 118.690 145.765 120.990 145.935 ;
        RECT 121.390 154.195 123.690 154.365 ;
        RECT 121.390 145.935 121.560 154.195 ;
        RECT 122.290 153.505 122.790 153.675 ;
        RECT 122.060 146.795 122.230 153.335 ;
        RECT 122.850 146.795 123.020 153.335 ;
        RECT 122.050 146.225 123.050 146.625 ;
        RECT 123.520 145.935 123.690 154.195 ;
        RECT 124.530 153.800 124.700 167.830 ;
        RECT 124.935 167.780 125.775 167.830 ;
        RECT 125.130 165.115 125.580 167.425 ;
        RECT 125.130 154.205 125.580 156.515 ;
        RECT 124.960 153.800 125.750 153.850 ;
        RECT 126.010 153.800 126.180 167.830 ;
        RECT 149.955 167.830 151.605 168.000 ;
        RECT 136.015 167.285 138.315 167.455 ;
        RECT 133.315 158.285 135.615 158.455 ;
        RECT 133.315 157.350 133.485 158.285 ;
        RECT 134.215 157.595 134.715 157.765 ;
        RECT 133.985 157.350 134.155 157.380 ;
        RECT 133.260 156.370 134.155 157.350 ;
        RECT 133.315 155.435 133.485 156.370 ;
        RECT 133.985 156.340 134.155 156.370 ;
        RECT 134.775 156.340 134.945 157.380 ;
        RECT 133.800 155.955 134.715 156.125 ;
        RECT 133.800 155.750 134.635 155.955 ;
        RECT 135.445 155.435 135.615 158.285 ;
        RECT 133.315 155.265 135.615 155.435 ;
        RECT 136.015 155.435 136.185 167.285 ;
        RECT 136.675 166.575 137.675 167.025 ;
        RECT 136.685 156.340 136.855 166.380 ;
        RECT 137.475 156.340 137.645 166.380 ;
        RECT 136.915 155.955 137.415 156.125 ;
        RECT 138.145 155.435 138.315 167.285 ;
        RECT 144.115 167.285 146.415 167.455 ;
        RECT 138.715 158.285 141.015 158.455 ;
        RECT 138.715 157.350 138.885 158.285 ;
        RECT 139.615 157.595 140.115 157.765 ;
        RECT 139.385 157.350 139.555 157.380 ;
        RECT 138.660 156.370 139.555 157.350 ;
        RECT 136.015 155.265 138.315 155.435 ;
        RECT 138.715 155.435 138.885 156.370 ;
        RECT 139.385 156.340 139.555 156.370 ;
        RECT 140.175 156.340 140.345 157.380 ;
        RECT 139.200 155.955 140.115 156.125 ;
        RECT 139.200 155.750 140.035 155.955 ;
        RECT 140.845 155.435 141.015 158.285 ;
        RECT 141.415 158.285 143.715 158.455 ;
        RECT 141.415 157.350 141.585 158.285 ;
        RECT 142.315 157.595 142.815 157.765 ;
        RECT 142.085 157.350 142.255 157.380 ;
        RECT 141.360 156.370 142.255 157.350 ;
        RECT 138.715 155.265 141.015 155.435 ;
        RECT 141.415 155.435 141.585 156.370 ;
        RECT 142.085 156.340 142.255 156.370 ;
        RECT 142.875 156.340 143.045 157.380 ;
        RECT 141.900 155.955 142.815 156.125 ;
        RECT 141.900 155.750 142.735 155.955 ;
        RECT 143.545 155.435 143.715 158.285 ;
        RECT 141.415 155.265 143.715 155.435 ;
        RECT 144.115 155.435 144.285 167.285 ;
        RECT 144.775 166.575 145.775 167.025 ;
        RECT 144.785 156.340 144.955 166.380 ;
        RECT 145.575 156.340 145.745 166.380 ;
        RECT 145.015 155.955 145.515 156.125 ;
        RECT 146.245 155.435 146.415 167.285 ;
        RECT 144.115 155.265 146.415 155.435 ;
        RECT 146.815 167.285 149.115 167.455 ;
        RECT 146.815 155.435 146.985 167.285 ;
        RECT 147.475 166.575 148.475 167.025 ;
        RECT 147.485 156.340 147.655 166.380 ;
        RECT 148.275 156.340 148.445 166.380 ;
        RECT 147.715 155.955 148.215 156.125 ;
        RECT 148.945 155.435 149.115 167.285 ;
        RECT 146.815 155.265 149.115 155.435 ;
        RECT 124.530 153.630 126.180 153.800 ;
        RECT 133.315 154.195 135.615 154.365 ;
        RECT 124.960 153.580 125.750 153.630 ;
        RECT 133.315 153.255 133.485 154.195 ;
        RECT 133.695 153.505 134.735 153.950 ;
        RECT 133.985 153.255 134.155 153.335 ;
        RECT 133.310 152.725 134.155 153.255 ;
        RECT 133.315 151.785 133.485 152.725 ;
        RECT 133.985 152.645 134.155 152.725 ;
        RECT 134.775 152.645 134.945 153.335 ;
        RECT 134.215 152.305 134.715 152.475 ;
        RECT 135.445 151.785 135.615 154.195 ;
        RECT 133.315 151.615 135.615 151.785 ;
        RECT 136.015 154.195 138.315 154.365 ;
        RECT 121.390 145.765 123.690 145.935 ;
        RECT 136.015 145.935 136.185 154.195 ;
        RECT 136.915 153.505 137.415 153.675 ;
        RECT 136.685 146.795 136.855 153.335 ;
        RECT 137.475 146.795 137.645 153.335 ;
        RECT 136.675 146.225 137.675 146.625 ;
        RECT 138.145 145.935 138.315 154.195 ;
        RECT 138.715 154.195 141.015 154.365 ;
        RECT 138.715 153.255 138.885 154.195 ;
        RECT 139.095 153.505 140.135 153.950 ;
        RECT 139.385 153.255 139.555 153.335 ;
        RECT 138.710 152.725 139.555 153.255 ;
        RECT 138.715 151.785 138.885 152.725 ;
        RECT 139.385 152.645 139.555 152.725 ;
        RECT 140.175 152.645 140.345 153.335 ;
        RECT 139.615 152.305 140.115 152.475 ;
        RECT 140.845 151.785 141.015 154.195 ;
        RECT 141.415 154.195 143.715 154.365 ;
        RECT 141.415 153.255 141.585 154.195 ;
        RECT 141.795 153.505 142.835 153.950 ;
        RECT 142.085 153.255 142.255 153.335 ;
        RECT 141.410 152.725 142.255 153.255 ;
        RECT 138.715 151.615 141.015 151.785 ;
        RECT 141.415 151.785 141.585 152.725 ;
        RECT 142.085 152.645 142.255 152.725 ;
        RECT 142.875 152.645 143.045 153.335 ;
        RECT 142.315 152.305 142.815 152.475 ;
        RECT 143.545 151.785 143.715 154.195 ;
        RECT 141.415 151.615 143.715 151.785 ;
        RECT 144.115 154.195 146.415 154.365 ;
        RECT 136.015 145.765 138.315 145.935 ;
        RECT 144.115 145.935 144.285 154.195 ;
        RECT 145.015 153.505 145.515 153.675 ;
        RECT 144.785 146.795 144.955 153.335 ;
        RECT 145.575 146.795 145.745 153.335 ;
        RECT 144.775 146.225 145.775 146.625 ;
        RECT 146.245 145.935 146.415 154.195 ;
        RECT 144.115 145.765 146.415 145.935 ;
        RECT 146.815 154.195 149.115 154.365 ;
        RECT 146.815 145.935 146.985 154.195 ;
        RECT 147.715 153.505 148.215 153.675 ;
        RECT 147.485 146.795 147.655 153.335 ;
        RECT 148.275 146.795 148.445 153.335 ;
        RECT 147.475 146.225 148.475 146.625 ;
        RECT 148.945 145.935 149.115 154.195 ;
        RECT 149.955 153.800 150.125 167.830 ;
        RECT 150.360 167.780 151.200 167.830 ;
        RECT 150.555 165.115 151.005 167.425 ;
        RECT 150.555 154.205 151.005 156.515 ;
        RECT 150.385 153.800 151.175 153.850 ;
        RECT 151.435 153.800 151.605 167.830 ;
        RECT 149.955 153.630 151.605 153.800 ;
        RECT 150.385 153.580 151.175 153.630 ;
        RECT 146.815 145.765 149.115 145.935 ;
        RECT 8.890 140.435 11.190 140.605 ;
        RECT 6.190 131.435 8.490 131.605 ;
        RECT 6.190 130.500 6.360 131.435 ;
        RECT 7.090 130.745 7.590 130.915 ;
        RECT 6.860 130.500 7.030 130.530 ;
        RECT 6.135 129.520 7.030 130.500 ;
        RECT 6.190 128.585 6.360 129.520 ;
        RECT 6.860 129.490 7.030 129.520 ;
        RECT 7.650 129.490 7.820 130.530 ;
        RECT 6.675 129.105 7.590 129.275 ;
        RECT 6.675 128.900 7.510 129.105 ;
        RECT 8.320 128.585 8.490 131.435 ;
        RECT 6.190 128.415 8.490 128.585 ;
        RECT 8.890 128.585 9.060 140.435 ;
        RECT 9.550 139.725 10.550 140.175 ;
        RECT 9.560 129.490 9.730 139.530 ;
        RECT 10.350 129.490 10.520 139.530 ;
        RECT 9.790 129.105 10.290 129.275 ;
        RECT 11.020 128.585 11.190 140.435 ;
        RECT 16.990 140.435 19.290 140.605 ;
        RECT 11.590 131.435 13.890 131.605 ;
        RECT 11.590 130.500 11.760 131.435 ;
        RECT 12.490 130.745 12.990 130.915 ;
        RECT 12.260 130.500 12.430 130.530 ;
        RECT 11.535 129.520 12.430 130.500 ;
        RECT 8.890 128.415 11.190 128.585 ;
        RECT 11.590 128.585 11.760 129.520 ;
        RECT 12.260 129.490 12.430 129.520 ;
        RECT 13.050 129.490 13.220 130.530 ;
        RECT 12.075 129.105 12.990 129.275 ;
        RECT 12.075 128.900 12.910 129.105 ;
        RECT 13.720 128.585 13.890 131.435 ;
        RECT 14.290 131.435 16.590 131.605 ;
        RECT 14.290 130.500 14.460 131.435 ;
        RECT 15.190 130.745 15.690 130.915 ;
        RECT 14.960 130.500 15.130 130.530 ;
        RECT 14.235 129.520 15.130 130.500 ;
        RECT 11.590 128.415 13.890 128.585 ;
        RECT 14.290 128.585 14.460 129.520 ;
        RECT 14.960 129.490 15.130 129.520 ;
        RECT 15.750 129.490 15.920 130.530 ;
        RECT 14.775 129.105 15.690 129.275 ;
        RECT 14.775 128.900 15.610 129.105 ;
        RECT 16.420 128.585 16.590 131.435 ;
        RECT 14.290 128.415 16.590 128.585 ;
        RECT 16.990 128.585 17.160 140.435 ;
        RECT 17.650 139.725 18.650 140.175 ;
        RECT 17.660 129.490 17.830 139.530 ;
        RECT 18.450 129.490 18.620 139.530 ;
        RECT 17.890 129.105 18.390 129.275 ;
        RECT 19.120 128.585 19.290 140.435 ;
        RECT 16.990 128.415 19.290 128.585 ;
        RECT 19.690 140.435 21.990 140.605 ;
        RECT 19.690 128.585 19.860 140.435 ;
        RECT 20.350 139.725 21.350 140.175 ;
        RECT 20.360 129.490 20.530 139.530 ;
        RECT 21.150 129.490 21.320 139.530 ;
        RECT 20.590 129.105 21.090 129.275 ;
        RECT 21.820 128.585 21.990 140.435 ;
        RECT 22.885 140.435 25.185 140.605 ;
        RECT 22.885 139.450 23.055 140.435 ;
        RECT 23.785 139.745 24.285 139.915 ;
        RECT 23.555 139.450 23.725 139.530 ;
        RECT 24.345 139.525 24.515 139.530 ;
        RECT 22.885 138.575 23.725 139.450 ;
        RECT 22.885 137.585 23.055 138.575 ;
        RECT 23.555 138.490 23.725 138.575 ;
        RECT 24.295 138.495 24.770 139.525 ;
        RECT 24.345 138.490 24.515 138.495 ;
        RECT 23.545 137.850 24.520 138.300 ;
        RECT 25.015 137.585 25.185 140.435 ;
        RECT 22.885 137.415 25.185 137.585 ;
        RECT 25.585 140.435 27.885 140.605 ;
        RECT 25.585 137.585 25.755 140.435 ;
        RECT 26.485 139.745 26.985 139.915 ;
        RECT 26.255 139.525 26.425 139.530 ;
        RECT 25.980 138.495 26.475 139.525 ;
        RECT 27.045 139.500 27.215 139.530 ;
        RECT 27.715 139.500 27.885 140.435 ;
        RECT 28.285 140.435 30.585 140.605 ;
        RECT 28.285 139.500 28.455 140.435 ;
        RECT 29.185 139.745 29.685 139.915 ;
        RECT 28.955 139.500 29.125 139.530 ;
        RECT 26.970 138.570 27.890 139.500 ;
        RECT 26.255 138.490 26.425 138.495 ;
        RECT 27.045 138.490 27.215 138.570 ;
        RECT 26.245 137.850 27.220 138.300 ;
        RECT 27.715 137.585 27.885 138.570 ;
        RECT 28.230 138.520 29.125 139.500 ;
        RECT 25.585 137.415 27.885 137.585 ;
        RECT 28.285 137.585 28.455 138.520 ;
        RECT 28.955 138.490 29.125 138.520 ;
        RECT 29.745 138.490 29.915 139.530 ;
        RECT 28.770 138.105 29.685 138.275 ;
        RECT 28.770 137.900 29.605 138.105 ;
        RECT 30.415 137.585 30.585 140.435 ;
        RECT 28.285 137.415 30.585 137.585 ;
        RECT 34.315 140.435 36.615 140.605 ;
        RECT 22.885 136.345 25.185 136.515 ;
        RECT 22.885 133.935 23.055 136.345 ;
        RECT 23.545 135.675 24.520 136.100 ;
        RECT 25.015 136.035 25.185 136.345 ;
        RECT 25.585 136.345 27.885 136.515 ;
        RECT 25.585 136.035 25.755 136.345 ;
        RECT 23.785 135.655 24.285 135.675 ;
        RECT 23.555 135.480 23.725 135.485 ;
        RECT 24.345 135.480 24.515 135.485 ;
        RECT 23.455 134.800 23.825 135.480 ;
        RECT 24.245 134.800 24.615 135.480 ;
        RECT 23.555 134.795 23.725 134.800 ;
        RECT 24.345 134.795 24.515 134.800 ;
        RECT 23.785 134.455 24.285 134.625 ;
        RECT 25.015 134.245 25.755 136.035 ;
        RECT 26.245 135.675 27.220 136.100 ;
        RECT 26.485 135.655 26.985 135.675 ;
        RECT 26.255 135.480 26.425 135.485 ;
        RECT 26.155 134.800 26.525 135.480 ;
        RECT 27.045 135.405 27.215 135.485 ;
        RECT 27.715 135.405 27.885 136.345 ;
        RECT 28.285 136.345 30.585 136.515 ;
        RECT 28.285 135.405 28.455 136.345 ;
        RECT 28.665 135.655 29.705 136.100 ;
        RECT 28.955 135.405 29.125 135.485 ;
        RECT 26.970 134.825 27.890 135.405 ;
        RECT 28.280 134.875 29.125 135.405 ;
        RECT 26.255 134.795 26.425 134.800 ;
        RECT 27.045 134.795 27.215 134.825 ;
        RECT 26.485 134.455 26.985 134.625 ;
        RECT 25.015 133.935 25.185 134.245 ;
        RECT 22.885 133.765 25.185 133.935 ;
        RECT 25.585 133.935 25.755 134.245 ;
        RECT 27.715 133.935 27.885 134.825 ;
        RECT 25.585 133.765 27.885 133.935 ;
        RECT 28.285 133.935 28.455 134.875 ;
        RECT 28.955 134.795 29.125 134.875 ;
        RECT 29.745 134.795 29.915 135.485 ;
        RECT 29.185 134.455 29.685 134.625 ;
        RECT 30.415 133.935 30.585 136.345 ;
        RECT 28.285 133.765 30.585 133.935 ;
        RECT 31.615 131.435 33.915 131.605 ;
        RECT 31.615 130.500 31.785 131.435 ;
        RECT 32.515 130.745 33.015 130.915 ;
        RECT 32.285 130.500 32.455 130.530 ;
        RECT 31.560 129.520 32.455 130.500 ;
        RECT 19.690 128.415 21.990 128.585 ;
        RECT 31.615 128.585 31.785 129.520 ;
        RECT 32.285 129.490 32.455 129.520 ;
        RECT 33.075 129.490 33.245 130.530 ;
        RECT 32.100 129.105 33.015 129.275 ;
        RECT 32.100 128.900 32.935 129.105 ;
        RECT 33.745 128.585 33.915 131.435 ;
        RECT 31.615 128.415 33.915 128.585 ;
        RECT 34.315 128.585 34.485 140.435 ;
        RECT 34.975 139.725 35.975 140.175 ;
        RECT 34.985 129.490 35.155 139.530 ;
        RECT 35.775 129.490 35.945 139.530 ;
        RECT 35.215 129.105 35.715 129.275 ;
        RECT 36.445 128.585 36.615 140.435 ;
        RECT 42.415 140.435 44.715 140.605 ;
        RECT 37.015 131.435 39.315 131.605 ;
        RECT 37.015 130.500 37.185 131.435 ;
        RECT 37.915 130.745 38.415 130.915 ;
        RECT 37.685 130.500 37.855 130.530 ;
        RECT 36.960 129.520 37.855 130.500 ;
        RECT 34.315 128.415 36.615 128.585 ;
        RECT 37.015 128.585 37.185 129.520 ;
        RECT 37.685 129.490 37.855 129.520 ;
        RECT 38.475 129.490 38.645 130.530 ;
        RECT 37.500 129.105 38.415 129.275 ;
        RECT 37.500 128.900 38.335 129.105 ;
        RECT 39.145 128.585 39.315 131.435 ;
        RECT 39.715 131.435 42.015 131.605 ;
        RECT 39.715 130.500 39.885 131.435 ;
        RECT 40.615 130.745 41.115 130.915 ;
        RECT 40.385 130.500 40.555 130.530 ;
        RECT 39.660 129.520 40.555 130.500 ;
        RECT 37.015 128.415 39.315 128.585 ;
        RECT 39.715 128.585 39.885 129.520 ;
        RECT 40.385 129.490 40.555 129.520 ;
        RECT 41.175 129.490 41.345 130.530 ;
        RECT 40.200 129.105 41.115 129.275 ;
        RECT 40.200 128.900 41.035 129.105 ;
        RECT 41.845 128.585 42.015 131.435 ;
        RECT 39.715 128.415 42.015 128.585 ;
        RECT 42.415 128.585 42.585 140.435 ;
        RECT 43.075 139.725 44.075 140.175 ;
        RECT 43.085 129.490 43.255 139.530 ;
        RECT 43.875 129.490 44.045 139.530 ;
        RECT 43.315 129.105 43.815 129.275 ;
        RECT 44.545 128.585 44.715 140.435 ;
        RECT 42.415 128.415 44.715 128.585 ;
        RECT 45.115 140.435 47.415 140.605 ;
        RECT 45.115 128.585 45.285 140.435 ;
        RECT 45.775 139.725 46.775 140.175 ;
        RECT 45.785 129.490 45.955 139.530 ;
        RECT 46.575 129.490 46.745 139.530 ;
        RECT 46.015 129.105 46.515 129.275 ;
        RECT 47.245 128.585 47.415 140.435 ;
        RECT 59.740 140.435 62.040 140.605 ;
        RECT 57.040 131.435 59.340 131.605 ;
        RECT 57.040 130.500 57.210 131.435 ;
        RECT 57.940 130.745 58.440 130.915 ;
        RECT 57.710 130.500 57.880 130.530 ;
        RECT 56.985 129.520 57.880 130.500 ;
        RECT 45.115 128.415 47.415 128.585 ;
        RECT 57.040 128.585 57.210 129.520 ;
        RECT 57.710 129.490 57.880 129.520 ;
        RECT 58.500 129.490 58.670 130.530 ;
        RECT 57.525 129.105 58.440 129.275 ;
        RECT 57.525 128.900 58.360 129.105 ;
        RECT 59.170 128.585 59.340 131.435 ;
        RECT 57.040 128.415 59.340 128.585 ;
        RECT 59.740 128.585 59.910 140.435 ;
        RECT 60.400 139.725 61.400 140.175 ;
        RECT 60.410 129.490 60.580 139.530 ;
        RECT 61.200 129.490 61.370 139.530 ;
        RECT 60.640 129.105 61.140 129.275 ;
        RECT 61.870 128.585 62.040 140.435 ;
        RECT 67.840 140.435 70.140 140.605 ;
        RECT 62.440 131.435 64.740 131.605 ;
        RECT 62.440 130.500 62.610 131.435 ;
        RECT 63.340 130.745 63.840 130.915 ;
        RECT 63.110 130.500 63.280 130.530 ;
        RECT 62.385 129.520 63.280 130.500 ;
        RECT 59.740 128.415 62.040 128.585 ;
        RECT 62.440 128.585 62.610 129.520 ;
        RECT 63.110 129.490 63.280 129.520 ;
        RECT 63.900 129.490 64.070 130.530 ;
        RECT 62.925 129.105 63.840 129.275 ;
        RECT 62.925 128.900 63.760 129.105 ;
        RECT 64.570 128.585 64.740 131.435 ;
        RECT 65.140 131.435 67.440 131.605 ;
        RECT 65.140 130.500 65.310 131.435 ;
        RECT 66.040 130.745 66.540 130.915 ;
        RECT 65.810 130.500 65.980 130.530 ;
        RECT 65.085 129.520 65.980 130.500 ;
        RECT 62.440 128.415 64.740 128.585 ;
        RECT 65.140 128.585 65.310 129.520 ;
        RECT 65.810 129.490 65.980 129.520 ;
        RECT 66.600 129.490 66.770 130.530 ;
        RECT 65.625 129.105 66.540 129.275 ;
        RECT 65.625 128.900 66.460 129.105 ;
        RECT 67.270 128.585 67.440 131.435 ;
        RECT 65.140 128.415 67.440 128.585 ;
        RECT 67.840 128.585 68.010 140.435 ;
        RECT 68.500 139.725 69.500 140.175 ;
        RECT 68.510 129.490 68.680 139.530 ;
        RECT 69.300 129.490 69.470 139.530 ;
        RECT 68.740 129.105 69.240 129.275 ;
        RECT 69.970 128.585 70.140 140.435 ;
        RECT 67.840 128.415 70.140 128.585 ;
        RECT 70.540 140.435 72.840 140.605 ;
        RECT 70.540 128.585 70.710 140.435 ;
        RECT 71.200 139.725 72.200 140.175 ;
        RECT 71.210 129.490 71.380 139.530 ;
        RECT 72.000 129.490 72.170 139.530 ;
        RECT 71.440 129.105 71.940 129.275 ;
        RECT 72.670 128.585 72.840 140.435 ;
        RECT 73.735 140.435 76.035 140.605 ;
        RECT 73.735 139.450 73.905 140.435 ;
        RECT 74.635 139.745 75.135 139.915 ;
        RECT 74.405 139.450 74.575 139.530 ;
        RECT 75.195 139.525 75.365 139.530 ;
        RECT 73.735 138.575 74.575 139.450 ;
        RECT 73.735 137.585 73.905 138.575 ;
        RECT 74.405 138.490 74.575 138.575 ;
        RECT 75.145 138.495 75.620 139.525 ;
        RECT 75.195 138.490 75.365 138.495 ;
        RECT 74.395 137.850 75.370 138.300 ;
        RECT 75.865 137.585 76.035 140.435 ;
        RECT 73.735 137.415 76.035 137.585 ;
        RECT 76.435 140.435 78.735 140.605 ;
        RECT 76.435 137.585 76.605 140.435 ;
        RECT 77.335 139.745 77.835 139.915 ;
        RECT 77.105 139.525 77.275 139.530 ;
        RECT 76.830 138.495 77.325 139.525 ;
        RECT 77.895 139.500 78.065 139.530 ;
        RECT 78.565 139.500 78.735 140.435 ;
        RECT 79.135 140.435 81.435 140.605 ;
        RECT 79.135 139.500 79.305 140.435 ;
        RECT 80.035 139.745 80.535 139.915 ;
        RECT 79.805 139.500 79.975 139.530 ;
        RECT 77.820 138.570 78.740 139.500 ;
        RECT 77.105 138.490 77.275 138.495 ;
        RECT 77.895 138.490 78.065 138.570 ;
        RECT 77.095 137.850 78.070 138.300 ;
        RECT 78.565 137.585 78.735 138.570 ;
        RECT 79.080 138.520 79.975 139.500 ;
        RECT 76.435 137.415 78.735 137.585 ;
        RECT 79.135 137.585 79.305 138.520 ;
        RECT 79.805 138.490 79.975 138.520 ;
        RECT 80.595 138.490 80.765 139.530 ;
        RECT 79.620 138.105 80.535 138.275 ;
        RECT 79.620 137.900 80.455 138.105 ;
        RECT 81.265 137.585 81.435 140.435 ;
        RECT 79.135 137.415 81.435 137.585 ;
        RECT 85.165 140.435 87.465 140.605 ;
        RECT 73.735 136.345 76.035 136.515 ;
        RECT 73.735 133.935 73.905 136.345 ;
        RECT 74.395 135.675 75.370 136.100 ;
        RECT 75.865 136.035 76.035 136.345 ;
        RECT 76.435 136.345 78.735 136.515 ;
        RECT 76.435 136.035 76.605 136.345 ;
        RECT 74.635 135.655 75.135 135.675 ;
        RECT 74.405 135.480 74.575 135.485 ;
        RECT 75.195 135.480 75.365 135.485 ;
        RECT 74.305 134.800 74.675 135.480 ;
        RECT 75.095 134.800 75.465 135.480 ;
        RECT 74.405 134.795 74.575 134.800 ;
        RECT 75.195 134.795 75.365 134.800 ;
        RECT 74.635 134.455 75.135 134.625 ;
        RECT 75.865 134.245 76.605 136.035 ;
        RECT 77.095 135.675 78.070 136.100 ;
        RECT 77.335 135.655 77.835 135.675 ;
        RECT 77.105 135.480 77.275 135.485 ;
        RECT 77.005 134.800 77.375 135.480 ;
        RECT 77.895 135.405 78.065 135.485 ;
        RECT 78.565 135.405 78.735 136.345 ;
        RECT 79.135 136.345 81.435 136.515 ;
        RECT 79.135 135.405 79.305 136.345 ;
        RECT 79.515 135.655 80.555 136.100 ;
        RECT 79.805 135.405 79.975 135.485 ;
        RECT 77.820 134.825 78.740 135.405 ;
        RECT 79.130 134.875 79.975 135.405 ;
        RECT 77.105 134.795 77.275 134.800 ;
        RECT 77.895 134.795 78.065 134.825 ;
        RECT 77.335 134.455 77.835 134.625 ;
        RECT 75.865 133.935 76.035 134.245 ;
        RECT 73.735 133.765 76.035 133.935 ;
        RECT 76.435 133.935 76.605 134.245 ;
        RECT 78.565 133.935 78.735 134.825 ;
        RECT 76.435 133.765 78.735 133.935 ;
        RECT 79.135 133.935 79.305 134.875 ;
        RECT 79.805 134.795 79.975 134.875 ;
        RECT 80.595 134.795 80.765 135.485 ;
        RECT 80.035 134.455 80.535 134.625 ;
        RECT 81.265 133.935 81.435 136.345 ;
        RECT 79.135 133.765 81.435 133.935 ;
        RECT 82.465 131.435 84.765 131.605 ;
        RECT 82.465 130.500 82.635 131.435 ;
        RECT 83.365 130.745 83.865 130.915 ;
        RECT 83.135 130.500 83.305 130.530 ;
        RECT 82.410 129.520 83.305 130.500 ;
        RECT 70.540 128.415 72.840 128.585 ;
        RECT 82.465 128.585 82.635 129.520 ;
        RECT 83.135 129.490 83.305 129.520 ;
        RECT 83.925 129.490 84.095 130.530 ;
        RECT 82.950 129.105 83.865 129.275 ;
        RECT 82.950 128.900 83.785 129.105 ;
        RECT 84.595 128.585 84.765 131.435 ;
        RECT 82.465 128.415 84.765 128.585 ;
        RECT 85.165 128.585 85.335 140.435 ;
        RECT 85.825 139.725 86.825 140.175 ;
        RECT 85.835 129.490 86.005 139.530 ;
        RECT 86.625 129.490 86.795 139.530 ;
        RECT 86.065 129.105 86.565 129.275 ;
        RECT 87.295 128.585 87.465 140.435 ;
        RECT 93.265 140.435 95.565 140.605 ;
        RECT 87.865 131.435 90.165 131.605 ;
        RECT 87.865 130.500 88.035 131.435 ;
        RECT 88.765 130.745 89.265 130.915 ;
        RECT 88.535 130.500 88.705 130.530 ;
        RECT 87.810 129.520 88.705 130.500 ;
        RECT 85.165 128.415 87.465 128.585 ;
        RECT 87.865 128.585 88.035 129.520 ;
        RECT 88.535 129.490 88.705 129.520 ;
        RECT 89.325 129.490 89.495 130.530 ;
        RECT 88.350 129.105 89.265 129.275 ;
        RECT 88.350 128.900 89.185 129.105 ;
        RECT 89.995 128.585 90.165 131.435 ;
        RECT 90.565 131.435 92.865 131.605 ;
        RECT 90.565 130.500 90.735 131.435 ;
        RECT 91.465 130.745 91.965 130.915 ;
        RECT 91.235 130.500 91.405 130.530 ;
        RECT 90.510 129.520 91.405 130.500 ;
        RECT 87.865 128.415 90.165 128.585 ;
        RECT 90.565 128.585 90.735 129.520 ;
        RECT 91.235 129.490 91.405 129.520 ;
        RECT 92.025 129.490 92.195 130.530 ;
        RECT 91.050 129.105 91.965 129.275 ;
        RECT 91.050 128.900 91.885 129.105 ;
        RECT 92.695 128.585 92.865 131.435 ;
        RECT 90.565 128.415 92.865 128.585 ;
        RECT 93.265 128.585 93.435 140.435 ;
        RECT 93.925 139.725 94.925 140.175 ;
        RECT 93.935 129.490 94.105 139.530 ;
        RECT 94.725 129.490 94.895 139.530 ;
        RECT 94.165 129.105 94.665 129.275 ;
        RECT 95.395 128.585 95.565 140.435 ;
        RECT 93.265 128.415 95.565 128.585 ;
        RECT 95.965 140.435 98.265 140.605 ;
        RECT 95.965 128.585 96.135 140.435 ;
        RECT 96.625 139.725 97.625 140.175 ;
        RECT 96.635 129.490 96.805 139.530 ;
        RECT 97.425 129.490 97.595 139.530 ;
        RECT 96.865 129.105 97.365 129.275 ;
        RECT 98.095 128.585 98.265 140.435 ;
        RECT 110.590 140.435 112.890 140.605 ;
        RECT 107.890 131.435 110.190 131.605 ;
        RECT 107.890 130.500 108.060 131.435 ;
        RECT 108.790 130.745 109.290 130.915 ;
        RECT 108.560 130.500 108.730 130.530 ;
        RECT 107.835 129.520 108.730 130.500 ;
        RECT 95.965 128.415 98.265 128.585 ;
        RECT 107.890 128.585 108.060 129.520 ;
        RECT 108.560 129.490 108.730 129.520 ;
        RECT 109.350 129.490 109.520 130.530 ;
        RECT 108.375 129.105 109.290 129.275 ;
        RECT 108.375 128.900 109.210 129.105 ;
        RECT 110.020 128.585 110.190 131.435 ;
        RECT 107.890 128.415 110.190 128.585 ;
        RECT 110.590 128.585 110.760 140.435 ;
        RECT 111.250 139.725 112.250 140.175 ;
        RECT 111.260 129.490 111.430 139.530 ;
        RECT 112.050 129.490 112.220 139.530 ;
        RECT 111.490 129.105 111.990 129.275 ;
        RECT 112.720 128.585 112.890 140.435 ;
        RECT 118.690 140.435 120.990 140.605 ;
        RECT 113.290 131.435 115.590 131.605 ;
        RECT 113.290 130.500 113.460 131.435 ;
        RECT 114.190 130.745 114.690 130.915 ;
        RECT 113.960 130.500 114.130 130.530 ;
        RECT 113.235 129.520 114.130 130.500 ;
        RECT 110.590 128.415 112.890 128.585 ;
        RECT 113.290 128.585 113.460 129.520 ;
        RECT 113.960 129.490 114.130 129.520 ;
        RECT 114.750 129.490 114.920 130.530 ;
        RECT 113.775 129.105 114.690 129.275 ;
        RECT 113.775 128.900 114.610 129.105 ;
        RECT 115.420 128.585 115.590 131.435 ;
        RECT 115.990 131.435 118.290 131.605 ;
        RECT 115.990 130.500 116.160 131.435 ;
        RECT 116.890 130.745 117.390 130.915 ;
        RECT 116.660 130.500 116.830 130.530 ;
        RECT 115.935 129.520 116.830 130.500 ;
        RECT 113.290 128.415 115.590 128.585 ;
        RECT 115.990 128.585 116.160 129.520 ;
        RECT 116.660 129.490 116.830 129.520 ;
        RECT 117.450 129.490 117.620 130.530 ;
        RECT 116.475 129.105 117.390 129.275 ;
        RECT 116.475 128.900 117.310 129.105 ;
        RECT 118.120 128.585 118.290 131.435 ;
        RECT 115.990 128.415 118.290 128.585 ;
        RECT 118.690 128.585 118.860 140.435 ;
        RECT 119.350 139.725 120.350 140.175 ;
        RECT 119.360 129.490 119.530 139.530 ;
        RECT 120.150 129.490 120.320 139.530 ;
        RECT 119.590 129.105 120.090 129.275 ;
        RECT 120.820 128.585 120.990 140.435 ;
        RECT 118.690 128.415 120.990 128.585 ;
        RECT 121.390 140.435 123.690 140.605 ;
        RECT 121.390 128.585 121.560 140.435 ;
        RECT 122.050 139.725 123.050 140.175 ;
        RECT 122.060 129.490 122.230 139.530 ;
        RECT 122.850 129.490 123.020 139.530 ;
        RECT 122.290 129.105 122.790 129.275 ;
        RECT 123.520 128.585 123.690 140.435 ;
        RECT 124.585 140.435 126.885 140.605 ;
        RECT 124.585 139.450 124.755 140.435 ;
        RECT 125.485 139.745 125.985 139.915 ;
        RECT 125.255 139.450 125.425 139.530 ;
        RECT 126.045 139.525 126.215 139.530 ;
        RECT 124.585 138.575 125.425 139.450 ;
        RECT 124.585 137.585 124.755 138.575 ;
        RECT 125.255 138.490 125.425 138.575 ;
        RECT 125.995 138.495 126.470 139.525 ;
        RECT 126.045 138.490 126.215 138.495 ;
        RECT 125.245 137.850 126.220 138.300 ;
        RECT 126.715 137.585 126.885 140.435 ;
        RECT 124.585 137.415 126.885 137.585 ;
        RECT 127.285 140.435 129.585 140.605 ;
        RECT 127.285 137.585 127.455 140.435 ;
        RECT 128.185 139.745 128.685 139.915 ;
        RECT 127.955 139.525 128.125 139.530 ;
        RECT 127.680 138.495 128.175 139.525 ;
        RECT 128.745 139.500 128.915 139.530 ;
        RECT 129.415 139.500 129.585 140.435 ;
        RECT 129.985 140.435 132.285 140.605 ;
        RECT 129.985 139.500 130.155 140.435 ;
        RECT 130.885 139.745 131.385 139.915 ;
        RECT 130.655 139.500 130.825 139.530 ;
        RECT 128.670 138.570 129.590 139.500 ;
        RECT 127.955 138.490 128.125 138.495 ;
        RECT 128.745 138.490 128.915 138.570 ;
        RECT 127.945 137.850 128.920 138.300 ;
        RECT 129.415 137.585 129.585 138.570 ;
        RECT 129.930 138.520 130.825 139.500 ;
        RECT 127.285 137.415 129.585 137.585 ;
        RECT 129.985 137.585 130.155 138.520 ;
        RECT 130.655 138.490 130.825 138.520 ;
        RECT 131.445 138.490 131.615 139.530 ;
        RECT 130.470 138.105 131.385 138.275 ;
        RECT 130.470 137.900 131.305 138.105 ;
        RECT 132.115 137.585 132.285 140.435 ;
        RECT 129.985 137.415 132.285 137.585 ;
        RECT 136.015 140.435 138.315 140.605 ;
        RECT 124.585 136.345 126.885 136.515 ;
        RECT 124.585 133.935 124.755 136.345 ;
        RECT 125.245 135.675 126.220 136.100 ;
        RECT 126.715 136.035 126.885 136.345 ;
        RECT 127.285 136.345 129.585 136.515 ;
        RECT 127.285 136.035 127.455 136.345 ;
        RECT 125.485 135.655 125.985 135.675 ;
        RECT 125.255 135.480 125.425 135.485 ;
        RECT 126.045 135.480 126.215 135.485 ;
        RECT 125.155 134.800 125.525 135.480 ;
        RECT 125.945 134.800 126.315 135.480 ;
        RECT 125.255 134.795 125.425 134.800 ;
        RECT 126.045 134.795 126.215 134.800 ;
        RECT 125.485 134.455 125.985 134.625 ;
        RECT 126.715 134.245 127.455 136.035 ;
        RECT 127.945 135.675 128.920 136.100 ;
        RECT 128.185 135.655 128.685 135.675 ;
        RECT 127.955 135.480 128.125 135.485 ;
        RECT 127.855 134.800 128.225 135.480 ;
        RECT 128.745 135.405 128.915 135.485 ;
        RECT 129.415 135.405 129.585 136.345 ;
        RECT 129.985 136.345 132.285 136.515 ;
        RECT 129.985 135.405 130.155 136.345 ;
        RECT 130.365 135.655 131.405 136.100 ;
        RECT 130.655 135.405 130.825 135.485 ;
        RECT 128.670 134.825 129.590 135.405 ;
        RECT 129.980 134.875 130.825 135.405 ;
        RECT 127.955 134.795 128.125 134.800 ;
        RECT 128.745 134.795 128.915 134.825 ;
        RECT 128.185 134.455 128.685 134.625 ;
        RECT 126.715 133.935 126.885 134.245 ;
        RECT 124.585 133.765 126.885 133.935 ;
        RECT 127.285 133.935 127.455 134.245 ;
        RECT 129.415 133.935 129.585 134.825 ;
        RECT 127.285 133.765 129.585 133.935 ;
        RECT 129.985 133.935 130.155 134.875 ;
        RECT 130.655 134.795 130.825 134.875 ;
        RECT 131.445 134.795 131.615 135.485 ;
        RECT 130.885 134.455 131.385 134.625 ;
        RECT 132.115 133.935 132.285 136.345 ;
        RECT 129.985 133.765 132.285 133.935 ;
        RECT 133.315 131.435 135.615 131.605 ;
        RECT 133.315 130.500 133.485 131.435 ;
        RECT 134.215 130.745 134.715 130.915 ;
        RECT 133.985 130.500 134.155 130.530 ;
        RECT 133.260 129.520 134.155 130.500 ;
        RECT 121.390 128.415 123.690 128.585 ;
        RECT 133.315 128.585 133.485 129.520 ;
        RECT 133.985 129.490 134.155 129.520 ;
        RECT 134.775 129.490 134.945 130.530 ;
        RECT 133.800 129.105 134.715 129.275 ;
        RECT 133.800 128.900 134.635 129.105 ;
        RECT 135.445 128.585 135.615 131.435 ;
        RECT 133.315 128.415 135.615 128.585 ;
        RECT 136.015 128.585 136.185 140.435 ;
        RECT 136.675 139.725 137.675 140.175 ;
        RECT 136.685 129.490 136.855 139.530 ;
        RECT 137.475 129.490 137.645 139.530 ;
        RECT 136.915 129.105 137.415 129.275 ;
        RECT 138.145 128.585 138.315 140.435 ;
        RECT 144.115 140.435 146.415 140.605 ;
        RECT 138.715 131.435 141.015 131.605 ;
        RECT 138.715 130.500 138.885 131.435 ;
        RECT 139.615 130.745 140.115 130.915 ;
        RECT 139.385 130.500 139.555 130.530 ;
        RECT 138.660 129.520 139.555 130.500 ;
        RECT 136.015 128.415 138.315 128.585 ;
        RECT 138.715 128.585 138.885 129.520 ;
        RECT 139.385 129.490 139.555 129.520 ;
        RECT 140.175 129.490 140.345 130.530 ;
        RECT 139.200 129.105 140.115 129.275 ;
        RECT 139.200 128.900 140.035 129.105 ;
        RECT 140.845 128.585 141.015 131.435 ;
        RECT 141.415 131.435 143.715 131.605 ;
        RECT 141.415 130.500 141.585 131.435 ;
        RECT 142.315 130.745 142.815 130.915 ;
        RECT 142.085 130.500 142.255 130.530 ;
        RECT 141.360 129.520 142.255 130.500 ;
        RECT 138.715 128.415 141.015 128.585 ;
        RECT 141.415 128.585 141.585 129.520 ;
        RECT 142.085 129.490 142.255 129.520 ;
        RECT 142.875 129.490 143.045 130.530 ;
        RECT 141.900 129.105 142.815 129.275 ;
        RECT 141.900 128.900 142.735 129.105 ;
        RECT 143.545 128.585 143.715 131.435 ;
        RECT 141.415 128.415 143.715 128.585 ;
        RECT 144.115 128.585 144.285 140.435 ;
        RECT 144.775 139.725 145.775 140.175 ;
        RECT 144.785 129.490 144.955 139.530 ;
        RECT 145.575 129.490 145.745 139.530 ;
        RECT 145.015 129.105 145.515 129.275 ;
        RECT 146.245 128.585 146.415 140.435 ;
        RECT 144.115 128.415 146.415 128.585 ;
        RECT 146.815 140.435 149.115 140.605 ;
        RECT 146.815 128.585 146.985 140.435 ;
        RECT 147.475 139.725 148.475 140.175 ;
        RECT 147.485 129.490 147.655 139.530 ;
        RECT 148.275 129.490 148.445 139.530 ;
        RECT 147.715 129.105 148.215 129.275 ;
        RECT 148.945 128.585 149.115 140.435 ;
        RECT 146.815 128.415 149.115 128.585 ;
        RECT 6.190 127.345 8.490 127.515 ;
        RECT 6.190 126.405 6.360 127.345 ;
        RECT 6.570 126.655 7.610 127.100 ;
        RECT 6.860 126.405 7.030 126.485 ;
        RECT 6.185 125.875 7.030 126.405 ;
        RECT 6.190 124.935 6.360 125.875 ;
        RECT 6.860 125.795 7.030 125.875 ;
        RECT 7.650 125.795 7.820 126.485 ;
        RECT 7.090 125.455 7.590 125.625 ;
        RECT 8.320 124.935 8.490 127.345 ;
        RECT 6.190 124.765 8.490 124.935 ;
        RECT 8.890 127.345 11.190 127.515 ;
        RECT 8.890 119.085 9.060 127.345 ;
        RECT 9.790 126.655 10.290 126.825 ;
        RECT 9.560 119.945 9.730 126.485 ;
        RECT 10.350 119.945 10.520 126.485 ;
        RECT 9.550 119.375 10.550 119.775 ;
        RECT 11.020 119.085 11.190 127.345 ;
        RECT 11.590 127.345 13.890 127.515 ;
        RECT 11.590 126.405 11.760 127.345 ;
        RECT 11.970 126.655 13.010 127.100 ;
        RECT 12.260 126.405 12.430 126.485 ;
        RECT 11.585 125.875 12.430 126.405 ;
        RECT 11.590 124.935 11.760 125.875 ;
        RECT 12.260 125.795 12.430 125.875 ;
        RECT 13.050 125.795 13.220 126.485 ;
        RECT 12.490 125.455 12.990 125.625 ;
        RECT 13.720 124.935 13.890 127.345 ;
        RECT 14.290 127.345 16.590 127.515 ;
        RECT 14.290 126.405 14.460 127.345 ;
        RECT 14.670 126.655 15.710 127.100 ;
        RECT 14.960 126.405 15.130 126.485 ;
        RECT 14.285 125.875 15.130 126.405 ;
        RECT 11.590 124.765 13.890 124.935 ;
        RECT 14.290 124.935 14.460 125.875 ;
        RECT 14.960 125.795 15.130 125.875 ;
        RECT 15.750 125.795 15.920 126.485 ;
        RECT 15.190 125.455 15.690 125.625 ;
        RECT 16.420 124.935 16.590 127.345 ;
        RECT 14.290 124.765 16.590 124.935 ;
        RECT 16.990 127.345 19.290 127.515 ;
        RECT 8.890 118.915 11.190 119.085 ;
        RECT 16.990 119.085 17.160 127.345 ;
        RECT 17.890 126.655 18.390 126.825 ;
        RECT 17.660 119.945 17.830 126.485 ;
        RECT 18.450 119.945 18.620 126.485 ;
        RECT 17.650 119.375 18.650 119.775 ;
        RECT 19.120 119.085 19.290 127.345 ;
        RECT 16.990 118.915 19.290 119.085 ;
        RECT 19.690 127.345 21.990 127.515 ;
        RECT 19.690 119.085 19.860 127.345 ;
        RECT 20.590 126.655 21.090 126.825 ;
        RECT 20.360 119.945 20.530 126.485 ;
        RECT 21.150 119.945 21.320 126.485 ;
        RECT 20.350 119.375 21.350 119.775 ;
        RECT 21.820 119.085 21.990 127.345 ;
        RECT 31.615 127.345 33.915 127.515 ;
        RECT 31.615 126.405 31.785 127.345 ;
        RECT 31.995 126.655 33.035 127.100 ;
        RECT 32.285 126.405 32.455 126.485 ;
        RECT 31.610 125.875 32.455 126.405 ;
        RECT 31.615 124.935 31.785 125.875 ;
        RECT 32.285 125.795 32.455 125.875 ;
        RECT 33.075 125.795 33.245 126.485 ;
        RECT 32.515 125.455 33.015 125.625 ;
        RECT 33.745 124.935 33.915 127.345 ;
        RECT 31.615 124.765 33.915 124.935 ;
        RECT 34.315 127.345 36.615 127.515 ;
        RECT 19.690 118.915 21.990 119.085 ;
        RECT 34.315 119.085 34.485 127.345 ;
        RECT 35.215 126.655 35.715 126.825 ;
        RECT 34.985 119.945 35.155 126.485 ;
        RECT 35.775 119.945 35.945 126.485 ;
        RECT 34.975 119.375 35.975 119.775 ;
        RECT 36.445 119.085 36.615 127.345 ;
        RECT 37.015 127.345 39.315 127.515 ;
        RECT 37.015 126.405 37.185 127.345 ;
        RECT 37.395 126.655 38.435 127.100 ;
        RECT 37.685 126.405 37.855 126.485 ;
        RECT 37.010 125.875 37.855 126.405 ;
        RECT 37.015 124.935 37.185 125.875 ;
        RECT 37.685 125.795 37.855 125.875 ;
        RECT 38.475 125.795 38.645 126.485 ;
        RECT 37.915 125.455 38.415 125.625 ;
        RECT 39.145 124.935 39.315 127.345 ;
        RECT 39.715 127.345 42.015 127.515 ;
        RECT 39.715 126.405 39.885 127.345 ;
        RECT 40.095 126.655 41.135 127.100 ;
        RECT 40.385 126.405 40.555 126.485 ;
        RECT 39.710 125.875 40.555 126.405 ;
        RECT 37.015 124.765 39.315 124.935 ;
        RECT 39.715 124.935 39.885 125.875 ;
        RECT 40.385 125.795 40.555 125.875 ;
        RECT 41.175 125.795 41.345 126.485 ;
        RECT 40.615 125.455 41.115 125.625 ;
        RECT 41.845 124.935 42.015 127.345 ;
        RECT 39.715 124.765 42.015 124.935 ;
        RECT 42.415 127.345 44.715 127.515 ;
        RECT 34.315 118.915 36.615 119.085 ;
        RECT 42.415 119.085 42.585 127.345 ;
        RECT 43.315 126.655 43.815 126.825 ;
        RECT 43.085 119.945 43.255 126.485 ;
        RECT 43.875 119.945 44.045 126.485 ;
        RECT 43.075 119.375 44.075 119.775 ;
        RECT 44.545 119.085 44.715 127.345 ;
        RECT 42.415 118.915 44.715 119.085 ;
        RECT 45.115 127.345 47.415 127.515 ;
        RECT 45.115 119.085 45.285 127.345 ;
        RECT 46.015 126.655 46.515 126.825 ;
        RECT 45.785 119.945 45.955 126.485 ;
        RECT 46.575 119.945 46.745 126.485 ;
        RECT 45.775 119.375 46.775 119.775 ;
        RECT 47.245 119.085 47.415 127.345 ;
        RECT 57.040 127.345 59.340 127.515 ;
        RECT 57.040 126.405 57.210 127.345 ;
        RECT 57.420 126.655 58.460 127.100 ;
        RECT 57.710 126.405 57.880 126.485 ;
        RECT 57.035 125.875 57.880 126.405 ;
        RECT 57.040 124.935 57.210 125.875 ;
        RECT 57.710 125.795 57.880 125.875 ;
        RECT 58.500 125.795 58.670 126.485 ;
        RECT 57.940 125.455 58.440 125.625 ;
        RECT 59.170 124.935 59.340 127.345 ;
        RECT 57.040 124.765 59.340 124.935 ;
        RECT 59.740 127.345 62.040 127.515 ;
        RECT 45.115 118.915 47.415 119.085 ;
        RECT 59.740 119.085 59.910 127.345 ;
        RECT 60.640 126.655 61.140 126.825 ;
        RECT 60.410 119.945 60.580 126.485 ;
        RECT 61.200 119.945 61.370 126.485 ;
        RECT 60.400 119.375 61.400 119.775 ;
        RECT 61.870 119.085 62.040 127.345 ;
        RECT 62.440 127.345 64.740 127.515 ;
        RECT 62.440 126.405 62.610 127.345 ;
        RECT 62.820 126.655 63.860 127.100 ;
        RECT 63.110 126.405 63.280 126.485 ;
        RECT 62.435 125.875 63.280 126.405 ;
        RECT 62.440 124.935 62.610 125.875 ;
        RECT 63.110 125.795 63.280 125.875 ;
        RECT 63.900 125.795 64.070 126.485 ;
        RECT 63.340 125.455 63.840 125.625 ;
        RECT 64.570 124.935 64.740 127.345 ;
        RECT 65.140 127.345 67.440 127.515 ;
        RECT 65.140 126.405 65.310 127.345 ;
        RECT 65.520 126.655 66.560 127.100 ;
        RECT 65.810 126.405 65.980 126.485 ;
        RECT 65.135 125.875 65.980 126.405 ;
        RECT 62.440 124.765 64.740 124.935 ;
        RECT 65.140 124.935 65.310 125.875 ;
        RECT 65.810 125.795 65.980 125.875 ;
        RECT 66.600 125.795 66.770 126.485 ;
        RECT 66.040 125.455 66.540 125.625 ;
        RECT 67.270 124.935 67.440 127.345 ;
        RECT 65.140 124.765 67.440 124.935 ;
        RECT 67.840 127.345 70.140 127.515 ;
        RECT 59.740 118.915 62.040 119.085 ;
        RECT 67.840 119.085 68.010 127.345 ;
        RECT 68.740 126.655 69.240 126.825 ;
        RECT 68.510 119.945 68.680 126.485 ;
        RECT 69.300 119.945 69.470 126.485 ;
        RECT 68.500 119.375 69.500 119.775 ;
        RECT 69.970 119.085 70.140 127.345 ;
        RECT 67.840 118.915 70.140 119.085 ;
        RECT 70.540 127.345 72.840 127.515 ;
        RECT 70.540 119.085 70.710 127.345 ;
        RECT 71.440 126.655 71.940 126.825 ;
        RECT 71.210 119.945 71.380 126.485 ;
        RECT 72.000 119.945 72.170 126.485 ;
        RECT 71.200 119.375 72.200 119.775 ;
        RECT 72.670 119.085 72.840 127.345 ;
        RECT 82.465 127.345 84.765 127.515 ;
        RECT 82.465 126.405 82.635 127.345 ;
        RECT 82.845 126.655 83.885 127.100 ;
        RECT 83.135 126.405 83.305 126.485 ;
        RECT 82.460 125.875 83.305 126.405 ;
        RECT 82.465 124.935 82.635 125.875 ;
        RECT 83.135 125.795 83.305 125.875 ;
        RECT 83.925 125.795 84.095 126.485 ;
        RECT 83.365 125.455 83.865 125.625 ;
        RECT 84.595 124.935 84.765 127.345 ;
        RECT 82.465 124.765 84.765 124.935 ;
        RECT 85.165 127.345 87.465 127.515 ;
        RECT 70.540 118.915 72.840 119.085 ;
        RECT 85.165 119.085 85.335 127.345 ;
        RECT 86.065 126.655 86.565 126.825 ;
        RECT 85.835 119.945 86.005 126.485 ;
        RECT 86.625 119.945 86.795 126.485 ;
        RECT 85.825 119.375 86.825 119.775 ;
        RECT 87.295 119.085 87.465 127.345 ;
        RECT 87.865 127.345 90.165 127.515 ;
        RECT 87.865 126.405 88.035 127.345 ;
        RECT 88.245 126.655 89.285 127.100 ;
        RECT 88.535 126.405 88.705 126.485 ;
        RECT 87.860 125.875 88.705 126.405 ;
        RECT 87.865 124.935 88.035 125.875 ;
        RECT 88.535 125.795 88.705 125.875 ;
        RECT 89.325 125.795 89.495 126.485 ;
        RECT 88.765 125.455 89.265 125.625 ;
        RECT 89.995 124.935 90.165 127.345 ;
        RECT 90.565 127.345 92.865 127.515 ;
        RECT 90.565 126.405 90.735 127.345 ;
        RECT 90.945 126.655 91.985 127.100 ;
        RECT 91.235 126.405 91.405 126.485 ;
        RECT 90.560 125.875 91.405 126.405 ;
        RECT 87.865 124.765 90.165 124.935 ;
        RECT 90.565 124.935 90.735 125.875 ;
        RECT 91.235 125.795 91.405 125.875 ;
        RECT 92.025 125.795 92.195 126.485 ;
        RECT 91.465 125.455 91.965 125.625 ;
        RECT 92.695 124.935 92.865 127.345 ;
        RECT 90.565 124.765 92.865 124.935 ;
        RECT 93.265 127.345 95.565 127.515 ;
        RECT 85.165 118.915 87.465 119.085 ;
        RECT 93.265 119.085 93.435 127.345 ;
        RECT 94.165 126.655 94.665 126.825 ;
        RECT 93.935 119.945 94.105 126.485 ;
        RECT 94.725 119.945 94.895 126.485 ;
        RECT 93.925 119.375 94.925 119.775 ;
        RECT 95.395 119.085 95.565 127.345 ;
        RECT 93.265 118.915 95.565 119.085 ;
        RECT 95.965 127.345 98.265 127.515 ;
        RECT 95.965 119.085 96.135 127.345 ;
        RECT 96.865 126.655 97.365 126.825 ;
        RECT 96.635 119.945 96.805 126.485 ;
        RECT 97.425 119.945 97.595 126.485 ;
        RECT 96.625 119.375 97.625 119.775 ;
        RECT 98.095 119.085 98.265 127.345 ;
        RECT 107.890 127.345 110.190 127.515 ;
        RECT 107.890 126.405 108.060 127.345 ;
        RECT 108.270 126.655 109.310 127.100 ;
        RECT 108.560 126.405 108.730 126.485 ;
        RECT 107.885 125.875 108.730 126.405 ;
        RECT 107.890 124.935 108.060 125.875 ;
        RECT 108.560 125.795 108.730 125.875 ;
        RECT 109.350 125.795 109.520 126.485 ;
        RECT 108.790 125.455 109.290 125.625 ;
        RECT 110.020 124.935 110.190 127.345 ;
        RECT 107.890 124.765 110.190 124.935 ;
        RECT 110.590 127.345 112.890 127.515 ;
        RECT 95.965 118.915 98.265 119.085 ;
        RECT 110.590 119.085 110.760 127.345 ;
        RECT 111.490 126.655 111.990 126.825 ;
        RECT 111.260 119.945 111.430 126.485 ;
        RECT 112.050 119.945 112.220 126.485 ;
        RECT 111.250 119.375 112.250 119.775 ;
        RECT 112.720 119.085 112.890 127.345 ;
        RECT 113.290 127.345 115.590 127.515 ;
        RECT 113.290 126.405 113.460 127.345 ;
        RECT 113.670 126.655 114.710 127.100 ;
        RECT 113.960 126.405 114.130 126.485 ;
        RECT 113.285 125.875 114.130 126.405 ;
        RECT 113.290 124.935 113.460 125.875 ;
        RECT 113.960 125.795 114.130 125.875 ;
        RECT 114.750 125.795 114.920 126.485 ;
        RECT 114.190 125.455 114.690 125.625 ;
        RECT 115.420 124.935 115.590 127.345 ;
        RECT 115.990 127.345 118.290 127.515 ;
        RECT 115.990 126.405 116.160 127.345 ;
        RECT 116.370 126.655 117.410 127.100 ;
        RECT 116.660 126.405 116.830 126.485 ;
        RECT 115.985 125.875 116.830 126.405 ;
        RECT 113.290 124.765 115.590 124.935 ;
        RECT 115.990 124.935 116.160 125.875 ;
        RECT 116.660 125.795 116.830 125.875 ;
        RECT 117.450 125.795 117.620 126.485 ;
        RECT 116.890 125.455 117.390 125.625 ;
        RECT 118.120 124.935 118.290 127.345 ;
        RECT 115.990 124.765 118.290 124.935 ;
        RECT 118.690 127.345 120.990 127.515 ;
        RECT 110.590 118.915 112.890 119.085 ;
        RECT 118.690 119.085 118.860 127.345 ;
        RECT 119.590 126.655 120.090 126.825 ;
        RECT 119.360 119.945 119.530 126.485 ;
        RECT 120.150 119.945 120.320 126.485 ;
        RECT 119.350 119.375 120.350 119.775 ;
        RECT 120.820 119.085 120.990 127.345 ;
        RECT 118.690 118.915 120.990 119.085 ;
        RECT 121.390 127.345 123.690 127.515 ;
        RECT 121.390 119.085 121.560 127.345 ;
        RECT 122.290 126.655 122.790 126.825 ;
        RECT 122.060 119.945 122.230 126.485 ;
        RECT 122.850 119.945 123.020 126.485 ;
        RECT 122.050 119.375 123.050 119.775 ;
        RECT 123.520 119.085 123.690 127.345 ;
        RECT 133.315 127.345 135.615 127.515 ;
        RECT 133.315 126.405 133.485 127.345 ;
        RECT 133.695 126.655 134.735 127.100 ;
        RECT 133.985 126.405 134.155 126.485 ;
        RECT 133.310 125.875 134.155 126.405 ;
        RECT 133.315 124.935 133.485 125.875 ;
        RECT 133.985 125.795 134.155 125.875 ;
        RECT 134.775 125.795 134.945 126.485 ;
        RECT 134.215 125.455 134.715 125.625 ;
        RECT 135.445 124.935 135.615 127.345 ;
        RECT 133.315 124.765 135.615 124.935 ;
        RECT 136.015 127.345 138.315 127.515 ;
        RECT 121.390 118.915 123.690 119.085 ;
        RECT 136.015 119.085 136.185 127.345 ;
        RECT 136.915 126.655 137.415 126.825 ;
        RECT 136.685 119.945 136.855 126.485 ;
        RECT 137.475 119.945 137.645 126.485 ;
        RECT 136.675 119.375 137.675 119.775 ;
        RECT 138.145 119.085 138.315 127.345 ;
        RECT 138.715 127.345 141.015 127.515 ;
        RECT 138.715 126.405 138.885 127.345 ;
        RECT 139.095 126.655 140.135 127.100 ;
        RECT 139.385 126.405 139.555 126.485 ;
        RECT 138.710 125.875 139.555 126.405 ;
        RECT 138.715 124.935 138.885 125.875 ;
        RECT 139.385 125.795 139.555 125.875 ;
        RECT 140.175 125.795 140.345 126.485 ;
        RECT 139.615 125.455 140.115 125.625 ;
        RECT 140.845 124.935 141.015 127.345 ;
        RECT 141.415 127.345 143.715 127.515 ;
        RECT 141.415 126.405 141.585 127.345 ;
        RECT 141.795 126.655 142.835 127.100 ;
        RECT 142.085 126.405 142.255 126.485 ;
        RECT 141.410 125.875 142.255 126.405 ;
        RECT 138.715 124.765 141.015 124.935 ;
        RECT 141.415 124.935 141.585 125.875 ;
        RECT 142.085 125.795 142.255 125.875 ;
        RECT 142.875 125.795 143.045 126.485 ;
        RECT 142.315 125.455 142.815 125.625 ;
        RECT 143.545 124.935 143.715 127.345 ;
        RECT 141.415 124.765 143.715 124.935 ;
        RECT 144.115 127.345 146.415 127.515 ;
        RECT 136.015 118.915 138.315 119.085 ;
        RECT 144.115 119.085 144.285 127.345 ;
        RECT 145.015 126.655 145.515 126.825 ;
        RECT 144.785 119.945 144.955 126.485 ;
        RECT 145.575 119.945 145.745 126.485 ;
        RECT 144.775 119.375 145.775 119.775 ;
        RECT 146.245 119.085 146.415 127.345 ;
        RECT 144.115 118.915 146.415 119.085 ;
        RECT 146.815 127.345 149.115 127.515 ;
        RECT 146.815 119.085 146.985 127.345 ;
        RECT 147.715 126.655 148.215 126.825 ;
        RECT 147.485 119.945 147.655 126.485 ;
        RECT 148.275 119.945 148.445 126.485 ;
        RECT 147.475 119.375 148.475 119.775 ;
        RECT 148.945 119.085 149.115 127.345 ;
        RECT 146.815 118.915 149.115 119.085 ;
        RECT 8.890 117.860 11.190 118.030 ;
        RECT 6.190 108.860 8.490 109.030 ;
        RECT 6.190 107.925 6.360 108.860 ;
        RECT 7.090 108.170 7.590 108.340 ;
        RECT 6.860 107.925 7.030 107.955 ;
        RECT 6.135 106.945 7.030 107.925 ;
        RECT 6.190 106.010 6.360 106.945 ;
        RECT 6.860 106.915 7.030 106.945 ;
        RECT 7.650 106.915 7.820 107.955 ;
        RECT 6.675 106.530 7.590 106.700 ;
        RECT 6.675 106.325 7.510 106.530 ;
        RECT 8.320 106.010 8.490 108.860 ;
        RECT 6.190 105.840 8.490 106.010 ;
        RECT 8.890 106.010 9.060 117.860 ;
        RECT 9.550 117.150 10.550 117.600 ;
        RECT 9.560 106.915 9.730 116.955 ;
        RECT 10.350 106.915 10.520 116.955 ;
        RECT 9.790 106.530 10.290 106.700 ;
        RECT 11.020 106.010 11.190 117.860 ;
        RECT 16.990 117.860 19.290 118.030 ;
        RECT 11.590 108.860 13.890 109.030 ;
        RECT 11.590 107.925 11.760 108.860 ;
        RECT 12.490 108.170 12.990 108.340 ;
        RECT 12.260 107.925 12.430 107.955 ;
        RECT 11.535 106.945 12.430 107.925 ;
        RECT 8.890 105.840 11.190 106.010 ;
        RECT 11.590 106.010 11.760 106.945 ;
        RECT 12.260 106.915 12.430 106.945 ;
        RECT 13.050 106.915 13.220 107.955 ;
        RECT 12.075 106.530 12.990 106.700 ;
        RECT 12.075 106.325 12.910 106.530 ;
        RECT 13.720 106.010 13.890 108.860 ;
        RECT 14.290 108.860 16.590 109.030 ;
        RECT 14.290 107.925 14.460 108.860 ;
        RECT 15.190 108.170 15.690 108.340 ;
        RECT 14.960 107.925 15.130 107.955 ;
        RECT 14.235 106.945 15.130 107.925 ;
        RECT 11.590 105.840 13.890 106.010 ;
        RECT 14.290 106.010 14.460 106.945 ;
        RECT 14.960 106.915 15.130 106.945 ;
        RECT 15.750 106.915 15.920 107.955 ;
        RECT 14.775 106.530 15.690 106.700 ;
        RECT 14.775 106.325 15.610 106.530 ;
        RECT 16.420 106.010 16.590 108.860 ;
        RECT 14.290 105.840 16.590 106.010 ;
        RECT 16.990 106.010 17.160 117.860 ;
        RECT 17.650 117.150 18.650 117.600 ;
        RECT 17.660 106.915 17.830 116.955 ;
        RECT 18.450 106.915 18.620 116.955 ;
        RECT 17.890 106.530 18.390 106.700 ;
        RECT 19.120 106.010 19.290 117.860 ;
        RECT 16.990 105.840 19.290 106.010 ;
        RECT 19.690 117.860 21.990 118.030 ;
        RECT 19.690 106.010 19.860 117.860 ;
        RECT 20.350 117.150 21.350 117.600 ;
        RECT 20.360 106.915 20.530 116.955 ;
        RECT 21.150 106.915 21.320 116.955 ;
        RECT 20.590 106.530 21.090 106.700 ;
        RECT 21.820 106.010 21.990 117.860 ;
        RECT 34.315 117.860 36.615 118.030 ;
        RECT 31.615 108.860 33.915 109.030 ;
        RECT 31.615 107.925 31.785 108.860 ;
        RECT 32.515 108.170 33.015 108.340 ;
        RECT 32.285 107.925 32.455 107.955 ;
        RECT 31.560 106.945 32.455 107.925 ;
        RECT 19.690 105.840 21.990 106.010 ;
        RECT 31.615 106.010 31.785 106.945 ;
        RECT 32.285 106.915 32.455 106.945 ;
        RECT 33.075 106.915 33.245 107.955 ;
        RECT 32.100 106.530 33.015 106.700 ;
        RECT 32.100 106.325 32.935 106.530 ;
        RECT 33.745 106.010 33.915 108.860 ;
        RECT 31.615 105.840 33.915 106.010 ;
        RECT 34.315 106.010 34.485 117.860 ;
        RECT 34.975 117.150 35.975 117.600 ;
        RECT 34.985 106.915 35.155 116.955 ;
        RECT 35.775 106.915 35.945 116.955 ;
        RECT 35.215 106.530 35.715 106.700 ;
        RECT 36.445 106.010 36.615 117.860 ;
        RECT 42.415 117.860 44.715 118.030 ;
        RECT 37.015 108.860 39.315 109.030 ;
        RECT 37.015 107.925 37.185 108.860 ;
        RECT 37.915 108.170 38.415 108.340 ;
        RECT 37.685 107.925 37.855 107.955 ;
        RECT 36.960 106.945 37.855 107.925 ;
        RECT 34.315 105.840 36.615 106.010 ;
        RECT 37.015 106.010 37.185 106.945 ;
        RECT 37.685 106.915 37.855 106.945 ;
        RECT 38.475 106.915 38.645 107.955 ;
        RECT 37.500 106.530 38.415 106.700 ;
        RECT 37.500 106.325 38.335 106.530 ;
        RECT 39.145 106.010 39.315 108.860 ;
        RECT 39.715 108.860 42.015 109.030 ;
        RECT 39.715 107.925 39.885 108.860 ;
        RECT 40.615 108.170 41.115 108.340 ;
        RECT 40.385 107.925 40.555 107.955 ;
        RECT 39.660 106.945 40.555 107.925 ;
        RECT 37.015 105.840 39.315 106.010 ;
        RECT 39.715 106.010 39.885 106.945 ;
        RECT 40.385 106.915 40.555 106.945 ;
        RECT 41.175 106.915 41.345 107.955 ;
        RECT 40.200 106.530 41.115 106.700 ;
        RECT 40.200 106.325 41.035 106.530 ;
        RECT 41.845 106.010 42.015 108.860 ;
        RECT 39.715 105.840 42.015 106.010 ;
        RECT 42.415 106.010 42.585 117.860 ;
        RECT 43.075 117.150 44.075 117.600 ;
        RECT 43.085 106.915 43.255 116.955 ;
        RECT 43.875 106.915 44.045 116.955 ;
        RECT 43.315 106.530 43.815 106.700 ;
        RECT 44.545 106.010 44.715 117.860 ;
        RECT 42.415 105.840 44.715 106.010 ;
        RECT 45.115 117.860 47.415 118.030 ;
        RECT 45.115 106.010 45.285 117.860 ;
        RECT 45.775 117.150 46.775 117.600 ;
        RECT 45.785 106.915 45.955 116.955 ;
        RECT 46.575 106.915 46.745 116.955 ;
        RECT 46.015 106.530 46.515 106.700 ;
        RECT 47.245 106.010 47.415 117.860 ;
        RECT 59.740 117.860 62.040 118.030 ;
        RECT 57.040 108.860 59.340 109.030 ;
        RECT 57.040 107.925 57.210 108.860 ;
        RECT 57.940 108.170 58.440 108.340 ;
        RECT 57.710 107.925 57.880 107.955 ;
        RECT 56.985 106.945 57.880 107.925 ;
        RECT 45.115 105.840 47.415 106.010 ;
        RECT 57.040 106.010 57.210 106.945 ;
        RECT 57.710 106.915 57.880 106.945 ;
        RECT 58.500 106.915 58.670 107.955 ;
        RECT 57.525 106.530 58.440 106.700 ;
        RECT 57.525 106.325 58.360 106.530 ;
        RECT 59.170 106.010 59.340 108.860 ;
        RECT 57.040 105.840 59.340 106.010 ;
        RECT 59.740 106.010 59.910 117.860 ;
        RECT 60.400 117.150 61.400 117.600 ;
        RECT 60.410 106.915 60.580 116.955 ;
        RECT 61.200 106.915 61.370 116.955 ;
        RECT 60.640 106.530 61.140 106.700 ;
        RECT 61.870 106.010 62.040 117.860 ;
        RECT 67.840 117.860 70.140 118.030 ;
        RECT 62.440 108.860 64.740 109.030 ;
        RECT 62.440 107.925 62.610 108.860 ;
        RECT 63.340 108.170 63.840 108.340 ;
        RECT 63.110 107.925 63.280 107.955 ;
        RECT 62.385 106.945 63.280 107.925 ;
        RECT 59.740 105.840 62.040 106.010 ;
        RECT 62.440 106.010 62.610 106.945 ;
        RECT 63.110 106.915 63.280 106.945 ;
        RECT 63.900 106.915 64.070 107.955 ;
        RECT 62.925 106.530 63.840 106.700 ;
        RECT 62.925 106.325 63.760 106.530 ;
        RECT 64.570 106.010 64.740 108.860 ;
        RECT 65.140 108.860 67.440 109.030 ;
        RECT 65.140 107.925 65.310 108.860 ;
        RECT 66.040 108.170 66.540 108.340 ;
        RECT 65.810 107.925 65.980 107.955 ;
        RECT 65.085 106.945 65.980 107.925 ;
        RECT 62.440 105.840 64.740 106.010 ;
        RECT 65.140 106.010 65.310 106.945 ;
        RECT 65.810 106.915 65.980 106.945 ;
        RECT 66.600 106.915 66.770 107.955 ;
        RECT 65.625 106.530 66.540 106.700 ;
        RECT 65.625 106.325 66.460 106.530 ;
        RECT 67.270 106.010 67.440 108.860 ;
        RECT 65.140 105.840 67.440 106.010 ;
        RECT 67.840 106.010 68.010 117.860 ;
        RECT 68.500 117.150 69.500 117.600 ;
        RECT 68.510 106.915 68.680 116.955 ;
        RECT 69.300 106.915 69.470 116.955 ;
        RECT 68.740 106.530 69.240 106.700 ;
        RECT 69.970 106.010 70.140 117.860 ;
        RECT 67.840 105.840 70.140 106.010 ;
        RECT 70.540 117.860 72.840 118.030 ;
        RECT 70.540 106.010 70.710 117.860 ;
        RECT 71.200 117.150 72.200 117.600 ;
        RECT 71.210 106.915 71.380 116.955 ;
        RECT 72.000 106.915 72.170 116.955 ;
        RECT 71.440 106.530 71.940 106.700 ;
        RECT 72.670 106.010 72.840 117.860 ;
        RECT 85.165 117.860 87.465 118.030 ;
        RECT 82.465 108.860 84.765 109.030 ;
        RECT 82.465 107.925 82.635 108.860 ;
        RECT 83.365 108.170 83.865 108.340 ;
        RECT 83.135 107.925 83.305 107.955 ;
        RECT 82.410 106.945 83.305 107.925 ;
        RECT 70.540 105.840 72.840 106.010 ;
        RECT 82.465 106.010 82.635 106.945 ;
        RECT 83.135 106.915 83.305 106.945 ;
        RECT 83.925 106.915 84.095 107.955 ;
        RECT 82.950 106.530 83.865 106.700 ;
        RECT 82.950 106.325 83.785 106.530 ;
        RECT 84.595 106.010 84.765 108.860 ;
        RECT 82.465 105.840 84.765 106.010 ;
        RECT 85.165 106.010 85.335 117.860 ;
        RECT 85.825 117.150 86.825 117.600 ;
        RECT 85.835 106.915 86.005 116.955 ;
        RECT 86.625 106.915 86.795 116.955 ;
        RECT 86.065 106.530 86.565 106.700 ;
        RECT 87.295 106.010 87.465 117.860 ;
        RECT 93.265 117.860 95.565 118.030 ;
        RECT 87.865 108.860 90.165 109.030 ;
        RECT 87.865 107.925 88.035 108.860 ;
        RECT 88.765 108.170 89.265 108.340 ;
        RECT 88.535 107.925 88.705 107.955 ;
        RECT 87.810 106.945 88.705 107.925 ;
        RECT 85.165 105.840 87.465 106.010 ;
        RECT 87.865 106.010 88.035 106.945 ;
        RECT 88.535 106.915 88.705 106.945 ;
        RECT 89.325 106.915 89.495 107.955 ;
        RECT 88.350 106.530 89.265 106.700 ;
        RECT 88.350 106.325 89.185 106.530 ;
        RECT 89.995 106.010 90.165 108.860 ;
        RECT 90.565 108.860 92.865 109.030 ;
        RECT 90.565 107.925 90.735 108.860 ;
        RECT 91.465 108.170 91.965 108.340 ;
        RECT 91.235 107.925 91.405 107.955 ;
        RECT 90.510 106.945 91.405 107.925 ;
        RECT 87.865 105.840 90.165 106.010 ;
        RECT 90.565 106.010 90.735 106.945 ;
        RECT 91.235 106.915 91.405 106.945 ;
        RECT 92.025 106.915 92.195 107.955 ;
        RECT 91.050 106.530 91.965 106.700 ;
        RECT 91.050 106.325 91.885 106.530 ;
        RECT 92.695 106.010 92.865 108.860 ;
        RECT 90.565 105.840 92.865 106.010 ;
        RECT 93.265 106.010 93.435 117.860 ;
        RECT 93.925 117.150 94.925 117.600 ;
        RECT 93.935 106.915 94.105 116.955 ;
        RECT 94.725 106.915 94.895 116.955 ;
        RECT 94.165 106.530 94.665 106.700 ;
        RECT 95.395 106.010 95.565 117.860 ;
        RECT 93.265 105.840 95.565 106.010 ;
        RECT 95.965 117.860 98.265 118.030 ;
        RECT 95.965 106.010 96.135 117.860 ;
        RECT 96.625 117.150 97.625 117.600 ;
        RECT 96.635 106.915 96.805 116.955 ;
        RECT 97.425 106.915 97.595 116.955 ;
        RECT 96.865 106.530 97.365 106.700 ;
        RECT 98.095 106.010 98.265 117.860 ;
        RECT 110.590 117.860 112.890 118.030 ;
        RECT 107.890 108.860 110.190 109.030 ;
        RECT 107.890 107.925 108.060 108.860 ;
        RECT 108.790 108.170 109.290 108.340 ;
        RECT 108.560 107.925 108.730 107.955 ;
        RECT 107.835 106.945 108.730 107.925 ;
        RECT 95.965 105.840 98.265 106.010 ;
        RECT 107.890 106.010 108.060 106.945 ;
        RECT 108.560 106.915 108.730 106.945 ;
        RECT 109.350 106.915 109.520 107.955 ;
        RECT 108.375 106.530 109.290 106.700 ;
        RECT 108.375 106.325 109.210 106.530 ;
        RECT 110.020 106.010 110.190 108.860 ;
        RECT 107.890 105.840 110.190 106.010 ;
        RECT 110.590 106.010 110.760 117.860 ;
        RECT 111.250 117.150 112.250 117.600 ;
        RECT 111.260 106.915 111.430 116.955 ;
        RECT 112.050 106.915 112.220 116.955 ;
        RECT 111.490 106.530 111.990 106.700 ;
        RECT 112.720 106.010 112.890 117.860 ;
        RECT 118.690 117.860 120.990 118.030 ;
        RECT 113.290 108.860 115.590 109.030 ;
        RECT 113.290 107.925 113.460 108.860 ;
        RECT 114.190 108.170 114.690 108.340 ;
        RECT 113.960 107.925 114.130 107.955 ;
        RECT 113.235 106.945 114.130 107.925 ;
        RECT 110.590 105.840 112.890 106.010 ;
        RECT 113.290 106.010 113.460 106.945 ;
        RECT 113.960 106.915 114.130 106.945 ;
        RECT 114.750 106.915 114.920 107.955 ;
        RECT 113.775 106.530 114.690 106.700 ;
        RECT 113.775 106.325 114.610 106.530 ;
        RECT 115.420 106.010 115.590 108.860 ;
        RECT 115.990 108.860 118.290 109.030 ;
        RECT 115.990 107.925 116.160 108.860 ;
        RECT 116.890 108.170 117.390 108.340 ;
        RECT 116.660 107.925 116.830 107.955 ;
        RECT 115.935 106.945 116.830 107.925 ;
        RECT 113.290 105.840 115.590 106.010 ;
        RECT 115.990 106.010 116.160 106.945 ;
        RECT 116.660 106.915 116.830 106.945 ;
        RECT 117.450 106.915 117.620 107.955 ;
        RECT 116.475 106.530 117.390 106.700 ;
        RECT 116.475 106.325 117.310 106.530 ;
        RECT 118.120 106.010 118.290 108.860 ;
        RECT 115.990 105.840 118.290 106.010 ;
        RECT 118.690 106.010 118.860 117.860 ;
        RECT 119.350 117.150 120.350 117.600 ;
        RECT 119.360 106.915 119.530 116.955 ;
        RECT 120.150 106.915 120.320 116.955 ;
        RECT 119.590 106.530 120.090 106.700 ;
        RECT 120.820 106.010 120.990 117.860 ;
        RECT 118.690 105.840 120.990 106.010 ;
        RECT 121.390 117.860 123.690 118.030 ;
        RECT 121.390 106.010 121.560 117.860 ;
        RECT 122.050 117.150 123.050 117.600 ;
        RECT 122.060 106.915 122.230 116.955 ;
        RECT 122.850 106.915 123.020 116.955 ;
        RECT 122.290 106.530 122.790 106.700 ;
        RECT 123.520 106.010 123.690 117.860 ;
        RECT 136.015 117.860 138.315 118.030 ;
        RECT 133.315 108.860 135.615 109.030 ;
        RECT 133.315 107.925 133.485 108.860 ;
        RECT 134.215 108.170 134.715 108.340 ;
        RECT 133.985 107.925 134.155 107.955 ;
        RECT 133.260 106.945 134.155 107.925 ;
        RECT 121.390 105.840 123.690 106.010 ;
        RECT 133.315 106.010 133.485 106.945 ;
        RECT 133.985 106.915 134.155 106.945 ;
        RECT 134.775 106.915 134.945 107.955 ;
        RECT 133.800 106.530 134.715 106.700 ;
        RECT 133.800 106.325 134.635 106.530 ;
        RECT 135.445 106.010 135.615 108.860 ;
        RECT 133.315 105.840 135.615 106.010 ;
        RECT 136.015 106.010 136.185 117.860 ;
        RECT 136.675 117.150 137.675 117.600 ;
        RECT 136.685 106.915 136.855 116.955 ;
        RECT 137.475 106.915 137.645 116.955 ;
        RECT 136.915 106.530 137.415 106.700 ;
        RECT 138.145 106.010 138.315 117.860 ;
        RECT 144.115 117.860 146.415 118.030 ;
        RECT 138.715 108.860 141.015 109.030 ;
        RECT 138.715 107.925 138.885 108.860 ;
        RECT 139.615 108.170 140.115 108.340 ;
        RECT 139.385 107.925 139.555 107.955 ;
        RECT 138.660 106.945 139.555 107.925 ;
        RECT 136.015 105.840 138.315 106.010 ;
        RECT 138.715 106.010 138.885 106.945 ;
        RECT 139.385 106.915 139.555 106.945 ;
        RECT 140.175 106.915 140.345 107.955 ;
        RECT 139.200 106.530 140.115 106.700 ;
        RECT 139.200 106.325 140.035 106.530 ;
        RECT 140.845 106.010 141.015 108.860 ;
        RECT 141.415 108.860 143.715 109.030 ;
        RECT 141.415 107.925 141.585 108.860 ;
        RECT 142.315 108.170 142.815 108.340 ;
        RECT 142.085 107.925 142.255 107.955 ;
        RECT 141.360 106.945 142.255 107.925 ;
        RECT 138.715 105.840 141.015 106.010 ;
        RECT 141.415 106.010 141.585 106.945 ;
        RECT 142.085 106.915 142.255 106.945 ;
        RECT 142.875 106.915 143.045 107.955 ;
        RECT 141.900 106.530 142.815 106.700 ;
        RECT 141.900 106.325 142.735 106.530 ;
        RECT 143.545 106.010 143.715 108.860 ;
        RECT 141.415 105.840 143.715 106.010 ;
        RECT 144.115 106.010 144.285 117.860 ;
        RECT 144.775 117.150 145.775 117.600 ;
        RECT 144.785 106.915 144.955 116.955 ;
        RECT 145.575 106.915 145.745 116.955 ;
        RECT 145.015 106.530 145.515 106.700 ;
        RECT 146.245 106.010 146.415 117.860 ;
        RECT 144.115 105.840 146.415 106.010 ;
        RECT 146.815 117.860 149.115 118.030 ;
        RECT 146.815 106.010 146.985 117.860 ;
        RECT 147.475 117.150 148.475 117.600 ;
        RECT 147.485 106.915 147.655 116.955 ;
        RECT 148.275 106.915 148.445 116.955 ;
        RECT 147.715 106.530 148.215 106.700 ;
        RECT 148.945 106.010 149.115 117.860 ;
        RECT 146.815 105.840 149.115 106.010 ;
        RECT 6.190 104.770 8.490 104.940 ;
        RECT 6.190 103.830 6.360 104.770 ;
        RECT 6.570 104.080 7.610 104.525 ;
        RECT 6.860 103.830 7.030 103.910 ;
        RECT 6.185 103.300 7.030 103.830 ;
        RECT 6.190 102.360 6.360 103.300 ;
        RECT 6.860 103.220 7.030 103.300 ;
        RECT 7.650 103.220 7.820 103.910 ;
        RECT 7.090 102.880 7.590 103.050 ;
        RECT 8.320 102.360 8.490 104.770 ;
        RECT 6.190 102.190 8.490 102.360 ;
        RECT 8.890 104.770 11.190 104.940 ;
        RECT 8.890 96.510 9.060 104.770 ;
        RECT 9.790 104.080 10.290 104.250 ;
        RECT 9.560 97.370 9.730 103.910 ;
        RECT 10.350 97.370 10.520 103.910 ;
        RECT 9.550 96.800 10.550 97.200 ;
        RECT 11.020 96.510 11.190 104.770 ;
        RECT 11.590 104.770 13.890 104.940 ;
        RECT 11.590 103.830 11.760 104.770 ;
        RECT 11.970 104.080 13.010 104.525 ;
        RECT 12.260 103.830 12.430 103.910 ;
        RECT 11.585 103.300 12.430 103.830 ;
        RECT 11.590 102.360 11.760 103.300 ;
        RECT 12.260 103.220 12.430 103.300 ;
        RECT 13.050 103.220 13.220 103.910 ;
        RECT 12.490 102.880 12.990 103.050 ;
        RECT 13.720 102.360 13.890 104.770 ;
        RECT 14.290 104.770 16.590 104.940 ;
        RECT 14.290 103.830 14.460 104.770 ;
        RECT 14.670 104.080 15.710 104.525 ;
        RECT 14.960 103.830 15.130 103.910 ;
        RECT 14.285 103.300 15.130 103.830 ;
        RECT 11.590 102.190 13.890 102.360 ;
        RECT 14.290 102.360 14.460 103.300 ;
        RECT 14.960 103.220 15.130 103.300 ;
        RECT 15.750 103.220 15.920 103.910 ;
        RECT 15.190 102.880 15.690 103.050 ;
        RECT 16.420 102.360 16.590 104.770 ;
        RECT 14.290 102.190 16.590 102.360 ;
        RECT 16.990 104.770 19.290 104.940 ;
        RECT 8.890 96.340 11.190 96.510 ;
        RECT 16.990 96.510 17.160 104.770 ;
        RECT 17.890 104.080 18.390 104.250 ;
        RECT 17.660 97.370 17.830 103.910 ;
        RECT 18.450 97.370 18.620 103.910 ;
        RECT 17.650 96.800 18.650 97.200 ;
        RECT 19.120 96.510 19.290 104.770 ;
        RECT 16.990 96.340 19.290 96.510 ;
        RECT 19.690 104.770 21.990 104.940 ;
        RECT 19.690 96.510 19.860 104.770 ;
        RECT 20.590 104.080 21.090 104.250 ;
        RECT 20.360 97.370 20.530 103.910 ;
        RECT 21.150 97.370 21.320 103.910 ;
        RECT 20.350 96.800 21.350 97.200 ;
        RECT 21.820 96.510 21.990 104.770 ;
        RECT 31.615 104.770 33.915 104.940 ;
        RECT 31.615 103.830 31.785 104.770 ;
        RECT 31.995 104.080 33.035 104.525 ;
        RECT 32.285 103.830 32.455 103.910 ;
        RECT 31.610 103.300 32.455 103.830 ;
        RECT 31.615 102.360 31.785 103.300 ;
        RECT 32.285 103.220 32.455 103.300 ;
        RECT 33.075 103.220 33.245 103.910 ;
        RECT 32.515 102.880 33.015 103.050 ;
        RECT 33.745 102.360 33.915 104.770 ;
        RECT 31.615 102.190 33.915 102.360 ;
        RECT 34.315 104.770 36.615 104.940 ;
        RECT 19.690 96.340 21.990 96.510 ;
        RECT 34.315 96.510 34.485 104.770 ;
        RECT 35.215 104.080 35.715 104.250 ;
        RECT 34.985 97.370 35.155 103.910 ;
        RECT 35.775 97.370 35.945 103.910 ;
        RECT 34.975 96.800 35.975 97.200 ;
        RECT 36.445 96.510 36.615 104.770 ;
        RECT 37.015 104.770 39.315 104.940 ;
        RECT 37.015 103.830 37.185 104.770 ;
        RECT 37.395 104.080 38.435 104.525 ;
        RECT 37.685 103.830 37.855 103.910 ;
        RECT 37.010 103.300 37.855 103.830 ;
        RECT 37.015 102.360 37.185 103.300 ;
        RECT 37.685 103.220 37.855 103.300 ;
        RECT 38.475 103.220 38.645 103.910 ;
        RECT 37.915 102.880 38.415 103.050 ;
        RECT 39.145 102.360 39.315 104.770 ;
        RECT 39.715 104.770 42.015 104.940 ;
        RECT 39.715 103.830 39.885 104.770 ;
        RECT 40.095 104.080 41.135 104.525 ;
        RECT 40.385 103.830 40.555 103.910 ;
        RECT 39.710 103.300 40.555 103.830 ;
        RECT 37.015 102.190 39.315 102.360 ;
        RECT 39.715 102.360 39.885 103.300 ;
        RECT 40.385 103.220 40.555 103.300 ;
        RECT 41.175 103.220 41.345 103.910 ;
        RECT 40.615 102.880 41.115 103.050 ;
        RECT 41.845 102.360 42.015 104.770 ;
        RECT 39.715 102.190 42.015 102.360 ;
        RECT 42.415 104.770 44.715 104.940 ;
        RECT 34.315 96.340 36.615 96.510 ;
        RECT 42.415 96.510 42.585 104.770 ;
        RECT 43.315 104.080 43.815 104.250 ;
        RECT 43.085 97.370 43.255 103.910 ;
        RECT 43.875 97.370 44.045 103.910 ;
        RECT 43.075 96.800 44.075 97.200 ;
        RECT 44.545 96.510 44.715 104.770 ;
        RECT 42.415 96.340 44.715 96.510 ;
        RECT 45.115 104.770 47.415 104.940 ;
        RECT 45.115 96.510 45.285 104.770 ;
        RECT 46.015 104.080 46.515 104.250 ;
        RECT 45.785 97.370 45.955 103.910 ;
        RECT 46.575 97.370 46.745 103.910 ;
        RECT 45.775 96.800 46.775 97.200 ;
        RECT 47.245 96.510 47.415 104.770 ;
        RECT 57.040 104.770 59.340 104.940 ;
        RECT 57.040 103.830 57.210 104.770 ;
        RECT 57.420 104.080 58.460 104.525 ;
        RECT 57.710 103.830 57.880 103.910 ;
        RECT 57.035 103.300 57.880 103.830 ;
        RECT 57.040 102.360 57.210 103.300 ;
        RECT 57.710 103.220 57.880 103.300 ;
        RECT 58.500 103.220 58.670 103.910 ;
        RECT 57.940 102.880 58.440 103.050 ;
        RECT 59.170 102.360 59.340 104.770 ;
        RECT 57.040 102.190 59.340 102.360 ;
        RECT 59.740 104.770 62.040 104.940 ;
        RECT 45.115 96.340 47.415 96.510 ;
        RECT 59.740 96.510 59.910 104.770 ;
        RECT 60.640 104.080 61.140 104.250 ;
        RECT 60.410 97.370 60.580 103.910 ;
        RECT 61.200 97.370 61.370 103.910 ;
        RECT 60.400 96.800 61.400 97.200 ;
        RECT 61.870 96.510 62.040 104.770 ;
        RECT 62.440 104.770 64.740 104.940 ;
        RECT 62.440 103.830 62.610 104.770 ;
        RECT 62.820 104.080 63.860 104.525 ;
        RECT 63.110 103.830 63.280 103.910 ;
        RECT 62.435 103.300 63.280 103.830 ;
        RECT 62.440 102.360 62.610 103.300 ;
        RECT 63.110 103.220 63.280 103.300 ;
        RECT 63.900 103.220 64.070 103.910 ;
        RECT 63.340 102.880 63.840 103.050 ;
        RECT 64.570 102.360 64.740 104.770 ;
        RECT 65.140 104.770 67.440 104.940 ;
        RECT 65.140 103.830 65.310 104.770 ;
        RECT 65.520 104.080 66.560 104.525 ;
        RECT 65.810 103.830 65.980 103.910 ;
        RECT 65.135 103.300 65.980 103.830 ;
        RECT 62.440 102.190 64.740 102.360 ;
        RECT 65.140 102.360 65.310 103.300 ;
        RECT 65.810 103.220 65.980 103.300 ;
        RECT 66.600 103.220 66.770 103.910 ;
        RECT 66.040 102.880 66.540 103.050 ;
        RECT 67.270 102.360 67.440 104.770 ;
        RECT 65.140 102.190 67.440 102.360 ;
        RECT 67.840 104.770 70.140 104.940 ;
        RECT 59.740 96.340 62.040 96.510 ;
        RECT 67.840 96.510 68.010 104.770 ;
        RECT 68.740 104.080 69.240 104.250 ;
        RECT 68.510 97.370 68.680 103.910 ;
        RECT 69.300 97.370 69.470 103.910 ;
        RECT 68.500 96.800 69.500 97.200 ;
        RECT 69.970 96.510 70.140 104.770 ;
        RECT 67.840 96.340 70.140 96.510 ;
        RECT 70.540 104.770 72.840 104.940 ;
        RECT 70.540 96.510 70.710 104.770 ;
        RECT 71.440 104.080 71.940 104.250 ;
        RECT 71.210 97.370 71.380 103.910 ;
        RECT 72.000 97.370 72.170 103.910 ;
        RECT 71.200 96.800 72.200 97.200 ;
        RECT 72.670 96.510 72.840 104.770 ;
        RECT 82.465 104.770 84.765 104.940 ;
        RECT 82.465 103.830 82.635 104.770 ;
        RECT 82.845 104.080 83.885 104.525 ;
        RECT 83.135 103.830 83.305 103.910 ;
        RECT 82.460 103.300 83.305 103.830 ;
        RECT 82.465 102.360 82.635 103.300 ;
        RECT 83.135 103.220 83.305 103.300 ;
        RECT 83.925 103.220 84.095 103.910 ;
        RECT 83.365 102.880 83.865 103.050 ;
        RECT 84.595 102.360 84.765 104.770 ;
        RECT 82.465 102.190 84.765 102.360 ;
        RECT 85.165 104.770 87.465 104.940 ;
        RECT 70.540 96.340 72.840 96.510 ;
        RECT 85.165 96.510 85.335 104.770 ;
        RECT 86.065 104.080 86.565 104.250 ;
        RECT 85.835 97.370 86.005 103.910 ;
        RECT 86.625 97.370 86.795 103.910 ;
        RECT 85.825 96.800 86.825 97.200 ;
        RECT 87.295 96.510 87.465 104.770 ;
        RECT 87.865 104.770 90.165 104.940 ;
        RECT 87.865 103.830 88.035 104.770 ;
        RECT 88.245 104.080 89.285 104.525 ;
        RECT 88.535 103.830 88.705 103.910 ;
        RECT 87.860 103.300 88.705 103.830 ;
        RECT 87.865 102.360 88.035 103.300 ;
        RECT 88.535 103.220 88.705 103.300 ;
        RECT 89.325 103.220 89.495 103.910 ;
        RECT 88.765 102.880 89.265 103.050 ;
        RECT 89.995 102.360 90.165 104.770 ;
        RECT 90.565 104.770 92.865 104.940 ;
        RECT 90.565 103.830 90.735 104.770 ;
        RECT 90.945 104.080 91.985 104.525 ;
        RECT 91.235 103.830 91.405 103.910 ;
        RECT 90.560 103.300 91.405 103.830 ;
        RECT 87.865 102.190 90.165 102.360 ;
        RECT 90.565 102.360 90.735 103.300 ;
        RECT 91.235 103.220 91.405 103.300 ;
        RECT 92.025 103.220 92.195 103.910 ;
        RECT 91.465 102.880 91.965 103.050 ;
        RECT 92.695 102.360 92.865 104.770 ;
        RECT 90.565 102.190 92.865 102.360 ;
        RECT 93.265 104.770 95.565 104.940 ;
        RECT 85.165 96.340 87.465 96.510 ;
        RECT 93.265 96.510 93.435 104.770 ;
        RECT 94.165 104.080 94.665 104.250 ;
        RECT 93.935 97.370 94.105 103.910 ;
        RECT 94.725 97.370 94.895 103.910 ;
        RECT 93.925 96.800 94.925 97.200 ;
        RECT 95.395 96.510 95.565 104.770 ;
        RECT 93.265 96.340 95.565 96.510 ;
        RECT 95.965 104.770 98.265 104.940 ;
        RECT 95.965 96.510 96.135 104.770 ;
        RECT 96.865 104.080 97.365 104.250 ;
        RECT 96.635 97.370 96.805 103.910 ;
        RECT 97.425 97.370 97.595 103.910 ;
        RECT 96.625 96.800 97.625 97.200 ;
        RECT 98.095 96.510 98.265 104.770 ;
        RECT 107.890 104.770 110.190 104.940 ;
        RECT 107.890 103.830 108.060 104.770 ;
        RECT 108.270 104.080 109.310 104.525 ;
        RECT 108.560 103.830 108.730 103.910 ;
        RECT 107.885 103.300 108.730 103.830 ;
        RECT 107.890 102.360 108.060 103.300 ;
        RECT 108.560 103.220 108.730 103.300 ;
        RECT 109.350 103.220 109.520 103.910 ;
        RECT 108.790 102.880 109.290 103.050 ;
        RECT 110.020 102.360 110.190 104.770 ;
        RECT 107.890 102.190 110.190 102.360 ;
        RECT 110.590 104.770 112.890 104.940 ;
        RECT 95.965 96.340 98.265 96.510 ;
        RECT 110.590 96.510 110.760 104.770 ;
        RECT 111.490 104.080 111.990 104.250 ;
        RECT 111.260 97.370 111.430 103.910 ;
        RECT 112.050 97.370 112.220 103.910 ;
        RECT 111.250 96.800 112.250 97.200 ;
        RECT 112.720 96.510 112.890 104.770 ;
        RECT 113.290 104.770 115.590 104.940 ;
        RECT 113.290 103.830 113.460 104.770 ;
        RECT 113.670 104.080 114.710 104.525 ;
        RECT 113.960 103.830 114.130 103.910 ;
        RECT 113.285 103.300 114.130 103.830 ;
        RECT 113.290 102.360 113.460 103.300 ;
        RECT 113.960 103.220 114.130 103.300 ;
        RECT 114.750 103.220 114.920 103.910 ;
        RECT 114.190 102.880 114.690 103.050 ;
        RECT 115.420 102.360 115.590 104.770 ;
        RECT 115.990 104.770 118.290 104.940 ;
        RECT 115.990 103.830 116.160 104.770 ;
        RECT 116.370 104.080 117.410 104.525 ;
        RECT 116.660 103.830 116.830 103.910 ;
        RECT 115.985 103.300 116.830 103.830 ;
        RECT 113.290 102.190 115.590 102.360 ;
        RECT 115.990 102.360 116.160 103.300 ;
        RECT 116.660 103.220 116.830 103.300 ;
        RECT 117.450 103.220 117.620 103.910 ;
        RECT 116.890 102.880 117.390 103.050 ;
        RECT 118.120 102.360 118.290 104.770 ;
        RECT 115.990 102.190 118.290 102.360 ;
        RECT 118.690 104.770 120.990 104.940 ;
        RECT 110.590 96.340 112.890 96.510 ;
        RECT 118.690 96.510 118.860 104.770 ;
        RECT 119.590 104.080 120.090 104.250 ;
        RECT 119.360 97.370 119.530 103.910 ;
        RECT 120.150 97.370 120.320 103.910 ;
        RECT 119.350 96.800 120.350 97.200 ;
        RECT 120.820 96.510 120.990 104.770 ;
        RECT 118.690 96.340 120.990 96.510 ;
        RECT 121.390 104.770 123.690 104.940 ;
        RECT 121.390 96.510 121.560 104.770 ;
        RECT 122.290 104.080 122.790 104.250 ;
        RECT 122.060 97.370 122.230 103.910 ;
        RECT 122.850 97.370 123.020 103.910 ;
        RECT 122.050 96.800 123.050 97.200 ;
        RECT 123.520 96.510 123.690 104.770 ;
        RECT 133.315 104.770 135.615 104.940 ;
        RECT 133.315 103.830 133.485 104.770 ;
        RECT 133.695 104.080 134.735 104.525 ;
        RECT 133.985 103.830 134.155 103.910 ;
        RECT 133.310 103.300 134.155 103.830 ;
        RECT 133.315 102.360 133.485 103.300 ;
        RECT 133.985 103.220 134.155 103.300 ;
        RECT 134.775 103.220 134.945 103.910 ;
        RECT 134.215 102.880 134.715 103.050 ;
        RECT 135.445 102.360 135.615 104.770 ;
        RECT 133.315 102.190 135.615 102.360 ;
        RECT 136.015 104.770 138.315 104.940 ;
        RECT 121.390 96.340 123.690 96.510 ;
        RECT 136.015 96.510 136.185 104.770 ;
        RECT 136.915 104.080 137.415 104.250 ;
        RECT 136.685 97.370 136.855 103.910 ;
        RECT 137.475 97.370 137.645 103.910 ;
        RECT 136.675 96.800 137.675 97.200 ;
        RECT 138.145 96.510 138.315 104.770 ;
        RECT 138.715 104.770 141.015 104.940 ;
        RECT 138.715 103.830 138.885 104.770 ;
        RECT 139.095 104.080 140.135 104.525 ;
        RECT 139.385 103.830 139.555 103.910 ;
        RECT 138.710 103.300 139.555 103.830 ;
        RECT 138.715 102.360 138.885 103.300 ;
        RECT 139.385 103.220 139.555 103.300 ;
        RECT 140.175 103.220 140.345 103.910 ;
        RECT 139.615 102.880 140.115 103.050 ;
        RECT 140.845 102.360 141.015 104.770 ;
        RECT 141.415 104.770 143.715 104.940 ;
        RECT 141.415 103.830 141.585 104.770 ;
        RECT 141.795 104.080 142.835 104.525 ;
        RECT 142.085 103.830 142.255 103.910 ;
        RECT 141.410 103.300 142.255 103.830 ;
        RECT 138.715 102.190 141.015 102.360 ;
        RECT 141.415 102.360 141.585 103.300 ;
        RECT 142.085 103.220 142.255 103.300 ;
        RECT 142.875 103.220 143.045 103.910 ;
        RECT 142.315 102.880 142.815 103.050 ;
        RECT 143.545 102.360 143.715 104.770 ;
        RECT 141.415 102.190 143.715 102.360 ;
        RECT 144.115 104.770 146.415 104.940 ;
        RECT 136.015 96.340 138.315 96.510 ;
        RECT 144.115 96.510 144.285 104.770 ;
        RECT 145.015 104.080 145.515 104.250 ;
        RECT 144.785 97.370 144.955 103.910 ;
        RECT 145.575 97.370 145.745 103.910 ;
        RECT 144.775 96.800 145.775 97.200 ;
        RECT 146.245 96.510 146.415 104.770 ;
        RECT 144.115 96.340 146.415 96.510 ;
        RECT 146.815 104.770 149.115 104.940 ;
        RECT 146.815 96.510 146.985 104.770 ;
        RECT 147.715 104.080 148.215 104.250 ;
        RECT 147.485 97.370 147.655 103.910 ;
        RECT 148.275 97.370 148.445 103.910 ;
        RECT 147.475 96.800 148.475 97.200 ;
        RECT 148.945 96.510 149.115 104.770 ;
        RECT 146.815 96.340 149.115 96.510 ;
        RECT 23.235 96.000 24.075 96.050 ;
        RECT 48.660 96.000 49.500 96.050 ;
        RECT 74.085 96.000 74.925 96.050 ;
        RECT 99.510 96.000 100.350 96.050 ;
        RECT 124.935 96.000 125.775 96.050 ;
        RECT 150.360 96.000 151.200 96.050 ;
        RECT 22.830 95.830 24.480 96.000 ;
        RECT 8.890 95.285 11.190 95.455 ;
        RECT 6.190 86.285 8.490 86.455 ;
        RECT 6.190 85.350 6.360 86.285 ;
        RECT 7.090 85.595 7.590 85.765 ;
        RECT 6.860 85.350 7.030 85.380 ;
        RECT 6.135 84.370 7.030 85.350 ;
        RECT 6.190 83.435 6.360 84.370 ;
        RECT 6.860 84.340 7.030 84.370 ;
        RECT 7.650 84.340 7.820 85.380 ;
        RECT 6.675 83.955 7.590 84.125 ;
        RECT 6.675 83.750 7.510 83.955 ;
        RECT 8.320 83.435 8.490 86.285 ;
        RECT 6.190 83.265 8.490 83.435 ;
        RECT 8.890 83.435 9.060 95.285 ;
        RECT 9.550 94.575 10.550 95.025 ;
        RECT 9.560 84.340 9.730 94.380 ;
        RECT 10.350 84.340 10.520 94.380 ;
        RECT 9.790 83.955 10.290 84.125 ;
        RECT 11.020 83.435 11.190 95.285 ;
        RECT 16.990 95.285 19.290 95.455 ;
        RECT 11.590 86.285 13.890 86.455 ;
        RECT 11.590 85.350 11.760 86.285 ;
        RECT 12.490 85.595 12.990 85.765 ;
        RECT 12.260 85.350 12.430 85.380 ;
        RECT 11.535 84.370 12.430 85.350 ;
        RECT 8.890 83.265 11.190 83.435 ;
        RECT 11.590 83.435 11.760 84.370 ;
        RECT 12.260 84.340 12.430 84.370 ;
        RECT 13.050 84.340 13.220 85.380 ;
        RECT 12.075 83.955 12.990 84.125 ;
        RECT 12.075 83.750 12.910 83.955 ;
        RECT 13.720 83.435 13.890 86.285 ;
        RECT 14.290 86.285 16.590 86.455 ;
        RECT 14.290 85.350 14.460 86.285 ;
        RECT 15.190 85.595 15.690 85.765 ;
        RECT 14.960 85.350 15.130 85.380 ;
        RECT 14.235 84.370 15.130 85.350 ;
        RECT 11.590 83.265 13.890 83.435 ;
        RECT 14.290 83.435 14.460 84.370 ;
        RECT 14.960 84.340 15.130 84.370 ;
        RECT 15.750 84.340 15.920 85.380 ;
        RECT 14.775 83.955 15.690 84.125 ;
        RECT 14.775 83.750 15.610 83.955 ;
        RECT 16.420 83.435 16.590 86.285 ;
        RECT 14.290 83.265 16.590 83.435 ;
        RECT 16.990 83.435 17.160 95.285 ;
        RECT 17.650 94.575 18.650 95.025 ;
        RECT 17.660 84.340 17.830 94.380 ;
        RECT 18.450 84.340 18.620 94.380 ;
        RECT 17.890 83.955 18.390 84.125 ;
        RECT 19.120 83.435 19.290 95.285 ;
        RECT 16.990 83.265 19.290 83.435 ;
        RECT 19.690 95.285 21.990 95.455 ;
        RECT 19.690 83.435 19.860 95.285 ;
        RECT 20.350 94.575 21.350 95.025 ;
        RECT 20.360 84.340 20.530 94.380 ;
        RECT 21.150 84.340 21.320 94.380 ;
        RECT 20.590 83.955 21.090 84.125 ;
        RECT 21.820 83.435 21.990 95.285 ;
        RECT 19.690 83.265 21.990 83.435 ;
        RECT 6.190 82.195 8.490 82.365 ;
        RECT 6.190 81.255 6.360 82.195 ;
        RECT 6.570 81.505 7.610 81.950 ;
        RECT 6.860 81.255 7.030 81.335 ;
        RECT 6.185 80.725 7.030 81.255 ;
        RECT 6.190 79.785 6.360 80.725 ;
        RECT 6.860 80.645 7.030 80.725 ;
        RECT 7.650 80.645 7.820 81.335 ;
        RECT 7.090 80.305 7.590 80.475 ;
        RECT 8.320 79.785 8.490 82.195 ;
        RECT 6.190 79.615 8.490 79.785 ;
        RECT 8.890 82.195 11.190 82.365 ;
        RECT 8.890 73.935 9.060 82.195 ;
        RECT 9.790 81.505 10.290 81.675 ;
        RECT 9.560 74.795 9.730 81.335 ;
        RECT 10.350 74.795 10.520 81.335 ;
        RECT 9.550 74.225 10.550 74.625 ;
        RECT 11.020 73.935 11.190 82.195 ;
        RECT 11.590 82.195 13.890 82.365 ;
        RECT 11.590 81.255 11.760 82.195 ;
        RECT 11.970 81.505 13.010 81.950 ;
        RECT 12.260 81.255 12.430 81.335 ;
        RECT 11.585 80.725 12.430 81.255 ;
        RECT 11.590 79.785 11.760 80.725 ;
        RECT 12.260 80.645 12.430 80.725 ;
        RECT 13.050 80.645 13.220 81.335 ;
        RECT 12.490 80.305 12.990 80.475 ;
        RECT 13.720 79.785 13.890 82.195 ;
        RECT 14.290 82.195 16.590 82.365 ;
        RECT 14.290 81.255 14.460 82.195 ;
        RECT 14.670 81.505 15.710 81.950 ;
        RECT 14.960 81.255 15.130 81.335 ;
        RECT 14.285 80.725 15.130 81.255 ;
        RECT 11.590 79.615 13.890 79.785 ;
        RECT 14.290 79.785 14.460 80.725 ;
        RECT 14.960 80.645 15.130 80.725 ;
        RECT 15.750 80.645 15.920 81.335 ;
        RECT 15.190 80.305 15.690 80.475 ;
        RECT 16.420 79.785 16.590 82.195 ;
        RECT 14.290 79.615 16.590 79.785 ;
        RECT 16.990 82.195 19.290 82.365 ;
        RECT 8.890 73.765 11.190 73.935 ;
        RECT 16.990 73.935 17.160 82.195 ;
        RECT 17.890 81.505 18.390 81.675 ;
        RECT 17.660 74.795 17.830 81.335 ;
        RECT 18.450 74.795 18.620 81.335 ;
        RECT 17.650 74.225 18.650 74.625 ;
        RECT 19.120 73.935 19.290 82.195 ;
        RECT 16.990 73.765 19.290 73.935 ;
        RECT 19.690 82.195 21.990 82.365 ;
        RECT 19.690 73.935 19.860 82.195 ;
        RECT 20.590 81.505 21.090 81.675 ;
        RECT 20.360 74.795 20.530 81.335 ;
        RECT 21.150 74.795 21.320 81.335 ;
        RECT 20.350 74.225 21.350 74.625 ;
        RECT 21.820 73.935 21.990 82.195 ;
        RECT 22.830 81.800 23.000 95.830 ;
        RECT 23.235 95.780 24.075 95.830 ;
        RECT 23.430 93.115 23.880 95.425 ;
        RECT 23.430 82.205 23.880 84.515 ;
        RECT 23.260 81.800 24.050 81.850 ;
        RECT 24.310 81.800 24.480 95.830 ;
        RECT 48.255 95.830 49.905 96.000 ;
        RECT 34.315 95.285 36.615 95.455 ;
        RECT 31.615 86.285 33.915 86.455 ;
        RECT 31.615 85.350 31.785 86.285 ;
        RECT 32.515 85.595 33.015 85.765 ;
        RECT 32.285 85.350 32.455 85.380 ;
        RECT 31.560 84.370 32.455 85.350 ;
        RECT 31.615 83.435 31.785 84.370 ;
        RECT 32.285 84.340 32.455 84.370 ;
        RECT 33.075 84.340 33.245 85.380 ;
        RECT 32.100 83.955 33.015 84.125 ;
        RECT 32.100 83.750 32.935 83.955 ;
        RECT 33.745 83.435 33.915 86.285 ;
        RECT 31.615 83.265 33.915 83.435 ;
        RECT 34.315 83.435 34.485 95.285 ;
        RECT 34.975 94.575 35.975 95.025 ;
        RECT 34.985 84.340 35.155 94.380 ;
        RECT 35.775 84.340 35.945 94.380 ;
        RECT 35.215 83.955 35.715 84.125 ;
        RECT 36.445 83.435 36.615 95.285 ;
        RECT 42.415 95.285 44.715 95.455 ;
        RECT 37.015 86.285 39.315 86.455 ;
        RECT 37.015 85.350 37.185 86.285 ;
        RECT 37.915 85.595 38.415 85.765 ;
        RECT 37.685 85.350 37.855 85.380 ;
        RECT 36.960 84.370 37.855 85.350 ;
        RECT 34.315 83.265 36.615 83.435 ;
        RECT 37.015 83.435 37.185 84.370 ;
        RECT 37.685 84.340 37.855 84.370 ;
        RECT 38.475 84.340 38.645 85.380 ;
        RECT 37.500 83.955 38.415 84.125 ;
        RECT 37.500 83.750 38.335 83.955 ;
        RECT 39.145 83.435 39.315 86.285 ;
        RECT 39.715 86.285 42.015 86.455 ;
        RECT 39.715 85.350 39.885 86.285 ;
        RECT 40.615 85.595 41.115 85.765 ;
        RECT 40.385 85.350 40.555 85.380 ;
        RECT 39.660 84.370 40.555 85.350 ;
        RECT 37.015 83.265 39.315 83.435 ;
        RECT 39.715 83.435 39.885 84.370 ;
        RECT 40.385 84.340 40.555 84.370 ;
        RECT 41.175 84.340 41.345 85.380 ;
        RECT 40.200 83.955 41.115 84.125 ;
        RECT 40.200 83.750 41.035 83.955 ;
        RECT 41.845 83.435 42.015 86.285 ;
        RECT 39.715 83.265 42.015 83.435 ;
        RECT 42.415 83.435 42.585 95.285 ;
        RECT 43.075 94.575 44.075 95.025 ;
        RECT 43.085 84.340 43.255 94.380 ;
        RECT 43.875 84.340 44.045 94.380 ;
        RECT 43.315 83.955 43.815 84.125 ;
        RECT 44.545 83.435 44.715 95.285 ;
        RECT 42.415 83.265 44.715 83.435 ;
        RECT 45.115 95.285 47.415 95.455 ;
        RECT 45.115 83.435 45.285 95.285 ;
        RECT 45.775 94.575 46.775 95.025 ;
        RECT 45.785 84.340 45.955 94.380 ;
        RECT 46.575 84.340 46.745 94.380 ;
        RECT 46.015 83.955 46.515 84.125 ;
        RECT 47.245 83.435 47.415 95.285 ;
        RECT 45.115 83.265 47.415 83.435 ;
        RECT 22.830 81.630 24.480 81.800 ;
        RECT 31.615 82.195 33.915 82.365 ;
        RECT 23.260 81.580 24.050 81.630 ;
        RECT 31.615 81.255 31.785 82.195 ;
        RECT 31.995 81.505 33.035 81.950 ;
        RECT 32.285 81.255 32.455 81.335 ;
        RECT 31.610 80.725 32.455 81.255 ;
        RECT 31.615 79.785 31.785 80.725 ;
        RECT 32.285 80.645 32.455 80.725 ;
        RECT 33.075 80.645 33.245 81.335 ;
        RECT 32.515 80.305 33.015 80.475 ;
        RECT 33.745 79.785 33.915 82.195 ;
        RECT 31.615 79.615 33.915 79.785 ;
        RECT 34.315 82.195 36.615 82.365 ;
        RECT 19.690 73.765 21.990 73.935 ;
        RECT 34.315 73.935 34.485 82.195 ;
        RECT 35.215 81.505 35.715 81.675 ;
        RECT 34.985 74.795 35.155 81.335 ;
        RECT 35.775 74.795 35.945 81.335 ;
        RECT 34.975 74.225 35.975 74.625 ;
        RECT 36.445 73.935 36.615 82.195 ;
        RECT 37.015 82.195 39.315 82.365 ;
        RECT 37.015 81.255 37.185 82.195 ;
        RECT 37.395 81.505 38.435 81.950 ;
        RECT 37.685 81.255 37.855 81.335 ;
        RECT 37.010 80.725 37.855 81.255 ;
        RECT 37.015 79.785 37.185 80.725 ;
        RECT 37.685 80.645 37.855 80.725 ;
        RECT 38.475 80.645 38.645 81.335 ;
        RECT 37.915 80.305 38.415 80.475 ;
        RECT 39.145 79.785 39.315 82.195 ;
        RECT 39.715 82.195 42.015 82.365 ;
        RECT 39.715 81.255 39.885 82.195 ;
        RECT 40.095 81.505 41.135 81.950 ;
        RECT 40.385 81.255 40.555 81.335 ;
        RECT 39.710 80.725 40.555 81.255 ;
        RECT 37.015 79.615 39.315 79.785 ;
        RECT 39.715 79.785 39.885 80.725 ;
        RECT 40.385 80.645 40.555 80.725 ;
        RECT 41.175 80.645 41.345 81.335 ;
        RECT 40.615 80.305 41.115 80.475 ;
        RECT 41.845 79.785 42.015 82.195 ;
        RECT 39.715 79.615 42.015 79.785 ;
        RECT 42.415 82.195 44.715 82.365 ;
        RECT 34.315 73.765 36.615 73.935 ;
        RECT 42.415 73.935 42.585 82.195 ;
        RECT 43.315 81.505 43.815 81.675 ;
        RECT 43.085 74.795 43.255 81.335 ;
        RECT 43.875 74.795 44.045 81.335 ;
        RECT 43.075 74.225 44.075 74.625 ;
        RECT 44.545 73.935 44.715 82.195 ;
        RECT 42.415 73.765 44.715 73.935 ;
        RECT 45.115 82.195 47.415 82.365 ;
        RECT 45.115 73.935 45.285 82.195 ;
        RECT 46.015 81.505 46.515 81.675 ;
        RECT 45.785 74.795 45.955 81.335 ;
        RECT 46.575 74.795 46.745 81.335 ;
        RECT 45.775 74.225 46.775 74.625 ;
        RECT 47.245 73.935 47.415 82.195 ;
        RECT 48.255 81.800 48.425 95.830 ;
        RECT 48.660 95.780 49.500 95.830 ;
        RECT 48.855 93.115 49.305 95.425 ;
        RECT 48.855 82.205 49.305 84.515 ;
        RECT 48.685 81.800 49.475 81.850 ;
        RECT 49.735 81.800 49.905 95.830 ;
        RECT 73.680 95.830 75.330 96.000 ;
        RECT 59.740 95.285 62.040 95.455 ;
        RECT 57.040 86.285 59.340 86.455 ;
        RECT 57.040 85.350 57.210 86.285 ;
        RECT 57.940 85.595 58.440 85.765 ;
        RECT 57.710 85.350 57.880 85.380 ;
        RECT 56.985 84.370 57.880 85.350 ;
        RECT 57.040 83.435 57.210 84.370 ;
        RECT 57.710 84.340 57.880 84.370 ;
        RECT 58.500 84.340 58.670 85.380 ;
        RECT 57.525 83.955 58.440 84.125 ;
        RECT 57.525 83.750 58.360 83.955 ;
        RECT 59.170 83.435 59.340 86.285 ;
        RECT 57.040 83.265 59.340 83.435 ;
        RECT 59.740 83.435 59.910 95.285 ;
        RECT 60.400 94.575 61.400 95.025 ;
        RECT 60.410 84.340 60.580 94.380 ;
        RECT 61.200 84.340 61.370 94.380 ;
        RECT 60.640 83.955 61.140 84.125 ;
        RECT 61.870 83.435 62.040 95.285 ;
        RECT 67.840 95.285 70.140 95.455 ;
        RECT 62.440 86.285 64.740 86.455 ;
        RECT 62.440 85.350 62.610 86.285 ;
        RECT 63.340 85.595 63.840 85.765 ;
        RECT 63.110 85.350 63.280 85.380 ;
        RECT 62.385 84.370 63.280 85.350 ;
        RECT 59.740 83.265 62.040 83.435 ;
        RECT 62.440 83.435 62.610 84.370 ;
        RECT 63.110 84.340 63.280 84.370 ;
        RECT 63.900 84.340 64.070 85.380 ;
        RECT 62.925 83.955 63.840 84.125 ;
        RECT 62.925 83.750 63.760 83.955 ;
        RECT 64.570 83.435 64.740 86.285 ;
        RECT 65.140 86.285 67.440 86.455 ;
        RECT 65.140 85.350 65.310 86.285 ;
        RECT 66.040 85.595 66.540 85.765 ;
        RECT 65.810 85.350 65.980 85.380 ;
        RECT 65.085 84.370 65.980 85.350 ;
        RECT 62.440 83.265 64.740 83.435 ;
        RECT 65.140 83.435 65.310 84.370 ;
        RECT 65.810 84.340 65.980 84.370 ;
        RECT 66.600 84.340 66.770 85.380 ;
        RECT 65.625 83.955 66.540 84.125 ;
        RECT 65.625 83.750 66.460 83.955 ;
        RECT 67.270 83.435 67.440 86.285 ;
        RECT 65.140 83.265 67.440 83.435 ;
        RECT 67.840 83.435 68.010 95.285 ;
        RECT 68.500 94.575 69.500 95.025 ;
        RECT 68.510 84.340 68.680 94.380 ;
        RECT 69.300 84.340 69.470 94.380 ;
        RECT 68.740 83.955 69.240 84.125 ;
        RECT 69.970 83.435 70.140 95.285 ;
        RECT 67.840 83.265 70.140 83.435 ;
        RECT 70.540 95.285 72.840 95.455 ;
        RECT 70.540 83.435 70.710 95.285 ;
        RECT 71.200 94.575 72.200 95.025 ;
        RECT 71.210 84.340 71.380 94.380 ;
        RECT 72.000 84.340 72.170 94.380 ;
        RECT 71.440 83.955 71.940 84.125 ;
        RECT 72.670 83.435 72.840 95.285 ;
        RECT 70.540 83.265 72.840 83.435 ;
        RECT 48.255 81.630 49.905 81.800 ;
        RECT 57.040 82.195 59.340 82.365 ;
        RECT 48.685 81.580 49.475 81.630 ;
        RECT 57.040 81.255 57.210 82.195 ;
        RECT 57.420 81.505 58.460 81.950 ;
        RECT 57.710 81.255 57.880 81.335 ;
        RECT 57.035 80.725 57.880 81.255 ;
        RECT 57.040 79.785 57.210 80.725 ;
        RECT 57.710 80.645 57.880 80.725 ;
        RECT 58.500 80.645 58.670 81.335 ;
        RECT 57.940 80.305 58.440 80.475 ;
        RECT 59.170 79.785 59.340 82.195 ;
        RECT 57.040 79.615 59.340 79.785 ;
        RECT 59.740 82.195 62.040 82.365 ;
        RECT 45.115 73.765 47.415 73.935 ;
        RECT 59.740 73.935 59.910 82.195 ;
        RECT 60.640 81.505 61.140 81.675 ;
        RECT 60.410 74.795 60.580 81.335 ;
        RECT 61.200 74.795 61.370 81.335 ;
        RECT 60.400 74.225 61.400 74.625 ;
        RECT 61.870 73.935 62.040 82.195 ;
        RECT 62.440 82.195 64.740 82.365 ;
        RECT 62.440 81.255 62.610 82.195 ;
        RECT 62.820 81.505 63.860 81.950 ;
        RECT 63.110 81.255 63.280 81.335 ;
        RECT 62.435 80.725 63.280 81.255 ;
        RECT 62.440 79.785 62.610 80.725 ;
        RECT 63.110 80.645 63.280 80.725 ;
        RECT 63.900 80.645 64.070 81.335 ;
        RECT 63.340 80.305 63.840 80.475 ;
        RECT 64.570 79.785 64.740 82.195 ;
        RECT 65.140 82.195 67.440 82.365 ;
        RECT 65.140 81.255 65.310 82.195 ;
        RECT 65.520 81.505 66.560 81.950 ;
        RECT 65.810 81.255 65.980 81.335 ;
        RECT 65.135 80.725 65.980 81.255 ;
        RECT 62.440 79.615 64.740 79.785 ;
        RECT 65.140 79.785 65.310 80.725 ;
        RECT 65.810 80.645 65.980 80.725 ;
        RECT 66.600 80.645 66.770 81.335 ;
        RECT 66.040 80.305 66.540 80.475 ;
        RECT 67.270 79.785 67.440 82.195 ;
        RECT 65.140 79.615 67.440 79.785 ;
        RECT 67.840 82.195 70.140 82.365 ;
        RECT 59.740 73.765 62.040 73.935 ;
        RECT 67.840 73.935 68.010 82.195 ;
        RECT 68.740 81.505 69.240 81.675 ;
        RECT 68.510 74.795 68.680 81.335 ;
        RECT 69.300 74.795 69.470 81.335 ;
        RECT 68.500 74.225 69.500 74.625 ;
        RECT 69.970 73.935 70.140 82.195 ;
        RECT 67.840 73.765 70.140 73.935 ;
        RECT 70.540 82.195 72.840 82.365 ;
        RECT 70.540 73.935 70.710 82.195 ;
        RECT 71.440 81.505 71.940 81.675 ;
        RECT 71.210 74.795 71.380 81.335 ;
        RECT 72.000 74.795 72.170 81.335 ;
        RECT 71.200 74.225 72.200 74.625 ;
        RECT 72.670 73.935 72.840 82.195 ;
        RECT 73.680 81.800 73.850 95.830 ;
        RECT 74.085 95.780 74.925 95.830 ;
        RECT 74.280 93.115 74.730 95.425 ;
        RECT 74.280 82.205 74.730 84.515 ;
        RECT 74.110 81.800 74.900 81.850 ;
        RECT 75.160 81.800 75.330 95.830 ;
        RECT 99.105 95.830 100.755 96.000 ;
        RECT 85.165 95.285 87.465 95.455 ;
        RECT 82.465 86.285 84.765 86.455 ;
        RECT 82.465 85.350 82.635 86.285 ;
        RECT 83.365 85.595 83.865 85.765 ;
        RECT 83.135 85.350 83.305 85.380 ;
        RECT 82.410 84.370 83.305 85.350 ;
        RECT 82.465 83.435 82.635 84.370 ;
        RECT 83.135 84.340 83.305 84.370 ;
        RECT 83.925 84.340 84.095 85.380 ;
        RECT 82.950 83.955 83.865 84.125 ;
        RECT 82.950 83.750 83.785 83.955 ;
        RECT 84.595 83.435 84.765 86.285 ;
        RECT 82.465 83.265 84.765 83.435 ;
        RECT 85.165 83.435 85.335 95.285 ;
        RECT 85.825 94.575 86.825 95.025 ;
        RECT 85.835 84.340 86.005 94.380 ;
        RECT 86.625 84.340 86.795 94.380 ;
        RECT 86.065 83.955 86.565 84.125 ;
        RECT 87.295 83.435 87.465 95.285 ;
        RECT 93.265 95.285 95.565 95.455 ;
        RECT 87.865 86.285 90.165 86.455 ;
        RECT 87.865 85.350 88.035 86.285 ;
        RECT 88.765 85.595 89.265 85.765 ;
        RECT 88.535 85.350 88.705 85.380 ;
        RECT 87.810 84.370 88.705 85.350 ;
        RECT 85.165 83.265 87.465 83.435 ;
        RECT 87.865 83.435 88.035 84.370 ;
        RECT 88.535 84.340 88.705 84.370 ;
        RECT 89.325 84.340 89.495 85.380 ;
        RECT 88.350 83.955 89.265 84.125 ;
        RECT 88.350 83.750 89.185 83.955 ;
        RECT 89.995 83.435 90.165 86.285 ;
        RECT 90.565 86.285 92.865 86.455 ;
        RECT 90.565 85.350 90.735 86.285 ;
        RECT 91.465 85.595 91.965 85.765 ;
        RECT 91.235 85.350 91.405 85.380 ;
        RECT 90.510 84.370 91.405 85.350 ;
        RECT 87.865 83.265 90.165 83.435 ;
        RECT 90.565 83.435 90.735 84.370 ;
        RECT 91.235 84.340 91.405 84.370 ;
        RECT 92.025 84.340 92.195 85.380 ;
        RECT 91.050 83.955 91.965 84.125 ;
        RECT 91.050 83.750 91.885 83.955 ;
        RECT 92.695 83.435 92.865 86.285 ;
        RECT 90.565 83.265 92.865 83.435 ;
        RECT 93.265 83.435 93.435 95.285 ;
        RECT 93.925 94.575 94.925 95.025 ;
        RECT 93.935 84.340 94.105 94.380 ;
        RECT 94.725 84.340 94.895 94.380 ;
        RECT 94.165 83.955 94.665 84.125 ;
        RECT 95.395 83.435 95.565 95.285 ;
        RECT 93.265 83.265 95.565 83.435 ;
        RECT 95.965 95.285 98.265 95.455 ;
        RECT 95.965 83.435 96.135 95.285 ;
        RECT 96.625 94.575 97.625 95.025 ;
        RECT 96.635 84.340 96.805 94.380 ;
        RECT 97.425 84.340 97.595 94.380 ;
        RECT 96.865 83.955 97.365 84.125 ;
        RECT 98.095 83.435 98.265 95.285 ;
        RECT 95.965 83.265 98.265 83.435 ;
        RECT 73.680 81.630 75.330 81.800 ;
        RECT 82.465 82.195 84.765 82.365 ;
        RECT 74.110 81.580 74.900 81.630 ;
        RECT 82.465 81.255 82.635 82.195 ;
        RECT 82.845 81.505 83.885 81.950 ;
        RECT 83.135 81.255 83.305 81.335 ;
        RECT 82.460 80.725 83.305 81.255 ;
        RECT 82.465 79.785 82.635 80.725 ;
        RECT 83.135 80.645 83.305 80.725 ;
        RECT 83.925 80.645 84.095 81.335 ;
        RECT 83.365 80.305 83.865 80.475 ;
        RECT 84.595 79.785 84.765 82.195 ;
        RECT 82.465 79.615 84.765 79.785 ;
        RECT 85.165 82.195 87.465 82.365 ;
        RECT 70.540 73.765 72.840 73.935 ;
        RECT 85.165 73.935 85.335 82.195 ;
        RECT 86.065 81.505 86.565 81.675 ;
        RECT 85.835 74.795 86.005 81.335 ;
        RECT 86.625 74.795 86.795 81.335 ;
        RECT 85.825 74.225 86.825 74.625 ;
        RECT 87.295 73.935 87.465 82.195 ;
        RECT 87.865 82.195 90.165 82.365 ;
        RECT 87.865 81.255 88.035 82.195 ;
        RECT 88.245 81.505 89.285 81.950 ;
        RECT 88.535 81.255 88.705 81.335 ;
        RECT 87.860 80.725 88.705 81.255 ;
        RECT 87.865 79.785 88.035 80.725 ;
        RECT 88.535 80.645 88.705 80.725 ;
        RECT 89.325 80.645 89.495 81.335 ;
        RECT 88.765 80.305 89.265 80.475 ;
        RECT 89.995 79.785 90.165 82.195 ;
        RECT 90.565 82.195 92.865 82.365 ;
        RECT 90.565 81.255 90.735 82.195 ;
        RECT 90.945 81.505 91.985 81.950 ;
        RECT 91.235 81.255 91.405 81.335 ;
        RECT 90.560 80.725 91.405 81.255 ;
        RECT 87.865 79.615 90.165 79.785 ;
        RECT 90.565 79.785 90.735 80.725 ;
        RECT 91.235 80.645 91.405 80.725 ;
        RECT 92.025 80.645 92.195 81.335 ;
        RECT 91.465 80.305 91.965 80.475 ;
        RECT 92.695 79.785 92.865 82.195 ;
        RECT 90.565 79.615 92.865 79.785 ;
        RECT 93.265 82.195 95.565 82.365 ;
        RECT 85.165 73.765 87.465 73.935 ;
        RECT 93.265 73.935 93.435 82.195 ;
        RECT 94.165 81.505 94.665 81.675 ;
        RECT 93.935 74.795 94.105 81.335 ;
        RECT 94.725 74.795 94.895 81.335 ;
        RECT 93.925 74.225 94.925 74.625 ;
        RECT 95.395 73.935 95.565 82.195 ;
        RECT 93.265 73.765 95.565 73.935 ;
        RECT 95.965 82.195 98.265 82.365 ;
        RECT 95.965 73.935 96.135 82.195 ;
        RECT 96.865 81.505 97.365 81.675 ;
        RECT 96.635 74.795 96.805 81.335 ;
        RECT 97.425 74.795 97.595 81.335 ;
        RECT 96.625 74.225 97.625 74.625 ;
        RECT 98.095 73.935 98.265 82.195 ;
        RECT 99.105 81.800 99.275 95.830 ;
        RECT 99.510 95.780 100.350 95.830 ;
        RECT 99.705 93.115 100.155 95.425 ;
        RECT 99.705 82.205 100.155 84.515 ;
        RECT 99.535 81.800 100.325 81.850 ;
        RECT 100.585 81.800 100.755 95.830 ;
        RECT 124.530 95.830 126.180 96.000 ;
        RECT 110.590 95.285 112.890 95.455 ;
        RECT 107.890 86.285 110.190 86.455 ;
        RECT 107.890 85.350 108.060 86.285 ;
        RECT 108.790 85.595 109.290 85.765 ;
        RECT 108.560 85.350 108.730 85.380 ;
        RECT 107.835 84.370 108.730 85.350 ;
        RECT 107.890 83.435 108.060 84.370 ;
        RECT 108.560 84.340 108.730 84.370 ;
        RECT 109.350 84.340 109.520 85.380 ;
        RECT 108.375 83.955 109.290 84.125 ;
        RECT 108.375 83.750 109.210 83.955 ;
        RECT 110.020 83.435 110.190 86.285 ;
        RECT 107.890 83.265 110.190 83.435 ;
        RECT 110.590 83.435 110.760 95.285 ;
        RECT 111.250 94.575 112.250 95.025 ;
        RECT 111.260 84.340 111.430 94.380 ;
        RECT 112.050 84.340 112.220 94.380 ;
        RECT 111.490 83.955 111.990 84.125 ;
        RECT 112.720 83.435 112.890 95.285 ;
        RECT 118.690 95.285 120.990 95.455 ;
        RECT 113.290 86.285 115.590 86.455 ;
        RECT 113.290 85.350 113.460 86.285 ;
        RECT 114.190 85.595 114.690 85.765 ;
        RECT 113.960 85.350 114.130 85.380 ;
        RECT 113.235 84.370 114.130 85.350 ;
        RECT 110.590 83.265 112.890 83.435 ;
        RECT 113.290 83.435 113.460 84.370 ;
        RECT 113.960 84.340 114.130 84.370 ;
        RECT 114.750 84.340 114.920 85.380 ;
        RECT 113.775 83.955 114.690 84.125 ;
        RECT 113.775 83.750 114.610 83.955 ;
        RECT 115.420 83.435 115.590 86.285 ;
        RECT 115.990 86.285 118.290 86.455 ;
        RECT 115.990 85.350 116.160 86.285 ;
        RECT 116.890 85.595 117.390 85.765 ;
        RECT 116.660 85.350 116.830 85.380 ;
        RECT 115.935 84.370 116.830 85.350 ;
        RECT 113.290 83.265 115.590 83.435 ;
        RECT 115.990 83.435 116.160 84.370 ;
        RECT 116.660 84.340 116.830 84.370 ;
        RECT 117.450 84.340 117.620 85.380 ;
        RECT 116.475 83.955 117.390 84.125 ;
        RECT 116.475 83.750 117.310 83.955 ;
        RECT 118.120 83.435 118.290 86.285 ;
        RECT 115.990 83.265 118.290 83.435 ;
        RECT 118.690 83.435 118.860 95.285 ;
        RECT 119.350 94.575 120.350 95.025 ;
        RECT 119.360 84.340 119.530 94.380 ;
        RECT 120.150 84.340 120.320 94.380 ;
        RECT 119.590 83.955 120.090 84.125 ;
        RECT 120.820 83.435 120.990 95.285 ;
        RECT 118.690 83.265 120.990 83.435 ;
        RECT 121.390 95.285 123.690 95.455 ;
        RECT 121.390 83.435 121.560 95.285 ;
        RECT 122.050 94.575 123.050 95.025 ;
        RECT 122.060 84.340 122.230 94.380 ;
        RECT 122.850 84.340 123.020 94.380 ;
        RECT 122.290 83.955 122.790 84.125 ;
        RECT 123.520 83.435 123.690 95.285 ;
        RECT 121.390 83.265 123.690 83.435 ;
        RECT 99.105 81.630 100.755 81.800 ;
        RECT 107.890 82.195 110.190 82.365 ;
        RECT 99.535 81.580 100.325 81.630 ;
        RECT 107.890 81.255 108.060 82.195 ;
        RECT 108.270 81.505 109.310 81.950 ;
        RECT 108.560 81.255 108.730 81.335 ;
        RECT 107.885 80.725 108.730 81.255 ;
        RECT 107.890 79.785 108.060 80.725 ;
        RECT 108.560 80.645 108.730 80.725 ;
        RECT 109.350 80.645 109.520 81.335 ;
        RECT 108.790 80.305 109.290 80.475 ;
        RECT 110.020 79.785 110.190 82.195 ;
        RECT 107.890 79.615 110.190 79.785 ;
        RECT 110.590 82.195 112.890 82.365 ;
        RECT 95.965 73.765 98.265 73.935 ;
        RECT 110.590 73.935 110.760 82.195 ;
        RECT 111.490 81.505 111.990 81.675 ;
        RECT 111.260 74.795 111.430 81.335 ;
        RECT 112.050 74.795 112.220 81.335 ;
        RECT 111.250 74.225 112.250 74.625 ;
        RECT 112.720 73.935 112.890 82.195 ;
        RECT 113.290 82.195 115.590 82.365 ;
        RECT 113.290 81.255 113.460 82.195 ;
        RECT 113.670 81.505 114.710 81.950 ;
        RECT 113.960 81.255 114.130 81.335 ;
        RECT 113.285 80.725 114.130 81.255 ;
        RECT 113.290 79.785 113.460 80.725 ;
        RECT 113.960 80.645 114.130 80.725 ;
        RECT 114.750 80.645 114.920 81.335 ;
        RECT 114.190 80.305 114.690 80.475 ;
        RECT 115.420 79.785 115.590 82.195 ;
        RECT 115.990 82.195 118.290 82.365 ;
        RECT 115.990 81.255 116.160 82.195 ;
        RECT 116.370 81.505 117.410 81.950 ;
        RECT 116.660 81.255 116.830 81.335 ;
        RECT 115.985 80.725 116.830 81.255 ;
        RECT 113.290 79.615 115.590 79.785 ;
        RECT 115.990 79.785 116.160 80.725 ;
        RECT 116.660 80.645 116.830 80.725 ;
        RECT 117.450 80.645 117.620 81.335 ;
        RECT 116.890 80.305 117.390 80.475 ;
        RECT 118.120 79.785 118.290 82.195 ;
        RECT 115.990 79.615 118.290 79.785 ;
        RECT 118.690 82.195 120.990 82.365 ;
        RECT 110.590 73.765 112.890 73.935 ;
        RECT 118.690 73.935 118.860 82.195 ;
        RECT 119.590 81.505 120.090 81.675 ;
        RECT 119.360 74.795 119.530 81.335 ;
        RECT 120.150 74.795 120.320 81.335 ;
        RECT 119.350 74.225 120.350 74.625 ;
        RECT 120.820 73.935 120.990 82.195 ;
        RECT 118.690 73.765 120.990 73.935 ;
        RECT 121.390 82.195 123.690 82.365 ;
        RECT 121.390 73.935 121.560 82.195 ;
        RECT 122.290 81.505 122.790 81.675 ;
        RECT 122.060 74.795 122.230 81.335 ;
        RECT 122.850 74.795 123.020 81.335 ;
        RECT 122.050 74.225 123.050 74.625 ;
        RECT 123.520 73.935 123.690 82.195 ;
        RECT 124.530 81.800 124.700 95.830 ;
        RECT 124.935 95.780 125.775 95.830 ;
        RECT 125.130 93.115 125.580 95.425 ;
        RECT 125.130 82.205 125.580 84.515 ;
        RECT 124.960 81.800 125.750 81.850 ;
        RECT 126.010 81.800 126.180 95.830 ;
        RECT 149.955 95.830 151.605 96.000 ;
        RECT 136.015 95.285 138.315 95.455 ;
        RECT 133.315 86.285 135.615 86.455 ;
        RECT 133.315 85.350 133.485 86.285 ;
        RECT 134.215 85.595 134.715 85.765 ;
        RECT 133.985 85.350 134.155 85.380 ;
        RECT 133.260 84.370 134.155 85.350 ;
        RECT 133.315 83.435 133.485 84.370 ;
        RECT 133.985 84.340 134.155 84.370 ;
        RECT 134.775 84.340 134.945 85.380 ;
        RECT 133.800 83.955 134.715 84.125 ;
        RECT 133.800 83.750 134.635 83.955 ;
        RECT 135.445 83.435 135.615 86.285 ;
        RECT 133.315 83.265 135.615 83.435 ;
        RECT 136.015 83.435 136.185 95.285 ;
        RECT 136.675 94.575 137.675 95.025 ;
        RECT 136.685 84.340 136.855 94.380 ;
        RECT 137.475 84.340 137.645 94.380 ;
        RECT 136.915 83.955 137.415 84.125 ;
        RECT 138.145 83.435 138.315 95.285 ;
        RECT 144.115 95.285 146.415 95.455 ;
        RECT 138.715 86.285 141.015 86.455 ;
        RECT 138.715 85.350 138.885 86.285 ;
        RECT 139.615 85.595 140.115 85.765 ;
        RECT 139.385 85.350 139.555 85.380 ;
        RECT 138.660 84.370 139.555 85.350 ;
        RECT 136.015 83.265 138.315 83.435 ;
        RECT 138.715 83.435 138.885 84.370 ;
        RECT 139.385 84.340 139.555 84.370 ;
        RECT 140.175 84.340 140.345 85.380 ;
        RECT 139.200 83.955 140.115 84.125 ;
        RECT 139.200 83.750 140.035 83.955 ;
        RECT 140.845 83.435 141.015 86.285 ;
        RECT 141.415 86.285 143.715 86.455 ;
        RECT 141.415 85.350 141.585 86.285 ;
        RECT 142.315 85.595 142.815 85.765 ;
        RECT 142.085 85.350 142.255 85.380 ;
        RECT 141.360 84.370 142.255 85.350 ;
        RECT 138.715 83.265 141.015 83.435 ;
        RECT 141.415 83.435 141.585 84.370 ;
        RECT 142.085 84.340 142.255 84.370 ;
        RECT 142.875 84.340 143.045 85.380 ;
        RECT 141.900 83.955 142.815 84.125 ;
        RECT 141.900 83.750 142.735 83.955 ;
        RECT 143.545 83.435 143.715 86.285 ;
        RECT 141.415 83.265 143.715 83.435 ;
        RECT 144.115 83.435 144.285 95.285 ;
        RECT 144.775 94.575 145.775 95.025 ;
        RECT 144.785 84.340 144.955 94.380 ;
        RECT 145.575 84.340 145.745 94.380 ;
        RECT 145.015 83.955 145.515 84.125 ;
        RECT 146.245 83.435 146.415 95.285 ;
        RECT 144.115 83.265 146.415 83.435 ;
        RECT 146.815 95.285 149.115 95.455 ;
        RECT 146.815 83.435 146.985 95.285 ;
        RECT 147.475 94.575 148.475 95.025 ;
        RECT 147.485 84.340 147.655 94.380 ;
        RECT 148.275 84.340 148.445 94.380 ;
        RECT 147.715 83.955 148.215 84.125 ;
        RECT 148.945 83.435 149.115 95.285 ;
        RECT 146.815 83.265 149.115 83.435 ;
        RECT 124.530 81.630 126.180 81.800 ;
        RECT 133.315 82.195 135.615 82.365 ;
        RECT 124.960 81.580 125.750 81.630 ;
        RECT 133.315 81.255 133.485 82.195 ;
        RECT 133.695 81.505 134.735 81.950 ;
        RECT 133.985 81.255 134.155 81.335 ;
        RECT 133.310 80.725 134.155 81.255 ;
        RECT 133.315 79.785 133.485 80.725 ;
        RECT 133.985 80.645 134.155 80.725 ;
        RECT 134.775 80.645 134.945 81.335 ;
        RECT 134.215 80.305 134.715 80.475 ;
        RECT 135.445 79.785 135.615 82.195 ;
        RECT 133.315 79.615 135.615 79.785 ;
        RECT 136.015 82.195 138.315 82.365 ;
        RECT 121.390 73.765 123.690 73.935 ;
        RECT 136.015 73.935 136.185 82.195 ;
        RECT 136.915 81.505 137.415 81.675 ;
        RECT 136.685 74.795 136.855 81.335 ;
        RECT 137.475 74.795 137.645 81.335 ;
        RECT 136.675 74.225 137.675 74.625 ;
        RECT 138.145 73.935 138.315 82.195 ;
        RECT 138.715 82.195 141.015 82.365 ;
        RECT 138.715 81.255 138.885 82.195 ;
        RECT 139.095 81.505 140.135 81.950 ;
        RECT 139.385 81.255 139.555 81.335 ;
        RECT 138.710 80.725 139.555 81.255 ;
        RECT 138.715 79.785 138.885 80.725 ;
        RECT 139.385 80.645 139.555 80.725 ;
        RECT 140.175 80.645 140.345 81.335 ;
        RECT 139.615 80.305 140.115 80.475 ;
        RECT 140.845 79.785 141.015 82.195 ;
        RECT 141.415 82.195 143.715 82.365 ;
        RECT 141.415 81.255 141.585 82.195 ;
        RECT 141.795 81.505 142.835 81.950 ;
        RECT 142.085 81.255 142.255 81.335 ;
        RECT 141.410 80.725 142.255 81.255 ;
        RECT 138.715 79.615 141.015 79.785 ;
        RECT 141.415 79.785 141.585 80.725 ;
        RECT 142.085 80.645 142.255 80.725 ;
        RECT 142.875 80.645 143.045 81.335 ;
        RECT 142.315 80.305 142.815 80.475 ;
        RECT 143.545 79.785 143.715 82.195 ;
        RECT 141.415 79.615 143.715 79.785 ;
        RECT 144.115 82.195 146.415 82.365 ;
        RECT 136.015 73.765 138.315 73.935 ;
        RECT 144.115 73.935 144.285 82.195 ;
        RECT 145.015 81.505 145.515 81.675 ;
        RECT 144.785 74.795 144.955 81.335 ;
        RECT 145.575 74.795 145.745 81.335 ;
        RECT 144.775 74.225 145.775 74.625 ;
        RECT 146.245 73.935 146.415 82.195 ;
        RECT 144.115 73.765 146.415 73.935 ;
        RECT 146.815 82.195 149.115 82.365 ;
        RECT 146.815 73.935 146.985 82.195 ;
        RECT 147.715 81.505 148.215 81.675 ;
        RECT 147.485 74.795 147.655 81.335 ;
        RECT 148.275 74.795 148.445 81.335 ;
        RECT 147.475 74.225 148.475 74.625 ;
        RECT 148.945 73.935 149.115 82.195 ;
        RECT 149.955 81.800 150.125 95.830 ;
        RECT 150.360 95.780 151.200 95.830 ;
        RECT 150.555 93.115 151.005 95.425 ;
        RECT 150.555 82.205 151.005 84.515 ;
        RECT 150.385 81.800 151.175 81.850 ;
        RECT 151.435 81.800 151.605 95.830 ;
        RECT 149.955 81.630 151.605 81.800 ;
        RECT 150.385 81.580 151.175 81.630 ;
        RECT 146.815 73.765 149.115 73.935 ;
        RECT 8.890 68.435 11.190 68.605 ;
        RECT 6.190 59.435 8.490 59.605 ;
        RECT 6.190 58.500 6.360 59.435 ;
        RECT 7.090 58.745 7.590 58.915 ;
        RECT 6.860 58.500 7.030 58.530 ;
        RECT 6.135 57.520 7.030 58.500 ;
        RECT 6.190 56.585 6.360 57.520 ;
        RECT 6.860 57.490 7.030 57.520 ;
        RECT 7.650 57.490 7.820 58.530 ;
        RECT 6.675 57.105 7.590 57.275 ;
        RECT 6.675 56.900 7.510 57.105 ;
        RECT 8.320 56.585 8.490 59.435 ;
        RECT 6.190 56.415 8.490 56.585 ;
        RECT 8.890 56.585 9.060 68.435 ;
        RECT 9.550 67.725 10.550 68.175 ;
        RECT 9.560 57.490 9.730 67.530 ;
        RECT 10.350 57.490 10.520 67.530 ;
        RECT 9.790 57.105 10.290 57.275 ;
        RECT 11.020 56.585 11.190 68.435 ;
        RECT 16.990 68.435 19.290 68.605 ;
        RECT 11.590 59.435 13.890 59.605 ;
        RECT 11.590 58.500 11.760 59.435 ;
        RECT 12.490 58.745 12.990 58.915 ;
        RECT 12.260 58.500 12.430 58.530 ;
        RECT 11.535 57.520 12.430 58.500 ;
        RECT 8.890 56.415 11.190 56.585 ;
        RECT 11.590 56.585 11.760 57.520 ;
        RECT 12.260 57.490 12.430 57.520 ;
        RECT 13.050 57.490 13.220 58.530 ;
        RECT 12.075 57.105 12.990 57.275 ;
        RECT 12.075 56.900 12.910 57.105 ;
        RECT 13.720 56.585 13.890 59.435 ;
        RECT 14.290 59.435 16.590 59.605 ;
        RECT 14.290 58.500 14.460 59.435 ;
        RECT 15.190 58.745 15.690 58.915 ;
        RECT 14.960 58.500 15.130 58.530 ;
        RECT 14.235 57.520 15.130 58.500 ;
        RECT 11.590 56.415 13.890 56.585 ;
        RECT 14.290 56.585 14.460 57.520 ;
        RECT 14.960 57.490 15.130 57.520 ;
        RECT 15.750 57.490 15.920 58.530 ;
        RECT 14.775 57.105 15.690 57.275 ;
        RECT 14.775 56.900 15.610 57.105 ;
        RECT 16.420 56.585 16.590 59.435 ;
        RECT 14.290 56.415 16.590 56.585 ;
        RECT 16.990 56.585 17.160 68.435 ;
        RECT 17.650 67.725 18.650 68.175 ;
        RECT 17.660 57.490 17.830 67.530 ;
        RECT 18.450 57.490 18.620 67.530 ;
        RECT 17.890 57.105 18.390 57.275 ;
        RECT 19.120 56.585 19.290 68.435 ;
        RECT 16.990 56.415 19.290 56.585 ;
        RECT 19.690 68.435 21.990 68.605 ;
        RECT 19.690 56.585 19.860 68.435 ;
        RECT 20.350 67.725 21.350 68.175 ;
        RECT 20.360 57.490 20.530 67.530 ;
        RECT 21.150 57.490 21.320 67.530 ;
        RECT 20.590 57.105 21.090 57.275 ;
        RECT 21.820 56.585 21.990 68.435 ;
        RECT 22.885 68.435 25.185 68.605 ;
        RECT 22.885 67.450 23.055 68.435 ;
        RECT 23.785 67.745 24.285 67.915 ;
        RECT 23.555 67.450 23.725 67.530 ;
        RECT 24.345 67.525 24.515 67.530 ;
        RECT 22.885 66.575 23.725 67.450 ;
        RECT 22.885 65.585 23.055 66.575 ;
        RECT 23.555 66.490 23.725 66.575 ;
        RECT 24.295 66.495 24.770 67.525 ;
        RECT 24.345 66.490 24.515 66.495 ;
        RECT 23.545 65.850 24.520 66.300 ;
        RECT 25.015 65.585 25.185 68.435 ;
        RECT 22.885 65.415 25.185 65.585 ;
        RECT 25.585 68.435 27.885 68.605 ;
        RECT 25.585 65.585 25.755 68.435 ;
        RECT 26.485 67.745 26.985 67.915 ;
        RECT 26.255 67.525 26.425 67.530 ;
        RECT 25.980 66.495 26.475 67.525 ;
        RECT 27.045 67.500 27.215 67.530 ;
        RECT 27.715 67.500 27.885 68.435 ;
        RECT 28.285 68.435 30.585 68.605 ;
        RECT 28.285 67.500 28.455 68.435 ;
        RECT 29.185 67.745 29.685 67.915 ;
        RECT 28.955 67.500 29.125 67.530 ;
        RECT 26.970 66.570 27.890 67.500 ;
        RECT 26.255 66.490 26.425 66.495 ;
        RECT 27.045 66.490 27.215 66.570 ;
        RECT 26.245 65.850 27.220 66.300 ;
        RECT 27.715 65.585 27.885 66.570 ;
        RECT 28.230 66.520 29.125 67.500 ;
        RECT 25.585 65.415 27.885 65.585 ;
        RECT 28.285 65.585 28.455 66.520 ;
        RECT 28.955 66.490 29.125 66.520 ;
        RECT 29.745 66.490 29.915 67.530 ;
        RECT 28.770 66.105 29.685 66.275 ;
        RECT 28.770 65.900 29.605 66.105 ;
        RECT 30.415 65.585 30.585 68.435 ;
        RECT 28.285 65.415 30.585 65.585 ;
        RECT 34.315 68.435 36.615 68.605 ;
        RECT 22.885 64.345 25.185 64.515 ;
        RECT 22.885 61.935 23.055 64.345 ;
        RECT 23.545 63.675 24.520 64.100 ;
        RECT 25.015 64.035 25.185 64.345 ;
        RECT 25.585 64.345 27.885 64.515 ;
        RECT 25.585 64.035 25.755 64.345 ;
        RECT 23.785 63.655 24.285 63.675 ;
        RECT 23.555 63.480 23.725 63.485 ;
        RECT 24.345 63.480 24.515 63.485 ;
        RECT 23.455 62.800 23.825 63.480 ;
        RECT 24.245 62.800 24.615 63.480 ;
        RECT 23.555 62.795 23.725 62.800 ;
        RECT 24.345 62.795 24.515 62.800 ;
        RECT 23.785 62.455 24.285 62.625 ;
        RECT 25.015 62.245 25.755 64.035 ;
        RECT 26.245 63.675 27.220 64.100 ;
        RECT 26.485 63.655 26.985 63.675 ;
        RECT 26.255 63.480 26.425 63.485 ;
        RECT 26.155 62.800 26.525 63.480 ;
        RECT 27.045 63.405 27.215 63.485 ;
        RECT 27.715 63.405 27.885 64.345 ;
        RECT 28.285 64.345 30.585 64.515 ;
        RECT 28.285 63.405 28.455 64.345 ;
        RECT 28.665 63.655 29.705 64.100 ;
        RECT 28.955 63.405 29.125 63.485 ;
        RECT 26.970 62.825 27.890 63.405 ;
        RECT 28.280 62.875 29.125 63.405 ;
        RECT 26.255 62.795 26.425 62.800 ;
        RECT 27.045 62.795 27.215 62.825 ;
        RECT 26.485 62.455 26.985 62.625 ;
        RECT 25.015 61.935 25.185 62.245 ;
        RECT 22.885 61.765 25.185 61.935 ;
        RECT 25.585 61.935 25.755 62.245 ;
        RECT 27.715 61.935 27.885 62.825 ;
        RECT 25.585 61.765 27.885 61.935 ;
        RECT 28.285 61.935 28.455 62.875 ;
        RECT 28.955 62.795 29.125 62.875 ;
        RECT 29.745 62.795 29.915 63.485 ;
        RECT 29.185 62.455 29.685 62.625 ;
        RECT 30.415 61.935 30.585 64.345 ;
        RECT 28.285 61.765 30.585 61.935 ;
        RECT 31.615 59.435 33.915 59.605 ;
        RECT 31.615 58.500 31.785 59.435 ;
        RECT 32.515 58.745 33.015 58.915 ;
        RECT 32.285 58.500 32.455 58.530 ;
        RECT 31.560 57.520 32.455 58.500 ;
        RECT 19.690 56.415 21.990 56.585 ;
        RECT 31.615 56.585 31.785 57.520 ;
        RECT 32.285 57.490 32.455 57.520 ;
        RECT 33.075 57.490 33.245 58.530 ;
        RECT 32.100 57.105 33.015 57.275 ;
        RECT 32.100 56.900 32.935 57.105 ;
        RECT 33.745 56.585 33.915 59.435 ;
        RECT 31.615 56.415 33.915 56.585 ;
        RECT 34.315 56.585 34.485 68.435 ;
        RECT 34.975 67.725 35.975 68.175 ;
        RECT 34.985 57.490 35.155 67.530 ;
        RECT 35.775 57.490 35.945 67.530 ;
        RECT 35.215 57.105 35.715 57.275 ;
        RECT 36.445 56.585 36.615 68.435 ;
        RECT 42.415 68.435 44.715 68.605 ;
        RECT 37.015 59.435 39.315 59.605 ;
        RECT 37.015 58.500 37.185 59.435 ;
        RECT 37.915 58.745 38.415 58.915 ;
        RECT 37.685 58.500 37.855 58.530 ;
        RECT 36.960 57.520 37.855 58.500 ;
        RECT 34.315 56.415 36.615 56.585 ;
        RECT 37.015 56.585 37.185 57.520 ;
        RECT 37.685 57.490 37.855 57.520 ;
        RECT 38.475 57.490 38.645 58.530 ;
        RECT 37.500 57.105 38.415 57.275 ;
        RECT 37.500 56.900 38.335 57.105 ;
        RECT 39.145 56.585 39.315 59.435 ;
        RECT 39.715 59.435 42.015 59.605 ;
        RECT 39.715 58.500 39.885 59.435 ;
        RECT 40.615 58.745 41.115 58.915 ;
        RECT 40.385 58.500 40.555 58.530 ;
        RECT 39.660 57.520 40.555 58.500 ;
        RECT 37.015 56.415 39.315 56.585 ;
        RECT 39.715 56.585 39.885 57.520 ;
        RECT 40.385 57.490 40.555 57.520 ;
        RECT 41.175 57.490 41.345 58.530 ;
        RECT 40.200 57.105 41.115 57.275 ;
        RECT 40.200 56.900 41.035 57.105 ;
        RECT 41.845 56.585 42.015 59.435 ;
        RECT 39.715 56.415 42.015 56.585 ;
        RECT 42.415 56.585 42.585 68.435 ;
        RECT 43.075 67.725 44.075 68.175 ;
        RECT 43.085 57.490 43.255 67.530 ;
        RECT 43.875 57.490 44.045 67.530 ;
        RECT 43.315 57.105 43.815 57.275 ;
        RECT 44.545 56.585 44.715 68.435 ;
        RECT 42.415 56.415 44.715 56.585 ;
        RECT 45.115 68.435 47.415 68.605 ;
        RECT 45.115 56.585 45.285 68.435 ;
        RECT 45.775 67.725 46.775 68.175 ;
        RECT 45.785 57.490 45.955 67.530 ;
        RECT 46.575 57.490 46.745 67.530 ;
        RECT 46.015 57.105 46.515 57.275 ;
        RECT 47.245 56.585 47.415 68.435 ;
        RECT 59.740 68.435 62.040 68.605 ;
        RECT 57.040 59.435 59.340 59.605 ;
        RECT 57.040 58.500 57.210 59.435 ;
        RECT 57.940 58.745 58.440 58.915 ;
        RECT 57.710 58.500 57.880 58.530 ;
        RECT 56.985 57.520 57.880 58.500 ;
        RECT 45.115 56.415 47.415 56.585 ;
        RECT 57.040 56.585 57.210 57.520 ;
        RECT 57.710 57.490 57.880 57.520 ;
        RECT 58.500 57.490 58.670 58.530 ;
        RECT 57.525 57.105 58.440 57.275 ;
        RECT 57.525 56.900 58.360 57.105 ;
        RECT 59.170 56.585 59.340 59.435 ;
        RECT 57.040 56.415 59.340 56.585 ;
        RECT 59.740 56.585 59.910 68.435 ;
        RECT 60.400 67.725 61.400 68.175 ;
        RECT 60.410 57.490 60.580 67.530 ;
        RECT 61.200 57.490 61.370 67.530 ;
        RECT 60.640 57.105 61.140 57.275 ;
        RECT 61.870 56.585 62.040 68.435 ;
        RECT 67.840 68.435 70.140 68.605 ;
        RECT 62.440 59.435 64.740 59.605 ;
        RECT 62.440 58.500 62.610 59.435 ;
        RECT 63.340 58.745 63.840 58.915 ;
        RECT 63.110 58.500 63.280 58.530 ;
        RECT 62.385 57.520 63.280 58.500 ;
        RECT 59.740 56.415 62.040 56.585 ;
        RECT 62.440 56.585 62.610 57.520 ;
        RECT 63.110 57.490 63.280 57.520 ;
        RECT 63.900 57.490 64.070 58.530 ;
        RECT 62.925 57.105 63.840 57.275 ;
        RECT 62.925 56.900 63.760 57.105 ;
        RECT 64.570 56.585 64.740 59.435 ;
        RECT 65.140 59.435 67.440 59.605 ;
        RECT 65.140 58.500 65.310 59.435 ;
        RECT 66.040 58.745 66.540 58.915 ;
        RECT 65.810 58.500 65.980 58.530 ;
        RECT 65.085 57.520 65.980 58.500 ;
        RECT 62.440 56.415 64.740 56.585 ;
        RECT 65.140 56.585 65.310 57.520 ;
        RECT 65.810 57.490 65.980 57.520 ;
        RECT 66.600 57.490 66.770 58.530 ;
        RECT 65.625 57.105 66.540 57.275 ;
        RECT 65.625 56.900 66.460 57.105 ;
        RECT 67.270 56.585 67.440 59.435 ;
        RECT 65.140 56.415 67.440 56.585 ;
        RECT 67.840 56.585 68.010 68.435 ;
        RECT 68.500 67.725 69.500 68.175 ;
        RECT 68.510 57.490 68.680 67.530 ;
        RECT 69.300 57.490 69.470 67.530 ;
        RECT 68.740 57.105 69.240 57.275 ;
        RECT 69.970 56.585 70.140 68.435 ;
        RECT 67.840 56.415 70.140 56.585 ;
        RECT 70.540 68.435 72.840 68.605 ;
        RECT 70.540 56.585 70.710 68.435 ;
        RECT 71.200 67.725 72.200 68.175 ;
        RECT 71.210 57.490 71.380 67.530 ;
        RECT 72.000 57.490 72.170 67.530 ;
        RECT 71.440 57.105 71.940 57.275 ;
        RECT 72.670 56.585 72.840 68.435 ;
        RECT 73.735 68.435 76.035 68.605 ;
        RECT 73.735 67.450 73.905 68.435 ;
        RECT 74.635 67.745 75.135 67.915 ;
        RECT 74.405 67.450 74.575 67.530 ;
        RECT 75.195 67.525 75.365 67.530 ;
        RECT 73.735 66.575 74.575 67.450 ;
        RECT 73.735 65.585 73.905 66.575 ;
        RECT 74.405 66.490 74.575 66.575 ;
        RECT 75.145 66.495 75.620 67.525 ;
        RECT 75.195 66.490 75.365 66.495 ;
        RECT 74.395 65.850 75.370 66.300 ;
        RECT 75.865 65.585 76.035 68.435 ;
        RECT 73.735 65.415 76.035 65.585 ;
        RECT 76.435 68.435 78.735 68.605 ;
        RECT 76.435 65.585 76.605 68.435 ;
        RECT 77.335 67.745 77.835 67.915 ;
        RECT 77.105 67.525 77.275 67.530 ;
        RECT 76.830 66.495 77.325 67.525 ;
        RECT 77.895 67.500 78.065 67.530 ;
        RECT 78.565 67.500 78.735 68.435 ;
        RECT 79.135 68.435 81.435 68.605 ;
        RECT 79.135 67.500 79.305 68.435 ;
        RECT 80.035 67.745 80.535 67.915 ;
        RECT 79.805 67.500 79.975 67.530 ;
        RECT 77.820 66.570 78.740 67.500 ;
        RECT 77.105 66.490 77.275 66.495 ;
        RECT 77.895 66.490 78.065 66.570 ;
        RECT 77.095 65.850 78.070 66.300 ;
        RECT 78.565 65.585 78.735 66.570 ;
        RECT 79.080 66.520 79.975 67.500 ;
        RECT 76.435 65.415 78.735 65.585 ;
        RECT 79.135 65.585 79.305 66.520 ;
        RECT 79.805 66.490 79.975 66.520 ;
        RECT 80.595 66.490 80.765 67.530 ;
        RECT 79.620 66.105 80.535 66.275 ;
        RECT 79.620 65.900 80.455 66.105 ;
        RECT 81.265 65.585 81.435 68.435 ;
        RECT 79.135 65.415 81.435 65.585 ;
        RECT 85.165 68.435 87.465 68.605 ;
        RECT 73.735 64.345 76.035 64.515 ;
        RECT 73.735 61.935 73.905 64.345 ;
        RECT 74.395 63.675 75.370 64.100 ;
        RECT 75.865 64.035 76.035 64.345 ;
        RECT 76.435 64.345 78.735 64.515 ;
        RECT 76.435 64.035 76.605 64.345 ;
        RECT 74.635 63.655 75.135 63.675 ;
        RECT 74.405 63.480 74.575 63.485 ;
        RECT 75.195 63.480 75.365 63.485 ;
        RECT 74.305 62.800 74.675 63.480 ;
        RECT 75.095 62.800 75.465 63.480 ;
        RECT 74.405 62.795 74.575 62.800 ;
        RECT 75.195 62.795 75.365 62.800 ;
        RECT 74.635 62.455 75.135 62.625 ;
        RECT 75.865 62.245 76.605 64.035 ;
        RECT 77.095 63.675 78.070 64.100 ;
        RECT 77.335 63.655 77.835 63.675 ;
        RECT 77.105 63.480 77.275 63.485 ;
        RECT 77.005 62.800 77.375 63.480 ;
        RECT 77.895 63.405 78.065 63.485 ;
        RECT 78.565 63.405 78.735 64.345 ;
        RECT 79.135 64.345 81.435 64.515 ;
        RECT 79.135 63.405 79.305 64.345 ;
        RECT 79.515 63.655 80.555 64.100 ;
        RECT 79.805 63.405 79.975 63.485 ;
        RECT 77.820 62.825 78.740 63.405 ;
        RECT 79.130 62.875 79.975 63.405 ;
        RECT 77.105 62.795 77.275 62.800 ;
        RECT 77.895 62.795 78.065 62.825 ;
        RECT 77.335 62.455 77.835 62.625 ;
        RECT 75.865 61.935 76.035 62.245 ;
        RECT 73.735 61.765 76.035 61.935 ;
        RECT 76.435 61.935 76.605 62.245 ;
        RECT 78.565 61.935 78.735 62.825 ;
        RECT 76.435 61.765 78.735 61.935 ;
        RECT 79.135 61.935 79.305 62.875 ;
        RECT 79.805 62.795 79.975 62.875 ;
        RECT 80.595 62.795 80.765 63.485 ;
        RECT 80.035 62.455 80.535 62.625 ;
        RECT 81.265 61.935 81.435 64.345 ;
        RECT 79.135 61.765 81.435 61.935 ;
        RECT 82.465 59.435 84.765 59.605 ;
        RECT 82.465 58.500 82.635 59.435 ;
        RECT 83.365 58.745 83.865 58.915 ;
        RECT 83.135 58.500 83.305 58.530 ;
        RECT 82.410 57.520 83.305 58.500 ;
        RECT 70.540 56.415 72.840 56.585 ;
        RECT 82.465 56.585 82.635 57.520 ;
        RECT 83.135 57.490 83.305 57.520 ;
        RECT 83.925 57.490 84.095 58.530 ;
        RECT 82.950 57.105 83.865 57.275 ;
        RECT 82.950 56.900 83.785 57.105 ;
        RECT 84.595 56.585 84.765 59.435 ;
        RECT 82.465 56.415 84.765 56.585 ;
        RECT 85.165 56.585 85.335 68.435 ;
        RECT 85.825 67.725 86.825 68.175 ;
        RECT 85.835 57.490 86.005 67.530 ;
        RECT 86.625 57.490 86.795 67.530 ;
        RECT 86.065 57.105 86.565 57.275 ;
        RECT 87.295 56.585 87.465 68.435 ;
        RECT 93.265 68.435 95.565 68.605 ;
        RECT 87.865 59.435 90.165 59.605 ;
        RECT 87.865 58.500 88.035 59.435 ;
        RECT 88.765 58.745 89.265 58.915 ;
        RECT 88.535 58.500 88.705 58.530 ;
        RECT 87.810 57.520 88.705 58.500 ;
        RECT 85.165 56.415 87.465 56.585 ;
        RECT 87.865 56.585 88.035 57.520 ;
        RECT 88.535 57.490 88.705 57.520 ;
        RECT 89.325 57.490 89.495 58.530 ;
        RECT 88.350 57.105 89.265 57.275 ;
        RECT 88.350 56.900 89.185 57.105 ;
        RECT 89.995 56.585 90.165 59.435 ;
        RECT 90.565 59.435 92.865 59.605 ;
        RECT 90.565 58.500 90.735 59.435 ;
        RECT 91.465 58.745 91.965 58.915 ;
        RECT 91.235 58.500 91.405 58.530 ;
        RECT 90.510 57.520 91.405 58.500 ;
        RECT 87.865 56.415 90.165 56.585 ;
        RECT 90.565 56.585 90.735 57.520 ;
        RECT 91.235 57.490 91.405 57.520 ;
        RECT 92.025 57.490 92.195 58.530 ;
        RECT 91.050 57.105 91.965 57.275 ;
        RECT 91.050 56.900 91.885 57.105 ;
        RECT 92.695 56.585 92.865 59.435 ;
        RECT 90.565 56.415 92.865 56.585 ;
        RECT 93.265 56.585 93.435 68.435 ;
        RECT 93.925 67.725 94.925 68.175 ;
        RECT 93.935 57.490 94.105 67.530 ;
        RECT 94.725 57.490 94.895 67.530 ;
        RECT 94.165 57.105 94.665 57.275 ;
        RECT 95.395 56.585 95.565 68.435 ;
        RECT 93.265 56.415 95.565 56.585 ;
        RECT 95.965 68.435 98.265 68.605 ;
        RECT 95.965 56.585 96.135 68.435 ;
        RECT 96.625 67.725 97.625 68.175 ;
        RECT 96.635 57.490 96.805 67.530 ;
        RECT 97.425 57.490 97.595 67.530 ;
        RECT 96.865 57.105 97.365 57.275 ;
        RECT 98.095 56.585 98.265 68.435 ;
        RECT 110.590 68.435 112.890 68.605 ;
        RECT 107.890 59.435 110.190 59.605 ;
        RECT 107.890 58.500 108.060 59.435 ;
        RECT 108.790 58.745 109.290 58.915 ;
        RECT 108.560 58.500 108.730 58.530 ;
        RECT 107.835 57.520 108.730 58.500 ;
        RECT 95.965 56.415 98.265 56.585 ;
        RECT 107.890 56.585 108.060 57.520 ;
        RECT 108.560 57.490 108.730 57.520 ;
        RECT 109.350 57.490 109.520 58.530 ;
        RECT 108.375 57.105 109.290 57.275 ;
        RECT 108.375 56.900 109.210 57.105 ;
        RECT 110.020 56.585 110.190 59.435 ;
        RECT 107.890 56.415 110.190 56.585 ;
        RECT 110.590 56.585 110.760 68.435 ;
        RECT 111.250 67.725 112.250 68.175 ;
        RECT 111.260 57.490 111.430 67.530 ;
        RECT 112.050 57.490 112.220 67.530 ;
        RECT 111.490 57.105 111.990 57.275 ;
        RECT 112.720 56.585 112.890 68.435 ;
        RECT 118.690 68.435 120.990 68.605 ;
        RECT 113.290 59.435 115.590 59.605 ;
        RECT 113.290 58.500 113.460 59.435 ;
        RECT 114.190 58.745 114.690 58.915 ;
        RECT 113.960 58.500 114.130 58.530 ;
        RECT 113.235 57.520 114.130 58.500 ;
        RECT 110.590 56.415 112.890 56.585 ;
        RECT 113.290 56.585 113.460 57.520 ;
        RECT 113.960 57.490 114.130 57.520 ;
        RECT 114.750 57.490 114.920 58.530 ;
        RECT 113.775 57.105 114.690 57.275 ;
        RECT 113.775 56.900 114.610 57.105 ;
        RECT 115.420 56.585 115.590 59.435 ;
        RECT 115.990 59.435 118.290 59.605 ;
        RECT 115.990 58.500 116.160 59.435 ;
        RECT 116.890 58.745 117.390 58.915 ;
        RECT 116.660 58.500 116.830 58.530 ;
        RECT 115.935 57.520 116.830 58.500 ;
        RECT 113.290 56.415 115.590 56.585 ;
        RECT 115.990 56.585 116.160 57.520 ;
        RECT 116.660 57.490 116.830 57.520 ;
        RECT 117.450 57.490 117.620 58.530 ;
        RECT 116.475 57.105 117.390 57.275 ;
        RECT 116.475 56.900 117.310 57.105 ;
        RECT 118.120 56.585 118.290 59.435 ;
        RECT 115.990 56.415 118.290 56.585 ;
        RECT 118.690 56.585 118.860 68.435 ;
        RECT 119.350 67.725 120.350 68.175 ;
        RECT 119.360 57.490 119.530 67.530 ;
        RECT 120.150 57.490 120.320 67.530 ;
        RECT 119.590 57.105 120.090 57.275 ;
        RECT 120.820 56.585 120.990 68.435 ;
        RECT 118.690 56.415 120.990 56.585 ;
        RECT 121.390 68.435 123.690 68.605 ;
        RECT 121.390 56.585 121.560 68.435 ;
        RECT 122.050 67.725 123.050 68.175 ;
        RECT 122.060 57.490 122.230 67.530 ;
        RECT 122.850 57.490 123.020 67.530 ;
        RECT 122.290 57.105 122.790 57.275 ;
        RECT 123.520 56.585 123.690 68.435 ;
        RECT 124.585 68.435 126.885 68.605 ;
        RECT 124.585 67.450 124.755 68.435 ;
        RECT 125.485 67.745 125.985 67.915 ;
        RECT 125.255 67.450 125.425 67.530 ;
        RECT 126.045 67.525 126.215 67.530 ;
        RECT 124.585 66.575 125.425 67.450 ;
        RECT 124.585 65.585 124.755 66.575 ;
        RECT 125.255 66.490 125.425 66.575 ;
        RECT 125.995 66.495 126.470 67.525 ;
        RECT 126.045 66.490 126.215 66.495 ;
        RECT 125.245 65.850 126.220 66.300 ;
        RECT 126.715 65.585 126.885 68.435 ;
        RECT 124.585 65.415 126.885 65.585 ;
        RECT 127.285 68.435 129.585 68.605 ;
        RECT 127.285 65.585 127.455 68.435 ;
        RECT 128.185 67.745 128.685 67.915 ;
        RECT 127.955 67.525 128.125 67.530 ;
        RECT 127.680 66.495 128.175 67.525 ;
        RECT 128.745 67.500 128.915 67.530 ;
        RECT 129.415 67.500 129.585 68.435 ;
        RECT 129.985 68.435 132.285 68.605 ;
        RECT 129.985 67.500 130.155 68.435 ;
        RECT 130.885 67.745 131.385 67.915 ;
        RECT 130.655 67.500 130.825 67.530 ;
        RECT 128.670 66.570 129.590 67.500 ;
        RECT 127.955 66.490 128.125 66.495 ;
        RECT 128.745 66.490 128.915 66.570 ;
        RECT 127.945 65.850 128.920 66.300 ;
        RECT 129.415 65.585 129.585 66.570 ;
        RECT 129.930 66.520 130.825 67.500 ;
        RECT 127.285 65.415 129.585 65.585 ;
        RECT 129.985 65.585 130.155 66.520 ;
        RECT 130.655 66.490 130.825 66.520 ;
        RECT 131.445 66.490 131.615 67.530 ;
        RECT 130.470 66.105 131.385 66.275 ;
        RECT 130.470 65.900 131.305 66.105 ;
        RECT 132.115 65.585 132.285 68.435 ;
        RECT 129.985 65.415 132.285 65.585 ;
        RECT 136.015 68.435 138.315 68.605 ;
        RECT 124.585 64.345 126.885 64.515 ;
        RECT 124.585 61.935 124.755 64.345 ;
        RECT 125.245 63.675 126.220 64.100 ;
        RECT 126.715 64.035 126.885 64.345 ;
        RECT 127.285 64.345 129.585 64.515 ;
        RECT 127.285 64.035 127.455 64.345 ;
        RECT 125.485 63.655 125.985 63.675 ;
        RECT 125.255 63.480 125.425 63.485 ;
        RECT 126.045 63.480 126.215 63.485 ;
        RECT 125.155 62.800 125.525 63.480 ;
        RECT 125.945 62.800 126.315 63.480 ;
        RECT 125.255 62.795 125.425 62.800 ;
        RECT 126.045 62.795 126.215 62.800 ;
        RECT 125.485 62.455 125.985 62.625 ;
        RECT 126.715 62.245 127.455 64.035 ;
        RECT 127.945 63.675 128.920 64.100 ;
        RECT 128.185 63.655 128.685 63.675 ;
        RECT 127.955 63.480 128.125 63.485 ;
        RECT 127.855 62.800 128.225 63.480 ;
        RECT 128.745 63.405 128.915 63.485 ;
        RECT 129.415 63.405 129.585 64.345 ;
        RECT 129.985 64.345 132.285 64.515 ;
        RECT 129.985 63.405 130.155 64.345 ;
        RECT 130.365 63.655 131.405 64.100 ;
        RECT 130.655 63.405 130.825 63.485 ;
        RECT 128.670 62.825 129.590 63.405 ;
        RECT 129.980 62.875 130.825 63.405 ;
        RECT 127.955 62.795 128.125 62.800 ;
        RECT 128.745 62.795 128.915 62.825 ;
        RECT 128.185 62.455 128.685 62.625 ;
        RECT 126.715 61.935 126.885 62.245 ;
        RECT 124.585 61.765 126.885 61.935 ;
        RECT 127.285 61.935 127.455 62.245 ;
        RECT 129.415 61.935 129.585 62.825 ;
        RECT 127.285 61.765 129.585 61.935 ;
        RECT 129.985 61.935 130.155 62.875 ;
        RECT 130.655 62.795 130.825 62.875 ;
        RECT 131.445 62.795 131.615 63.485 ;
        RECT 130.885 62.455 131.385 62.625 ;
        RECT 132.115 61.935 132.285 64.345 ;
        RECT 129.985 61.765 132.285 61.935 ;
        RECT 133.315 59.435 135.615 59.605 ;
        RECT 133.315 58.500 133.485 59.435 ;
        RECT 134.215 58.745 134.715 58.915 ;
        RECT 133.985 58.500 134.155 58.530 ;
        RECT 133.260 57.520 134.155 58.500 ;
        RECT 121.390 56.415 123.690 56.585 ;
        RECT 133.315 56.585 133.485 57.520 ;
        RECT 133.985 57.490 134.155 57.520 ;
        RECT 134.775 57.490 134.945 58.530 ;
        RECT 133.800 57.105 134.715 57.275 ;
        RECT 133.800 56.900 134.635 57.105 ;
        RECT 135.445 56.585 135.615 59.435 ;
        RECT 133.315 56.415 135.615 56.585 ;
        RECT 136.015 56.585 136.185 68.435 ;
        RECT 136.675 67.725 137.675 68.175 ;
        RECT 136.685 57.490 136.855 67.530 ;
        RECT 137.475 57.490 137.645 67.530 ;
        RECT 136.915 57.105 137.415 57.275 ;
        RECT 138.145 56.585 138.315 68.435 ;
        RECT 144.115 68.435 146.415 68.605 ;
        RECT 138.715 59.435 141.015 59.605 ;
        RECT 138.715 58.500 138.885 59.435 ;
        RECT 139.615 58.745 140.115 58.915 ;
        RECT 139.385 58.500 139.555 58.530 ;
        RECT 138.660 57.520 139.555 58.500 ;
        RECT 136.015 56.415 138.315 56.585 ;
        RECT 138.715 56.585 138.885 57.520 ;
        RECT 139.385 57.490 139.555 57.520 ;
        RECT 140.175 57.490 140.345 58.530 ;
        RECT 139.200 57.105 140.115 57.275 ;
        RECT 139.200 56.900 140.035 57.105 ;
        RECT 140.845 56.585 141.015 59.435 ;
        RECT 141.415 59.435 143.715 59.605 ;
        RECT 141.415 58.500 141.585 59.435 ;
        RECT 142.315 58.745 142.815 58.915 ;
        RECT 142.085 58.500 142.255 58.530 ;
        RECT 141.360 57.520 142.255 58.500 ;
        RECT 138.715 56.415 141.015 56.585 ;
        RECT 141.415 56.585 141.585 57.520 ;
        RECT 142.085 57.490 142.255 57.520 ;
        RECT 142.875 57.490 143.045 58.530 ;
        RECT 141.900 57.105 142.815 57.275 ;
        RECT 141.900 56.900 142.735 57.105 ;
        RECT 143.545 56.585 143.715 59.435 ;
        RECT 141.415 56.415 143.715 56.585 ;
        RECT 144.115 56.585 144.285 68.435 ;
        RECT 144.775 67.725 145.775 68.175 ;
        RECT 144.785 57.490 144.955 67.530 ;
        RECT 145.575 57.490 145.745 67.530 ;
        RECT 145.015 57.105 145.515 57.275 ;
        RECT 146.245 56.585 146.415 68.435 ;
        RECT 144.115 56.415 146.415 56.585 ;
        RECT 146.815 68.435 149.115 68.605 ;
        RECT 146.815 56.585 146.985 68.435 ;
        RECT 147.475 67.725 148.475 68.175 ;
        RECT 147.485 57.490 147.655 67.530 ;
        RECT 148.275 57.490 148.445 67.530 ;
        RECT 147.715 57.105 148.215 57.275 ;
        RECT 148.945 56.585 149.115 68.435 ;
        RECT 146.815 56.415 149.115 56.585 ;
        RECT 6.190 55.345 8.490 55.515 ;
        RECT 6.190 54.405 6.360 55.345 ;
        RECT 6.570 54.655 7.610 55.100 ;
        RECT 6.860 54.405 7.030 54.485 ;
        RECT 6.185 53.875 7.030 54.405 ;
        RECT 6.190 52.935 6.360 53.875 ;
        RECT 6.860 53.795 7.030 53.875 ;
        RECT 7.650 53.795 7.820 54.485 ;
        RECT 7.090 53.455 7.590 53.625 ;
        RECT 8.320 52.935 8.490 55.345 ;
        RECT 6.190 52.765 8.490 52.935 ;
        RECT 8.890 55.345 11.190 55.515 ;
        RECT 8.890 47.085 9.060 55.345 ;
        RECT 9.790 54.655 10.290 54.825 ;
        RECT 9.560 47.945 9.730 54.485 ;
        RECT 10.350 47.945 10.520 54.485 ;
        RECT 9.550 47.375 10.550 47.775 ;
        RECT 11.020 47.085 11.190 55.345 ;
        RECT 11.590 55.345 13.890 55.515 ;
        RECT 11.590 54.405 11.760 55.345 ;
        RECT 11.970 54.655 13.010 55.100 ;
        RECT 12.260 54.405 12.430 54.485 ;
        RECT 11.585 53.875 12.430 54.405 ;
        RECT 11.590 52.935 11.760 53.875 ;
        RECT 12.260 53.795 12.430 53.875 ;
        RECT 13.050 53.795 13.220 54.485 ;
        RECT 12.490 53.455 12.990 53.625 ;
        RECT 13.720 52.935 13.890 55.345 ;
        RECT 14.290 55.345 16.590 55.515 ;
        RECT 14.290 54.405 14.460 55.345 ;
        RECT 14.670 54.655 15.710 55.100 ;
        RECT 14.960 54.405 15.130 54.485 ;
        RECT 14.285 53.875 15.130 54.405 ;
        RECT 11.590 52.765 13.890 52.935 ;
        RECT 14.290 52.935 14.460 53.875 ;
        RECT 14.960 53.795 15.130 53.875 ;
        RECT 15.750 53.795 15.920 54.485 ;
        RECT 15.190 53.455 15.690 53.625 ;
        RECT 16.420 52.935 16.590 55.345 ;
        RECT 14.290 52.765 16.590 52.935 ;
        RECT 16.990 55.345 19.290 55.515 ;
        RECT 8.890 46.915 11.190 47.085 ;
        RECT 16.990 47.085 17.160 55.345 ;
        RECT 17.890 54.655 18.390 54.825 ;
        RECT 17.660 47.945 17.830 54.485 ;
        RECT 18.450 47.945 18.620 54.485 ;
        RECT 17.650 47.375 18.650 47.775 ;
        RECT 19.120 47.085 19.290 55.345 ;
        RECT 16.990 46.915 19.290 47.085 ;
        RECT 19.690 55.345 21.990 55.515 ;
        RECT 19.690 47.085 19.860 55.345 ;
        RECT 20.590 54.655 21.090 54.825 ;
        RECT 20.360 47.945 20.530 54.485 ;
        RECT 21.150 47.945 21.320 54.485 ;
        RECT 20.350 47.375 21.350 47.775 ;
        RECT 21.820 47.085 21.990 55.345 ;
        RECT 31.615 55.345 33.915 55.515 ;
        RECT 31.615 54.405 31.785 55.345 ;
        RECT 31.995 54.655 33.035 55.100 ;
        RECT 32.285 54.405 32.455 54.485 ;
        RECT 31.610 53.875 32.455 54.405 ;
        RECT 31.615 52.935 31.785 53.875 ;
        RECT 32.285 53.795 32.455 53.875 ;
        RECT 33.075 53.795 33.245 54.485 ;
        RECT 32.515 53.455 33.015 53.625 ;
        RECT 33.745 52.935 33.915 55.345 ;
        RECT 31.615 52.765 33.915 52.935 ;
        RECT 34.315 55.345 36.615 55.515 ;
        RECT 19.690 46.915 21.990 47.085 ;
        RECT 34.315 47.085 34.485 55.345 ;
        RECT 35.215 54.655 35.715 54.825 ;
        RECT 34.985 47.945 35.155 54.485 ;
        RECT 35.775 47.945 35.945 54.485 ;
        RECT 34.975 47.375 35.975 47.775 ;
        RECT 36.445 47.085 36.615 55.345 ;
        RECT 37.015 55.345 39.315 55.515 ;
        RECT 37.015 54.405 37.185 55.345 ;
        RECT 37.395 54.655 38.435 55.100 ;
        RECT 37.685 54.405 37.855 54.485 ;
        RECT 37.010 53.875 37.855 54.405 ;
        RECT 37.015 52.935 37.185 53.875 ;
        RECT 37.685 53.795 37.855 53.875 ;
        RECT 38.475 53.795 38.645 54.485 ;
        RECT 37.915 53.455 38.415 53.625 ;
        RECT 39.145 52.935 39.315 55.345 ;
        RECT 39.715 55.345 42.015 55.515 ;
        RECT 39.715 54.405 39.885 55.345 ;
        RECT 40.095 54.655 41.135 55.100 ;
        RECT 40.385 54.405 40.555 54.485 ;
        RECT 39.710 53.875 40.555 54.405 ;
        RECT 37.015 52.765 39.315 52.935 ;
        RECT 39.715 52.935 39.885 53.875 ;
        RECT 40.385 53.795 40.555 53.875 ;
        RECT 41.175 53.795 41.345 54.485 ;
        RECT 40.615 53.455 41.115 53.625 ;
        RECT 41.845 52.935 42.015 55.345 ;
        RECT 39.715 52.765 42.015 52.935 ;
        RECT 42.415 55.345 44.715 55.515 ;
        RECT 34.315 46.915 36.615 47.085 ;
        RECT 42.415 47.085 42.585 55.345 ;
        RECT 43.315 54.655 43.815 54.825 ;
        RECT 43.085 47.945 43.255 54.485 ;
        RECT 43.875 47.945 44.045 54.485 ;
        RECT 43.075 47.375 44.075 47.775 ;
        RECT 44.545 47.085 44.715 55.345 ;
        RECT 42.415 46.915 44.715 47.085 ;
        RECT 45.115 55.345 47.415 55.515 ;
        RECT 45.115 47.085 45.285 55.345 ;
        RECT 46.015 54.655 46.515 54.825 ;
        RECT 45.785 47.945 45.955 54.485 ;
        RECT 46.575 47.945 46.745 54.485 ;
        RECT 45.775 47.375 46.775 47.775 ;
        RECT 47.245 47.085 47.415 55.345 ;
        RECT 57.040 55.345 59.340 55.515 ;
        RECT 57.040 54.405 57.210 55.345 ;
        RECT 57.420 54.655 58.460 55.100 ;
        RECT 57.710 54.405 57.880 54.485 ;
        RECT 57.035 53.875 57.880 54.405 ;
        RECT 57.040 52.935 57.210 53.875 ;
        RECT 57.710 53.795 57.880 53.875 ;
        RECT 58.500 53.795 58.670 54.485 ;
        RECT 57.940 53.455 58.440 53.625 ;
        RECT 59.170 52.935 59.340 55.345 ;
        RECT 57.040 52.765 59.340 52.935 ;
        RECT 59.740 55.345 62.040 55.515 ;
        RECT 45.115 46.915 47.415 47.085 ;
        RECT 59.740 47.085 59.910 55.345 ;
        RECT 60.640 54.655 61.140 54.825 ;
        RECT 60.410 47.945 60.580 54.485 ;
        RECT 61.200 47.945 61.370 54.485 ;
        RECT 60.400 47.375 61.400 47.775 ;
        RECT 61.870 47.085 62.040 55.345 ;
        RECT 62.440 55.345 64.740 55.515 ;
        RECT 62.440 54.405 62.610 55.345 ;
        RECT 62.820 54.655 63.860 55.100 ;
        RECT 63.110 54.405 63.280 54.485 ;
        RECT 62.435 53.875 63.280 54.405 ;
        RECT 62.440 52.935 62.610 53.875 ;
        RECT 63.110 53.795 63.280 53.875 ;
        RECT 63.900 53.795 64.070 54.485 ;
        RECT 63.340 53.455 63.840 53.625 ;
        RECT 64.570 52.935 64.740 55.345 ;
        RECT 65.140 55.345 67.440 55.515 ;
        RECT 65.140 54.405 65.310 55.345 ;
        RECT 65.520 54.655 66.560 55.100 ;
        RECT 65.810 54.405 65.980 54.485 ;
        RECT 65.135 53.875 65.980 54.405 ;
        RECT 62.440 52.765 64.740 52.935 ;
        RECT 65.140 52.935 65.310 53.875 ;
        RECT 65.810 53.795 65.980 53.875 ;
        RECT 66.600 53.795 66.770 54.485 ;
        RECT 66.040 53.455 66.540 53.625 ;
        RECT 67.270 52.935 67.440 55.345 ;
        RECT 65.140 52.765 67.440 52.935 ;
        RECT 67.840 55.345 70.140 55.515 ;
        RECT 59.740 46.915 62.040 47.085 ;
        RECT 67.840 47.085 68.010 55.345 ;
        RECT 68.740 54.655 69.240 54.825 ;
        RECT 68.510 47.945 68.680 54.485 ;
        RECT 69.300 47.945 69.470 54.485 ;
        RECT 68.500 47.375 69.500 47.775 ;
        RECT 69.970 47.085 70.140 55.345 ;
        RECT 67.840 46.915 70.140 47.085 ;
        RECT 70.540 55.345 72.840 55.515 ;
        RECT 70.540 47.085 70.710 55.345 ;
        RECT 71.440 54.655 71.940 54.825 ;
        RECT 71.210 47.945 71.380 54.485 ;
        RECT 72.000 47.945 72.170 54.485 ;
        RECT 71.200 47.375 72.200 47.775 ;
        RECT 72.670 47.085 72.840 55.345 ;
        RECT 82.465 55.345 84.765 55.515 ;
        RECT 82.465 54.405 82.635 55.345 ;
        RECT 82.845 54.655 83.885 55.100 ;
        RECT 83.135 54.405 83.305 54.485 ;
        RECT 82.460 53.875 83.305 54.405 ;
        RECT 82.465 52.935 82.635 53.875 ;
        RECT 83.135 53.795 83.305 53.875 ;
        RECT 83.925 53.795 84.095 54.485 ;
        RECT 83.365 53.455 83.865 53.625 ;
        RECT 84.595 52.935 84.765 55.345 ;
        RECT 82.465 52.765 84.765 52.935 ;
        RECT 85.165 55.345 87.465 55.515 ;
        RECT 70.540 46.915 72.840 47.085 ;
        RECT 85.165 47.085 85.335 55.345 ;
        RECT 86.065 54.655 86.565 54.825 ;
        RECT 85.835 47.945 86.005 54.485 ;
        RECT 86.625 47.945 86.795 54.485 ;
        RECT 85.825 47.375 86.825 47.775 ;
        RECT 87.295 47.085 87.465 55.345 ;
        RECT 87.865 55.345 90.165 55.515 ;
        RECT 87.865 54.405 88.035 55.345 ;
        RECT 88.245 54.655 89.285 55.100 ;
        RECT 88.535 54.405 88.705 54.485 ;
        RECT 87.860 53.875 88.705 54.405 ;
        RECT 87.865 52.935 88.035 53.875 ;
        RECT 88.535 53.795 88.705 53.875 ;
        RECT 89.325 53.795 89.495 54.485 ;
        RECT 88.765 53.455 89.265 53.625 ;
        RECT 89.995 52.935 90.165 55.345 ;
        RECT 90.565 55.345 92.865 55.515 ;
        RECT 90.565 54.405 90.735 55.345 ;
        RECT 90.945 54.655 91.985 55.100 ;
        RECT 91.235 54.405 91.405 54.485 ;
        RECT 90.560 53.875 91.405 54.405 ;
        RECT 87.865 52.765 90.165 52.935 ;
        RECT 90.565 52.935 90.735 53.875 ;
        RECT 91.235 53.795 91.405 53.875 ;
        RECT 92.025 53.795 92.195 54.485 ;
        RECT 91.465 53.455 91.965 53.625 ;
        RECT 92.695 52.935 92.865 55.345 ;
        RECT 90.565 52.765 92.865 52.935 ;
        RECT 93.265 55.345 95.565 55.515 ;
        RECT 85.165 46.915 87.465 47.085 ;
        RECT 93.265 47.085 93.435 55.345 ;
        RECT 94.165 54.655 94.665 54.825 ;
        RECT 93.935 47.945 94.105 54.485 ;
        RECT 94.725 47.945 94.895 54.485 ;
        RECT 93.925 47.375 94.925 47.775 ;
        RECT 95.395 47.085 95.565 55.345 ;
        RECT 93.265 46.915 95.565 47.085 ;
        RECT 95.965 55.345 98.265 55.515 ;
        RECT 95.965 47.085 96.135 55.345 ;
        RECT 96.865 54.655 97.365 54.825 ;
        RECT 96.635 47.945 96.805 54.485 ;
        RECT 97.425 47.945 97.595 54.485 ;
        RECT 96.625 47.375 97.625 47.775 ;
        RECT 98.095 47.085 98.265 55.345 ;
        RECT 107.890 55.345 110.190 55.515 ;
        RECT 107.890 54.405 108.060 55.345 ;
        RECT 108.270 54.655 109.310 55.100 ;
        RECT 108.560 54.405 108.730 54.485 ;
        RECT 107.885 53.875 108.730 54.405 ;
        RECT 107.890 52.935 108.060 53.875 ;
        RECT 108.560 53.795 108.730 53.875 ;
        RECT 109.350 53.795 109.520 54.485 ;
        RECT 108.790 53.455 109.290 53.625 ;
        RECT 110.020 52.935 110.190 55.345 ;
        RECT 107.890 52.765 110.190 52.935 ;
        RECT 110.590 55.345 112.890 55.515 ;
        RECT 95.965 46.915 98.265 47.085 ;
        RECT 110.590 47.085 110.760 55.345 ;
        RECT 111.490 54.655 111.990 54.825 ;
        RECT 111.260 47.945 111.430 54.485 ;
        RECT 112.050 47.945 112.220 54.485 ;
        RECT 111.250 47.375 112.250 47.775 ;
        RECT 112.720 47.085 112.890 55.345 ;
        RECT 113.290 55.345 115.590 55.515 ;
        RECT 113.290 54.405 113.460 55.345 ;
        RECT 113.670 54.655 114.710 55.100 ;
        RECT 113.960 54.405 114.130 54.485 ;
        RECT 113.285 53.875 114.130 54.405 ;
        RECT 113.290 52.935 113.460 53.875 ;
        RECT 113.960 53.795 114.130 53.875 ;
        RECT 114.750 53.795 114.920 54.485 ;
        RECT 114.190 53.455 114.690 53.625 ;
        RECT 115.420 52.935 115.590 55.345 ;
        RECT 115.990 55.345 118.290 55.515 ;
        RECT 115.990 54.405 116.160 55.345 ;
        RECT 116.370 54.655 117.410 55.100 ;
        RECT 116.660 54.405 116.830 54.485 ;
        RECT 115.985 53.875 116.830 54.405 ;
        RECT 113.290 52.765 115.590 52.935 ;
        RECT 115.990 52.935 116.160 53.875 ;
        RECT 116.660 53.795 116.830 53.875 ;
        RECT 117.450 53.795 117.620 54.485 ;
        RECT 116.890 53.455 117.390 53.625 ;
        RECT 118.120 52.935 118.290 55.345 ;
        RECT 115.990 52.765 118.290 52.935 ;
        RECT 118.690 55.345 120.990 55.515 ;
        RECT 110.590 46.915 112.890 47.085 ;
        RECT 118.690 47.085 118.860 55.345 ;
        RECT 119.590 54.655 120.090 54.825 ;
        RECT 119.360 47.945 119.530 54.485 ;
        RECT 120.150 47.945 120.320 54.485 ;
        RECT 119.350 47.375 120.350 47.775 ;
        RECT 120.820 47.085 120.990 55.345 ;
        RECT 118.690 46.915 120.990 47.085 ;
        RECT 121.390 55.345 123.690 55.515 ;
        RECT 121.390 47.085 121.560 55.345 ;
        RECT 122.290 54.655 122.790 54.825 ;
        RECT 122.060 47.945 122.230 54.485 ;
        RECT 122.850 47.945 123.020 54.485 ;
        RECT 122.050 47.375 123.050 47.775 ;
        RECT 123.520 47.085 123.690 55.345 ;
        RECT 133.315 55.345 135.615 55.515 ;
        RECT 133.315 54.405 133.485 55.345 ;
        RECT 133.695 54.655 134.735 55.100 ;
        RECT 133.985 54.405 134.155 54.485 ;
        RECT 133.310 53.875 134.155 54.405 ;
        RECT 133.315 52.935 133.485 53.875 ;
        RECT 133.985 53.795 134.155 53.875 ;
        RECT 134.775 53.795 134.945 54.485 ;
        RECT 134.215 53.455 134.715 53.625 ;
        RECT 135.445 52.935 135.615 55.345 ;
        RECT 133.315 52.765 135.615 52.935 ;
        RECT 136.015 55.345 138.315 55.515 ;
        RECT 121.390 46.915 123.690 47.085 ;
        RECT 136.015 47.085 136.185 55.345 ;
        RECT 136.915 54.655 137.415 54.825 ;
        RECT 136.685 47.945 136.855 54.485 ;
        RECT 137.475 47.945 137.645 54.485 ;
        RECT 136.675 47.375 137.675 47.775 ;
        RECT 138.145 47.085 138.315 55.345 ;
        RECT 138.715 55.345 141.015 55.515 ;
        RECT 138.715 54.405 138.885 55.345 ;
        RECT 139.095 54.655 140.135 55.100 ;
        RECT 139.385 54.405 139.555 54.485 ;
        RECT 138.710 53.875 139.555 54.405 ;
        RECT 138.715 52.935 138.885 53.875 ;
        RECT 139.385 53.795 139.555 53.875 ;
        RECT 140.175 53.795 140.345 54.485 ;
        RECT 139.615 53.455 140.115 53.625 ;
        RECT 140.845 52.935 141.015 55.345 ;
        RECT 141.415 55.345 143.715 55.515 ;
        RECT 141.415 54.405 141.585 55.345 ;
        RECT 141.795 54.655 142.835 55.100 ;
        RECT 142.085 54.405 142.255 54.485 ;
        RECT 141.410 53.875 142.255 54.405 ;
        RECT 138.715 52.765 141.015 52.935 ;
        RECT 141.415 52.935 141.585 53.875 ;
        RECT 142.085 53.795 142.255 53.875 ;
        RECT 142.875 53.795 143.045 54.485 ;
        RECT 142.315 53.455 142.815 53.625 ;
        RECT 143.545 52.935 143.715 55.345 ;
        RECT 141.415 52.765 143.715 52.935 ;
        RECT 144.115 55.345 146.415 55.515 ;
        RECT 136.015 46.915 138.315 47.085 ;
        RECT 144.115 47.085 144.285 55.345 ;
        RECT 145.015 54.655 145.515 54.825 ;
        RECT 144.785 47.945 144.955 54.485 ;
        RECT 145.575 47.945 145.745 54.485 ;
        RECT 144.775 47.375 145.775 47.775 ;
        RECT 146.245 47.085 146.415 55.345 ;
        RECT 144.115 46.915 146.415 47.085 ;
        RECT 146.815 55.345 149.115 55.515 ;
        RECT 146.815 47.085 146.985 55.345 ;
        RECT 147.715 54.655 148.215 54.825 ;
        RECT 147.485 47.945 147.655 54.485 ;
        RECT 148.275 47.945 148.445 54.485 ;
        RECT 147.475 47.375 148.475 47.775 ;
        RECT 148.945 47.085 149.115 55.345 ;
        RECT 146.815 46.915 149.115 47.085 ;
        RECT 8.890 45.860 11.190 46.030 ;
        RECT 6.190 36.860 8.490 37.030 ;
        RECT 6.190 35.925 6.360 36.860 ;
        RECT 7.090 36.170 7.590 36.340 ;
        RECT 6.860 35.925 7.030 35.955 ;
        RECT 6.135 34.945 7.030 35.925 ;
        RECT 6.190 34.010 6.360 34.945 ;
        RECT 6.860 34.915 7.030 34.945 ;
        RECT 7.650 34.915 7.820 35.955 ;
        RECT 6.675 34.530 7.590 34.700 ;
        RECT 6.675 34.325 7.510 34.530 ;
        RECT 8.320 34.010 8.490 36.860 ;
        RECT 6.190 33.840 8.490 34.010 ;
        RECT 8.890 34.010 9.060 45.860 ;
        RECT 9.550 45.150 10.550 45.600 ;
        RECT 9.560 34.915 9.730 44.955 ;
        RECT 10.350 34.915 10.520 44.955 ;
        RECT 9.790 34.530 10.290 34.700 ;
        RECT 11.020 34.010 11.190 45.860 ;
        RECT 16.990 45.860 19.290 46.030 ;
        RECT 11.590 36.860 13.890 37.030 ;
        RECT 11.590 35.925 11.760 36.860 ;
        RECT 12.490 36.170 12.990 36.340 ;
        RECT 12.260 35.925 12.430 35.955 ;
        RECT 11.535 34.945 12.430 35.925 ;
        RECT 8.890 33.840 11.190 34.010 ;
        RECT 11.590 34.010 11.760 34.945 ;
        RECT 12.260 34.915 12.430 34.945 ;
        RECT 13.050 34.915 13.220 35.955 ;
        RECT 12.075 34.530 12.990 34.700 ;
        RECT 12.075 34.325 12.910 34.530 ;
        RECT 13.720 34.010 13.890 36.860 ;
        RECT 14.290 36.860 16.590 37.030 ;
        RECT 14.290 35.925 14.460 36.860 ;
        RECT 15.190 36.170 15.690 36.340 ;
        RECT 14.960 35.925 15.130 35.955 ;
        RECT 14.235 34.945 15.130 35.925 ;
        RECT 11.590 33.840 13.890 34.010 ;
        RECT 14.290 34.010 14.460 34.945 ;
        RECT 14.960 34.915 15.130 34.945 ;
        RECT 15.750 34.915 15.920 35.955 ;
        RECT 14.775 34.530 15.690 34.700 ;
        RECT 14.775 34.325 15.610 34.530 ;
        RECT 16.420 34.010 16.590 36.860 ;
        RECT 14.290 33.840 16.590 34.010 ;
        RECT 16.990 34.010 17.160 45.860 ;
        RECT 17.650 45.150 18.650 45.600 ;
        RECT 17.660 34.915 17.830 44.955 ;
        RECT 18.450 34.915 18.620 44.955 ;
        RECT 17.890 34.530 18.390 34.700 ;
        RECT 19.120 34.010 19.290 45.860 ;
        RECT 16.990 33.840 19.290 34.010 ;
        RECT 19.690 45.860 21.990 46.030 ;
        RECT 19.690 34.010 19.860 45.860 ;
        RECT 20.350 45.150 21.350 45.600 ;
        RECT 20.360 34.915 20.530 44.955 ;
        RECT 21.150 34.915 21.320 44.955 ;
        RECT 20.590 34.530 21.090 34.700 ;
        RECT 21.820 34.010 21.990 45.860 ;
        RECT 34.315 45.860 36.615 46.030 ;
        RECT 31.615 36.860 33.915 37.030 ;
        RECT 31.615 35.925 31.785 36.860 ;
        RECT 32.515 36.170 33.015 36.340 ;
        RECT 32.285 35.925 32.455 35.955 ;
        RECT 31.560 34.945 32.455 35.925 ;
        RECT 19.690 33.840 21.990 34.010 ;
        RECT 31.615 34.010 31.785 34.945 ;
        RECT 32.285 34.915 32.455 34.945 ;
        RECT 33.075 34.915 33.245 35.955 ;
        RECT 32.100 34.530 33.015 34.700 ;
        RECT 32.100 34.325 32.935 34.530 ;
        RECT 33.745 34.010 33.915 36.860 ;
        RECT 31.615 33.840 33.915 34.010 ;
        RECT 34.315 34.010 34.485 45.860 ;
        RECT 34.975 45.150 35.975 45.600 ;
        RECT 34.985 34.915 35.155 44.955 ;
        RECT 35.775 34.915 35.945 44.955 ;
        RECT 35.215 34.530 35.715 34.700 ;
        RECT 36.445 34.010 36.615 45.860 ;
        RECT 42.415 45.860 44.715 46.030 ;
        RECT 37.015 36.860 39.315 37.030 ;
        RECT 37.015 35.925 37.185 36.860 ;
        RECT 37.915 36.170 38.415 36.340 ;
        RECT 37.685 35.925 37.855 35.955 ;
        RECT 36.960 34.945 37.855 35.925 ;
        RECT 34.315 33.840 36.615 34.010 ;
        RECT 37.015 34.010 37.185 34.945 ;
        RECT 37.685 34.915 37.855 34.945 ;
        RECT 38.475 34.915 38.645 35.955 ;
        RECT 37.500 34.530 38.415 34.700 ;
        RECT 37.500 34.325 38.335 34.530 ;
        RECT 39.145 34.010 39.315 36.860 ;
        RECT 39.715 36.860 42.015 37.030 ;
        RECT 39.715 35.925 39.885 36.860 ;
        RECT 40.615 36.170 41.115 36.340 ;
        RECT 40.385 35.925 40.555 35.955 ;
        RECT 39.660 34.945 40.555 35.925 ;
        RECT 37.015 33.840 39.315 34.010 ;
        RECT 39.715 34.010 39.885 34.945 ;
        RECT 40.385 34.915 40.555 34.945 ;
        RECT 41.175 34.915 41.345 35.955 ;
        RECT 40.200 34.530 41.115 34.700 ;
        RECT 40.200 34.325 41.035 34.530 ;
        RECT 41.845 34.010 42.015 36.860 ;
        RECT 39.715 33.840 42.015 34.010 ;
        RECT 42.415 34.010 42.585 45.860 ;
        RECT 43.075 45.150 44.075 45.600 ;
        RECT 43.085 34.915 43.255 44.955 ;
        RECT 43.875 34.915 44.045 44.955 ;
        RECT 43.315 34.530 43.815 34.700 ;
        RECT 44.545 34.010 44.715 45.860 ;
        RECT 42.415 33.840 44.715 34.010 ;
        RECT 45.115 45.860 47.415 46.030 ;
        RECT 45.115 34.010 45.285 45.860 ;
        RECT 45.775 45.150 46.775 45.600 ;
        RECT 45.785 34.915 45.955 44.955 ;
        RECT 46.575 34.915 46.745 44.955 ;
        RECT 46.015 34.530 46.515 34.700 ;
        RECT 47.245 34.010 47.415 45.860 ;
        RECT 59.740 45.860 62.040 46.030 ;
        RECT 57.040 36.860 59.340 37.030 ;
        RECT 57.040 35.925 57.210 36.860 ;
        RECT 57.940 36.170 58.440 36.340 ;
        RECT 57.710 35.925 57.880 35.955 ;
        RECT 56.985 34.945 57.880 35.925 ;
        RECT 45.115 33.840 47.415 34.010 ;
        RECT 57.040 34.010 57.210 34.945 ;
        RECT 57.710 34.915 57.880 34.945 ;
        RECT 58.500 34.915 58.670 35.955 ;
        RECT 57.525 34.530 58.440 34.700 ;
        RECT 57.525 34.325 58.360 34.530 ;
        RECT 59.170 34.010 59.340 36.860 ;
        RECT 57.040 33.840 59.340 34.010 ;
        RECT 59.740 34.010 59.910 45.860 ;
        RECT 60.400 45.150 61.400 45.600 ;
        RECT 60.410 34.915 60.580 44.955 ;
        RECT 61.200 34.915 61.370 44.955 ;
        RECT 60.640 34.530 61.140 34.700 ;
        RECT 61.870 34.010 62.040 45.860 ;
        RECT 67.840 45.860 70.140 46.030 ;
        RECT 62.440 36.860 64.740 37.030 ;
        RECT 62.440 35.925 62.610 36.860 ;
        RECT 63.340 36.170 63.840 36.340 ;
        RECT 63.110 35.925 63.280 35.955 ;
        RECT 62.385 34.945 63.280 35.925 ;
        RECT 59.740 33.840 62.040 34.010 ;
        RECT 62.440 34.010 62.610 34.945 ;
        RECT 63.110 34.915 63.280 34.945 ;
        RECT 63.900 34.915 64.070 35.955 ;
        RECT 62.925 34.530 63.840 34.700 ;
        RECT 62.925 34.325 63.760 34.530 ;
        RECT 64.570 34.010 64.740 36.860 ;
        RECT 65.140 36.860 67.440 37.030 ;
        RECT 65.140 35.925 65.310 36.860 ;
        RECT 66.040 36.170 66.540 36.340 ;
        RECT 65.810 35.925 65.980 35.955 ;
        RECT 65.085 34.945 65.980 35.925 ;
        RECT 62.440 33.840 64.740 34.010 ;
        RECT 65.140 34.010 65.310 34.945 ;
        RECT 65.810 34.915 65.980 34.945 ;
        RECT 66.600 34.915 66.770 35.955 ;
        RECT 65.625 34.530 66.540 34.700 ;
        RECT 65.625 34.325 66.460 34.530 ;
        RECT 67.270 34.010 67.440 36.860 ;
        RECT 65.140 33.840 67.440 34.010 ;
        RECT 67.840 34.010 68.010 45.860 ;
        RECT 68.500 45.150 69.500 45.600 ;
        RECT 68.510 34.915 68.680 44.955 ;
        RECT 69.300 34.915 69.470 44.955 ;
        RECT 68.740 34.530 69.240 34.700 ;
        RECT 69.970 34.010 70.140 45.860 ;
        RECT 67.840 33.840 70.140 34.010 ;
        RECT 70.540 45.860 72.840 46.030 ;
        RECT 70.540 34.010 70.710 45.860 ;
        RECT 71.200 45.150 72.200 45.600 ;
        RECT 71.210 34.915 71.380 44.955 ;
        RECT 72.000 34.915 72.170 44.955 ;
        RECT 71.440 34.530 71.940 34.700 ;
        RECT 72.670 34.010 72.840 45.860 ;
        RECT 85.165 45.860 87.465 46.030 ;
        RECT 82.465 36.860 84.765 37.030 ;
        RECT 82.465 35.925 82.635 36.860 ;
        RECT 83.365 36.170 83.865 36.340 ;
        RECT 83.135 35.925 83.305 35.955 ;
        RECT 82.410 34.945 83.305 35.925 ;
        RECT 70.540 33.840 72.840 34.010 ;
        RECT 82.465 34.010 82.635 34.945 ;
        RECT 83.135 34.915 83.305 34.945 ;
        RECT 83.925 34.915 84.095 35.955 ;
        RECT 82.950 34.530 83.865 34.700 ;
        RECT 82.950 34.325 83.785 34.530 ;
        RECT 84.595 34.010 84.765 36.860 ;
        RECT 82.465 33.840 84.765 34.010 ;
        RECT 85.165 34.010 85.335 45.860 ;
        RECT 85.825 45.150 86.825 45.600 ;
        RECT 85.835 34.915 86.005 44.955 ;
        RECT 86.625 34.915 86.795 44.955 ;
        RECT 86.065 34.530 86.565 34.700 ;
        RECT 87.295 34.010 87.465 45.860 ;
        RECT 93.265 45.860 95.565 46.030 ;
        RECT 87.865 36.860 90.165 37.030 ;
        RECT 87.865 35.925 88.035 36.860 ;
        RECT 88.765 36.170 89.265 36.340 ;
        RECT 88.535 35.925 88.705 35.955 ;
        RECT 87.810 34.945 88.705 35.925 ;
        RECT 85.165 33.840 87.465 34.010 ;
        RECT 87.865 34.010 88.035 34.945 ;
        RECT 88.535 34.915 88.705 34.945 ;
        RECT 89.325 34.915 89.495 35.955 ;
        RECT 88.350 34.530 89.265 34.700 ;
        RECT 88.350 34.325 89.185 34.530 ;
        RECT 89.995 34.010 90.165 36.860 ;
        RECT 90.565 36.860 92.865 37.030 ;
        RECT 90.565 35.925 90.735 36.860 ;
        RECT 91.465 36.170 91.965 36.340 ;
        RECT 91.235 35.925 91.405 35.955 ;
        RECT 90.510 34.945 91.405 35.925 ;
        RECT 87.865 33.840 90.165 34.010 ;
        RECT 90.565 34.010 90.735 34.945 ;
        RECT 91.235 34.915 91.405 34.945 ;
        RECT 92.025 34.915 92.195 35.955 ;
        RECT 91.050 34.530 91.965 34.700 ;
        RECT 91.050 34.325 91.885 34.530 ;
        RECT 92.695 34.010 92.865 36.860 ;
        RECT 90.565 33.840 92.865 34.010 ;
        RECT 93.265 34.010 93.435 45.860 ;
        RECT 93.925 45.150 94.925 45.600 ;
        RECT 93.935 34.915 94.105 44.955 ;
        RECT 94.725 34.915 94.895 44.955 ;
        RECT 94.165 34.530 94.665 34.700 ;
        RECT 95.395 34.010 95.565 45.860 ;
        RECT 93.265 33.840 95.565 34.010 ;
        RECT 95.965 45.860 98.265 46.030 ;
        RECT 95.965 34.010 96.135 45.860 ;
        RECT 96.625 45.150 97.625 45.600 ;
        RECT 96.635 34.915 96.805 44.955 ;
        RECT 97.425 34.915 97.595 44.955 ;
        RECT 96.865 34.530 97.365 34.700 ;
        RECT 98.095 34.010 98.265 45.860 ;
        RECT 110.590 45.860 112.890 46.030 ;
        RECT 107.890 36.860 110.190 37.030 ;
        RECT 107.890 35.925 108.060 36.860 ;
        RECT 108.790 36.170 109.290 36.340 ;
        RECT 108.560 35.925 108.730 35.955 ;
        RECT 107.835 34.945 108.730 35.925 ;
        RECT 95.965 33.840 98.265 34.010 ;
        RECT 107.890 34.010 108.060 34.945 ;
        RECT 108.560 34.915 108.730 34.945 ;
        RECT 109.350 34.915 109.520 35.955 ;
        RECT 108.375 34.530 109.290 34.700 ;
        RECT 108.375 34.325 109.210 34.530 ;
        RECT 110.020 34.010 110.190 36.860 ;
        RECT 107.890 33.840 110.190 34.010 ;
        RECT 110.590 34.010 110.760 45.860 ;
        RECT 111.250 45.150 112.250 45.600 ;
        RECT 111.260 34.915 111.430 44.955 ;
        RECT 112.050 34.915 112.220 44.955 ;
        RECT 111.490 34.530 111.990 34.700 ;
        RECT 112.720 34.010 112.890 45.860 ;
        RECT 118.690 45.860 120.990 46.030 ;
        RECT 113.290 36.860 115.590 37.030 ;
        RECT 113.290 35.925 113.460 36.860 ;
        RECT 114.190 36.170 114.690 36.340 ;
        RECT 113.960 35.925 114.130 35.955 ;
        RECT 113.235 34.945 114.130 35.925 ;
        RECT 110.590 33.840 112.890 34.010 ;
        RECT 113.290 34.010 113.460 34.945 ;
        RECT 113.960 34.915 114.130 34.945 ;
        RECT 114.750 34.915 114.920 35.955 ;
        RECT 113.775 34.530 114.690 34.700 ;
        RECT 113.775 34.325 114.610 34.530 ;
        RECT 115.420 34.010 115.590 36.860 ;
        RECT 115.990 36.860 118.290 37.030 ;
        RECT 115.990 35.925 116.160 36.860 ;
        RECT 116.890 36.170 117.390 36.340 ;
        RECT 116.660 35.925 116.830 35.955 ;
        RECT 115.935 34.945 116.830 35.925 ;
        RECT 113.290 33.840 115.590 34.010 ;
        RECT 115.990 34.010 116.160 34.945 ;
        RECT 116.660 34.915 116.830 34.945 ;
        RECT 117.450 34.915 117.620 35.955 ;
        RECT 116.475 34.530 117.390 34.700 ;
        RECT 116.475 34.325 117.310 34.530 ;
        RECT 118.120 34.010 118.290 36.860 ;
        RECT 115.990 33.840 118.290 34.010 ;
        RECT 118.690 34.010 118.860 45.860 ;
        RECT 119.350 45.150 120.350 45.600 ;
        RECT 119.360 34.915 119.530 44.955 ;
        RECT 120.150 34.915 120.320 44.955 ;
        RECT 119.590 34.530 120.090 34.700 ;
        RECT 120.820 34.010 120.990 45.860 ;
        RECT 118.690 33.840 120.990 34.010 ;
        RECT 121.390 45.860 123.690 46.030 ;
        RECT 121.390 34.010 121.560 45.860 ;
        RECT 122.050 45.150 123.050 45.600 ;
        RECT 122.060 34.915 122.230 44.955 ;
        RECT 122.850 34.915 123.020 44.955 ;
        RECT 122.290 34.530 122.790 34.700 ;
        RECT 123.520 34.010 123.690 45.860 ;
        RECT 136.015 45.860 138.315 46.030 ;
        RECT 133.315 36.860 135.615 37.030 ;
        RECT 133.315 35.925 133.485 36.860 ;
        RECT 134.215 36.170 134.715 36.340 ;
        RECT 133.985 35.925 134.155 35.955 ;
        RECT 133.260 34.945 134.155 35.925 ;
        RECT 121.390 33.840 123.690 34.010 ;
        RECT 133.315 34.010 133.485 34.945 ;
        RECT 133.985 34.915 134.155 34.945 ;
        RECT 134.775 34.915 134.945 35.955 ;
        RECT 133.800 34.530 134.715 34.700 ;
        RECT 133.800 34.325 134.635 34.530 ;
        RECT 135.445 34.010 135.615 36.860 ;
        RECT 133.315 33.840 135.615 34.010 ;
        RECT 136.015 34.010 136.185 45.860 ;
        RECT 136.675 45.150 137.675 45.600 ;
        RECT 136.685 34.915 136.855 44.955 ;
        RECT 137.475 34.915 137.645 44.955 ;
        RECT 136.915 34.530 137.415 34.700 ;
        RECT 138.145 34.010 138.315 45.860 ;
        RECT 144.115 45.860 146.415 46.030 ;
        RECT 138.715 36.860 141.015 37.030 ;
        RECT 138.715 35.925 138.885 36.860 ;
        RECT 139.615 36.170 140.115 36.340 ;
        RECT 139.385 35.925 139.555 35.955 ;
        RECT 138.660 34.945 139.555 35.925 ;
        RECT 136.015 33.840 138.315 34.010 ;
        RECT 138.715 34.010 138.885 34.945 ;
        RECT 139.385 34.915 139.555 34.945 ;
        RECT 140.175 34.915 140.345 35.955 ;
        RECT 139.200 34.530 140.115 34.700 ;
        RECT 139.200 34.325 140.035 34.530 ;
        RECT 140.845 34.010 141.015 36.860 ;
        RECT 141.415 36.860 143.715 37.030 ;
        RECT 141.415 35.925 141.585 36.860 ;
        RECT 142.315 36.170 142.815 36.340 ;
        RECT 142.085 35.925 142.255 35.955 ;
        RECT 141.360 34.945 142.255 35.925 ;
        RECT 138.715 33.840 141.015 34.010 ;
        RECT 141.415 34.010 141.585 34.945 ;
        RECT 142.085 34.915 142.255 34.945 ;
        RECT 142.875 34.915 143.045 35.955 ;
        RECT 141.900 34.530 142.815 34.700 ;
        RECT 141.900 34.325 142.735 34.530 ;
        RECT 143.545 34.010 143.715 36.860 ;
        RECT 141.415 33.840 143.715 34.010 ;
        RECT 144.115 34.010 144.285 45.860 ;
        RECT 144.775 45.150 145.775 45.600 ;
        RECT 144.785 34.915 144.955 44.955 ;
        RECT 145.575 34.915 145.745 44.955 ;
        RECT 145.015 34.530 145.515 34.700 ;
        RECT 146.245 34.010 146.415 45.860 ;
        RECT 144.115 33.840 146.415 34.010 ;
        RECT 146.815 45.860 149.115 46.030 ;
        RECT 146.815 34.010 146.985 45.860 ;
        RECT 147.475 45.150 148.475 45.600 ;
        RECT 147.485 34.915 147.655 44.955 ;
        RECT 148.275 34.915 148.445 44.955 ;
        RECT 147.715 34.530 148.215 34.700 ;
        RECT 148.945 34.010 149.115 45.860 ;
        RECT 146.815 33.840 149.115 34.010 ;
        RECT 6.190 32.770 8.490 32.940 ;
        RECT 6.190 31.830 6.360 32.770 ;
        RECT 6.570 32.080 7.610 32.525 ;
        RECT 6.860 31.830 7.030 31.910 ;
        RECT 6.185 31.300 7.030 31.830 ;
        RECT 6.190 30.360 6.360 31.300 ;
        RECT 6.860 31.220 7.030 31.300 ;
        RECT 7.650 31.220 7.820 31.910 ;
        RECT 7.090 30.880 7.590 31.050 ;
        RECT 8.320 30.360 8.490 32.770 ;
        RECT 6.190 30.190 8.490 30.360 ;
        RECT 8.890 32.770 11.190 32.940 ;
        RECT 8.890 24.510 9.060 32.770 ;
        RECT 9.790 32.080 10.290 32.250 ;
        RECT 9.560 25.370 9.730 31.910 ;
        RECT 10.350 25.370 10.520 31.910 ;
        RECT 9.550 24.800 10.550 25.200 ;
        RECT 11.020 24.510 11.190 32.770 ;
        RECT 11.590 32.770 13.890 32.940 ;
        RECT 11.590 31.830 11.760 32.770 ;
        RECT 11.970 32.080 13.010 32.525 ;
        RECT 12.260 31.830 12.430 31.910 ;
        RECT 11.585 31.300 12.430 31.830 ;
        RECT 11.590 30.360 11.760 31.300 ;
        RECT 12.260 31.220 12.430 31.300 ;
        RECT 13.050 31.220 13.220 31.910 ;
        RECT 12.490 30.880 12.990 31.050 ;
        RECT 13.720 30.360 13.890 32.770 ;
        RECT 14.290 32.770 16.590 32.940 ;
        RECT 14.290 31.830 14.460 32.770 ;
        RECT 14.670 32.080 15.710 32.525 ;
        RECT 14.960 31.830 15.130 31.910 ;
        RECT 14.285 31.300 15.130 31.830 ;
        RECT 11.590 30.190 13.890 30.360 ;
        RECT 14.290 30.360 14.460 31.300 ;
        RECT 14.960 31.220 15.130 31.300 ;
        RECT 15.750 31.220 15.920 31.910 ;
        RECT 15.190 30.880 15.690 31.050 ;
        RECT 16.420 30.360 16.590 32.770 ;
        RECT 14.290 30.190 16.590 30.360 ;
        RECT 16.990 32.770 19.290 32.940 ;
        RECT 8.890 24.340 11.190 24.510 ;
        RECT 16.990 24.510 17.160 32.770 ;
        RECT 17.890 32.080 18.390 32.250 ;
        RECT 17.660 25.370 17.830 31.910 ;
        RECT 18.450 25.370 18.620 31.910 ;
        RECT 17.650 24.800 18.650 25.200 ;
        RECT 19.120 24.510 19.290 32.770 ;
        RECT 16.990 24.340 19.290 24.510 ;
        RECT 19.690 32.770 21.990 32.940 ;
        RECT 19.690 24.510 19.860 32.770 ;
        RECT 20.590 32.080 21.090 32.250 ;
        RECT 20.360 25.370 20.530 31.910 ;
        RECT 21.150 25.370 21.320 31.910 ;
        RECT 20.350 24.800 21.350 25.200 ;
        RECT 21.820 24.510 21.990 32.770 ;
        RECT 31.615 32.770 33.915 32.940 ;
        RECT 31.615 31.830 31.785 32.770 ;
        RECT 31.995 32.080 33.035 32.525 ;
        RECT 32.285 31.830 32.455 31.910 ;
        RECT 31.610 31.300 32.455 31.830 ;
        RECT 31.615 30.360 31.785 31.300 ;
        RECT 32.285 31.220 32.455 31.300 ;
        RECT 33.075 31.220 33.245 31.910 ;
        RECT 32.515 30.880 33.015 31.050 ;
        RECT 33.745 30.360 33.915 32.770 ;
        RECT 31.615 30.190 33.915 30.360 ;
        RECT 34.315 32.770 36.615 32.940 ;
        RECT 19.690 24.340 21.990 24.510 ;
        RECT 34.315 24.510 34.485 32.770 ;
        RECT 35.215 32.080 35.715 32.250 ;
        RECT 34.985 25.370 35.155 31.910 ;
        RECT 35.775 25.370 35.945 31.910 ;
        RECT 34.975 24.800 35.975 25.200 ;
        RECT 36.445 24.510 36.615 32.770 ;
        RECT 37.015 32.770 39.315 32.940 ;
        RECT 37.015 31.830 37.185 32.770 ;
        RECT 37.395 32.080 38.435 32.525 ;
        RECT 37.685 31.830 37.855 31.910 ;
        RECT 37.010 31.300 37.855 31.830 ;
        RECT 37.015 30.360 37.185 31.300 ;
        RECT 37.685 31.220 37.855 31.300 ;
        RECT 38.475 31.220 38.645 31.910 ;
        RECT 37.915 30.880 38.415 31.050 ;
        RECT 39.145 30.360 39.315 32.770 ;
        RECT 39.715 32.770 42.015 32.940 ;
        RECT 39.715 31.830 39.885 32.770 ;
        RECT 40.095 32.080 41.135 32.525 ;
        RECT 40.385 31.830 40.555 31.910 ;
        RECT 39.710 31.300 40.555 31.830 ;
        RECT 37.015 30.190 39.315 30.360 ;
        RECT 39.715 30.360 39.885 31.300 ;
        RECT 40.385 31.220 40.555 31.300 ;
        RECT 41.175 31.220 41.345 31.910 ;
        RECT 40.615 30.880 41.115 31.050 ;
        RECT 41.845 30.360 42.015 32.770 ;
        RECT 39.715 30.190 42.015 30.360 ;
        RECT 42.415 32.770 44.715 32.940 ;
        RECT 34.315 24.340 36.615 24.510 ;
        RECT 42.415 24.510 42.585 32.770 ;
        RECT 43.315 32.080 43.815 32.250 ;
        RECT 43.085 25.370 43.255 31.910 ;
        RECT 43.875 25.370 44.045 31.910 ;
        RECT 43.075 24.800 44.075 25.200 ;
        RECT 44.545 24.510 44.715 32.770 ;
        RECT 42.415 24.340 44.715 24.510 ;
        RECT 45.115 32.770 47.415 32.940 ;
        RECT 45.115 24.510 45.285 32.770 ;
        RECT 46.015 32.080 46.515 32.250 ;
        RECT 45.785 25.370 45.955 31.910 ;
        RECT 46.575 25.370 46.745 31.910 ;
        RECT 45.775 24.800 46.775 25.200 ;
        RECT 47.245 24.510 47.415 32.770 ;
        RECT 57.040 32.770 59.340 32.940 ;
        RECT 57.040 31.830 57.210 32.770 ;
        RECT 57.420 32.080 58.460 32.525 ;
        RECT 57.710 31.830 57.880 31.910 ;
        RECT 57.035 31.300 57.880 31.830 ;
        RECT 57.040 30.360 57.210 31.300 ;
        RECT 57.710 31.220 57.880 31.300 ;
        RECT 58.500 31.220 58.670 31.910 ;
        RECT 57.940 30.880 58.440 31.050 ;
        RECT 59.170 30.360 59.340 32.770 ;
        RECT 57.040 30.190 59.340 30.360 ;
        RECT 59.740 32.770 62.040 32.940 ;
        RECT 45.115 24.340 47.415 24.510 ;
        RECT 59.740 24.510 59.910 32.770 ;
        RECT 60.640 32.080 61.140 32.250 ;
        RECT 60.410 25.370 60.580 31.910 ;
        RECT 61.200 25.370 61.370 31.910 ;
        RECT 60.400 24.800 61.400 25.200 ;
        RECT 61.870 24.510 62.040 32.770 ;
        RECT 62.440 32.770 64.740 32.940 ;
        RECT 62.440 31.830 62.610 32.770 ;
        RECT 62.820 32.080 63.860 32.525 ;
        RECT 63.110 31.830 63.280 31.910 ;
        RECT 62.435 31.300 63.280 31.830 ;
        RECT 62.440 30.360 62.610 31.300 ;
        RECT 63.110 31.220 63.280 31.300 ;
        RECT 63.900 31.220 64.070 31.910 ;
        RECT 63.340 30.880 63.840 31.050 ;
        RECT 64.570 30.360 64.740 32.770 ;
        RECT 65.140 32.770 67.440 32.940 ;
        RECT 65.140 31.830 65.310 32.770 ;
        RECT 65.520 32.080 66.560 32.525 ;
        RECT 65.810 31.830 65.980 31.910 ;
        RECT 65.135 31.300 65.980 31.830 ;
        RECT 62.440 30.190 64.740 30.360 ;
        RECT 65.140 30.360 65.310 31.300 ;
        RECT 65.810 31.220 65.980 31.300 ;
        RECT 66.600 31.220 66.770 31.910 ;
        RECT 66.040 30.880 66.540 31.050 ;
        RECT 67.270 30.360 67.440 32.770 ;
        RECT 65.140 30.190 67.440 30.360 ;
        RECT 67.840 32.770 70.140 32.940 ;
        RECT 59.740 24.340 62.040 24.510 ;
        RECT 67.840 24.510 68.010 32.770 ;
        RECT 68.740 32.080 69.240 32.250 ;
        RECT 68.510 25.370 68.680 31.910 ;
        RECT 69.300 25.370 69.470 31.910 ;
        RECT 68.500 24.800 69.500 25.200 ;
        RECT 69.970 24.510 70.140 32.770 ;
        RECT 67.840 24.340 70.140 24.510 ;
        RECT 70.540 32.770 72.840 32.940 ;
        RECT 70.540 24.510 70.710 32.770 ;
        RECT 71.440 32.080 71.940 32.250 ;
        RECT 71.210 25.370 71.380 31.910 ;
        RECT 72.000 25.370 72.170 31.910 ;
        RECT 71.200 24.800 72.200 25.200 ;
        RECT 72.670 24.510 72.840 32.770 ;
        RECT 82.465 32.770 84.765 32.940 ;
        RECT 82.465 31.830 82.635 32.770 ;
        RECT 82.845 32.080 83.885 32.525 ;
        RECT 83.135 31.830 83.305 31.910 ;
        RECT 82.460 31.300 83.305 31.830 ;
        RECT 82.465 30.360 82.635 31.300 ;
        RECT 83.135 31.220 83.305 31.300 ;
        RECT 83.925 31.220 84.095 31.910 ;
        RECT 83.365 30.880 83.865 31.050 ;
        RECT 84.595 30.360 84.765 32.770 ;
        RECT 82.465 30.190 84.765 30.360 ;
        RECT 85.165 32.770 87.465 32.940 ;
        RECT 70.540 24.340 72.840 24.510 ;
        RECT 85.165 24.510 85.335 32.770 ;
        RECT 86.065 32.080 86.565 32.250 ;
        RECT 85.835 25.370 86.005 31.910 ;
        RECT 86.625 25.370 86.795 31.910 ;
        RECT 85.825 24.800 86.825 25.200 ;
        RECT 87.295 24.510 87.465 32.770 ;
        RECT 87.865 32.770 90.165 32.940 ;
        RECT 87.865 31.830 88.035 32.770 ;
        RECT 88.245 32.080 89.285 32.525 ;
        RECT 88.535 31.830 88.705 31.910 ;
        RECT 87.860 31.300 88.705 31.830 ;
        RECT 87.865 30.360 88.035 31.300 ;
        RECT 88.535 31.220 88.705 31.300 ;
        RECT 89.325 31.220 89.495 31.910 ;
        RECT 88.765 30.880 89.265 31.050 ;
        RECT 89.995 30.360 90.165 32.770 ;
        RECT 90.565 32.770 92.865 32.940 ;
        RECT 90.565 31.830 90.735 32.770 ;
        RECT 90.945 32.080 91.985 32.525 ;
        RECT 91.235 31.830 91.405 31.910 ;
        RECT 90.560 31.300 91.405 31.830 ;
        RECT 87.865 30.190 90.165 30.360 ;
        RECT 90.565 30.360 90.735 31.300 ;
        RECT 91.235 31.220 91.405 31.300 ;
        RECT 92.025 31.220 92.195 31.910 ;
        RECT 91.465 30.880 91.965 31.050 ;
        RECT 92.695 30.360 92.865 32.770 ;
        RECT 90.565 30.190 92.865 30.360 ;
        RECT 93.265 32.770 95.565 32.940 ;
        RECT 85.165 24.340 87.465 24.510 ;
        RECT 93.265 24.510 93.435 32.770 ;
        RECT 94.165 32.080 94.665 32.250 ;
        RECT 93.935 25.370 94.105 31.910 ;
        RECT 94.725 25.370 94.895 31.910 ;
        RECT 93.925 24.800 94.925 25.200 ;
        RECT 95.395 24.510 95.565 32.770 ;
        RECT 93.265 24.340 95.565 24.510 ;
        RECT 95.965 32.770 98.265 32.940 ;
        RECT 95.965 24.510 96.135 32.770 ;
        RECT 96.865 32.080 97.365 32.250 ;
        RECT 96.635 25.370 96.805 31.910 ;
        RECT 97.425 25.370 97.595 31.910 ;
        RECT 96.625 24.800 97.625 25.200 ;
        RECT 98.095 24.510 98.265 32.770 ;
        RECT 107.890 32.770 110.190 32.940 ;
        RECT 107.890 31.830 108.060 32.770 ;
        RECT 108.270 32.080 109.310 32.525 ;
        RECT 108.560 31.830 108.730 31.910 ;
        RECT 107.885 31.300 108.730 31.830 ;
        RECT 107.890 30.360 108.060 31.300 ;
        RECT 108.560 31.220 108.730 31.300 ;
        RECT 109.350 31.220 109.520 31.910 ;
        RECT 108.790 30.880 109.290 31.050 ;
        RECT 110.020 30.360 110.190 32.770 ;
        RECT 107.890 30.190 110.190 30.360 ;
        RECT 110.590 32.770 112.890 32.940 ;
        RECT 95.965 24.340 98.265 24.510 ;
        RECT 110.590 24.510 110.760 32.770 ;
        RECT 111.490 32.080 111.990 32.250 ;
        RECT 111.260 25.370 111.430 31.910 ;
        RECT 112.050 25.370 112.220 31.910 ;
        RECT 111.250 24.800 112.250 25.200 ;
        RECT 112.720 24.510 112.890 32.770 ;
        RECT 113.290 32.770 115.590 32.940 ;
        RECT 113.290 31.830 113.460 32.770 ;
        RECT 113.670 32.080 114.710 32.525 ;
        RECT 113.960 31.830 114.130 31.910 ;
        RECT 113.285 31.300 114.130 31.830 ;
        RECT 113.290 30.360 113.460 31.300 ;
        RECT 113.960 31.220 114.130 31.300 ;
        RECT 114.750 31.220 114.920 31.910 ;
        RECT 114.190 30.880 114.690 31.050 ;
        RECT 115.420 30.360 115.590 32.770 ;
        RECT 115.990 32.770 118.290 32.940 ;
        RECT 115.990 31.830 116.160 32.770 ;
        RECT 116.370 32.080 117.410 32.525 ;
        RECT 116.660 31.830 116.830 31.910 ;
        RECT 115.985 31.300 116.830 31.830 ;
        RECT 113.290 30.190 115.590 30.360 ;
        RECT 115.990 30.360 116.160 31.300 ;
        RECT 116.660 31.220 116.830 31.300 ;
        RECT 117.450 31.220 117.620 31.910 ;
        RECT 116.890 30.880 117.390 31.050 ;
        RECT 118.120 30.360 118.290 32.770 ;
        RECT 115.990 30.190 118.290 30.360 ;
        RECT 118.690 32.770 120.990 32.940 ;
        RECT 110.590 24.340 112.890 24.510 ;
        RECT 118.690 24.510 118.860 32.770 ;
        RECT 119.590 32.080 120.090 32.250 ;
        RECT 119.360 25.370 119.530 31.910 ;
        RECT 120.150 25.370 120.320 31.910 ;
        RECT 119.350 24.800 120.350 25.200 ;
        RECT 120.820 24.510 120.990 32.770 ;
        RECT 118.690 24.340 120.990 24.510 ;
        RECT 121.390 32.770 123.690 32.940 ;
        RECT 121.390 24.510 121.560 32.770 ;
        RECT 122.290 32.080 122.790 32.250 ;
        RECT 122.060 25.370 122.230 31.910 ;
        RECT 122.850 25.370 123.020 31.910 ;
        RECT 122.050 24.800 123.050 25.200 ;
        RECT 123.520 24.510 123.690 32.770 ;
        RECT 133.315 32.770 135.615 32.940 ;
        RECT 133.315 31.830 133.485 32.770 ;
        RECT 133.695 32.080 134.735 32.525 ;
        RECT 133.985 31.830 134.155 31.910 ;
        RECT 133.310 31.300 134.155 31.830 ;
        RECT 133.315 30.360 133.485 31.300 ;
        RECT 133.985 31.220 134.155 31.300 ;
        RECT 134.775 31.220 134.945 31.910 ;
        RECT 134.215 30.880 134.715 31.050 ;
        RECT 135.445 30.360 135.615 32.770 ;
        RECT 133.315 30.190 135.615 30.360 ;
        RECT 136.015 32.770 138.315 32.940 ;
        RECT 121.390 24.340 123.690 24.510 ;
        RECT 136.015 24.510 136.185 32.770 ;
        RECT 136.915 32.080 137.415 32.250 ;
        RECT 136.685 25.370 136.855 31.910 ;
        RECT 137.475 25.370 137.645 31.910 ;
        RECT 136.675 24.800 137.675 25.200 ;
        RECT 138.145 24.510 138.315 32.770 ;
        RECT 138.715 32.770 141.015 32.940 ;
        RECT 138.715 31.830 138.885 32.770 ;
        RECT 139.095 32.080 140.135 32.525 ;
        RECT 139.385 31.830 139.555 31.910 ;
        RECT 138.710 31.300 139.555 31.830 ;
        RECT 138.715 30.360 138.885 31.300 ;
        RECT 139.385 31.220 139.555 31.300 ;
        RECT 140.175 31.220 140.345 31.910 ;
        RECT 139.615 30.880 140.115 31.050 ;
        RECT 140.845 30.360 141.015 32.770 ;
        RECT 141.415 32.770 143.715 32.940 ;
        RECT 141.415 31.830 141.585 32.770 ;
        RECT 141.795 32.080 142.835 32.525 ;
        RECT 142.085 31.830 142.255 31.910 ;
        RECT 141.410 31.300 142.255 31.830 ;
        RECT 138.715 30.190 141.015 30.360 ;
        RECT 141.415 30.360 141.585 31.300 ;
        RECT 142.085 31.220 142.255 31.300 ;
        RECT 142.875 31.220 143.045 31.910 ;
        RECT 142.315 30.880 142.815 31.050 ;
        RECT 143.545 30.360 143.715 32.770 ;
        RECT 141.415 30.190 143.715 30.360 ;
        RECT 144.115 32.770 146.415 32.940 ;
        RECT 136.015 24.340 138.315 24.510 ;
        RECT 144.115 24.510 144.285 32.770 ;
        RECT 145.015 32.080 145.515 32.250 ;
        RECT 144.785 25.370 144.955 31.910 ;
        RECT 145.575 25.370 145.745 31.910 ;
        RECT 144.775 24.800 145.775 25.200 ;
        RECT 146.245 24.510 146.415 32.770 ;
        RECT 144.115 24.340 146.415 24.510 ;
        RECT 146.815 32.770 149.115 32.940 ;
        RECT 146.815 24.510 146.985 32.770 ;
        RECT 147.715 32.080 148.215 32.250 ;
        RECT 147.485 25.370 147.655 31.910 ;
        RECT 148.275 25.370 148.445 31.910 ;
        RECT 147.475 24.800 148.475 25.200 ;
        RECT 148.945 24.510 149.115 32.770 ;
        RECT 146.815 24.340 149.115 24.510 ;
        RECT 23.235 24.000 24.075 24.050 ;
        RECT 48.660 24.000 49.500 24.050 ;
        RECT 74.085 24.000 74.925 24.050 ;
        RECT 99.510 24.000 100.350 24.050 ;
        RECT 124.935 24.000 125.775 24.050 ;
        RECT 150.360 24.000 151.200 24.050 ;
        RECT 22.830 23.830 24.480 24.000 ;
        RECT 8.890 23.285 11.190 23.455 ;
        RECT 6.190 14.285 8.490 14.455 ;
        RECT 6.190 13.350 6.360 14.285 ;
        RECT 7.090 13.595 7.590 13.765 ;
        RECT 6.860 13.350 7.030 13.380 ;
        RECT 6.135 12.370 7.030 13.350 ;
        RECT 6.190 11.435 6.360 12.370 ;
        RECT 6.860 12.340 7.030 12.370 ;
        RECT 7.650 12.340 7.820 13.380 ;
        RECT 6.675 11.955 7.590 12.125 ;
        RECT 6.675 11.750 7.510 11.955 ;
        RECT 8.320 11.435 8.490 14.285 ;
        RECT 6.190 11.265 8.490 11.435 ;
        RECT 8.890 11.435 9.060 23.285 ;
        RECT 9.550 22.575 10.550 23.025 ;
        RECT 9.560 12.340 9.730 22.380 ;
        RECT 10.350 12.340 10.520 22.380 ;
        RECT 9.790 11.955 10.290 12.125 ;
        RECT 11.020 11.435 11.190 23.285 ;
        RECT 16.990 23.285 19.290 23.455 ;
        RECT 11.590 14.285 13.890 14.455 ;
        RECT 11.590 13.350 11.760 14.285 ;
        RECT 12.490 13.595 12.990 13.765 ;
        RECT 12.260 13.350 12.430 13.380 ;
        RECT 11.535 12.370 12.430 13.350 ;
        RECT 8.890 11.265 11.190 11.435 ;
        RECT 11.590 11.435 11.760 12.370 ;
        RECT 12.260 12.340 12.430 12.370 ;
        RECT 13.050 12.340 13.220 13.380 ;
        RECT 12.075 11.955 12.990 12.125 ;
        RECT 12.075 11.750 12.910 11.955 ;
        RECT 13.720 11.435 13.890 14.285 ;
        RECT 14.290 14.285 16.590 14.455 ;
        RECT 14.290 13.350 14.460 14.285 ;
        RECT 15.190 13.595 15.690 13.765 ;
        RECT 14.960 13.350 15.130 13.380 ;
        RECT 14.235 12.370 15.130 13.350 ;
        RECT 11.590 11.265 13.890 11.435 ;
        RECT 14.290 11.435 14.460 12.370 ;
        RECT 14.960 12.340 15.130 12.370 ;
        RECT 15.750 12.340 15.920 13.380 ;
        RECT 14.775 11.955 15.690 12.125 ;
        RECT 14.775 11.750 15.610 11.955 ;
        RECT 16.420 11.435 16.590 14.285 ;
        RECT 14.290 11.265 16.590 11.435 ;
        RECT 16.990 11.435 17.160 23.285 ;
        RECT 17.650 22.575 18.650 23.025 ;
        RECT 17.660 12.340 17.830 22.380 ;
        RECT 18.450 12.340 18.620 22.380 ;
        RECT 17.890 11.955 18.390 12.125 ;
        RECT 19.120 11.435 19.290 23.285 ;
        RECT 16.990 11.265 19.290 11.435 ;
        RECT 19.690 23.285 21.990 23.455 ;
        RECT 19.690 11.435 19.860 23.285 ;
        RECT 20.350 22.575 21.350 23.025 ;
        RECT 20.360 12.340 20.530 22.380 ;
        RECT 21.150 12.340 21.320 22.380 ;
        RECT 20.590 11.955 21.090 12.125 ;
        RECT 21.820 11.435 21.990 23.285 ;
        RECT 19.690 11.265 21.990 11.435 ;
        RECT 6.190 10.195 8.490 10.365 ;
        RECT 6.190 9.255 6.360 10.195 ;
        RECT 6.570 9.505 7.610 9.950 ;
        RECT 6.860 9.255 7.030 9.335 ;
        RECT 6.185 8.725 7.030 9.255 ;
        RECT 6.190 7.785 6.360 8.725 ;
        RECT 6.860 8.645 7.030 8.725 ;
        RECT 7.650 8.645 7.820 9.335 ;
        RECT 7.090 8.305 7.590 8.475 ;
        RECT 8.320 7.785 8.490 10.195 ;
        RECT 6.190 7.615 8.490 7.785 ;
        RECT 8.890 10.195 11.190 10.365 ;
        RECT 8.890 1.935 9.060 10.195 ;
        RECT 9.790 9.505 10.290 9.675 ;
        RECT 9.560 2.795 9.730 9.335 ;
        RECT 10.350 2.795 10.520 9.335 ;
        RECT 9.550 2.225 10.550 2.625 ;
        RECT 11.020 1.935 11.190 10.195 ;
        RECT 11.590 10.195 13.890 10.365 ;
        RECT 11.590 9.255 11.760 10.195 ;
        RECT 11.970 9.505 13.010 9.950 ;
        RECT 12.260 9.255 12.430 9.335 ;
        RECT 11.585 8.725 12.430 9.255 ;
        RECT 11.590 7.785 11.760 8.725 ;
        RECT 12.260 8.645 12.430 8.725 ;
        RECT 13.050 8.645 13.220 9.335 ;
        RECT 12.490 8.305 12.990 8.475 ;
        RECT 13.720 7.785 13.890 10.195 ;
        RECT 14.290 10.195 16.590 10.365 ;
        RECT 14.290 9.255 14.460 10.195 ;
        RECT 14.670 9.505 15.710 9.950 ;
        RECT 14.960 9.255 15.130 9.335 ;
        RECT 14.285 8.725 15.130 9.255 ;
        RECT 11.590 7.615 13.890 7.785 ;
        RECT 14.290 7.785 14.460 8.725 ;
        RECT 14.960 8.645 15.130 8.725 ;
        RECT 15.750 8.645 15.920 9.335 ;
        RECT 15.190 8.305 15.690 8.475 ;
        RECT 16.420 7.785 16.590 10.195 ;
        RECT 14.290 7.615 16.590 7.785 ;
        RECT 16.990 10.195 19.290 10.365 ;
        RECT 8.890 1.765 11.190 1.935 ;
        RECT 16.990 1.935 17.160 10.195 ;
        RECT 17.890 9.505 18.390 9.675 ;
        RECT 17.660 2.795 17.830 9.335 ;
        RECT 18.450 2.795 18.620 9.335 ;
        RECT 17.650 2.225 18.650 2.625 ;
        RECT 19.120 1.935 19.290 10.195 ;
        RECT 16.990 1.765 19.290 1.935 ;
        RECT 19.690 10.195 21.990 10.365 ;
        RECT 19.690 1.935 19.860 10.195 ;
        RECT 20.590 9.505 21.090 9.675 ;
        RECT 20.360 2.795 20.530 9.335 ;
        RECT 21.150 2.795 21.320 9.335 ;
        RECT 20.350 2.225 21.350 2.625 ;
        RECT 21.820 1.935 21.990 10.195 ;
        RECT 22.830 9.800 23.000 23.830 ;
        RECT 23.235 23.780 24.075 23.830 ;
        RECT 23.430 21.115 23.880 23.425 ;
        RECT 23.430 10.205 23.880 12.515 ;
        RECT 23.260 9.800 24.050 9.850 ;
        RECT 24.310 9.800 24.480 23.830 ;
        RECT 48.255 23.830 49.905 24.000 ;
        RECT 34.315 23.285 36.615 23.455 ;
        RECT 31.615 14.285 33.915 14.455 ;
        RECT 31.615 13.350 31.785 14.285 ;
        RECT 32.515 13.595 33.015 13.765 ;
        RECT 32.285 13.350 32.455 13.380 ;
        RECT 31.560 12.370 32.455 13.350 ;
        RECT 31.615 11.435 31.785 12.370 ;
        RECT 32.285 12.340 32.455 12.370 ;
        RECT 33.075 12.340 33.245 13.380 ;
        RECT 32.100 11.955 33.015 12.125 ;
        RECT 32.100 11.750 32.935 11.955 ;
        RECT 33.745 11.435 33.915 14.285 ;
        RECT 31.615 11.265 33.915 11.435 ;
        RECT 34.315 11.435 34.485 23.285 ;
        RECT 34.975 22.575 35.975 23.025 ;
        RECT 34.985 12.340 35.155 22.380 ;
        RECT 35.775 12.340 35.945 22.380 ;
        RECT 35.215 11.955 35.715 12.125 ;
        RECT 36.445 11.435 36.615 23.285 ;
        RECT 42.415 23.285 44.715 23.455 ;
        RECT 37.015 14.285 39.315 14.455 ;
        RECT 37.015 13.350 37.185 14.285 ;
        RECT 37.915 13.595 38.415 13.765 ;
        RECT 37.685 13.350 37.855 13.380 ;
        RECT 36.960 12.370 37.855 13.350 ;
        RECT 34.315 11.265 36.615 11.435 ;
        RECT 37.015 11.435 37.185 12.370 ;
        RECT 37.685 12.340 37.855 12.370 ;
        RECT 38.475 12.340 38.645 13.380 ;
        RECT 37.500 11.955 38.415 12.125 ;
        RECT 37.500 11.750 38.335 11.955 ;
        RECT 39.145 11.435 39.315 14.285 ;
        RECT 39.715 14.285 42.015 14.455 ;
        RECT 39.715 13.350 39.885 14.285 ;
        RECT 40.615 13.595 41.115 13.765 ;
        RECT 40.385 13.350 40.555 13.380 ;
        RECT 39.660 12.370 40.555 13.350 ;
        RECT 37.015 11.265 39.315 11.435 ;
        RECT 39.715 11.435 39.885 12.370 ;
        RECT 40.385 12.340 40.555 12.370 ;
        RECT 41.175 12.340 41.345 13.380 ;
        RECT 40.200 11.955 41.115 12.125 ;
        RECT 40.200 11.750 41.035 11.955 ;
        RECT 41.845 11.435 42.015 14.285 ;
        RECT 39.715 11.265 42.015 11.435 ;
        RECT 42.415 11.435 42.585 23.285 ;
        RECT 43.075 22.575 44.075 23.025 ;
        RECT 43.085 12.340 43.255 22.380 ;
        RECT 43.875 12.340 44.045 22.380 ;
        RECT 43.315 11.955 43.815 12.125 ;
        RECT 44.545 11.435 44.715 23.285 ;
        RECT 42.415 11.265 44.715 11.435 ;
        RECT 45.115 23.285 47.415 23.455 ;
        RECT 45.115 11.435 45.285 23.285 ;
        RECT 45.775 22.575 46.775 23.025 ;
        RECT 45.785 12.340 45.955 22.380 ;
        RECT 46.575 12.340 46.745 22.380 ;
        RECT 46.015 11.955 46.515 12.125 ;
        RECT 47.245 11.435 47.415 23.285 ;
        RECT 45.115 11.265 47.415 11.435 ;
        RECT 22.830 9.630 24.480 9.800 ;
        RECT 31.615 10.195 33.915 10.365 ;
        RECT 23.260 9.580 24.050 9.630 ;
        RECT 31.615 9.255 31.785 10.195 ;
        RECT 31.995 9.505 33.035 9.950 ;
        RECT 32.285 9.255 32.455 9.335 ;
        RECT 31.610 8.725 32.455 9.255 ;
        RECT 31.615 7.785 31.785 8.725 ;
        RECT 32.285 8.645 32.455 8.725 ;
        RECT 33.075 8.645 33.245 9.335 ;
        RECT 32.515 8.305 33.015 8.475 ;
        RECT 33.745 7.785 33.915 10.195 ;
        RECT 31.615 7.615 33.915 7.785 ;
        RECT 34.315 10.195 36.615 10.365 ;
        RECT 19.690 1.765 21.990 1.935 ;
        RECT 34.315 1.935 34.485 10.195 ;
        RECT 35.215 9.505 35.715 9.675 ;
        RECT 34.985 2.795 35.155 9.335 ;
        RECT 35.775 2.795 35.945 9.335 ;
        RECT 34.975 2.225 35.975 2.625 ;
        RECT 36.445 1.935 36.615 10.195 ;
        RECT 37.015 10.195 39.315 10.365 ;
        RECT 37.015 9.255 37.185 10.195 ;
        RECT 37.395 9.505 38.435 9.950 ;
        RECT 37.685 9.255 37.855 9.335 ;
        RECT 37.010 8.725 37.855 9.255 ;
        RECT 37.015 7.785 37.185 8.725 ;
        RECT 37.685 8.645 37.855 8.725 ;
        RECT 38.475 8.645 38.645 9.335 ;
        RECT 37.915 8.305 38.415 8.475 ;
        RECT 39.145 7.785 39.315 10.195 ;
        RECT 39.715 10.195 42.015 10.365 ;
        RECT 39.715 9.255 39.885 10.195 ;
        RECT 40.095 9.505 41.135 9.950 ;
        RECT 40.385 9.255 40.555 9.335 ;
        RECT 39.710 8.725 40.555 9.255 ;
        RECT 37.015 7.615 39.315 7.785 ;
        RECT 39.715 7.785 39.885 8.725 ;
        RECT 40.385 8.645 40.555 8.725 ;
        RECT 41.175 8.645 41.345 9.335 ;
        RECT 40.615 8.305 41.115 8.475 ;
        RECT 41.845 7.785 42.015 10.195 ;
        RECT 39.715 7.615 42.015 7.785 ;
        RECT 42.415 10.195 44.715 10.365 ;
        RECT 34.315 1.765 36.615 1.935 ;
        RECT 42.415 1.935 42.585 10.195 ;
        RECT 43.315 9.505 43.815 9.675 ;
        RECT 43.085 2.795 43.255 9.335 ;
        RECT 43.875 2.795 44.045 9.335 ;
        RECT 43.075 2.225 44.075 2.625 ;
        RECT 44.545 1.935 44.715 10.195 ;
        RECT 42.415 1.765 44.715 1.935 ;
        RECT 45.115 10.195 47.415 10.365 ;
        RECT 45.115 1.935 45.285 10.195 ;
        RECT 46.015 9.505 46.515 9.675 ;
        RECT 45.785 2.795 45.955 9.335 ;
        RECT 46.575 2.795 46.745 9.335 ;
        RECT 45.775 2.225 46.775 2.625 ;
        RECT 47.245 1.935 47.415 10.195 ;
        RECT 48.255 9.800 48.425 23.830 ;
        RECT 48.660 23.780 49.500 23.830 ;
        RECT 48.855 21.115 49.305 23.425 ;
        RECT 48.855 10.205 49.305 12.515 ;
        RECT 48.685 9.800 49.475 9.850 ;
        RECT 49.735 9.800 49.905 23.830 ;
        RECT 73.680 23.830 75.330 24.000 ;
        RECT 59.740 23.285 62.040 23.455 ;
        RECT 57.040 14.285 59.340 14.455 ;
        RECT 57.040 13.350 57.210 14.285 ;
        RECT 57.940 13.595 58.440 13.765 ;
        RECT 57.710 13.350 57.880 13.380 ;
        RECT 56.985 12.370 57.880 13.350 ;
        RECT 57.040 11.435 57.210 12.370 ;
        RECT 57.710 12.340 57.880 12.370 ;
        RECT 58.500 12.340 58.670 13.380 ;
        RECT 57.525 11.955 58.440 12.125 ;
        RECT 57.525 11.750 58.360 11.955 ;
        RECT 59.170 11.435 59.340 14.285 ;
        RECT 57.040 11.265 59.340 11.435 ;
        RECT 59.740 11.435 59.910 23.285 ;
        RECT 60.400 22.575 61.400 23.025 ;
        RECT 60.410 12.340 60.580 22.380 ;
        RECT 61.200 12.340 61.370 22.380 ;
        RECT 60.640 11.955 61.140 12.125 ;
        RECT 61.870 11.435 62.040 23.285 ;
        RECT 67.840 23.285 70.140 23.455 ;
        RECT 62.440 14.285 64.740 14.455 ;
        RECT 62.440 13.350 62.610 14.285 ;
        RECT 63.340 13.595 63.840 13.765 ;
        RECT 63.110 13.350 63.280 13.380 ;
        RECT 62.385 12.370 63.280 13.350 ;
        RECT 59.740 11.265 62.040 11.435 ;
        RECT 62.440 11.435 62.610 12.370 ;
        RECT 63.110 12.340 63.280 12.370 ;
        RECT 63.900 12.340 64.070 13.380 ;
        RECT 62.925 11.955 63.840 12.125 ;
        RECT 62.925 11.750 63.760 11.955 ;
        RECT 64.570 11.435 64.740 14.285 ;
        RECT 65.140 14.285 67.440 14.455 ;
        RECT 65.140 13.350 65.310 14.285 ;
        RECT 66.040 13.595 66.540 13.765 ;
        RECT 65.810 13.350 65.980 13.380 ;
        RECT 65.085 12.370 65.980 13.350 ;
        RECT 62.440 11.265 64.740 11.435 ;
        RECT 65.140 11.435 65.310 12.370 ;
        RECT 65.810 12.340 65.980 12.370 ;
        RECT 66.600 12.340 66.770 13.380 ;
        RECT 65.625 11.955 66.540 12.125 ;
        RECT 65.625 11.750 66.460 11.955 ;
        RECT 67.270 11.435 67.440 14.285 ;
        RECT 65.140 11.265 67.440 11.435 ;
        RECT 67.840 11.435 68.010 23.285 ;
        RECT 68.500 22.575 69.500 23.025 ;
        RECT 68.510 12.340 68.680 22.380 ;
        RECT 69.300 12.340 69.470 22.380 ;
        RECT 68.740 11.955 69.240 12.125 ;
        RECT 69.970 11.435 70.140 23.285 ;
        RECT 67.840 11.265 70.140 11.435 ;
        RECT 70.540 23.285 72.840 23.455 ;
        RECT 70.540 11.435 70.710 23.285 ;
        RECT 71.200 22.575 72.200 23.025 ;
        RECT 71.210 12.340 71.380 22.380 ;
        RECT 72.000 12.340 72.170 22.380 ;
        RECT 71.440 11.955 71.940 12.125 ;
        RECT 72.670 11.435 72.840 23.285 ;
        RECT 70.540 11.265 72.840 11.435 ;
        RECT 48.255 9.630 49.905 9.800 ;
        RECT 57.040 10.195 59.340 10.365 ;
        RECT 48.685 9.580 49.475 9.630 ;
        RECT 57.040 9.255 57.210 10.195 ;
        RECT 57.420 9.505 58.460 9.950 ;
        RECT 57.710 9.255 57.880 9.335 ;
        RECT 57.035 8.725 57.880 9.255 ;
        RECT 57.040 7.785 57.210 8.725 ;
        RECT 57.710 8.645 57.880 8.725 ;
        RECT 58.500 8.645 58.670 9.335 ;
        RECT 57.940 8.305 58.440 8.475 ;
        RECT 59.170 7.785 59.340 10.195 ;
        RECT 57.040 7.615 59.340 7.785 ;
        RECT 59.740 10.195 62.040 10.365 ;
        RECT 45.115 1.765 47.415 1.935 ;
        RECT 59.740 1.935 59.910 10.195 ;
        RECT 60.640 9.505 61.140 9.675 ;
        RECT 60.410 2.795 60.580 9.335 ;
        RECT 61.200 2.795 61.370 9.335 ;
        RECT 60.400 2.225 61.400 2.625 ;
        RECT 61.870 1.935 62.040 10.195 ;
        RECT 62.440 10.195 64.740 10.365 ;
        RECT 62.440 9.255 62.610 10.195 ;
        RECT 62.820 9.505 63.860 9.950 ;
        RECT 63.110 9.255 63.280 9.335 ;
        RECT 62.435 8.725 63.280 9.255 ;
        RECT 62.440 7.785 62.610 8.725 ;
        RECT 63.110 8.645 63.280 8.725 ;
        RECT 63.900 8.645 64.070 9.335 ;
        RECT 63.340 8.305 63.840 8.475 ;
        RECT 64.570 7.785 64.740 10.195 ;
        RECT 65.140 10.195 67.440 10.365 ;
        RECT 65.140 9.255 65.310 10.195 ;
        RECT 65.520 9.505 66.560 9.950 ;
        RECT 65.810 9.255 65.980 9.335 ;
        RECT 65.135 8.725 65.980 9.255 ;
        RECT 62.440 7.615 64.740 7.785 ;
        RECT 65.140 7.785 65.310 8.725 ;
        RECT 65.810 8.645 65.980 8.725 ;
        RECT 66.600 8.645 66.770 9.335 ;
        RECT 66.040 8.305 66.540 8.475 ;
        RECT 67.270 7.785 67.440 10.195 ;
        RECT 65.140 7.615 67.440 7.785 ;
        RECT 67.840 10.195 70.140 10.365 ;
        RECT 59.740 1.765 62.040 1.935 ;
        RECT 67.840 1.935 68.010 10.195 ;
        RECT 68.740 9.505 69.240 9.675 ;
        RECT 68.510 2.795 68.680 9.335 ;
        RECT 69.300 2.795 69.470 9.335 ;
        RECT 68.500 2.225 69.500 2.625 ;
        RECT 69.970 1.935 70.140 10.195 ;
        RECT 67.840 1.765 70.140 1.935 ;
        RECT 70.540 10.195 72.840 10.365 ;
        RECT 70.540 1.935 70.710 10.195 ;
        RECT 71.440 9.505 71.940 9.675 ;
        RECT 71.210 2.795 71.380 9.335 ;
        RECT 72.000 2.795 72.170 9.335 ;
        RECT 71.200 2.225 72.200 2.625 ;
        RECT 72.670 1.935 72.840 10.195 ;
        RECT 73.680 9.800 73.850 23.830 ;
        RECT 74.085 23.780 74.925 23.830 ;
        RECT 74.280 21.115 74.730 23.425 ;
        RECT 74.280 10.205 74.730 12.515 ;
        RECT 74.110 9.800 74.900 9.850 ;
        RECT 75.160 9.800 75.330 23.830 ;
        RECT 99.105 23.830 100.755 24.000 ;
        RECT 85.165 23.285 87.465 23.455 ;
        RECT 82.465 14.285 84.765 14.455 ;
        RECT 82.465 13.350 82.635 14.285 ;
        RECT 83.365 13.595 83.865 13.765 ;
        RECT 83.135 13.350 83.305 13.380 ;
        RECT 82.410 12.370 83.305 13.350 ;
        RECT 82.465 11.435 82.635 12.370 ;
        RECT 83.135 12.340 83.305 12.370 ;
        RECT 83.925 12.340 84.095 13.380 ;
        RECT 82.950 11.955 83.865 12.125 ;
        RECT 82.950 11.750 83.785 11.955 ;
        RECT 84.595 11.435 84.765 14.285 ;
        RECT 82.465 11.265 84.765 11.435 ;
        RECT 85.165 11.435 85.335 23.285 ;
        RECT 85.825 22.575 86.825 23.025 ;
        RECT 85.835 12.340 86.005 22.380 ;
        RECT 86.625 12.340 86.795 22.380 ;
        RECT 86.065 11.955 86.565 12.125 ;
        RECT 87.295 11.435 87.465 23.285 ;
        RECT 93.265 23.285 95.565 23.455 ;
        RECT 87.865 14.285 90.165 14.455 ;
        RECT 87.865 13.350 88.035 14.285 ;
        RECT 88.765 13.595 89.265 13.765 ;
        RECT 88.535 13.350 88.705 13.380 ;
        RECT 87.810 12.370 88.705 13.350 ;
        RECT 85.165 11.265 87.465 11.435 ;
        RECT 87.865 11.435 88.035 12.370 ;
        RECT 88.535 12.340 88.705 12.370 ;
        RECT 89.325 12.340 89.495 13.380 ;
        RECT 88.350 11.955 89.265 12.125 ;
        RECT 88.350 11.750 89.185 11.955 ;
        RECT 89.995 11.435 90.165 14.285 ;
        RECT 90.565 14.285 92.865 14.455 ;
        RECT 90.565 13.350 90.735 14.285 ;
        RECT 91.465 13.595 91.965 13.765 ;
        RECT 91.235 13.350 91.405 13.380 ;
        RECT 90.510 12.370 91.405 13.350 ;
        RECT 87.865 11.265 90.165 11.435 ;
        RECT 90.565 11.435 90.735 12.370 ;
        RECT 91.235 12.340 91.405 12.370 ;
        RECT 92.025 12.340 92.195 13.380 ;
        RECT 91.050 11.955 91.965 12.125 ;
        RECT 91.050 11.750 91.885 11.955 ;
        RECT 92.695 11.435 92.865 14.285 ;
        RECT 90.565 11.265 92.865 11.435 ;
        RECT 93.265 11.435 93.435 23.285 ;
        RECT 93.925 22.575 94.925 23.025 ;
        RECT 93.935 12.340 94.105 22.380 ;
        RECT 94.725 12.340 94.895 22.380 ;
        RECT 94.165 11.955 94.665 12.125 ;
        RECT 95.395 11.435 95.565 23.285 ;
        RECT 93.265 11.265 95.565 11.435 ;
        RECT 95.965 23.285 98.265 23.455 ;
        RECT 95.965 11.435 96.135 23.285 ;
        RECT 96.625 22.575 97.625 23.025 ;
        RECT 96.635 12.340 96.805 22.380 ;
        RECT 97.425 12.340 97.595 22.380 ;
        RECT 96.865 11.955 97.365 12.125 ;
        RECT 98.095 11.435 98.265 23.285 ;
        RECT 95.965 11.265 98.265 11.435 ;
        RECT 73.680 9.630 75.330 9.800 ;
        RECT 82.465 10.195 84.765 10.365 ;
        RECT 74.110 9.580 74.900 9.630 ;
        RECT 82.465 9.255 82.635 10.195 ;
        RECT 82.845 9.505 83.885 9.950 ;
        RECT 83.135 9.255 83.305 9.335 ;
        RECT 82.460 8.725 83.305 9.255 ;
        RECT 82.465 7.785 82.635 8.725 ;
        RECT 83.135 8.645 83.305 8.725 ;
        RECT 83.925 8.645 84.095 9.335 ;
        RECT 83.365 8.305 83.865 8.475 ;
        RECT 84.595 7.785 84.765 10.195 ;
        RECT 82.465 7.615 84.765 7.785 ;
        RECT 85.165 10.195 87.465 10.365 ;
        RECT 70.540 1.765 72.840 1.935 ;
        RECT 85.165 1.935 85.335 10.195 ;
        RECT 86.065 9.505 86.565 9.675 ;
        RECT 85.835 2.795 86.005 9.335 ;
        RECT 86.625 2.795 86.795 9.335 ;
        RECT 85.825 2.225 86.825 2.625 ;
        RECT 87.295 1.935 87.465 10.195 ;
        RECT 87.865 10.195 90.165 10.365 ;
        RECT 87.865 9.255 88.035 10.195 ;
        RECT 88.245 9.505 89.285 9.950 ;
        RECT 88.535 9.255 88.705 9.335 ;
        RECT 87.860 8.725 88.705 9.255 ;
        RECT 87.865 7.785 88.035 8.725 ;
        RECT 88.535 8.645 88.705 8.725 ;
        RECT 89.325 8.645 89.495 9.335 ;
        RECT 88.765 8.305 89.265 8.475 ;
        RECT 89.995 7.785 90.165 10.195 ;
        RECT 90.565 10.195 92.865 10.365 ;
        RECT 90.565 9.255 90.735 10.195 ;
        RECT 90.945 9.505 91.985 9.950 ;
        RECT 91.235 9.255 91.405 9.335 ;
        RECT 90.560 8.725 91.405 9.255 ;
        RECT 87.865 7.615 90.165 7.785 ;
        RECT 90.565 7.785 90.735 8.725 ;
        RECT 91.235 8.645 91.405 8.725 ;
        RECT 92.025 8.645 92.195 9.335 ;
        RECT 91.465 8.305 91.965 8.475 ;
        RECT 92.695 7.785 92.865 10.195 ;
        RECT 90.565 7.615 92.865 7.785 ;
        RECT 93.265 10.195 95.565 10.365 ;
        RECT 85.165 1.765 87.465 1.935 ;
        RECT 93.265 1.935 93.435 10.195 ;
        RECT 94.165 9.505 94.665 9.675 ;
        RECT 93.935 2.795 94.105 9.335 ;
        RECT 94.725 2.795 94.895 9.335 ;
        RECT 93.925 2.225 94.925 2.625 ;
        RECT 95.395 1.935 95.565 10.195 ;
        RECT 93.265 1.765 95.565 1.935 ;
        RECT 95.965 10.195 98.265 10.365 ;
        RECT 95.965 1.935 96.135 10.195 ;
        RECT 96.865 9.505 97.365 9.675 ;
        RECT 96.635 2.795 96.805 9.335 ;
        RECT 97.425 2.795 97.595 9.335 ;
        RECT 96.625 2.225 97.625 2.625 ;
        RECT 98.095 1.935 98.265 10.195 ;
        RECT 99.105 9.800 99.275 23.830 ;
        RECT 99.510 23.780 100.350 23.830 ;
        RECT 99.705 21.115 100.155 23.425 ;
        RECT 99.705 10.205 100.155 12.515 ;
        RECT 99.535 9.800 100.325 9.850 ;
        RECT 100.585 9.800 100.755 23.830 ;
        RECT 124.530 23.830 126.180 24.000 ;
        RECT 110.590 23.285 112.890 23.455 ;
        RECT 107.890 14.285 110.190 14.455 ;
        RECT 107.890 13.350 108.060 14.285 ;
        RECT 108.790 13.595 109.290 13.765 ;
        RECT 108.560 13.350 108.730 13.380 ;
        RECT 107.835 12.370 108.730 13.350 ;
        RECT 107.890 11.435 108.060 12.370 ;
        RECT 108.560 12.340 108.730 12.370 ;
        RECT 109.350 12.340 109.520 13.380 ;
        RECT 108.375 11.955 109.290 12.125 ;
        RECT 108.375 11.750 109.210 11.955 ;
        RECT 110.020 11.435 110.190 14.285 ;
        RECT 107.890 11.265 110.190 11.435 ;
        RECT 110.590 11.435 110.760 23.285 ;
        RECT 111.250 22.575 112.250 23.025 ;
        RECT 111.260 12.340 111.430 22.380 ;
        RECT 112.050 12.340 112.220 22.380 ;
        RECT 111.490 11.955 111.990 12.125 ;
        RECT 112.720 11.435 112.890 23.285 ;
        RECT 118.690 23.285 120.990 23.455 ;
        RECT 113.290 14.285 115.590 14.455 ;
        RECT 113.290 13.350 113.460 14.285 ;
        RECT 114.190 13.595 114.690 13.765 ;
        RECT 113.960 13.350 114.130 13.380 ;
        RECT 113.235 12.370 114.130 13.350 ;
        RECT 110.590 11.265 112.890 11.435 ;
        RECT 113.290 11.435 113.460 12.370 ;
        RECT 113.960 12.340 114.130 12.370 ;
        RECT 114.750 12.340 114.920 13.380 ;
        RECT 113.775 11.955 114.690 12.125 ;
        RECT 113.775 11.750 114.610 11.955 ;
        RECT 115.420 11.435 115.590 14.285 ;
        RECT 115.990 14.285 118.290 14.455 ;
        RECT 115.990 13.350 116.160 14.285 ;
        RECT 116.890 13.595 117.390 13.765 ;
        RECT 116.660 13.350 116.830 13.380 ;
        RECT 115.935 12.370 116.830 13.350 ;
        RECT 113.290 11.265 115.590 11.435 ;
        RECT 115.990 11.435 116.160 12.370 ;
        RECT 116.660 12.340 116.830 12.370 ;
        RECT 117.450 12.340 117.620 13.380 ;
        RECT 116.475 11.955 117.390 12.125 ;
        RECT 116.475 11.750 117.310 11.955 ;
        RECT 118.120 11.435 118.290 14.285 ;
        RECT 115.990 11.265 118.290 11.435 ;
        RECT 118.690 11.435 118.860 23.285 ;
        RECT 119.350 22.575 120.350 23.025 ;
        RECT 119.360 12.340 119.530 22.380 ;
        RECT 120.150 12.340 120.320 22.380 ;
        RECT 119.590 11.955 120.090 12.125 ;
        RECT 120.820 11.435 120.990 23.285 ;
        RECT 118.690 11.265 120.990 11.435 ;
        RECT 121.390 23.285 123.690 23.455 ;
        RECT 121.390 11.435 121.560 23.285 ;
        RECT 122.050 22.575 123.050 23.025 ;
        RECT 122.060 12.340 122.230 22.380 ;
        RECT 122.850 12.340 123.020 22.380 ;
        RECT 122.290 11.955 122.790 12.125 ;
        RECT 123.520 11.435 123.690 23.285 ;
        RECT 121.390 11.265 123.690 11.435 ;
        RECT 99.105 9.630 100.755 9.800 ;
        RECT 107.890 10.195 110.190 10.365 ;
        RECT 99.535 9.580 100.325 9.630 ;
        RECT 107.890 9.255 108.060 10.195 ;
        RECT 108.270 9.505 109.310 9.950 ;
        RECT 108.560 9.255 108.730 9.335 ;
        RECT 107.885 8.725 108.730 9.255 ;
        RECT 107.890 7.785 108.060 8.725 ;
        RECT 108.560 8.645 108.730 8.725 ;
        RECT 109.350 8.645 109.520 9.335 ;
        RECT 108.790 8.305 109.290 8.475 ;
        RECT 110.020 7.785 110.190 10.195 ;
        RECT 107.890 7.615 110.190 7.785 ;
        RECT 110.590 10.195 112.890 10.365 ;
        RECT 95.965 1.765 98.265 1.935 ;
        RECT 110.590 1.935 110.760 10.195 ;
        RECT 111.490 9.505 111.990 9.675 ;
        RECT 111.260 2.795 111.430 9.335 ;
        RECT 112.050 2.795 112.220 9.335 ;
        RECT 111.250 2.225 112.250 2.625 ;
        RECT 112.720 1.935 112.890 10.195 ;
        RECT 113.290 10.195 115.590 10.365 ;
        RECT 113.290 9.255 113.460 10.195 ;
        RECT 113.670 9.505 114.710 9.950 ;
        RECT 113.960 9.255 114.130 9.335 ;
        RECT 113.285 8.725 114.130 9.255 ;
        RECT 113.290 7.785 113.460 8.725 ;
        RECT 113.960 8.645 114.130 8.725 ;
        RECT 114.750 8.645 114.920 9.335 ;
        RECT 114.190 8.305 114.690 8.475 ;
        RECT 115.420 7.785 115.590 10.195 ;
        RECT 115.990 10.195 118.290 10.365 ;
        RECT 115.990 9.255 116.160 10.195 ;
        RECT 116.370 9.505 117.410 9.950 ;
        RECT 116.660 9.255 116.830 9.335 ;
        RECT 115.985 8.725 116.830 9.255 ;
        RECT 113.290 7.615 115.590 7.785 ;
        RECT 115.990 7.785 116.160 8.725 ;
        RECT 116.660 8.645 116.830 8.725 ;
        RECT 117.450 8.645 117.620 9.335 ;
        RECT 116.890 8.305 117.390 8.475 ;
        RECT 118.120 7.785 118.290 10.195 ;
        RECT 115.990 7.615 118.290 7.785 ;
        RECT 118.690 10.195 120.990 10.365 ;
        RECT 110.590 1.765 112.890 1.935 ;
        RECT 118.690 1.935 118.860 10.195 ;
        RECT 119.590 9.505 120.090 9.675 ;
        RECT 119.360 2.795 119.530 9.335 ;
        RECT 120.150 2.795 120.320 9.335 ;
        RECT 119.350 2.225 120.350 2.625 ;
        RECT 120.820 1.935 120.990 10.195 ;
        RECT 118.690 1.765 120.990 1.935 ;
        RECT 121.390 10.195 123.690 10.365 ;
        RECT 121.390 1.935 121.560 10.195 ;
        RECT 122.290 9.505 122.790 9.675 ;
        RECT 122.060 2.795 122.230 9.335 ;
        RECT 122.850 2.795 123.020 9.335 ;
        RECT 122.050 2.225 123.050 2.625 ;
        RECT 123.520 1.935 123.690 10.195 ;
        RECT 124.530 9.800 124.700 23.830 ;
        RECT 124.935 23.780 125.775 23.830 ;
        RECT 125.130 21.115 125.580 23.425 ;
        RECT 125.130 10.205 125.580 12.515 ;
        RECT 124.960 9.800 125.750 9.850 ;
        RECT 126.010 9.800 126.180 23.830 ;
        RECT 149.955 23.830 151.605 24.000 ;
        RECT 136.015 23.285 138.315 23.455 ;
        RECT 133.315 14.285 135.615 14.455 ;
        RECT 133.315 13.350 133.485 14.285 ;
        RECT 134.215 13.595 134.715 13.765 ;
        RECT 133.985 13.350 134.155 13.380 ;
        RECT 133.260 12.370 134.155 13.350 ;
        RECT 133.315 11.435 133.485 12.370 ;
        RECT 133.985 12.340 134.155 12.370 ;
        RECT 134.775 12.340 134.945 13.380 ;
        RECT 133.800 11.955 134.715 12.125 ;
        RECT 133.800 11.750 134.635 11.955 ;
        RECT 135.445 11.435 135.615 14.285 ;
        RECT 133.315 11.265 135.615 11.435 ;
        RECT 136.015 11.435 136.185 23.285 ;
        RECT 136.675 22.575 137.675 23.025 ;
        RECT 136.685 12.340 136.855 22.380 ;
        RECT 137.475 12.340 137.645 22.380 ;
        RECT 136.915 11.955 137.415 12.125 ;
        RECT 138.145 11.435 138.315 23.285 ;
        RECT 144.115 23.285 146.415 23.455 ;
        RECT 138.715 14.285 141.015 14.455 ;
        RECT 138.715 13.350 138.885 14.285 ;
        RECT 139.615 13.595 140.115 13.765 ;
        RECT 139.385 13.350 139.555 13.380 ;
        RECT 138.660 12.370 139.555 13.350 ;
        RECT 136.015 11.265 138.315 11.435 ;
        RECT 138.715 11.435 138.885 12.370 ;
        RECT 139.385 12.340 139.555 12.370 ;
        RECT 140.175 12.340 140.345 13.380 ;
        RECT 139.200 11.955 140.115 12.125 ;
        RECT 139.200 11.750 140.035 11.955 ;
        RECT 140.845 11.435 141.015 14.285 ;
        RECT 141.415 14.285 143.715 14.455 ;
        RECT 141.415 13.350 141.585 14.285 ;
        RECT 142.315 13.595 142.815 13.765 ;
        RECT 142.085 13.350 142.255 13.380 ;
        RECT 141.360 12.370 142.255 13.350 ;
        RECT 138.715 11.265 141.015 11.435 ;
        RECT 141.415 11.435 141.585 12.370 ;
        RECT 142.085 12.340 142.255 12.370 ;
        RECT 142.875 12.340 143.045 13.380 ;
        RECT 141.900 11.955 142.815 12.125 ;
        RECT 141.900 11.750 142.735 11.955 ;
        RECT 143.545 11.435 143.715 14.285 ;
        RECT 141.415 11.265 143.715 11.435 ;
        RECT 144.115 11.435 144.285 23.285 ;
        RECT 144.775 22.575 145.775 23.025 ;
        RECT 144.785 12.340 144.955 22.380 ;
        RECT 145.575 12.340 145.745 22.380 ;
        RECT 145.015 11.955 145.515 12.125 ;
        RECT 146.245 11.435 146.415 23.285 ;
        RECT 144.115 11.265 146.415 11.435 ;
        RECT 146.815 23.285 149.115 23.455 ;
        RECT 146.815 11.435 146.985 23.285 ;
        RECT 147.475 22.575 148.475 23.025 ;
        RECT 147.485 12.340 147.655 22.380 ;
        RECT 148.275 12.340 148.445 22.380 ;
        RECT 147.715 11.955 148.215 12.125 ;
        RECT 148.945 11.435 149.115 23.285 ;
        RECT 146.815 11.265 149.115 11.435 ;
        RECT 124.530 9.630 126.180 9.800 ;
        RECT 133.315 10.195 135.615 10.365 ;
        RECT 124.960 9.580 125.750 9.630 ;
        RECT 133.315 9.255 133.485 10.195 ;
        RECT 133.695 9.505 134.735 9.950 ;
        RECT 133.985 9.255 134.155 9.335 ;
        RECT 133.310 8.725 134.155 9.255 ;
        RECT 133.315 7.785 133.485 8.725 ;
        RECT 133.985 8.645 134.155 8.725 ;
        RECT 134.775 8.645 134.945 9.335 ;
        RECT 134.215 8.305 134.715 8.475 ;
        RECT 135.445 7.785 135.615 10.195 ;
        RECT 133.315 7.615 135.615 7.785 ;
        RECT 136.015 10.195 138.315 10.365 ;
        RECT 121.390 1.765 123.690 1.935 ;
        RECT 136.015 1.935 136.185 10.195 ;
        RECT 136.915 9.505 137.415 9.675 ;
        RECT 136.685 2.795 136.855 9.335 ;
        RECT 137.475 2.795 137.645 9.335 ;
        RECT 136.675 2.225 137.675 2.625 ;
        RECT 138.145 1.935 138.315 10.195 ;
        RECT 138.715 10.195 141.015 10.365 ;
        RECT 138.715 9.255 138.885 10.195 ;
        RECT 139.095 9.505 140.135 9.950 ;
        RECT 139.385 9.255 139.555 9.335 ;
        RECT 138.710 8.725 139.555 9.255 ;
        RECT 138.715 7.785 138.885 8.725 ;
        RECT 139.385 8.645 139.555 8.725 ;
        RECT 140.175 8.645 140.345 9.335 ;
        RECT 139.615 8.305 140.115 8.475 ;
        RECT 140.845 7.785 141.015 10.195 ;
        RECT 141.415 10.195 143.715 10.365 ;
        RECT 141.415 9.255 141.585 10.195 ;
        RECT 141.795 9.505 142.835 9.950 ;
        RECT 142.085 9.255 142.255 9.335 ;
        RECT 141.410 8.725 142.255 9.255 ;
        RECT 138.715 7.615 141.015 7.785 ;
        RECT 141.415 7.785 141.585 8.725 ;
        RECT 142.085 8.645 142.255 8.725 ;
        RECT 142.875 8.645 143.045 9.335 ;
        RECT 142.315 8.305 142.815 8.475 ;
        RECT 143.545 7.785 143.715 10.195 ;
        RECT 141.415 7.615 143.715 7.785 ;
        RECT 144.115 10.195 146.415 10.365 ;
        RECT 136.015 1.765 138.315 1.935 ;
        RECT 144.115 1.935 144.285 10.195 ;
        RECT 145.015 9.505 145.515 9.675 ;
        RECT 144.785 2.795 144.955 9.335 ;
        RECT 145.575 2.795 145.745 9.335 ;
        RECT 144.775 2.225 145.775 2.625 ;
        RECT 146.245 1.935 146.415 10.195 ;
        RECT 144.115 1.765 146.415 1.935 ;
        RECT 146.815 10.195 149.115 10.365 ;
        RECT 146.815 1.935 146.985 10.195 ;
        RECT 147.715 9.505 148.215 9.675 ;
        RECT 147.485 2.795 147.655 9.335 ;
        RECT 148.275 2.795 148.445 9.335 ;
        RECT 147.475 2.225 148.475 2.625 ;
        RECT 148.945 1.935 149.115 10.195 ;
        RECT 149.955 9.800 150.125 23.830 ;
        RECT 150.360 23.780 151.200 23.830 ;
        RECT 150.555 21.115 151.005 23.425 ;
        RECT 150.555 10.205 151.005 12.515 ;
        RECT 150.385 9.800 151.175 9.850 ;
        RECT 151.435 9.800 151.605 23.830 ;
        RECT 149.955 9.630 151.605 9.800 ;
        RECT 150.385 9.580 151.175 9.630 ;
        RECT 146.815 1.765 149.115 1.935 ;
      LAYER met1 ;
        RECT 35.200 225.300 36.200 225.330 ;
        RECT 86.050 225.300 87.050 225.330 ;
        RECT 136.900 225.300 137.900 225.330 ;
        RECT 2.560 224.300 157.545 225.300 ;
        RECT 35.200 224.270 36.200 224.300 ;
        RECT 86.050 224.270 87.050 224.300 ;
        RECT 136.900 224.270 137.900 224.300 ;
        RECT 33.200 223.550 34.200 223.580 ;
        RECT 84.050 223.550 85.050 223.580 ;
        RECT 134.900 223.550 135.900 223.580 ;
        RECT 2.560 222.550 157.545 223.550 ;
        RECT 33.200 222.520 34.200 222.550 ;
        RECT 84.050 222.520 85.050 222.550 ;
        RECT 134.900 222.520 135.900 222.550 ;
        RECT 31.200 221.800 32.200 221.830 ;
        RECT 82.050 221.800 83.050 221.830 ;
        RECT 132.900 221.800 133.900 221.830 ;
        RECT 2.560 220.800 157.545 221.800 ;
        RECT 31.200 220.770 32.200 220.800 ;
        RECT 82.050 220.770 83.050 220.800 ;
        RECT 132.900 220.770 133.900 220.800 ;
        RECT 9.775 220.050 10.775 220.080 ;
        RECT 60.625 220.050 61.625 220.080 ;
        RECT 111.475 220.050 112.475 220.080 ;
        RECT 128.775 220.050 129.775 220.080 ;
        RECT 2.560 219.050 157.545 220.050 ;
        RECT 9.775 219.020 10.775 219.050 ;
        RECT 60.625 219.020 61.625 219.050 ;
        RECT 111.475 219.020 112.475 219.050 ;
        RECT 128.775 219.020 129.775 219.050 ;
        RECT 7.775 218.300 8.775 218.330 ;
        RECT 58.625 218.300 59.625 218.330 ;
        RECT 109.475 218.300 110.475 218.330 ;
        RECT 125.075 218.300 126.075 218.330 ;
        RECT 2.560 217.300 157.545 218.300 ;
        RECT 7.775 217.270 8.775 217.300 ;
        RECT 58.625 217.270 59.625 217.300 ;
        RECT 109.475 217.270 110.475 217.300 ;
        RECT 125.075 217.270 126.075 217.300 ;
        RECT 5.775 216.550 6.775 216.580 ;
        RECT 56.625 216.550 57.625 216.580 ;
        RECT 107.475 216.550 108.475 216.580 ;
        RECT 121.425 216.550 122.425 216.580 ;
        RECT 2.580 215.550 157.545 216.550 ;
        RECT 5.775 215.520 6.775 215.550 ;
        RECT 56.625 215.520 57.625 215.550 ;
        RECT 107.475 215.520 108.475 215.550 ;
        RECT 121.425 215.520 122.425 215.550 ;
        RECT 7.500 213.550 153.425 214.550 ;
        RECT 11.725 212.175 12.725 212.205 ;
        RECT 15.400 212.175 16.400 212.205 ;
        RECT 37.150 212.175 38.150 212.205 ;
        RECT 40.825 212.175 41.825 212.205 ;
        RECT 9.550 211.725 10.550 212.175 ;
        RECT 9.810 211.715 10.270 211.725 ;
        RECT 8.790 209.120 9.160 210.225 ;
        RECT 9.530 206.500 9.760 211.510 ;
        RECT 10.320 206.500 10.550 211.510 ;
        RECT 11.725 211.145 13.650 212.175 ;
        RECT 10.920 210.175 11.290 210.225 ;
        RECT 10.920 209.120 12.025 210.175 ;
        RECT 7.110 202.715 7.570 202.945 ;
        RECT 6.830 202.500 7.060 202.510 ;
        RECT 7.620 202.500 7.850 202.510 ;
        RECT 6.085 201.520 7.130 202.500 ;
        RECT 7.550 201.520 7.920 202.500 ;
        RECT 9.460 201.520 9.830 206.500 ;
        RECT 10.250 201.520 10.620 206.500 ;
        RECT 11.025 204.425 12.025 209.120 ;
        RECT 12.650 206.075 13.650 211.145 ;
        RECT 14.450 211.145 16.400 212.175 ;
        RECT 17.650 211.725 18.650 212.175 ;
        RECT 20.350 211.725 21.350 212.175 ;
        RECT 27.270 211.975 28.270 212.125 ;
        RECT 17.910 211.715 18.370 211.725 ;
        RECT 20.610 211.715 21.070 211.725 ;
        RECT 23.805 211.715 24.265 211.945 ;
        RECT 26.505 211.715 26.965 211.945 ;
        RECT 27.120 211.525 28.270 211.975 ;
        RECT 29.205 211.715 29.665 211.945 ;
        RECT 34.975 211.725 35.975 212.175 ;
        RECT 35.235 211.715 35.695 211.725 ;
        RECT 14.450 206.820 15.450 211.145 ;
        RECT 16.890 210.175 17.260 210.225 ;
        RECT 16.175 209.120 17.260 210.175 ;
        RECT 12.650 205.075 15.480 206.075 ;
        RECT 16.175 204.425 17.175 209.120 ;
        RECT 17.630 206.500 17.860 211.510 ;
        RECT 18.420 206.500 18.650 211.510 ;
        RECT 19.020 209.120 19.390 210.225 ;
        RECT 19.590 209.120 19.960 210.225 ;
        RECT 20.330 206.500 20.560 211.510 ;
        RECT 21.120 206.500 21.350 211.510 ;
        RECT 23.525 210.510 23.755 211.510 ;
        RECT 24.295 210.495 26.475 211.525 ;
        RECT 26.970 211.500 28.270 211.525 ;
        RECT 28.925 211.500 29.155 211.510 ;
        RECT 29.715 211.500 29.945 211.510 ;
        RECT 26.970 210.975 29.225 211.500 ;
        RECT 26.970 210.570 27.890 210.975 ;
        RECT 27.015 210.510 27.245 210.570 ;
        RECT 28.180 210.520 29.225 210.975 ;
        RECT 29.645 210.520 30.015 211.500 ;
        RECT 28.925 210.510 29.155 210.520 ;
        RECT 29.715 210.510 29.945 210.520 ;
        RECT 21.720 209.120 22.090 210.225 ;
        RECT 23.520 207.625 24.520 210.355 ;
        RECT 26.245 207.625 27.245 210.325 ;
        RECT 28.670 209.850 29.705 210.325 ;
        RECT 34.215 209.120 34.585 210.225 ;
        RECT 28.665 207.605 29.705 208.100 ;
        RECT 23.205 206.800 23.850 207.480 ;
        RECT 24.245 206.800 26.525 207.480 ;
        RECT 27.015 207.405 27.245 207.465 ;
        RECT 28.925 207.455 29.155 207.465 ;
        RECT 29.715 207.455 29.945 207.465 ;
        RECT 26.970 207.250 27.890 207.405 ;
        RECT 28.180 207.250 29.225 207.455 ;
        RECT 26.970 206.825 29.225 207.250 ;
        RECT 29.645 206.825 30.015 207.455 ;
        RECT 27.015 206.815 28.270 206.825 ;
        RECT 28.925 206.815 29.155 206.825 ;
        RECT 29.715 206.815 29.945 206.825 ;
        RECT 27.020 206.800 28.270 206.815 ;
        RECT 11.025 203.425 17.175 204.425 ;
        RECT 12.510 202.715 12.970 202.945 ;
        RECT 15.210 202.715 15.670 202.945 ;
        RECT 12.230 202.500 12.460 202.510 ;
        RECT 13.020 202.500 13.250 202.510 ;
        RECT 14.930 202.500 15.160 202.510 ;
        RECT 15.720 202.500 15.950 202.510 ;
        RECT 11.485 201.520 12.530 202.500 ;
        RECT 12.950 201.520 13.320 202.500 ;
        RECT 14.185 201.520 15.230 202.500 ;
        RECT 15.650 201.520 16.020 202.500 ;
        RECT 17.560 201.520 17.930 206.500 ;
        RECT 18.350 201.520 18.720 206.500 ;
        RECT 20.260 201.520 20.630 206.500 ;
        RECT 21.050 201.520 21.420 206.500 ;
        RECT 23.805 206.425 24.265 206.655 ;
        RECT 26.505 206.425 26.965 206.655 ;
        RECT 27.115 206.250 28.270 206.800 ;
        RECT 29.205 206.425 29.665 206.655 ;
        RECT 34.955 206.500 35.185 211.510 ;
        RECT 35.745 206.500 35.975 211.510 ;
        RECT 37.150 211.145 39.075 212.175 ;
        RECT 36.345 210.175 36.715 210.225 ;
        RECT 36.345 209.120 37.450 210.175 ;
        RECT 27.115 206.200 28.175 206.250 ;
        RECT 6.830 201.510 7.060 201.520 ;
        RECT 7.620 201.510 7.850 201.520 ;
        RECT 9.530 201.510 9.760 201.520 ;
        RECT 10.320 201.510 10.550 201.520 ;
        RECT 12.230 201.510 12.460 201.520 ;
        RECT 13.020 201.510 13.250 201.520 ;
        RECT 14.930 201.510 15.160 201.520 ;
        RECT 15.720 201.510 15.950 201.520 ;
        RECT 17.630 201.510 17.860 201.520 ;
        RECT 18.420 201.510 18.650 201.520 ;
        RECT 20.330 201.510 20.560 201.520 ;
        RECT 21.120 201.510 21.350 201.520 ;
        RECT 6.575 200.850 7.610 201.325 ;
        RECT 9.810 201.075 10.270 201.305 ;
        RECT 11.975 200.850 13.010 201.325 ;
        RECT 14.675 200.850 15.710 201.325 ;
        RECT 17.910 201.075 18.370 201.305 ;
        RECT 20.610 201.075 21.070 201.305 ;
        RECT 3.950 200.475 4.950 200.530 ;
        RECT 24.820 200.510 25.925 205.180 ;
        RECT 32.535 202.715 32.995 202.945 ;
        RECT 32.255 202.500 32.485 202.510 ;
        RECT 33.045 202.500 33.275 202.510 ;
        RECT 31.510 201.520 32.555 202.500 ;
        RECT 32.975 201.520 33.345 202.500 ;
        RECT 34.885 201.520 35.255 206.500 ;
        RECT 35.675 201.520 36.045 206.500 ;
        RECT 36.450 204.425 37.450 209.120 ;
        RECT 38.075 206.075 39.075 211.145 ;
        RECT 39.875 211.145 41.825 212.175 ;
        RECT 43.075 211.725 44.075 212.175 ;
        RECT 45.775 211.725 46.775 212.175 ;
        RECT 43.335 211.715 43.795 211.725 ;
        RECT 46.035 211.715 46.495 211.725 ;
        RECT 39.875 206.820 40.875 211.145 ;
        RECT 42.315 210.175 42.685 210.225 ;
        RECT 41.600 209.120 42.685 210.175 ;
        RECT 38.075 205.075 40.905 206.075 ;
        RECT 41.600 204.425 42.600 209.120 ;
        RECT 43.055 206.500 43.285 211.510 ;
        RECT 43.845 206.500 44.075 211.510 ;
        RECT 44.445 209.120 44.815 210.225 ;
        RECT 45.015 209.120 45.385 210.225 ;
        RECT 45.755 206.500 45.985 211.510 ;
        RECT 46.545 206.500 46.775 211.510 ;
        RECT 47.145 209.120 47.515 210.225 ;
        RECT 36.450 203.425 42.600 204.425 ;
        RECT 37.935 202.715 38.395 202.945 ;
        RECT 40.635 202.715 41.095 202.945 ;
        RECT 37.655 202.500 37.885 202.510 ;
        RECT 38.445 202.500 38.675 202.510 ;
        RECT 40.355 202.500 40.585 202.510 ;
        RECT 41.145 202.500 41.375 202.510 ;
        RECT 36.910 201.520 37.955 202.500 ;
        RECT 38.375 201.520 38.745 202.500 ;
        RECT 39.610 201.520 40.655 202.500 ;
        RECT 41.075 201.520 41.445 202.500 ;
        RECT 42.985 201.520 43.355 206.500 ;
        RECT 43.775 201.520 44.145 206.500 ;
        RECT 45.685 201.520 46.055 206.500 ;
        RECT 46.475 201.520 46.845 206.500 ;
        RECT 32.255 201.510 32.485 201.520 ;
        RECT 33.045 201.510 33.275 201.520 ;
        RECT 34.955 201.510 35.185 201.520 ;
        RECT 35.745 201.510 35.975 201.520 ;
        RECT 37.655 201.510 37.885 201.520 ;
        RECT 38.445 201.510 38.675 201.520 ;
        RECT 40.355 201.510 40.585 201.520 ;
        RECT 41.145 201.510 41.375 201.520 ;
        RECT 43.055 201.510 43.285 201.520 ;
        RECT 43.845 201.510 44.075 201.520 ;
        RECT 45.755 201.510 45.985 201.520 ;
        RECT 46.545 201.510 46.775 201.520 ;
        RECT 32.000 200.850 33.035 201.325 ;
        RECT 35.235 201.075 35.695 201.305 ;
        RECT 37.400 200.850 38.435 201.325 ;
        RECT 40.100 200.850 41.135 201.325 ;
        RECT 43.335 201.075 43.795 201.305 ;
        RECT 46.035 201.075 46.495 201.305 ;
        RECT 29.375 200.510 30.375 200.530 ;
        RECT 3.920 199.475 4.980 200.475 ;
        RECT 3.950 196.250 4.950 199.475 ;
        RECT 24.820 199.405 30.430 200.510 ;
        RECT 50.725 200.475 51.725 213.550 ;
        RECT 62.575 212.175 63.575 212.205 ;
        RECT 66.250 212.175 67.250 212.205 ;
        RECT 88.000 212.175 89.000 212.205 ;
        RECT 91.675 212.175 92.675 212.205 ;
        RECT 60.400 211.725 61.400 212.175 ;
        RECT 60.660 211.715 61.120 211.725 ;
        RECT 59.640 209.120 60.010 210.225 ;
        RECT 60.380 206.500 60.610 211.510 ;
        RECT 61.170 206.500 61.400 211.510 ;
        RECT 62.575 211.145 64.500 212.175 ;
        RECT 61.770 210.175 62.140 210.225 ;
        RECT 61.770 209.120 62.875 210.175 ;
        RECT 57.960 202.715 58.420 202.945 ;
        RECT 57.680 202.500 57.910 202.510 ;
        RECT 58.470 202.500 58.700 202.510 ;
        RECT 56.935 201.520 57.980 202.500 ;
        RECT 58.400 201.520 58.770 202.500 ;
        RECT 60.310 201.520 60.680 206.500 ;
        RECT 61.100 201.520 61.470 206.500 ;
        RECT 61.875 204.425 62.875 209.120 ;
        RECT 63.500 206.075 64.500 211.145 ;
        RECT 65.300 211.145 67.250 212.175 ;
        RECT 68.500 211.725 69.500 212.175 ;
        RECT 71.200 211.725 72.200 212.175 ;
        RECT 78.120 211.975 79.120 212.125 ;
        RECT 68.760 211.715 69.220 211.725 ;
        RECT 71.460 211.715 71.920 211.725 ;
        RECT 74.655 211.715 75.115 211.945 ;
        RECT 77.355 211.715 77.815 211.945 ;
        RECT 77.970 211.525 79.120 211.975 ;
        RECT 80.055 211.715 80.515 211.945 ;
        RECT 85.825 211.725 86.825 212.175 ;
        RECT 86.085 211.715 86.545 211.725 ;
        RECT 65.300 206.820 66.300 211.145 ;
        RECT 67.740 210.175 68.110 210.225 ;
        RECT 67.025 209.120 68.110 210.175 ;
        RECT 63.500 205.075 66.330 206.075 ;
        RECT 67.025 204.425 68.025 209.120 ;
        RECT 68.480 206.500 68.710 211.510 ;
        RECT 69.270 206.500 69.500 211.510 ;
        RECT 69.870 209.120 70.240 210.225 ;
        RECT 70.440 209.120 70.810 210.225 ;
        RECT 71.180 206.500 71.410 211.510 ;
        RECT 71.970 206.500 72.200 211.510 ;
        RECT 74.375 210.510 74.605 211.510 ;
        RECT 75.145 210.495 77.325 211.525 ;
        RECT 77.820 211.500 79.120 211.525 ;
        RECT 79.775 211.500 80.005 211.510 ;
        RECT 80.565 211.500 80.795 211.510 ;
        RECT 77.820 210.975 80.075 211.500 ;
        RECT 77.820 210.570 78.740 210.975 ;
        RECT 77.865 210.510 78.095 210.570 ;
        RECT 79.030 210.520 80.075 210.975 ;
        RECT 80.495 210.520 80.865 211.500 ;
        RECT 79.775 210.510 80.005 210.520 ;
        RECT 80.565 210.510 80.795 210.520 ;
        RECT 72.570 209.120 72.940 210.225 ;
        RECT 74.370 207.625 75.370 210.355 ;
        RECT 77.095 207.625 78.095 210.325 ;
        RECT 79.520 209.850 80.555 210.325 ;
        RECT 85.065 209.120 85.435 210.225 ;
        RECT 79.515 207.605 80.555 208.100 ;
        RECT 74.055 206.800 74.700 207.480 ;
        RECT 75.095 206.800 77.375 207.480 ;
        RECT 77.865 207.405 78.095 207.465 ;
        RECT 79.775 207.455 80.005 207.465 ;
        RECT 80.565 207.455 80.795 207.465 ;
        RECT 77.820 207.250 78.740 207.405 ;
        RECT 79.030 207.250 80.075 207.455 ;
        RECT 77.820 206.825 80.075 207.250 ;
        RECT 80.495 206.825 80.865 207.455 ;
        RECT 77.865 206.815 79.120 206.825 ;
        RECT 79.775 206.815 80.005 206.825 ;
        RECT 80.565 206.815 80.795 206.825 ;
        RECT 77.870 206.800 79.120 206.815 ;
        RECT 61.875 203.425 68.025 204.425 ;
        RECT 63.360 202.715 63.820 202.945 ;
        RECT 66.060 202.715 66.520 202.945 ;
        RECT 63.080 202.500 63.310 202.510 ;
        RECT 63.870 202.500 64.100 202.510 ;
        RECT 65.780 202.500 66.010 202.510 ;
        RECT 66.570 202.500 66.800 202.510 ;
        RECT 62.335 201.520 63.380 202.500 ;
        RECT 63.800 201.520 64.170 202.500 ;
        RECT 65.035 201.520 66.080 202.500 ;
        RECT 66.500 201.520 66.870 202.500 ;
        RECT 68.410 201.520 68.780 206.500 ;
        RECT 69.200 201.520 69.570 206.500 ;
        RECT 71.110 201.520 71.480 206.500 ;
        RECT 71.900 201.520 72.270 206.500 ;
        RECT 74.655 206.425 75.115 206.655 ;
        RECT 77.355 206.425 77.815 206.655 ;
        RECT 77.965 206.250 79.120 206.800 ;
        RECT 80.055 206.425 80.515 206.655 ;
        RECT 85.805 206.500 86.035 211.510 ;
        RECT 86.595 206.500 86.825 211.510 ;
        RECT 88.000 211.145 89.925 212.175 ;
        RECT 87.195 210.175 87.565 210.225 ;
        RECT 87.195 209.120 88.300 210.175 ;
        RECT 77.965 206.200 79.025 206.250 ;
        RECT 57.680 201.510 57.910 201.520 ;
        RECT 58.470 201.510 58.700 201.520 ;
        RECT 60.380 201.510 60.610 201.520 ;
        RECT 61.170 201.510 61.400 201.520 ;
        RECT 63.080 201.510 63.310 201.520 ;
        RECT 63.870 201.510 64.100 201.520 ;
        RECT 65.780 201.510 66.010 201.520 ;
        RECT 66.570 201.510 66.800 201.520 ;
        RECT 68.480 201.510 68.710 201.520 ;
        RECT 69.270 201.510 69.500 201.520 ;
        RECT 71.180 201.510 71.410 201.520 ;
        RECT 71.970 201.510 72.200 201.520 ;
        RECT 57.425 200.850 58.460 201.325 ;
        RECT 60.660 201.075 61.120 201.305 ;
        RECT 62.825 200.850 63.860 201.325 ;
        RECT 65.525 200.850 66.560 201.325 ;
        RECT 68.760 201.075 69.220 201.305 ;
        RECT 71.460 201.075 71.920 201.305 ;
        RECT 54.800 200.475 55.800 200.530 ;
        RECT 75.670 200.510 76.775 205.180 ;
        RECT 83.385 202.715 83.845 202.945 ;
        RECT 83.105 202.500 83.335 202.510 ;
        RECT 83.895 202.500 84.125 202.510 ;
        RECT 82.360 201.520 83.405 202.500 ;
        RECT 83.825 201.520 84.195 202.500 ;
        RECT 85.735 201.520 86.105 206.500 ;
        RECT 86.525 201.520 86.895 206.500 ;
        RECT 87.300 204.425 88.300 209.120 ;
        RECT 88.925 206.075 89.925 211.145 ;
        RECT 90.725 211.145 92.675 212.175 ;
        RECT 93.925 211.725 94.925 212.175 ;
        RECT 96.625 211.725 97.625 212.175 ;
        RECT 94.185 211.715 94.645 211.725 ;
        RECT 96.885 211.715 97.345 211.725 ;
        RECT 90.725 206.820 91.725 211.145 ;
        RECT 93.165 210.175 93.535 210.225 ;
        RECT 92.450 209.120 93.535 210.175 ;
        RECT 88.925 205.075 91.755 206.075 ;
        RECT 92.450 204.425 93.450 209.120 ;
        RECT 93.905 206.500 94.135 211.510 ;
        RECT 94.695 206.500 94.925 211.510 ;
        RECT 95.295 209.120 95.665 210.225 ;
        RECT 95.865 209.120 96.235 210.225 ;
        RECT 96.605 206.500 96.835 211.510 ;
        RECT 97.395 206.500 97.625 211.510 ;
        RECT 97.995 209.120 98.365 210.225 ;
        RECT 87.300 203.425 93.450 204.425 ;
        RECT 88.785 202.715 89.245 202.945 ;
        RECT 91.485 202.715 91.945 202.945 ;
        RECT 88.505 202.500 88.735 202.510 ;
        RECT 89.295 202.500 89.525 202.510 ;
        RECT 91.205 202.500 91.435 202.510 ;
        RECT 91.995 202.500 92.225 202.510 ;
        RECT 87.760 201.520 88.805 202.500 ;
        RECT 89.225 201.520 89.595 202.500 ;
        RECT 90.460 201.520 91.505 202.500 ;
        RECT 91.925 201.520 92.295 202.500 ;
        RECT 93.835 201.520 94.205 206.500 ;
        RECT 94.625 201.520 94.995 206.500 ;
        RECT 96.535 201.520 96.905 206.500 ;
        RECT 97.325 201.520 97.695 206.500 ;
        RECT 83.105 201.510 83.335 201.520 ;
        RECT 83.895 201.510 84.125 201.520 ;
        RECT 85.805 201.510 86.035 201.520 ;
        RECT 86.595 201.510 86.825 201.520 ;
        RECT 88.505 201.510 88.735 201.520 ;
        RECT 89.295 201.510 89.525 201.520 ;
        RECT 91.205 201.510 91.435 201.520 ;
        RECT 91.995 201.510 92.225 201.520 ;
        RECT 93.905 201.510 94.135 201.520 ;
        RECT 94.695 201.510 94.925 201.520 ;
        RECT 96.605 201.510 96.835 201.520 ;
        RECT 97.395 201.510 97.625 201.520 ;
        RECT 82.850 200.850 83.885 201.325 ;
        RECT 86.085 201.075 86.545 201.305 ;
        RECT 88.250 200.850 89.285 201.325 ;
        RECT 90.950 200.850 91.985 201.325 ;
        RECT 94.185 201.075 94.645 201.305 ;
        RECT 96.885 201.075 97.345 201.305 ;
        RECT 80.225 200.510 81.225 200.530 ;
        RECT 50.695 199.475 51.755 200.475 ;
        RECT 54.770 199.475 55.830 200.475 ;
        RECT 6.570 198.605 7.610 199.100 ;
        RECT 9.810 198.625 10.270 198.855 ;
        RECT 11.970 198.605 13.010 199.100 ;
        RECT 14.670 198.605 15.710 199.100 ;
        RECT 17.910 198.625 18.370 198.855 ;
        RECT 20.610 198.625 21.070 198.855 ;
        RECT 6.830 198.455 7.060 198.465 ;
        RECT 7.620 198.455 7.850 198.465 ;
        RECT 9.530 198.455 9.760 198.465 ;
        RECT 10.320 198.455 10.550 198.465 ;
        RECT 12.230 198.455 12.460 198.465 ;
        RECT 13.020 198.455 13.250 198.465 ;
        RECT 14.930 198.455 15.160 198.465 ;
        RECT 15.720 198.455 15.950 198.465 ;
        RECT 17.630 198.455 17.860 198.465 ;
        RECT 18.420 198.455 18.650 198.465 ;
        RECT 20.330 198.455 20.560 198.465 ;
        RECT 21.120 198.455 21.350 198.465 ;
        RECT 6.085 197.825 7.130 198.455 ;
        RECT 7.550 197.825 7.920 198.455 ;
        RECT 6.830 197.815 7.060 197.825 ;
        RECT 7.620 197.815 7.850 197.825 ;
        RECT 7.110 197.425 7.570 197.655 ;
        RECT 1.900 195.250 4.950 196.250 ;
        RECT 9.460 195.275 9.830 198.455 ;
        RECT 10.250 195.275 10.620 198.455 ;
        RECT 11.485 197.825 12.530 198.455 ;
        RECT 12.950 197.825 13.320 198.455 ;
        RECT 14.185 197.825 15.230 198.455 ;
        RECT 15.650 197.825 16.020 198.455 ;
        RECT 12.230 197.815 12.460 197.825 ;
        RECT 13.020 197.815 13.250 197.825 ;
        RECT 14.930 197.815 15.160 197.825 ;
        RECT 15.720 197.815 15.950 197.825 ;
        RECT 12.510 197.425 12.970 197.655 ;
        RECT 15.210 197.425 15.670 197.655 ;
        RECT 17.560 195.275 17.930 198.455 ;
        RECT 18.350 195.275 18.720 198.455 ;
        RECT 20.260 195.275 20.630 198.455 ;
        RECT 21.050 195.275 21.420 198.455 ;
        RECT 29.375 196.250 30.375 199.405 ;
        RECT 31.995 198.605 33.035 199.100 ;
        RECT 35.235 198.625 35.695 198.855 ;
        RECT 37.395 198.605 38.435 199.100 ;
        RECT 40.095 198.605 41.135 199.100 ;
        RECT 43.335 198.625 43.795 198.855 ;
        RECT 46.035 198.625 46.495 198.855 ;
        RECT 32.255 198.455 32.485 198.465 ;
        RECT 33.045 198.455 33.275 198.465 ;
        RECT 34.955 198.455 35.185 198.465 ;
        RECT 35.745 198.455 35.975 198.465 ;
        RECT 37.655 198.455 37.885 198.465 ;
        RECT 38.445 198.455 38.675 198.465 ;
        RECT 40.355 198.455 40.585 198.465 ;
        RECT 41.145 198.455 41.375 198.465 ;
        RECT 43.055 198.455 43.285 198.465 ;
        RECT 43.845 198.455 44.075 198.465 ;
        RECT 45.755 198.455 45.985 198.465 ;
        RECT 46.545 198.455 46.775 198.465 ;
        RECT 31.510 197.825 32.555 198.455 ;
        RECT 32.975 197.825 33.345 198.455 ;
        RECT 32.255 197.815 32.485 197.825 ;
        RECT 33.045 197.815 33.275 197.825 ;
        RECT 32.535 197.425 32.995 197.655 ;
        RECT 1.900 177.900 2.900 195.250 ;
        RECT 3.905 194.430 5.020 194.485 ;
        RECT 3.875 193.315 5.050 194.430 ;
        RECT 8.790 193.320 9.160 194.435 ;
        RECT 1.870 176.900 2.930 177.900 ;
        RECT 1.900 155.325 2.900 176.900 ;
        RECT 3.905 171.855 5.020 193.315 ;
        RECT 9.530 191.965 9.760 195.275 ;
        RECT 10.320 191.965 10.550 195.275 ;
        RECT 10.920 193.320 11.290 194.435 ;
        RECT 16.890 193.320 17.260 194.435 ;
        RECT 17.630 191.965 17.860 195.275 ;
        RECT 18.420 191.965 18.650 195.275 ;
        RECT 19.020 193.320 19.390 194.435 ;
        RECT 19.590 193.320 19.960 194.435 ;
        RECT 20.330 191.965 20.560 195.275 ;
        RECT 21.120 191.965 21.350 195.275 ;
        RECT 27.325 195.250 30.375 196.250 ;
        RECT 34.885 195.275 35.255 198.455 ;
        RECT 35.675 195.275 36.045 198.455 ;
        RECT 36.910 197.825 37.955 198.455 ;
        RECT 38.375 197.825 38.745 198.455 ;
        RECT 39.610 197.825 40.655 198.455 ;
        RECT 41.075 197.825 41.445 198.455 ;
        RECT 37.655 197.815 37.885 197.825 ;
        RECT 38.445 197.815 38.675 197.825 ;
        RECT 40.355 197.815 40.585 197.825 ;
        RECT 41.145 197.815 41.375 197.825 ;
        RECT 37.935 197.425 38.395 197.655 ;
        RECT 40.635 197.425 41.095 197.655 ;
        RECT 42.985 195.275 43.355 198.455 ;
        RECT 43.775 195.275 44.145 198.455 ;
        RECT 45.685 195.275 46.055 198.455 ;
        RECT 46.475 195.275 46.845 198.455 ;
        RECT 54.800 196.250 55.800 199.475 ;
        RECT 75.670 199.405 81.280 200.510 ;
        RECT 101.575 200.475 102.575 213.550 ;
        RECT 113.425 212.175 114.425 212.205 ;
        RECT 117.100 212.175 118.100 212.205 ;
        RECT 138.850 212.175 139.850 212.205 ;
        RECT 142.525 212.175 143.525 212.205 ;
        RECT 111.250 211.725 112.250 212.175 ;
        RECT 111.510 211.715 111.970 211.725 ;
        RECT 110.490 209.120 110.860 210.225 ;
        RECT 111.230 206.500 111.460 211.510 ;
        RECT 112.020 206.500 112.250 211.510 ;
        RECT 113.425 211.145 115.350 212.175 ;
        RECT 112.620 210.175 112.990 210.225 ;
        RECT 112.620 209.120 113.725 210.175 ;
        RECT 108.810 202.715 109.270 202.945 ;
        RECT 108.530 202.500 108.760 202.510 ;
        RECT 109.320 202.500 109.550 202.510 ;
        RECT 107.785 201.520 108.830 202.500 ;
        RECT 109.250 201.520 109.620 202.500 ;
        RECT 111.160 201.520 111.530 206.500 ;
        RECT 111.950 201.520 112.320 206.500 ;
        RECT 112.725 204.425 113.725 209.120 ;
        RECT 114.350 206.075 115.350 211.145 ;
        RECT 116.150 211.145 118.100 212.175 ;
        RECT 119.350 211.725 120.350 212.175 ;
        RECT 122.050 211.725 123.050 212.175 ;
        RECT 128.970 211.975 129.970 212.125 ;
        RECT 119.610 211.715 120.070 211.725 ;
        RECT 122.310 211.715 122.770 211.725 ;
        RECT 125.505 211.715 125.965 211.945 ;
        RECT 128.205 211.715 128.665 211.945 ;
        RECT 128.820 211.525 129.970 211.975 ;
        RECT 130.905 211.715 131.365 211.945 ;
        RECT 136.675 211.725 137.675 212.175 ;
        RECT 136.935 211.715 137.395 211.725 ;
        RECT 116.150 206.820 117.150 211.145 ;
        RECT 118.590 210.175 118.960 210.225 ;
        RECT 117.875 209.120 118.960 210.175 ;
        RECT 114.350 205.075 117.180 206.075 ;
        RECT 117.875 204.425 118.875 209.120 ;
        RECT 119.330 206.500 119.560 211.510 ;
        RECT 120.120 206.500 120.350 211.510 ;
        RECT 120.720 209.120 121.090 210.225 ;
        RECT 121.290 209.120 121.660 210.225 ;
        RECT 122.030 206.500 122.260 211.510 ;
        RECT 122.820 206.500 123.050 211.510 ;
        RECT 125.225 210.510 125.455 211.510 ;
        RECT 125.995 210.495 128.175 211.525 ;
        RECT 128.670 211.500 129.970 211.525 ;
        RECT 130.625 211.500 130.855 211.510 ;
        RECT 131.415 211.500 131.645 211.510 ;
        RECT 128.670 210.975 130.925 211.500 ;
        RECT 128.670 210.570 129.590 210.975 ;
        RECT 128.715 210.510 128.945 210.570 ;
        RECT 129.880 210.520 130.925 210.975 ;
        RECT 131.345 210.520 131.715 211.500 ;
        RECT 130.625 210.510 130.855 210.520 ;
        RECT 131.415 210.510 131.645 210.520 ;
        RECT 123.420 209.120 123.790 210.225 ;
        RECT 125.220 207.625 126.220 210.355 ;
        RECT 127.945 207.625 128.945 210.325 ;
        RECT 130.370 209.850 131.405 210.325 ;
        RECT 135.915 209.120 136.285 210.225 ;
        RECT 130.365 207.605 131.405 208.100 ;
        RECT 124.905 206.800 125.550 207.480 ;
        RECT 125.945 206.800 128.225 207.480 ;
        RECT 128.715 207.405 128.945 207.465 ;
        RECT 130.625 207.455 130.855 207.465 ;
        RECT 131.415 207.455 131.645 207.465 ;
        RECT 128.670 207.250 129.590 207.405 ;
        RECT 129.880 207.250 130.925 207.455 ;
        RECT 128.670 206.825 130.925 207.250 ;
        RECT 131.345 206.825 131.715 207.455 ;
        RECT 128.715 206.815 129.970 206.825 ;
        RECT 130.625 206.815 130.855 206.825 ;
        RECT 131.415 206.815 131.645 206.825 ;
        RECT 128.720 206.800 129.970 206.815 ;
        RECT 112.725 203.425 118.875 204.425 ;
        RECT 114.210 202.715 114.670 202.945 ;
        RECT 116.910 202.715 117.370 202.945 ;
        RECT 113.930 202.500 114.160 202.510 ;
        RECT 114.720 202.500 114.950 202.510 ;
        RECT 116.630 202.500 116.860 202.510 ;
        RECT 117.420 202.500 117.650 202.510 ;
        RECT 113.185 201.520 114.230 202.500 ;
        RECT 114.650 201.520 115.020 202.500 ;
        RECT 115.885 201.520 116.930 202.500 ;
        RECT 117.350 201.520 117.720 202.500 ;
        RECT 119.260 201.520 119.630 206.500 ;
        RECT 120.050 201.520 120.420 206.500 ;
        RECT 121.960 201.520 122.330 206.500 ;
        RECT 122.750 201.520 123.120 206.500 ;
        RECT 125.505 206.425 125.965 206.655 ;
        RECT 128.205 206.425 128.665 206.655 ;
        RECT 128.815 206.250 129.970 206.800 ;
        RECT 130.905 206.425 131.365 206.655 ;
        RECT 136.655 206.500 136.885 211.510 ;
        RECT 137.445 206.500 137.675 211.510 ;
        RECT 138.850 211.145 140.775 212.175 ;
        RECT 138.045 210.175 138.415 210.225 ;
        RECT 138.045 209.120 139.150 210.175 ;
        RECT 128.815 206.200 129.875 206.250 ;
        RECT 108.530 201.510 108.760 201.520 ;
        RECT 109.320 201.510 109.550 201.520 ;
        RECT 111.230 201.510 111.460 201.520 ;
        RECT 112.020 201.510 112.250 201.520 ;
        RECT 113.930 201.510 114.160 201.520 ;
        RECT 114.720 201.510 114.950 201.520 ;
        RECT 116.630 201.510 116.860 201.520 ;
        RECT 117.420 201.510 117.650 201.520 ;
        RECT 119.330 201.510 119.560 201.520 ;
        RECT 120.120 201.510 120.350 201.520 ;
        RECT 122.030 201.510 122.260 201.520 ;
        RECT 122.820 201.510 123.050 201.520 ;
        RECT 108.275 200.850 109.310 201.325 ;
        RECT 111.510 201.075 111.970 201.305 ;
        RECT 113.675 200.850 114.710 201.325 ;
        RECT 116.375 200.850 117.410 201.325 ;
        RECT 119.610 201.075 120.070 201.305 ;
        RECT 122.310 201.075 122.770 201.305 ;
        RECT 105.650 200.475 106.650 200.530 ;
        RECT 126.520 200.510 127.625 205.180 ;
        RECT 134.235 202.715 134.695 202.945 ;
        RECT 133.955 202.500 134.185 202.510 ;
        RECT 134.745 202.500 134.975 202.510 ;
        RECT 133.210 201.520 134.255 202.500 ;
        RECT 134.675 201.520 135.045 202.500 ;
        RECT 136.585 201.520 136.955 206.500 ;
        RECT 137.375 201.520 137.745 206.500 ;
        RECT 138.150 204.425 139.150 209.120 ;
        RECT 139.775 206.075 140.775 211.145 ;
        RECT 141.575 211.145 143.525 212.175 ;
        RECT 144.775 211.725 145.775 212.175 ;
        RECT 147.475 211.725 148.475 212.175 ;
        RECT 145.035 211.715 145.495 211.725 ;
        RECT 147.735 211.715 148.195 211.725 ;
        RECT 141.575 206.820 142.575 211.145 ;
        RECT 144.015 210.175 144.385 210.225 ;
        RECT 143.300 209.120 144.385 210.175 ;
        RECT 139.775 205.075 142.605 206.075 ;
        RECT 143.300 204.425 144.300 209.120 ;
        RECT 144.755 206.500 144.985 211.510 ;
        RECT 145.545 206.500 145.775 211.510 ;
        RECT 146.145 209.120 146.515 210.225 ;
        RECT 146.715 209.120 147.085 210.225 ;
        RECT 147.455 206.500 147.685 211.510 ;
        RECT 148.245 206.500 148.475 211.510 ;
        RECT 148.845 209.120 149.215 210.225 ;
        RECT 138.150 203.425 144.300 204.425 ;
        RECT 139.635 202.715 140.095 202.945 ;
        RECT 142.335 202.715 142.795 202.945 ;
        RECT 139.355 202.500 139.585 202.510 ;
        RECT 140.145 202.500 140.375 202.510 ;
        RECT 142.055 202.500 142.285 202.510 ;
        RECT 142.845 202.500 143.075 202.510 ;
        RECT 138.610 201.520 139.655 202.500 ;
        RECT 140.075 201.520 140.445 202.500 ;
        RECT 141.310 201.520 142.355 202.500 ;
        RECT 142.775 201.520 143.145 202.500 ;
        RECT 144.685 201.520 145.055 206.500 ;
        RECT 145.475 201.520 145.845 206.500 ;
        RECT 147.385 201.520 147.755 206.500 ;
        RECT 148.175 201.520 148.545 206.500 ;
        RECT 133.955 201.510 134.185 201.520 ;
        RECT 134.745 201.510 134.975 201.520 ;
        RECT 136.655 201.510 136.885 201.520 ;
        RECT 137.445 201.510 137.675 201.520 ;
        RECT 139.355 201.510 139.585 201.520 ;
        RECT 140.145 201.510 140.375 201.520 ;
        RECT 142.055 201.510 142.285 201.520 ;
        RECT 142.845 201.510 143.075 201.520 ;
        RECT 144.755 201.510 144.985 201.520 ;
        RECT 145.545 201.510 145.775 201.520 ;
        RECT 147.455 201.510 147.685 201.520 ;
        RECT 148.245 201.510 148.475 201.520 ;
        RECT 133.700 200.850 134.735 201.325 ;
        RECT 136.935 201.075 137.395 201.305 ;
        RECT 139.100 200.850 140.135 201.325 ;
        RECT 141.800 200.850 142.835 201.325 ;
        RECT 145.035 201.075 145.495 201.305 ;
        RECT 147.735 201.075 148.195 201.305 ;
        RECT 131.075 200.510 132.075 200.530 ;
        RECT 101.545 199.475 102.605 200.475 ;
        RECT 105.620 199.475 106.680 200.475 ;
        RECT 57.420 198.605 58.460 199.100 ;
        RECT 60.660 198.625 61.120 198.855 ;
        RECT 62.820 198.605 63.860 199.100 ;
        RECT 65.520 198.605 66.560 199.100 ;
        RECT 68.760 198.625 69.220 198.855 ;
        RECT 71.460 198.625 71.920 198.855 ;
        RECT 57.680 198.455 57.910 198.465 ;
        RECT 58.470 198.455 58.700 198.465 ;
        RECT 60.380 198.455 60.610 198.465 ;
        RECT 61.170 198.455 61.400 198.465 ;
        RECT 63.080 198.455 63.310 198.465 ;
        RECT 63.870 198.455 64.100 198.465 ;
        RECT 65.780 198.455 66.010 198.465 ;
        RECT 66.570 198.455 66.800 198.465 ;
        RECT 68.480 198.455 68.710 198.465 ;
        RECT 69.270 198.455 69.500 198.465 ;
        RECT 71.180 198.455 71.410 198.465 ;
        RECT 71.970 198.455 72.200 198.465 ;
        RECT 56.935 197.825 57.980 198.455 ;
        RECT 58.400 197.825 58.770 198.455 ;
        RECT 57.680 197.815 57.910 197.825 ;
        RECT 58.470 197.815 58.700 197.825 ;
        RECT 57.960 197.425 58.420 197.655 ;
        RECT 21.720 193.320 22.090 194.435 ;
        RECT 9.810 191.775 10.270 191.805 ;
        RECT 17.910 191.775 18.370 191.805 ;
        RECT 20.610 191.775 21.070 191.805 ;
        RECT 9.550 191.375 10.550 191.775 ;
        RECT 17.650 191.375 18.650 191.775 ;
        RECT 20.350 191.375 21.350 191.775 ;
        RECT 11.725 189.600 12.725 189.630 ;
        RECT 15.400 189.600 16.400 189.630 ;
        RECT 9.550 189.150 10.550 189.600 ;
        RECT 9.810 189.140 10.270 189.150 ;
        RECT 8.790 186.545 9.160 187.650 ;
        RECT 9.530 183.925 9.760 188.935 ;
        RECT 10.320 183.925 10.550 188.935 ;
        RECT 11.725 188.570 13.650 189.600 ;
        RECT 10.920 187.600 11.290 187.650 ;
        RECT 10.920 186.545 12.025 187.600 ;
        RECT 7.110 180.140 7.570 180.370 ;
        RECT 6.830 179.925 7.060 179.935 ;
        RECT 7.620 179.925 7.850 179.935 ;
        RECT 6.085 178.945 7.130 179.925 ;
        RECT 7.550 178.945 7.920 179.925 ;
        RECT 9.460 178.945 9.830 183.925 ;
        RECT 10.250 178.945 10.620 183.925 ;
        RECT 11.025 181.850 12.025 186.545 ;
        RECT 12.650 183.500 13.650 188.570 ;
        RECT 14.450 188.570 16.400 189.600 ;
        RECT 17.650 189.150 18.650 189.600 ;
        RECT 20.350 189.150 21.350 189.600 ;
        RECT 17.910 189.140 18.370 189.150 ;
        RECT 20.610 189.140 21.070 189.150 ;
        RECT 14.450 184.245 15.450 188.570 ;
        RECT 16.890 187.600 17.260 187.650 ;
        RECT 16.175 186.545 17.260 187.600 ;
        RECT 12.650 182.500 15.480 183.500 ;
        RECT 16.175 181.850 17.175 186.545 ;
        RECT 17.630 183.925 17.860 188.935 ;
        RECT 18.420 183.925 18.650 188.935 ;
        RECT 19.020 186.545 19.390 187.650 ;
        RECT 19.590 186.545 19.960 187.650 ;
        RECT 20.330 183.925 20.560 188.935 ;
        RECT 21.120 183.925 21.350 188.935 ;
        RECT 21.720 186.545 22.090 187.650 ;
        RECT 11.025 180.850 17.175 181.850 ;
        RECT 12.510 180.140 12.970 180.370 ;
        RECT 15.210 180.140 15.670 180.370 ;
        RECT 12.230 179.925 12.460 179.935 ;
        RECT 13.020 179.925 13.250 179.935 ;
        RECT 14.930 179.925 15.160 179.935 ;
        RECT 15.720 179.925 15.950 179.935 ;
        RECT 11.485 178.945 12.530 179.925 ;
        RECT 12.950 178.945 13.320 179.925 ;
        RECT 14.185 178.945 15.230 179.925 ;
        RECT 15.650 178.945 16.020 179.925 ;
        RECT 17.560 178.945 17.930 183.925 ;
        RECT 18.350 178.945 18.720 183.925 ;
        RECT 20.260 178.945 20.630 183.925 ;
        RECT 21.050 178.945 21.420 183.925 ;
        RECT 6.830 178.935 7.060 178.945 ;
        RECT 7.620 178.935 7.850 178.945 ;
        RECT 9.530 178.935 9.760 178.945 ;
        RECT 10.320 178.935 10.550 178.945 ;
        RECT 12.230 178.935 12.460 178.945 ;
        RECT 13.020 178.935 13.250 178.945 ;
        RECT 14.930 178.935 15.160 178.945 ;
        RECT 15.720 178.935 15.950 178.945 ;
        RECT 17.630 178.935 17.860 178.945 ;
        RECT 18.420 178.935 18.650 178.945 ;
        RECT 20.330 178.935 20.560 178.945 ;
        RECT 21.120 178.935 21.350 178.945 ;
        RECT 6.575 178.275 7.610 178.750 ;
        RECT 9.810 178.500 10.270 178.730 ;
        RECT 11.975 178.275 13.010 178.750 ;
        RECT 14.675 178.275 15.710 178.750 ;
        RECT 17.910 178.500 18.370 178.730 ;
        RECT 20.610 178.500 21.070 178.730 ;
        RECT 27.325 177.900 28.325 195.250 ;
        RECT 29.330 194.430 30.445 194.485 ;
        RECT 29.300 193.315 30.475 194.430 ;
        RECT 34.215 193.320 34.585 194.435 ;
        RECT 27.295 176.900 28.355 177.900 ;
        RECT 6.570 176.030 7.610 176.525 ;
        RECT 9.810 176.050 10.270 176.280 ;
        RECT 11.970 176.030 13.010 176.525 ;
        RECT 14.670 176.030 15.710 176.525 ;
        RECT 17.910 176.050 18.370 176.280 ;
        RECT 20.610 176.050 21.070 176.280 ;
        RECT 6.830 175.880 7.060 175.890 ;
        RECT 7.620 175.880 7.850 175.890 ;
        RECT 9.530 175.880 9.760 175.890 ;
        RECT 10.320 175.880 10.550 175.890 ;
        RECT 12.230 175.880 12.460 175.890 ;
        RECT 13.020 175.880 13.250 175.890 ;
        RECT 14.930 175.880 15.160 175.890 ;
        RECT 15.720 175.880 15.950 175.890 ;
        RECT 17.630 175.880 17.860 175.890 ;
        RECT 18.420 175.880 18.650 175.890 ;
        RECT 20.330 175.880 20.560 175.890 ;
        RECT 21.120 175.880 21.350 175.890 ;
        RECT 6.085 175.250 7.130 175.880 ;
        RECT 7.550 175.250 7.920 175.880 ;
        RECT 6.830 175.240 7.060 175.250 ;
        RECT 7.620 175.240 7.850 175.250 ;
        RECT 7.110 174.850 7.570 175.080 ;
        RECT 9.460 172.700 9.830 175.880 ;
        RECT 10.250 172.700 10.620 175.880 ;
        RECT 11.485 175.250 12.530 175.880 ;
        RECT 12.950 175.250 13.320 175.880 ;
        RECT 14.185 175.250 15.230 175.880 ;
        RECT 15.650 175.250 16.020 175.880 ;
        RECT 12.230 175.240 12.460 175.250 ;
        RECT 13.020 175.240 13.250 175.250 ;
        RECT 14.930 175.240 15.160 175.250 ;
        RECT 15.720 175.240 15.950 175.250 ;
        RECT 12.510 174.850 12.970 175.080 ;
        RECT 15.210 174.850 15.670 175.080 ;
        RECT 17.560 172.700 17.930 175.880 ;
        RECT 18.350 172.700 18.720 175.880 ;
        RECT 20.260 172.700 20.630 175.880 ;
        RECT 21.050 172.700 21.420 175.880 ;
        RECT 3.875 170.740 5.050 171.855 ;
        RECT 8.790 170.745 9.160 171.860 ;
        RECT 1.870 154.325 2.930 155.325 ;
        RECT 1.900 154.295 2.900 154.325 ;
        RECT 3.905 149.285 5.020 170.740 ;
        RECT 9.530 169.390 9.760 172.700 ;
        RECT 10.320 169.390 10.550 172.700 ;
        RECT 10.920 170.745 11.290 171.860 ;
        RECT 16.890 170.745 17.260 171.860 ;
        RECT 17.630 169.390 17.860 172.700 ;
        RECT 18.420 169.390 18.650 172.700 ;
        RECT 19.020 170.745 19.390 171.860 ;
        RECT 19.590 170.745 19.960 171.860 ;
        RECT 20.330 169.390 20.560 172.700 ;
        RECT 21.120 169.390 21.350 172.700 ;
        RECT 21.720 170.745 22.090 171.860 ;
        RECT 23.085 170.745 24.260 171.860 ;
        RECT 9.810 169.200 10.270 169.230 ;
        RECT 17.910 169.200 18.370 169.230 ;
        RECT 20.610 169.200 21.070 169.230 ;
        RECT 9.550 168.800 10.550 169.200 ;
        RECT 17.650 168.800 18.650 169.200 ;
        RECT 20.350 168.800 21.350 169.200 ;
        RECT 23.115 167.770 24.230 170.745 ;
        RECT 11.725 167.025 12.725 167.055 ;
        RECT 15.400 167.025 16.400 167.055 ;
        RECT 9.550 166.575 10.550 167.025 ;
        RECT 9.810 166.565 10.270 166.575 ;
        RECT 8.790 163.970 9.160 165.075 ;
        RECT 9.530 161.350 9.760 166.360 ;
        RECT 10.320 161.350 10.550 166.360 ;
        RECT 11.725 165.995 13.650 167.025 ;
        RECT 10.920 165.025 11.290 165.075 ;
        RECT 10.920 163.970 12.025 165.025 ;
        RECT 7.110 157.565 7.570 157.795 ;
        RECT 6.830 157.350 7.060 157.360 ;
        RECT 7.620 157.350 7.850 157.360 ;
        RECT 6.085 156.370 7.130 157.350 ;
        RECT 7.550 156.370 7.920 157.350 ;
        RECT 9.460 156.370 9.830 161.350 ;
        RECT 10.250 156.370 10.620 161.350 ;
        RECT 11.025 159.275 12.025 163.970 ;
        RECT 12.650 160.925 13.650 165.995 ;
        RECT 14.450 165.995 16.400 167.025 ;
        RECT 17.650 166.575 18.650 167.025 ;
        RECT 20.350 166.575 21.350 167.025 ;
        RECT 17.910 166.565 18.370 166.575 ;
        RECT 20.610 166.565 21.070 166.575 ;
        RECT 14.450 161.670 15.450 165.995 ;
        RECT 16.890 165.025 17.260 165.075 ;
        RECT 16.175 163.970 17.260 165.025 ;
        RECT 12.650 159.925 15.480 160.925 ;
        RECT 16.175 159.275 17.175 163.970 ;
        RECT 17.630 161.350 17.860 166.360 ;
        RECT 18.420 161.350 18.650 166.360 ;
        RECT 19.020 163.970 19.390 165.075 ;
        RECT 19.590 163.970 19.960 165.075 ;
        RECT 20.330 161.350 20.560 166.360 ;
        RECT 21.120 161.350 21.350 166.360 ;
        RECT 23.430 165.115 23.880 167.425 ;
        RECT 21.720 163.970 22.090 165.075 ;
        RECT 11.025 158.275 17.175 159.275 ;
        RECT 12.510 157.565 12.970 157.795 ;
        RECT 15.210 157.565 15.670 157.795 ;
        RECT 12.230 157.350 12.460 157.360 ;
        RECT 13.020 157.350 13.250 157.360 ;
        RECT 14.930 157.350 15.160 157.360 ;
        RECT 15.720 157.350 15.950 157.360 ;
        RECT 11.485 156.370 12.530 157.350 ;
        RECT 12.950 156.370 13.320 157.350 ;
        RECT 14.185 156.370 15.230 157.350 ;
        RECT 15.650 156.370 16.020 157.350 ;
        RECT 17.560 156.370 17.930 161.350 ;
        RECT 18.350 156.370 18.720 161.350 ;
        RECT 20.260 156.370 20.630 161.350 ;
        RECT 21.050 156.370 21.420 161.350 ;
        RECT 6.830 156.360 7.060 156.370 ;
        RECT 7.620 156.360 7.850 156.370 ;
        RECT 9.530 156.360 9.760 156.370 ;
        RECT 10.320 156.360 10.550 156.370 ;
        RECT 12.230 156.360 12.460 156.370 ;
        RECT 13.020 156.360 13.250 156.370 ;
        RECT 14.930 156.360 15.160 156.370 ;
        RECT 15.720 156.360 15.950 156.370 ;
        RECT 17.630 156.360 17.860 156.370 ;
        RECT 18.420 156.360 18.650 156.370 ;
        RECT 20.330 156.360 20.560 156.370 ;
        RECT 21.120 156.360 21.350 156.370 ;
        RECT 6.575 155.700 7.610 156.175 ;
        RECT 9.810 155.925 10.270 156.155 ;
        RECT 11.975 155.700 13.010 156.175 ;
        RECT 14.675 155.700 15.710 156.175 ;
        RECT 17.910 155.925 18.370 156.155 ;
        RECT 20.610 155.925 21.070 156.155 ;
        RECT 23.430 154.205 23.880 156.515 ;
        RECT 27.325 155.325 28.325 176.900 ;
        RECT 29.330 171.855 30.445 193.315 ;
        RECT 34.955 191.965 35.185 195.275 ;
        RECT 35.745 191.965 35.975 195.275 ;
        RECT 36.345 193.320 36.715 194.435 ;
        RECT 42.315 193.320 42.685 194.435 ;
        RECT 43.055 191.965 43.285 195.275 ;
        RECT 43.845 191.965 44.075 195.275 ;
        RECT 44.445 193.320 44.815 194.435 ;
        RECT 45.015 193.320 45.385 194.435 ;
        RECT 45.755 191.965 45.985 195.275 ;
        RECT 46.545 191.965 46.775 195.275 ;
        RECT 52.750 195.250 55.800 196.250 ;
        RECT 60.310 195.275 60.680 198.455 ;
        RECT 61.100 195.275 61.470 198.455 ;
        RECT 62.335 197.825 63.380 198.455 ;
        RECT 63.800 197.825 64.170 198.455 ;
        RECT 65.035 197.825 66.080 198.455 ;
        RECT 66.500 197.825 66.870 198.455 ;
        RECT 63.080 197.815 63.310 197.825 ;
        RECT 63.870 197.815 64.100 197.825 ;
        RECT 65.780 197.815 66.010 197.825 ;
        RECT 66.570 197.815 66.800 197.825 ;
        RECT 63.360 197.425 63.820 197.655 ;
        RECT 66.060 197.425 66.520 197.655 ;
        RECT 68.410 195.275 68.780 198.455 ;
        RECT 69.200 195.275 69.570 198.455 ;
        RECT 71.110 195.275 71.480 198.455 ;
        RECT 71.900 195.275 72.270 198.455 ;
        RECT 80.225 196.250 81.225 199.405 ;
        RECT 82.845 198.605 83.885 199.100 ;
        RECT 86.085 198.625 86.545 198.855 ;
        RECT 88.245 198.605 89.285 199.100 ;
        RECT 90.945 198.605 91.985 199.100 ;
        RECT 94.185 198.625 94.645 198.855 ;
        RECT 96.885 198.625 97.345 198.855 ;
        RECT 83.105 198.455 83.335 198.465 ;
        RECT 83.895 198.455 84.125 198.465 ;
        RECT 85.805 198.455 86.035 198.465 ;
        RECT 86.595 198.455 86.825 198.465 ;
        RECT 88.505 198.455 88.735 198.465 ;
        RECT 89.295 198.455 89.525 198.465 ;
        RECT 91.205 198.455 91.435 198.465 ;
        RECT 91.995 198.455 92.225 198.465 ;
        RECT 93.905 198.455 94.135 198.465 ;
        RECT 94.695 198.455 94.925 198.465 ;
        RECT 96.605 198.455 96.835 198.465 ;
        RECT 97.395 198.455 97.625 198.465 ;
        RECT 82.360 197.825 83.405 198.455 ;
        RECT 83.825 197.825 84.195 198.455 ;
        RECT 83.105 197.815 83.335 197.825 ;
        RECT 83.895 197.815 84.125 197.825 ;
        RECT 83.385 197.425 83.845 197.655 ;
        RECT 47.145 193.320 47.515 194.435 ;
        RECT 35.235 191.775 35.695 191.805 ;
        RECT 43.335 191.775 43.795 191.805 ;
        RECT 46.035 191.775 46.495 191.805 ;
        RECT 34.975 191.375 35.975 191.775 ;
        RECT 43.075 191.375 44.075 191.775 ;
        RECT 45.775 191.375 46.775 191.775 ;
        RECT 37.150 189.600 38.150 189.630 ;
        RECT 40.825 189.600 41.825 189.630 ;
        RECT 34.975 189.150 35.975 189.600 ;
        RECT 35.235 189.140 35.695 189.150 ;
        RECT 34.215 186.545 34.585 187.650 ;
        RECT 34.955 183.925 35.185 188.935 ;
        RECT 35.745 183.925 35.975 188.935 ;
        RECT 37.150 188.570 39.075 189.600 ;
        RECT 36.345 187.600 36.715 187.650 ;
        RECT 36.345 186.545 37.450 187.600 ;
        RECT 32.535 180.140 32.995 180.370 ;
        RECT 32.255 179.925 32.485 179.935 ;
        RECT 33.045 179.925 33.275 179.935 ;
        RECT 31.510 178.945 32.555 179.925 ;
        RECT 32.975 178.945 33.345 179.925 ;
        RECT 34.885 178.945 35.255 183.925 ;
        RECT 35.675 178.945 36.045 183.925 ;
        RECT 36.450 181.850 37.450 186.545 ;
        RECT 38.075 183.500 39.075 188.570 ;
        RECT 39.875 188.570 41.825 189.600 ;
        RECT 43.075 189.150 44.075 189.600 ;
        RECT 45.775 189.150 46.775 189.600 ;
        RECT 43.335 189.140 43.795 189.150 ;
        RECT 46.035 189.140 46.495 189.150 ;
        RECT 39.875 184.245 40.875 188.570 ;
        RECT 42.315 187.600 42.685 187.650 ;
        RECT 41.600 186.545 42.685 187.600 ;
        RECT 38.075 182.500 40.905 183.500 ;
        RECT 41.600 181.850 42.600 186.545 ;
        RECT 43.055 183.925 43.285 188.935 ;
        RECT 43.845 183.925 44.075 188.935 ;
        RECT 44.445 186.545 44.815 187.650 ;
        RECT 45.015 186.545 45.385 187.650 ;
        RECT 45.755 183.925 45.985 188.935 ;
        RECT 46.545 183.925 46.775 188.935 ;
        RECT 47.145 186.545 47.515 187.650 ;
        RECT 36.450 180.850 42.600 181.850 ;
        RECT 37.935 180.140 38.395 180.370 ;
        RECT 40.635 180.140 41.095 180.370 ;
        RECT 37.655 179.925 37.885 179.935 ;
        RECT 38.445 179.925 38.675 179.935 ;
        RECT 40.355 179.925 40.585 179.935 ;
        RECT 41.145 179.925 41.375 179.935 ;
        RECT 36.910 178.945 37.955 179.925 ;
        RECT 38.375 178.945 38.745 179.925 ;
        RECT 39.610 178.945 40.655 179.925 ;
        RECT 41.075 178.945 41.445 179.925 ;
        RECT 42.985 178.945 43.355 183.925 ;
        RECT 43.775 178.945 44.145 183.925 ;
        RECT 45.685 178.945 46.055 183.925 ;
        RECT 46.475 178.945 46.845 183.925 ;
        RECT 32.255 178.935 32.485 178.945 ;
        RECT 33.045 178.935 33.275 178.945 ;
        RECT 34.955 178.935 35.185 178.945 ;
        RECT 35.745 178.935 35.975 178.945 ;
        RECT 37.655 178.935 37.885 178.945 ;
        RECT 38.445 178.935 38.675 178.945 ;
        RECT 40.355 178.935 40.585 178.945 ;
        RECT 41.145 178.935 41.375 178.945 ;
        RECT 43.055 178.935 43.285 178.945 ;
        RECT 43.845 178.935 44.075 178.945 ;
        RECT 45.755 178.935 45.985 178.945 ;
        RECT 46.545 178.935 46.775 178.945 ;
        RECT 32.000 178.275 33.035 178.750 ;
        RECT 35.235 178.500 35.695 178.730 ;
        RECT 37.400 178.275 38.435 178.750 ;
        RECT 40.100 178.275 41.135 178.750 ;
        RECT 43.335 178.500 43.795 178.730 ;
        RECT 46.035 178.500 46.495 178.730 ;
        RECT 52.750 177.900 53.750 195.250 ;
        RECT 54.755 194.430 55.870 194.485 ;
        RECT 54.725 193.315 55.900 194.430 ;
        RECT 59.640 193.320 60.010 194.435 ;
        RECT 52.720 176.900 53.780 177.900 ;
        RECT 31.995 176.030 33.035 176.525 ;
        RECT 35.235 176.050 35.695 176.280 ;
        RECT 37.395 176.030 38.435 176.525 ;
        RECT 40.095 176.030 41.135 176.525 ;
        RECT 43.335 176.050 43.795 176.280 ;
        RECT 46.035 176.050 46.495 176.280 ;
        RECT 32.255 175.880 32.485 175.890 ;
        RECT 33.045 175.880 33.275 175.890 ;
        RECT 34.955 175.880 35.185 175.890 ;
        RECT 35.745 175.880 35.975 175.890 ;
        RECT 37.655 175.880 37.885 175.890 ;
        RECT 38.445 175.880 38.675 175.890 ;
        RECT 40.355 175.880 40.585 175.890 ;
        RECT 41.145 175.880 41.375 175.890 ;
        RECT 43.055 175.880 43.285 175.890 ;
        RECT 43.845 175.880 44.075 175.890 ;
        RECT 45.755 175.880 45.985 175.890 ;
        RECT 46.545 175.880 46.775 175.890 ;
        RECT 31.510 175.250 32.555 175.880 ;
        RECT 32.975 175.250 33.345 175.880 ;
        RECT 32.255 175.240 32.485 175.250 ;
        RECT 33.045 175.240 33.275 175.250 ;
        RECT 32.535 174.850 32.995 175.080 ;
        RECT 34.885 172.700 35.255 175.880 ;
        RECT 35.675 172.700 36.045 175.880 ;
        RECT 36.910 175.250 37.955 175.880 ;
        RECT 38.375 175.250 38.745 175.880 ;
        RECT 39.610 175.250 40.655 175.880 ;
        RECT 41.075 175.250 41.445 175.880 ;
        RECT 37.655 175.240 37.885 175.250 ;
        RECT 38.445 175.240 38.675 175.250 ;
        RECT 40.355 175.240 40.585 175.250 ;
        RECT 41.145 175.240 41.375 175.250 ;
        RECT 37.935 174.850 38.395 175.080 ;
        RECT 40.635 174.850 41.095 175.080 ;
        RECT 42.985 172.700 43.355 175.880 ;
        RECT 43.775 172.700 44.145 175.880 ;
        RECT 45.685 172.700 46.055 175.880 ;
        RECT 46.475 172.700 46.845 175.880 ;
        RECT 29.300 170.740 30.475 171.855 ;
        RECT 34.215 170.745 34.585 171.860 ;
        RECT 27.295 154.325 28.355 155.325 ;
        RECT 27.325 154.295 28.325 154.325 ;
        RECT 6.570 153.455 7.610 153.950 ;
        RECT 9.810 153.475 10.270 153.705 ;
        RECT 11.970 153.455 13.010 153.950 ;
        RECT 14.670 153.455 15.710 153.950 ;
        RECT 17.910 153.475 18.370 153.705 ;
        RECT 20.610 153.475 21.070 153.705 ;
        RECT 6.830 153.305 7.060 153.315 ;
        RECT 7.620 153.305 7.850 153.315 ;
        RECT 9.530 153.305 9.760 153.315 ;
        RECT 10.320 153.305 10.550 153.315 ;
        RECT 12.230 153.305 12.460 153.315 ;
        RECT 13.020 153.305 13.250 153.315 ;
        RECT 14.930 153.305 15.160 153.315 ;
        RECT 15.720 153.305 15.950 153.315 ;
        RECT 17.630 153.305 17.860 153.315 ;
        RECT 18.420 153.305 18.650 153.315 ;
        RECT 20.330 153.305 20.560 153.315 ;
        RECT 21.120 153.305 21.350 153.315 ;
        RECT 6.085 152.675 7.130 153.305 ;
        RECT 7.550 152.675 7.920 153.305 ;
        RECT 6.830 152.665 7.060 152.675 ;
        RECT 7.620 152.665 7.850 152.675 ;
        RECT 7.110 152.275 7.570 152.505 ;
        RECT 9.460 150.125 9.830 153.305 ;
        RECT 10.250 150.125 10.620 153.305 ;
        RECT 11.485 152.675 12.530 153.305 ;
        RECT 12.950 152.675 13.320 153.305 ;
        RECT 14.185 152.675 15.230 153.305 ;
        RECT 15.650 152.675 16.020 153.305 ;
        RECT 12.230 152.665 12.460 152.675 ;
        RECT 13.020 152.665 13.250 152.675 ;
        RECT 14.930 152.665 15.160 152.675 ;
        RECT 15.720 152.665 15.950 152.675 ;
        RECT 12.510 152.275 12.970 152.505 ;
        RECT 15.210 152.275 15.670 152.505 ;
        RECT 17.560 150.125 17.930 153.305 ;
        RECT 18.350 150.125 18.720 153.305 ;
        RECT 20.260 150.125 20.630 153.305 ;
        RECT 21.050 150.125 21.420 153.305 ;
        RECT 3.860 148.170 5.060 149.285 ;
        RECT 8.790 148.170 9.160 149.285 ;
        RECT 3.905 148.140 5.020 148.170 ;
        RECT 9.530 146.815 9.760 150.125 ;
        RECT 10.320 146.815 10.550 150.125 ;
        RECT 10.920 148.170 11.290 149.285 ;
        RECT 16.890 148.170 17.260 149.285 ;
        RECT 17.630 146.815 17.860 150.125 ;
        RECT 18.420 146.815 18.650 150.125 ;
        RECT 19.020 148.170 19.390 149.285 ;
        RECT 19.590 148.170 19.960 149.285 ;
        RECT 20.330 146.815 20.560 150.125 ;
        RECT 21.120 146.815 21.350 150.125 ;
        RECT 21.720 148.170 22.090 149.285 ;
        RECT 23.090 148.140 24.205 153.855 ;
        RECT 29.330 149.285 30.445 170.740 ;
        RECT 34.955 169.390 35.185 172.700 ;
        RECT 35.745 169.390 35.975 172.700 ;
        RECT 36.345 170.745 36.715 171.860 ;
        RECT 42.315 170.745 42.685 171.860 ;
        RECT 43.055 169.390 43.285 172.700 ;
        RECT 43.845 169.390 44.075 172.700 ;
        RECT 44.445 170.745 44.815 171.860 ;
        RECT 45.015 170.745 45.385 171.860 ;
        RECT 45.755 169.390 45.985 172.700 ;
        RECT 46.545 169.390 46.775 172.700 ;
        RECT 47.145 170.745 47.515 171.860 ;
        RECT 48.510 170.745 49.685 171.860 ;
        RECT 35.235 169.200 35.695 169.230 ;
        RECT 43.335 169.200 43.795 169.230 ;
        RECT 46.035 169.200 46.495 169.230 ;
        RECT 34.975 168.800 35.975 169.200 ;
        RECT 43.075 168.800 44.075 169.200 ;
        RECT 45.775 168.800 46.775 169.200 ;
        RECT 48.540 167.770 49.655 170.745 ;
        RECT 37.150 167.025 38.150 167.055 ;
        RECT 40.825 167.025 41.825 167.055 ;
        RECT 34.975 166.575 35.975 167.025 ;
        RECT 35.235 166.565 35.695 166.575 ;
        RECT 34.215 163.970 34.585 165.075 ;
        RECT 34.955 161.350 35.185 166.360 ;
        RECT 35.745 161.350 35.975 166.360 ;
        RECT 37.150 165.995 39.075 167.025 ;
        RECT 36.345 165.025 36.715 165.075 ;
        RECT 36.345 163.970 37.450 165.025 ;
        RECT 32.535 157.565 32.995 157.795 ;
        RECT 32.255 157.350 32.485 157.360 ;
        RECT 33.045 157.350 33.275 157.360 ;
        RECT 31.510 156.370 32.555 157.350 ;
        RECT 32.975 156.370 33.345 157.350 ;
        RECT 34.885 156.370 35.255 161.350 ;
        RECT 35.675 156.370 36.045 161.350 ;
        RECT 36.450 159.275 37.450 163.970 ;
        RECT 38.075 160.925 39.075 165.995 ;
        RECT 39.875 165.995 41.825 167.025 ;
        RECT 43.075 166.575 44.075 167.025 ;
        RECT 45.775 166.575 46.775 167.025 ;
        RECT 43.335 166.565 43.795 166.575 ;
        RECT 46.035 166.565 46.495 166.575 ;
        RECT 39.875 161.670 40.875 165.995 ;
        RECT 42.315 165.025 42.685 165.075 ;
        RECT 41.600 163.970 42.685 165.025 ;
        RECT 38.075 159.925 40.905 160.925 ;
        RECT 41.600 159.275 42.600 163.970 ;
        RECT 43.055 161.350 43.285 166.360 ;
        RECT 43.845 161.350 44.075 166.360 ;
        RECT 44.445 163.970 44.815 165.075 ;
        RECT 45.015 163.970 45.385 165.075 ;
        RECT 45.755 161.350 45.985 166.360 ;
        RECT 46.545 161.350 46.775 166.360 ;
        RECT 48.855 165.115 49.305 167.425 ;
        RECT 47.145 163.970 47.515 165.075 ;
        RECT 36.450 158.275 42.600 159.275 ;
        RECT 37.935 157.565 38.395 157.795 ;
        RECT 40.635 157.565 41.095 157.795 ;
        RECT 37.655 157.350 37.885 157.360 ;
        RECT 38.445 157.350 38.675 157.360 ;
        RECT 40.355 157.350 40.585 157.360 ;
        RECT 41.145 157.350 41.375 157.360 ;
        RECT 36.910 156.370 37.955 157.350 ;
        RECT 38.375 156.370 38.745 157.350 ;
        RECT 39.610 156.370 40.655 157.350 ;
        RECT 41.075 156.370 41.445 157.350 ;
        RECT 42.985 156.370 43.355 161.350 ;
        RECT 43.775 156.370 44.145 161.350 ;
        RECT 45.685 156.370 46.055 161.350 ;
        RECT 46.475 156.370 46.845 161.350 ;
        RECT 32.255 156.360 32.485 156.370 ;
        RECT 33.045 156.360 33.275 156.370 ;
        RECT 34.955 156.360 35.185 156.370 ;
        RECT 35.745 156.360 35.975 156.370 ;
        RECT 37.655 156.360 37.885 156.370 ;
        RECT 38.445 156.360 38.675 156.370 ;
        RECT 40.355 156.360 40.585 156.370 ;
        RECT 41.145 156.360 41.375 156.370 ;
        RECT 43.055 156.360 43.285 156.370 ;
        RECT 43.845 156.360 44.075 156.370 ;
        RECT 45.755 156.360 45.985 156.370 ;
        RECT 46.545 156.360 46.775 156.370 ;
        RECT 32.000 155.700 33.035 156.175 ;
        RECT 35.235 155.925 35.695 156.155 ;
        RECT 37.400 155.700 38.435 156.175 ;
        RECT 40.100 155.700 41.135 156.175 ;
        RECT 43.335 155.925 43.795 156.155 ;
        RECT 46.035 155.925 46.495 156.155 ;
        RECT 48.855 154.205 49.305 156.515 ;
        RECT 52.750 155.325 53.750 176.900 ;
        RECT 54.755 171.855 55.870 193.315 ;
        RECT 60.380 191.965 60.610 195.275 ;
        RECT 61.170 191.965 61.400 195.275 ;
        RECT 61.770 193.320 62.140 194.435 ;
        RECT 67.740 193.320 68.110 194.435 ;
        RECT 68.480 191.965 68.710 195.275 ;
        RECT 69.270 191.965 69.500 195.275 ;
        RECT 69.870 193.320 70.240 194.435 ;
        RECT 70.440 193.320 70.810 194.435 ;
        RECT 71.180 191.965 71.410 195.275 ;
        RECT 71.970 191.965 72.200 195.275 ;
        RECT 78.175 195.250 81.225 196.250 ;
        RECT 85.735 195.275 86.105 198.455 ;
        RECT 86.525 195.275 86.895 198.455 ;
        RECT 87.760 197.825 88.805 198.455 ;
        RECT 89.225 197.825 89.595 198.455 ;
        RECT 90.460 197.825 91.505 198.455 ;
        RECT 91.925 197.825 92.295 198.455 ;
        RECT 88.505 197.815 88.735 197.825 ;
        RECT 89.295 197.815 89.525 197.825 ;
        RECT 91.205 197.815 91.435 197.825 ;
        RECT 91.995 197.815 92.225 197.825 ;
        RECT 88.785 197.425 89.245 197.655 ;
        RECT 91.485 197.425 91.945 197.655 ;
        RECT 93.835 195.275 94.205 198.455 ;
        RECT 94.625 195.275 94.995 198.455 ;
        RECT 96.535 195.275 96.905 198.455 ;
        RECT 97.325 195.275 97.695 198.455 ;
        RECT 105.650 196.250 106.650 199.475 ;
        RECT 126.520 199.405 132.130 200.510 ;
        RECT 152.425 200.475 153.425 213.550 ;
        RECT 152.395 199.475 153.455 200.475 ;
        RECT 108.270 198.605 109.310 199.100 ;
        RECT 111.510 198.625 111.970 198.855 ;
        RECT 113.670 198.605 114.710 199.100 ;
        RECT 116.370 198.605 117.410 199.100 ;
        RECT 119.610 198.625 120.070 198.855 ;
        RECT 122.310 198.625 122.770 198.855 ;
        RECT 108.530 198.455 108.760 198.465 ;
        RECT 109.320 198.455 109.550 198.465 ;
        RECT 111.230 198.455 111.460 198.465 ;
        RECT 112.020 198.455 112.250 198.465 ;
        RECT 113.930 198.455 114.160 198.465 ;
        RECT 114.720 198.455 114.950 198.465 ;
        RECT 116.630 198.455 116.860 198.465 ;
        RECT 117.420 198.455 117.650 198.465 ;
        RECT 119.330 198.455 119.560 198.465 ;
        RECT 120.120 198.455 120.350 198.465 ;
        RECT 122.030 198.455 122.260 198.465 ;
        RECT 122.820 198.455 123.050 198.465 ;
        RECT 107.785 197.825 108.830 198.455 ;
        RECT 109.250 197.825 109.620 198.455 ;
        RECT 108.530 197.815 108.760 197.825 ;
        RECT 109.320 197.815 109.550 197.825 ;
        RECT 108.810 197.425 109.270 197.655 ;
        RECT 72.570 193.320 72.940 194.435 ;
        RECT 60.660 191.775 61.120 191.805 ;
        RECT 68.760 191.775 69.220 191.805 ;
        RECT 71.460 191.775 71.920 191.805 ;
        RECT 60.400 191.375 61.400 191.775 ;
        RECT 68.500 191.375 69.500 191.775 ;
        RECT 71.200 191.375 72.200 191.775 ;
        RECT 62.575 189.600 63.575 189.630 ;
        RECT 66.250 189.600 67.250 189.630 ;
        RECT 60.400 189.150 61.400 189.600 ;
        RECT 60.660 189.140 61.120 189.150 ;
        RECT 59.640 186.545 60.010 187.650 ;
        RECT 60.380 183.925 60.610 188.935 ;
        RECT 61.170 183.925 61.400 188.935 ;
        RECT 62.575 188.570 64.500 189.600 ;
        RECT 61.770 187.600 62.140 187.650 ;
        RECT 61.770 186.545 62.875 187.600 ;
        RECT 57.960 180.140 58.420 180.370 ;
        RECT 57.680 179.925 57.910 179.935 ;
        RECT 58.470 179.925 58.700 179.935 ;
        RECT 56.935 178.945 57.980 179.925 ;
        RECT 58.400 178.945 58.770 179.925 ;
        RECT 60.310 178.945 60.680 183.925 ;
        RECT 61.100 178.945 61.470 183.925 ;
        RECT 61.875 181.850 62.875 186.545 ;
        RECT 63.500 183.500 64.500 188.570 ;
        RECT 65.300 188.570 67.250 189.600 ;
        RECT 68.500 189.150 69.500 189.600 ;
        RECT 71.200 189.150 72.200 189.600 ;
        RECT 68.760 189.140 69.220 189.150 ;
        RECT 71.460 189.140 71.920 189.150 ;
        RECT 65.300 184.245 66.300 188.570 ;
        RECT 67.740 187.600 68.110 187.650 ;
        RECT 67.025 186.545 68.110 187.600 ;
        RECT 63.500 182.500 66.330 183.500 ;
        RECT 67.025 181.850 68.025 186.545 ;
        RECT 68.480 183.925 68.710 188.935 ;
        RECT 69.270 183.925 69.500 188.935 ;
        RECT 69.870 186.545 70.240 187.650 ;
        RECT 70.440 186.545 70.810 187.650 ;
        RECT 71.180 183.925 71.410 188.935 ;
        RECT 71.970 183.925 72.200 188.935 ;
        RECT 72.570 186.545 72.940 187.650 ;
        RECT 61.875 180.850 68.025 181.850 ;
        RECT 63.360 180.140 63.820 180.370 ;
        RECT 66.060 180.140 66.520 180.370 ;
        RECT 63.080 179.925 63.310 179.935 ;
        RECT 63.870 179.925 64.100 179.935 ;
        RECT 65.780 179.925 66.010 179.935 ;
        RECT 66.570 179.925 66.800 179.935 ;
        RECT 62.335 178.945 63.380 179.925 ;
        RECT 63.800 178.945 64.170 179.925 ;
        RECT 65.035 178.945 66.080 179.925 ;
        RECT 66.500 178.945 66.870 179.925 ;
        RECT 68.410 178.945 68.780 183.925 ;
        RECT 69.200 178.945 69.570 183.925 ;
        RECT 71.110 178.945 71.480 183.925 ;
        RECT 71.900 178.945 72.270 183.925 ;
        RECT 57.680 178.935 57.910 178.945 ;
        RECT 58.470 178.935 58.700 178.945 ;
        RECT 60.380 178.935 60.610 178.945 ;
        RECT 61.170 178.935 61.400 178.945 ;
        RECT 63.080 178.935 63.310 178.945 ;
        RECT 63.870 178.935 64.100 178.945 ;
        RECT 65.780 178.935 66.010 178.945 ;
        RECT 66.570 178.935 66.800 178.945 ;
        RECT 68.480 178.935 68.710 178.945 ;
        RECT 69.270 178.935 69.500 178.945 ;
        RECT 71.180 178.935 71.410 178.945 ;
        RECT 71.970 178.935 72.200 178.945 ;
        RECT 57.425 178.275 58.460 178.750 ;
        RECT 60.660 178.500 61.120 178.730 ;
        RECT 62.825 178.275 63.860 178.750 ;
        RECT 65.525 178.275 66.560 178.750 ;
        RECT 68.760 178.500 69.220 178.730 ;
        RECT 71.460 178.500 71.920 178.730 ;
        RECT 78.175 177.900 79.175 195.250 ;
        RECT 80.180 194.430 81.295 194.485 ;
        RECT 80.150 193.315 81.325 194.430 ;
        RECT 85.065 193.320 85.435 194.435 ;
        RECT 78.145 176.900 79.205 177.900 ;
        RECT 57.420 176.030 58.460 176.525 ;
        RECT 60.660 176.050 61.120 176.280 ;
        RECT 62.820 176.030 63.860 176.525 ;
        RECT 65.520 176.030 66.560 176.525 ;
        RECT 68.760 176.050 69.220 176.280 ;
        RECT 71.460 176.050 71.920 176.280 ;
        RECT 57.680 175.880 57.910 175.890 ;
        RECT 58.470 175.880 58.700 175.890 ;
        RECT 60.380 175.880 60.610 175.890 ;
        RECT 61.170 175.880 61.400 175.890 ;
        RECT 63.080 175.880 63.310 175.890 ;
        RECT 63.870 175.880 64.100 175.890 ;
        RECT 65.780 175.880 66.010 175.890 ;
        RECT 66.570 175.880 66.800 175.890 ;
        RECT 68.480 175.880 68.710 175.890 ;
        RECT 69.270 175.880 69.500 175.890 ;
        RECT 71.180 175.880 71.410 175.890 ;
        RECT 71.970 175.880 72.200 175.890 ;
        RECT 56.935 175.250 57.980 175.880 ;
        RECT 58.400 175.250 58.770 175.880 ;
        RECT 57.680 175.240 57.910 175.250 ;
        RECT 58.470 175.240 58.700 175.250 ;
        RECT 57.960 174.850 58.420 175.080 ;
        RECT 60.310 172.700 60.680 175.880 ;
        RECT 61.100 172.700 61.470 175.880 ;
        RECT 62.335 175.250 63.380 175.880 ;
        RECT 63.800 175.250 64.170 175.880 ;
        RECT 65.035 175.250 66.080 175.880 ;
        RECT 66.500 175.250 66.870 175.880 ;
        RECT 63.080 175.240 63.310 175.250 ;
        RECT 63.870 175.240 64.100 175.250 ;
        RECT 65.780 175.240 66.010 175.250 ;
        RECT 66.570 175.240 66.800 175.250 ;
        RECT 63.360 174.850 63.820 175.080 ;
        RECT 66.060 174.850 66.520 175.080 ;
        RECT 68.410 172.700 68.780 175.880 ;
        RECT 69.200 172.700 69.570 175.880 ;
        RECT 71.110 172.700 71.480 175.880 ;
        RECT 71.900 172.700 72.270 175.880 ;
        RECT 54.725 170.740 55.900 171.855 ;
        RECT 59.640 170.745 60.010 171.860 ;
        RECT 52.720 154.325 53.780 155.325 ;
        RECT 52.750 154.295 53.750 154.325 ;
        RECT 31.995 153.455 33.035 153.950 ;
        RECT 35.235 153.475 35.695 153.705 ;
        RECT 37.395 153.455 38.435 153.950 ;
        RECT 40.095 153.455 41.135 153.950 ;
        RECT 43.335 153.475 43.795 153.705 ;
        RECT 46.035 153.475 46.495 153.705 ;
        RECT 32.255 153.305 32.485 153.315 ;
        RECT 33.045 153.305 33.275 153.315 ;
        RECT 34.955 153.305 35.185 153.315 ;
        RECT 35.745 153.305 35.975 153.315 ;
        RECT 37.655 153.305 37.885 153.315 ;
        RECT 38.445 153.305 38.675 153.315 ;
        RECT 40.355 153.305 40.585 153.315 ;
        RECT 41.145 153.305 41.375 153.315 ;
        RECT 43.055 153.305 43.285 153.315 ;
        RECT 43.845 153.305 44.075 153.315 ;
        RECT 45.755 153.305 45.985 153.315 ;
        RECT 46.545 153.305 46.775 153.315 ;
        RECT 31.510 152.675 32.555 153.305 ;
        RECT 32.975 152.675 33.345 153.305 ;
        RECT 32.255 152.665 32.485 152.675 ;
        RECT 33.045 152.665 33.275 152.675 ;
        RECT 32.535 152.275 32.995 152.505 ;
        RECT 34.885 150.125 35.255 153.305 ;
        RECT 35.675 150.125 36.045 153.305 ;
        RECT 36.910 152.675 37.955 153.305 ;
        RECT 38.375 152.675 38.745 153.305 ;
        RECT 39.610 152.675 40.655 153.305 ;
        RECT 41.075 152.675 41.445 153.305 ;
        RECT 37.655 152.665 37.885 152.675 ;
        RECT 38.445 152.665 38.675 152.675 ;
        RECT 40.355 152.665 40.585 152.675 ;
        RECT 41.145 152.665 41.375 152.675 ;
        RECT 37.935 152.275 38.395 152.505 ;
        RECT 40.635 152.275 41.095 152.505 ;
        RECT 42.985 150.125 43.355 153.305 ;
        RECT 43.775 150.125 44.145 153.305 ;
        RECT 45.685 150.125 46.055 153.305 ;
        RECT 46.475 150.125 46.845 153.305 ;
        RECT 29.285 148.170 30.485 149.285 ;
        RECT 34.215 148.170 34.585 149.285 ;
        RECT 29.330 148.140 30.445 148.170 ;
        RECT 34.955 146.815 35.185 150.125 ;
        RECT 35.745 146.815 35.975 150.125 ;
        RECT 36.345 148.170 36.715 149.285 ;
        RECT 42.315 148.170 42.685 149.285 ;
        RECT 43.055 146.815 43.285 150.125 ;
        RECT 43.845 146.815 44.075 150.125 ;
        RECT 44.445 148.170 44.815 149.285 ;
        RECT 45.015 148.170 45.385 149.285 ;
        RECT 45.755 146.815 45.985 150.125 ;
        RECT 46.545 146.815 46.775 150.125 ;
        RECT 47.145 148.170 47.515 149.285 ;
        RECT 48.515 148.140 49.630 153.855 ;
        RECT 54.755 149.285 55.870 170.740 ;
        RECT 60.380 169.390 60.610 172.700 ;
        RECT 61.170 169.390 61.400 172.700 ;
        RECT 61.770 170.745 62.140 171.860 ;
        RECT 67.740 170.745 68.110 171.860 ;
        RECT 68.480 169.390 68.710 172.700 ;
        RECT 69.270 169.390 69.500 172.700 ;
        RECT 69.870 170.745 70.240 171.860 ;
        RECT 70.440 170.745 70.810 171.860 ;
        RECT 71.180 169.390 71.410 172.700 ;
        RECT 71.970 169.390 72.200 172.700 ;
        RECT 72.570 170.745 72.940 171.860 ;
        RECT 73.935 170.745 75.110 171.860 ;
        RECT 60.660 169.200 61.120 169.230 ;
        RECT 68.760 169.200 69.220 169.230 ;
        RECT 71.460 169.200 71.920 169.230 ;
        RECT 60.400 168.800 61.400 169.200 ;
        RECT 68.500 168.800 69.500 169.200 ;
        RECT 71.200 168.800 72.200 169.200 ;
        RECT 73.965 167.770 75.080 170.745 ;
        RECT 62.575 167.025 63.575 167.055 ;
        RECT 66.250 167.025 67.250 167.055 ;
        RECT 60.400 166.575 61.400 167.025 ;
        RECT 60.660 166.565 61.120 166.575 ;
        RECT 59.640 163.970 60.010 165.075 ;
        RECT 60.380 161.350 60.610 166.360 ;
        RECT 61.170 161.350 61.400 166.360 ;
        RECT 62.575 165.995 64.500 167.025 ;
        RECT 61.770 165.025 62.140 165.075 ;
        RECT 61.770 163.970 62.875 165.025 ;
        RECT 57.960 157.565 58.420 157.795 ;
        RECT 57.680 157.350 57.910 157.360 ;
        RECT 58.470 157.350 58.700 157.360 ;
        RECT 56.935 156.370 57.980 157.350 ;
        RECT 58.400 156.370 58.770 157.350 ;
        RECT 60.310 156.370 60.680 161.350 ;
        RECT 61.100 156.370 61.470 161.350 ;
        RECT 61.875 159.275 62.875 163.970 ;
        RECT 63.500 160.925 64.500 165.995 ;
        RECT 65.300 165.995 67.250 167.025 ;
        RECT 68.500 166.575 69.500 167.025 ;
        RECT 71.200 166.575 72.200 167.025 ;
        RECT 68.760 166.565 69.220 166.575 ;
        RECT 71.460 166.565 71.920 166.575 ;
        RECT 65.300 161.670 66.300 165.995 ;
        RECT 67.740 165.025 68.110 165.075 ;
        RECT 67.025 163.970 68.110 165.025 ;
        RECT 63.500 159.925 66.330 160.925 ;
        RECT 67.025 159.275 68.025 163.970 ;
        RECT 68.480 161.350 68.710 166.360 ;
        RECT 69.270 161.350 69.500 166.360 ;
        RECT 69.870 163.970 70.240 165.075 ;
        RECT 70.440 163.970 70.810 165.075 ;
        RECT 71.180 161.350 71.410 166.360 ;
        RECT 71.970 161.350 72.200 166.360 ;
        RECT 74.280 165.115 74.730 167.425 ;
        RECT 72.570 163.970 72.940 165.075 ;
        RECT 61.875 158.275 68.025 159.275 ;
        RECT 63.360 157.565 63.820 157.795 ;
        RECT 66.060 157.565 66.520 157.795 ;
        RECT 63.080 157.350 63.310 157.360 ;
        RECT 63.870 157.350 64.100 157.360 ;
        RECT 65.780 157.350 66.010 157.360 ;
        RECT 66.570 157.350 66.800 157.360 ;
        RECT 62.335 156.370 63.380 157.350 ;
        RECT 63.800 156.370 64.170 157.350 ;
        RECT 65.035 156.370 66.080 157.350 ;
        RECT 66.500 156.370 66.870 157.350 ;
        RECT 68.410 156.370 68.780 161.350 ;
        RECT 69.200 156.370 69.570 161.350 ;
        RECT 71.110 156.370 71.480 161.350 ;
        RECT 71.900 156.370 72.270 161.350 ;
        RECT 57.680 156.360 57.910 156.370 ;
        RECT 58.470 156.360 58.700 156.370 ;
        RECT 60.380 156.360 60.610 156.370 ;
        RECT 61.170 156.360 61.400 156.370 ;
        RECT 63.080 156.360 63.310 156.370 ;
        RECT 63.870 156.360 64.100 156.370 ;
        RECT 65.780 156.360 66.010 156.370 ;
        RECT 66.570 156.360 66.800 156.370 ;
        RECT 68.480 156.360 68.710 156.370 ;
        RECT 69.270 156.360 69.500 156.370 ;
        RECT 71.180 156.360 71.410 156.370 ;
        RECT 71.970 156.360 72.200 156.370 ;
        RECT 57.425 155.700 58.460 156.175 ;
        RECT 60.660 155.925 61.120 156.155 ;
        RECT 62.825 155.700 63.860 156.175 ;
        RECT 65.525 155.700 66.560 156.175 ;
        RECT 68.760 155.925 69.220 156.155 ;
        RECT 71.460 155.925 71.920 156.155 ;
        RECT 74.280 154.205 74.730 156.515 ;
        RECT 78.175 155.325 79.175 176.900 ;
        RECT 80.180 171.855 81.295 193.315 ;
        RECT 85.805 191.965 86.035 195.275 ;
        RECT 86.595 191.965 86.825 195.275 ;
        RECT 87.195 193.320 87.565 194.435 ;
        RECT 93.165 193.320 93.535 194.435 ;
        RECT 93.905 191.965 94.135 195.275 ;
        RECT 94.695 191.965 94.925 195.275 ;
        RECT 95.295 193.320 95.665 194.435 ;
        RECT 95.865 193.320 96.235 194.435 ;
        RECT 96.605 191.965 96.835 195.275 ;
        RECT 97.395 191.965 97.625 195.275 ;
        RECT 103.600 195.250 106.650 196.250 ;
        RECT 111.160 195.275 111.530 198.455 ;
        RECT 111.950 195.275 112.320 198.455 ;
        RECT 113.185 197.825 114.230 198.455 ;
        RECT 114.650 197.825 115.020 198.455 ;
        RECT 115.885 197.825 116.930 198.455 ;
        RECT 117.350 197.825 117.720 198.455 ;
        RECT 113.930 197.815 114.160 197.825 ;
        RECT 114.720 197.815 114.950 197.825 ;
        RECT 116.630 197.815 116.860 197.825 ;
        RECT 117.420 197.815 117.650 197.825 ;
        RECT 114.210 197.425 114.670 197.655 ;
        RECT 116.910 197.425 117.370 197.655 ;
        RECT 119.260 195.275 119.630 198.455 ;
        RECT 120.050 195.275 120.420 198.455 ;
        RECT 121.960 195.275 122.330 198.455 ;
        RECT 122.750 195.275 123.120 198.455 ;
        RECT 131.075 196.250 132.075 199.405 ;
        RECT 133.695 198.605 134.735 199.100 ;
        RECT 136.935 198.625 137.395 198.855 ;
        RECT 139.095 198.605 140.135 199.100 ;
        RECT 141.795 198.605 142.835 199.100 ;
        RECT 145.035 198.625 145.495 198.855 ;
        RECT 147.735 198.625 148.195 198.855 ;
        RECT 133.955 198.455 134.185 198.465 ;
        RECT 134.745 198.455 134.975 198.465 ;
        RECT 136.655 198.455 136.885 198.465 ;
        RECT 137.445 198.455 137.675 198.465 ;
        RECT 139.355 198.455 139.585 198.465 ;
        RECT 140.145 198.455 140.375 198.465 ;
        RECT 142.055 198.455 142.285 198.465 ;
        RECT 142.845 198.455 143.075 198.465 ;
        RECT 144.755 198.455 144.985 198.465 ;
        RECT 145.545 198.455 145.775 198.465 ;
        RECT 147.455 198.455 147.685 198.465 ;
        RECT 148.245 198.455 148.475 198.465 ;
        RECT 133.210 197.825 134.255 198.455 ;
        RECT 134.675 197.825 135.045 198.455 ;
        RECT 133.955 197.815 134.185 197.825 ;
        RECT 134.745 197.815 134.975 197.825 ;
        RECT 134.235 197.425 134.695 197.655 ;
        RECT 97.995 193.320 98.365 194.435 ;
        RECT 86.085 191.775 86.545 191.805 ;
        RECT 94.185 191.775 94.645 191.805 ;
        RECT 96.885 191.775 97.345 191.805 ;
        RECT 85.825 191.375 86.825 191.775 ;
        RECT 93.925 191.375 94.925 191.775 ;
        RECT 96.625 191.375 97.625 191.775 ;
        RECT 88.000 189.600 89.000 189.630 ;
        RECT 91.675 189.600 92.675 189.630 ;
        RECT 85.825 189.150 86.825 189.600 ;
        RECT 86.085 189.140 86.545 189.150 ;
        RECT 85.065 186.545 85.435 187.650 ;
        RECT 85.805 183.925 86.035 188.935 ;
        RECT 86.595 183.925 86.825 188.935 ;
        RECT 88.000 188.570 89.925 189.600 ;
        RECT 87.195 187.600 87.565 187.650 ;
        RECT 87.195 186.545 88.300 187.600 ;
        RECT 83.385 180.140 83.845 180.370 ;
        RECT 83.105 179.925 83.335 179.935 ;
        RECT 83.895 179.925 84.125 179.935 ;
        RECT 82.360 178.945 83.405 179.925 ;
        RECT 83.825 178.945 84.195 179.925 ;
        RECT 85.735 178.945 86.105 183.925 ;
        RECT 86.525 178.945 86.895 183.925 ;
        RECT 87.300 181.850 88.300 186.545 ;
        RECT 88.925 183.500 89.925 188.570 ;
        RECT 90.725 188.570 92.675 189.600 ;
        RECT 93.925 189.150 94.925 189.600 ;
        RECT 96.625 189.150 97.625 189.600 ;
        RECT 94.185 189.140 94.645 189.150 ;
        RECT 96.885 189.140 97.345 189.150 ;
        RECT 90.725 184.245 91.725 188.570 ;
        RECT 93.165 187.600 93.535 187.650 ;
        RECT 92.450 186.545 93.535 187.600 ;
        RECT 88.925 182.500 91.755 183.500 ;
        RECT 92.450 181.850 93.450 186.545 ;
        RECT 93.905 183.925 94.135 188.935 ;
        RECT 94.695 183.925 94.925 188.935 ;
        RECT 95.295 186.545 95.665 187.650 ;
        RECT 95.865 186.545 96.235 187.650 ;
        RECT 96.605 183.925 96.835 188.935 ;
        RECT 97.395 183.925 97.625 188.935 ;
        RECT 97.995 186.545 98.365 187.650 ;
        RECT 87.300 180.850 93.450 181.850 ;
        RECT 88.785 180.140 89.245 180.370 ;
        RECT 91.485 180.140 91.945 180.370 ;
        RECT 88.505 179.925 88.735 179.935 ;
        RECT 89.295 179.925 89.525 179.935 ;
        RECT 91.205 179.925 91.435 179.935 ;
        RECT 91.995 179.925 92.225 179.935 ;
        RECT 87.760 178.945 88.805 179.925 ;
        RECT 89.225 178.945 89.595 179.925 ;
        RECT 90.460 178.945 91.505 179.925 ;
        RECT 91.925 178.945 92.295 179.925 ;
        RECT 93.835 178.945 94.205 183.925 ;
        RECT 94.625 178.945 94.995 183.925 ;
        RECT 96.535 178.945 96.905 183.925 ;
        RECT 97.325 178.945 97.695 183.925 ;
        RECT 83.105 178.935 83.335 178.945 ;
        RECT 83.895 178.935 84.125 178.945 ;
        RECT 85.805 178.935 86.035 178.945 ;
        RECT 86.595 178.935 86.825 178.945 ;
        RECT 88.505 178.935 88.735 178.945 ;
        RECT 89.295 178.935 89.525 178.945 ;
        RECT 91.205 178.935 91.435 178.945 ;
        RECT 91.995 178.935 92.225 178.945 ;
        RECT 93.905 178.935 94.135 178.945 ;
        RECT 94.695 178.935 94.925 178.945 ;
        RECT 96.605 178.935 96.835 178.945 ;
        RECT 97.395 178.935 97.625 178.945 ;
        RECT 82.850 178.275 83.885 178.750 ;
        RECT 86.085 178.500 86.545 178.730 ;
        RECT 88.250 178.275 89.285 178.750 ;
        RECT 90.950 178.275 91.985 178.750 ;
        RECT 94.185 178.500 94.645 178.730 ;
        RECT 96.885 178.500 97.345 178.730 ;
        RECT 103.600 177.900 104.600 195.250 ;
        RECT 105.605 194.430 106.720 194.485 ;
        RECT 105.575 193.315 106.750 194.430 ;
        RECT 110.490 193.320 110.860 194.435 ;
        RECT 103.570 176.900 104.630 177.900 ;
        RECT 82.845 176.030 83.885 176.525 ;
        RECT 86.085 176.050 86.545 176.280 ;
        RECT 88.245 176.030 89.285 176.525 ;
        RECT 90.945 176.030 91.985 176.525 ;
        RECT 94.185 176.050 94.645 176.280 ;
        RECT 96.885 176.050 97.345 176.280 ;
        RECT 83.105 175.880 83.335 175.890 ;
        RECT 83.895 175.880 84.125 175.890 ;
        RECT 85.805 175.880 86.035 175.890 ;
        RECT 86.595 175.880 86.825 175.890 ;
        RECT 88.505 175.880 88.735 175.890 ;
        RECT 89.295 175.880 89.525 175.890 ;
        RECT 91.205 175.880 91.435 175.890 ;
        RECT 91.995 175.880 92.225 175.890 ;
        RECT 93.905 175.880 94.135 175.890 ;
        RECT 94.695 175.880 94.925 175.890 ;
        RECT 96.605 175.880 96.835 175.890 ;
        RECT 97.395 175.880 97.625 175.890 ;
        RECT 82.360 175.250 83.405 175.880 ;
        RECT 83.825 175.250 84.195 175.880 ;
        RECT 83.105 175.240 83.335 175.250 ;
        RECT 83.895 175.240 84.125 175.250 ;
        RECT 83.385 174.850 83.845 175.080 ;
        RECT 85.735 172.700 86.105 175.880 ;
        RECT 86.525 172.700 86.895 175.880 ;
        RECT 87.760 175.250 88.805 175.880 ;
        RECT 89.225 175.250 89.595 175.880 ;
        RECT 90.460 175.250 91.505 175.880 ;
        RECT 91.925 175.250 92.295 175.880 ;
        RECT 88.505 175.240 88.735 175.250 ;
        RECT 89.295 175.240 89.525 175.250 ;
        RECT 91.205 175.240 91.435 175.250 ;
        RECT 91.995 175.240 92.225 175.250 ;
        RECT 88.785 174.850 89.245 175.080 ;
        RECT 91.485 174.850 91.945 175.080 ;
        RECT 93.835 172.700 94.205 175.880 ;
        RECT 94.625 172.700 94.995 175.880 ;
        RECT 96.535 172.700 96.905 175.880 ;
        RECT 97.325 172.700 97.695 175.880 ;
        RECT 80.150 170.740 81.325 171.855 ;
        RECT 85.065 170.745 85.435 171.860 ;
        RECT 78.145 154.325 79.205 155.325 ;
        RECT 78.175 154.295 79.175 154.325 ;
        RECT 57.420 153.455 58.460 153.950 ;
        RECT 60.660 153.475 61.120 153.705 ;
        RECT 62.820 153.455 63.860 153.950 ;
        RECT 65.520 153.455 66.560 153.950 ;
        RECT 68.760 153.475 69.220 153.705 ;
        RECT 71.460 153.475 71.920 153.705 ;
        RECT 57.680 153.305 57.910 153.315 ;
        RECT 58.470 153.305 58.700 153.315 ;
        RECT 60.380 153.305 60.610 153.315 ;
        RECT 61.170 153.305 61.400 153.315 ;
        RECT 63.080 153.305 63.310 153.315 ;
        RECT 63.870 153.305 64.100 153.315 ;
        RECT 65.780 153.305 66.010 153.315 ;
        RECT 66.570 153.305 66.800 153.315 ;
        RECT 68.480 153.305 68.710 153.315 ;
        RECT 69.270 153.305 69.500 153.315 ;
        RECT 71.180 153.305 71.410 153.315 ;
        RECT 71.970 153.305 72.200 153.315 ;
        RECT 56.935 152.675 57.980 153.305 ;
        RECT 58.400 152.675 58.770 153.305 ;
        RECT 57.680 152.665 57.910 152.675 ;
        RECT 58.470 152.665 58.700 152.675 ;
        RECT 57.960 152.275 58.420 152.505 ;
        RECT 60.310 150.125 60.680 153.305 ;
        RECT 61.100 150.125 61.470 153.305 ;
        RECT 62.335 152.675 63.380 153.305 ;
        RECT 63.800 152.675 64.170 153.305 ;
        RECT 65.035 152.675 66.080 153.305 ;
        RECT 66.500 152.675 66.870 153.305 ;
        RECT 63.080 152.665 63.310 152.675 ;
        RECT 63.870 152.665 64.100 152.675 ;
        RECT 65.780 152.665 66.010 152.675 ;
        RECT 66.570 152.665 66.800 152.675 ;
        RECT 63.360 152.275 63.820 152.505 ;
        RECT 66.060 152.275 66.520 152.505 ;
        RECT 68.410 150.125 68.780 153.305 ;
        RECT 69.200 150.125 69.570 153.305 ;
        RECT 71.110 150.125 71.480 153.305 ;
        RECT 71.900 150.125 72.270 153.305 ;
        RECT 54.710 148.170 55.910 149.285 ;
        RECT 59.640 148.170 60.010 149.285 ;
        RECT 54.755 148.140 55.870 148.170 ;
        RECT 60.380 146.815 60.610 150.125 ;
        RECT 61.170 146.815 61.400 150.125 ;
        RECT 61.770 148.170 62.140 149.285 ;
        RECT 67.740 148.170 68.110 149.285 ;
        RECT 68.480 146.815 68.710 150.125 ;
        RECT 69.270 146.815 69.500 150.125 ;
        RECT 69.870 148.170 70.240 149.285 ;
        RECT 70.440 148.170 70.810 149.285 ;
        RECT 71.180 146.815 71.410 150.125 ;
        RECT 71.970 146.815 72.200 150.125 ;
        RECT 72.570 148.170 72.940 149.285 ;
        RECT 73.940 148.140 75.055 153.855 ;
        RECT 80.180 149.285 81.295 170.740 ;
        RECT 85.805 169.390 86.035 172.700 ;
        RECT 86.595 169.390 86.825 172.700 ;
        RECT 87.195 170.745 87.565 171.860 ;
        RECT 93.165 170.745 93.535 171.860 ;
        RECT 93.905 169.390 94.135 172.700 ;
        RECT 94.695 169.390 94.925 172.700 ;
        RECT 95.295 170.745 95.665 171.860 ;
        RECT 95.865 170.745 96.235 171.860 ;
        RECT 96.605 169.390 96.835 172.700 ;
        RECT 97.395 169.390 97.625 172.700 ;
        RECT 97.995 170.745 98.365 171.860 ;
        RECT 99.360 170.745 100.535 171.860 ;
        RECT 86.085 169.200 86.545 169.230 ;
        RECT 94.185 169.200 94.645 169.230 ;
        RECT 96.885 169.200 97.345 169.230 ;
        RECT 85.825 168.800 86.825 169.200 ;
        RECT 93.925 168.800 94.925 169.200 ;
        RECT 96.625 168.800 97.625 169.200 ;
        RECT 99.390 167.770 100.505 170.745 ;
        RECT 88.000 167.025 89.000 167.055 ;
        RECT 91.675 167.025 92.675 167.055 ;
        RECT 85.825 166.575 86.825 167.025 ;
        RECT 86.085 166.565 86.545 166.575 ;
        RECT 85.065 163.970 85.435 165.075 ;
        RECT 85.805 161.350 86.035 166.360 ;
        RECT 86.595 161.350 86.825 166.360 ;
        RECT 88.000 165.995 89.925 167.025 ;
        RECT 87.195 165.025 87.565 165.075 ;
        RECT 87.195 163.970 88.300 165.025 ;
        RECT 83.385 157.565 83.845 157.795 ;
        RECT 83.105 157.350 83.335 157.360 ;
        RECT 83.895 157.350 84.125 157.360 ;
        RECT 82.360 156.370 83.405 157.350 ;
        RECT 83.825 156.370 84.195 157.350 ;
        RECT 85.735 156.370 86.105 161.350 ;
        RECT 86.525 156.370 86.895 161.350 ;
        RECT 87.300 159.275 88.300 163.970 ;
        RECT 88.925 160.925 89.925 165.995 ;
        RECT 90.725 165.995 92.675 167.025 ;
        RECT 93.925 166.575 94.925 167.025 ;
        RECT 96.625 166.575 97.625 167.025 ;
        RECT 94.185 166.565 94.645 166.575 ;
        RECT 96.885 166.565 97.345 166.575 ;
        RECT 90.725 161.670 91.725 165.995 ;
        RECT 93.165 165.025 93.535 165.075 ;
        RECT 92.450 163.970 93.535 165.025 ;
        RECT 88.925 159.925 91.755 160.925 ;
        RECT 92.450 159.275 93.450 163.970 ;
        RECT 93.905 161.350 94.135 166.360 ;
        RECT 94.695 161.350 94.925 166.360 ;
        RECT 95.295 163.970 95.665 165.075 ;
        RECT 95.865 163.970 96.235 165.075 ;
        RECT 96.605 161.350 96.835 166.360 ;
        RECT 97.395 161.350 97.625 166.360 ;
        RECT 99.705 165.115 100.155 167.425 ;
        RECT 97.995 163.970 98.365 165.075 ;
        RECT 87.300 158.275 93.450 159.275 ;
        RECT 88.785 157.565 89.245 157.795 ;
        RECT 91.485 157.565 91.945 157.795 ;
        RECT 88.505 157.350 88.735 157.360 ;
        RECT 89.295 157.350 89.525 157.360 ;
        RECT 91.205 157.350 91.435 157.360 ;
        RECT 91.995 157.350 92.225 157.360 ;
        RECT 87.760 156.370 88.805 157.350 ;
        RECT 89.225 156.370 89.595 157.350 ;
        RECT 90.460 156.370 91.505 157.350 ;
        RECT 91.925 156.370 92.295 157.350 ;
        RECT 93.835 156.370 94.205 161.350 ;
        RECT 94.625 156.370 94.995 161.350 ;
        RECT 96.535 156.370 96.905 161.350 ;
        RECT 97.325 156.370 97.695 161.350 ;
        RECT 83.105 156.360 83.335 156.370 ;
        RECT 83.895 156.360 84.125 156.370 ;
        RECT 85.805 156.360 86.035 156.370 ;
        RECT 86.595 156.360 86.825 156.370 ;
        RECT 88.505 156.360 88.735 156.370 ;
        RECT 89.295 156.360 89.525 156.370 ;
        RECT 91.205 156.360 91.435 156.370 ;
        RECT 91.995 156.360 92.225 156.370 ;
        RECT 93.905 156.360 94.135 156.370 ;
        RECT 94.695 156.360 94.925 156.370 ;
        RECT 96.605 156.360 96.835 156.370 ;
        RECT 97.395 156.360 97.625 156.370 ;
        RECT 82.850 155.700 83.885 156.175 ;
        RECT 86.085 155.925 86.545 156.155 ;
        RECT 88.250 155.700 89.285 156.175 ;
        RECT 90.950 155.700 91.985 156.175 ;
        RECT 94.185 155.925 94.645 156.155 ;
        RECT 96.885 155.925 97.345 156.155 ;
        RECT 99.705 154.205 100.155 156.515 ;
        RECT 103.600 155.325 104.600 176.900 ;
        RECT 105.605 171.855 106.720 193.315 ;
        RECT 111.230 191.965 111.460 195.275 ;
        RECT 112.020 191.965 112.250 195.275 ;
        RECT 112.620 193.320 112.990 194.435 ;
        RECT 118.590 193.320 118.960 194.435 ;
        RECT 119.330 191.965 119.560 195.275 ;
        RECT 120.120 191.965 120.350 195.275 ;
        RECT 120.720 193.320 121.090 194.435 ;
        RECT 121.290 193.320 121.660 194.435 ;
        RECT 122.030 191.965 122.260 195.275 ;
        RECT 122.820 191.965 123.050 195.275 ;
        RECT 129.025 195.250 132.075 196.250 ;
        RECT 136.585 195.275 136.955 198.455 ;
        RECT 137.375 195.275 137.745 198.455 ;
        RECT 138.610 197.825 139.655 198.455 ;
        RECT 140.075 197.825 140.445 198.455 ;
        RECT 141.310 197.825 142.355 198.455 ;
        RECT 142.775 197.825 143.145 198.455 ;
        RECT 139.355 197.815 139.585 197.825 ;
        RECT 140.145 197.815 140.375 197.825 ;
        RECT 142.055 197.815 142.285 197.825 ;
        RECT 142.845 197.815 143.075 197.825 ;
        RECT 139.635 197.425 140.095 197.655 ;
        RECT 142.335 197.425 142.795 197.655 ;
        RECT 144.685 195.275 145.055 198.455 ;
        RECT 145.475 195.275 145.845 198.455 ;
        RECT 147.385 195.275 147.755 198.455 ;
        RECT 148.175 195.275 148.545 198.455 ;
        RECT 123.420 193.320 123.790 194.435 ;
        RECT 111.510 191.775 111.970 191.805 ;
        RECT 119.610 191.775 120.070 191.805 ;
        RECT 122.310 191.775 122.770 191.805 ;
        RECT 111.250 191.375 112.250 191.775 ;
        RECT 119.350 191.375 120.350 191.775 ;
        RECT 122.050 191.375 123.050 191.775 ;
        RECT 113.425 189.600 114.425 189.630 ;
        RECT 117.100 189.600 118.100 189.630 ;
        RECT 111.250 189.150 112.250 189.600 ;
        RECT 111.510 189.140 111.970 189.150 ;
        RECT 110.490 186.545 110.860 187.650 ;
        RECT 111.230 183.925 111.460 188.935 ;
        RECT 112.020 183.925 112.250 188.935 ;
        RECT 113.425 188.570 115.350 189.600 ;
        RECT 112.620 187.600 112.990 187.650 ;
        RECT 112.620 186.545 113.725 187.600 ;
        RECT 108.810 180.140 109.270 180.370 ;
        RECT 108.530 179.925 108.760 179.935 ;
        RECT 109.320 179.925 109.550 179.935 ;
        RECT 107.785 178.945 108.830 179.925 ;
        RECT 109.250 178.945 109.620 179.925 ;
        RECT 111.160 178.945 111.530 183.925 ;
        RECT 111.950 178.945 112.320 183.925 ;
        RECT 112.725 181.850 113.725 186.545 ;
        RECT 114.350 183.500 115.350 188.570 ;
        RECT 116.150 188.570 118.100 189.600 ;
        RECT 119.350 189.150 120.350 189.600 ;
        RECT 122.050 189.150 123.050 189.600 ;
        RECT 119.610 189.140 120.070 189.150 ;
        RECT 122.310 189.140 122.770 189.150 ;
        RECT 116.150 184.245 117.150 188.570 ;
        RECT 118.590 187.600 118.960 187.650 ;
        RECT 117.875 186.545 118.960 187.600 ;
        RECT 114.350 182.500 117.180 183.500 ;
        RECT 117.875 181.850 118.875 186.545 ;
        RECT 119.330 183.925 119.560 188.935 ;
        RECT 120.120 183.925 120.350 188.935 ;
        RECT 120.720 186.545 121.090 187.650 ;
        RECT 121.290 186.545 121.660 187.650 ;
        RECT 122.030 183.925 122.260 188.935 ;
        RECT 122.820 183.925 123.050 188.935 ;
        RECT 123.420 186.545 123.790 187.650 ;
        RECT 112.725 180.850 118.875 181.850 ;
        RECT 114.210 180.140 114.670 180.370 ;
        RECT 116.910 180.140 117.370 180.370 ;
        RECT 113.930 179.925 114.160 179.935 ;
        RECT 114.720 179.925 114.950 179.935 ;
        RECT 116.630 179.925 116.860 179.935 ;
        RECT 117.420 179.925 117.650 179.935 ;
        RECT 113.185 178.945 114.230 179.925 ;
        RECT 114.650 178.945 115.020 179.925 ;
        RECT 115.885 178.945 116.930 179.925 ;
        RECT 117.350 178.945 117.720 179.925 ;
        RECT 119.260 178.945 119.630 183.925 ;
        RECT 120.050 178.945 120.420 183.925 ;
        RECT 121.960 178.945 122.330 183.925 ;
        RECT 122.750 178.945 123.120 183.925 ;
        RECT 108.530 178.935 108.760 178.945 ;
        RECT 109.320 178.935 109.550 178.945 ;
        RECT 111.230 178.935 111.460 178.945 ;
        RECT 112.020 178.935 112.250 178.945 ;
        RECT 113.930 178.935 114.160 178.945 ;
        RECT 114.720 178.935 114.950 178.945 ;
        RECT 116.630 178.935 116.860 178.945 ;
        RECT 117.420 178.935 117.650 178.945 ;
        RECT 119.330 178.935 119.560 178.945 ;
        RECT 120.120 178.935 120.350 178.945 ;
        RECT 122.030 178.935 122.260 178.945 ;
        RECT 122.820 178.935 123.050 178.945 ;
        RECT 108.275 178.275 109.310 178.750 ;
        RECT 111.510 178.500 111.970 178.730 ;
        RECT 113.675 178.275 114.710 178.750 ;
        RECT 116.375 178.275 117.410 178.750 ;
        RECT 119.610 178.500 120.070 178.730 ;
        RECT 122.310 178.500 122.770 178.730 ;
        RECT 129.025 177.900 130.025 195.250 ;
        RECT 131.030 194.430 132.145 194.485 ;
        RECT 131.000 193.315 132.175 194.430 ;
        RECT 135.915 193.320 136.285 194.435 ;
        RECT 128.995 176.900 130.055 177.900 ;
        RECT 108.270 176.030 109.310 176.525 ;
        RECT 111.510 176.050 111.970 176.280 ;
        RECT 113.670 176.030 114.710 176.525 ;
        RECT 116.370 176.030 117.410 176.525 ;
        RECT 119.610 176.050 120.070 176.280 ;
        RECT 122.310 176.050 122.770 176.280 ;
        RECT 108.530 175.880 108.760 175.890 ;
        RECT 109.320 175.880 109.550 175.890 ;
        RECT 111.230 175.880 111.460 175.890 ;
        RECT 112.020 175.880 112.250 175.890 ;
        RECT 113.930 175.880 114.160 175.890 ;
        RECT 114.720 175.880 114.950 175.890 ;
        RECT 116.630 175.880 116.860 175.890 ;
        RECT 117.420 175.880 117.650 175.890 ;
        RECT 119.330 175.880 119.560 175.890 ;
        RECT 120.120 175.880 120.350 175.890 ;
        RECT 122.030 175.880 122.260 175.890 ;
        RECT 122.820 175.880 123.050 175.890 ;
        RECT 107.785 175.250 108.830 175.880 ;
        RECT 109.250 175.250 109.620 175.880 ;
        RECT 108.530 175.240 108.760 175.250 ;
        RECT 109.320 175.240 109.550 175.250 ;
        RECT 108.810 174.850 109.270 175.080 ;
        RECT 111.160 172.700 111.530 175.880 ;
        RECT 111.950 172.700 112.320 175.880 ;
        RECT 113.185 175.250 114.230 175.880 ;
        RECT 114.650 175.250 115.020 175.880 ;
        RECT 115.885 175.250 116.930 175.880 ;
        RECT 117.350 175.250 117.720 175.880 ;
        RECT 113.930 175.240 114.160 175.250 ;
        RECT 114.720 175.240 114.950 175.250 ;
        RECT 116.630 175.240 116.860 175.250 ;
        RECT 117.420 175.240 117.650 175.250 ;
        RECT 114.210 174.850 114.670 175.080 ;
        RECT 116.910 174.850 117.370 175.080 ;
        RECT 119.260 172.700 119.630 175.880 ;
        RECT 120.050 172.700 120.420 175.880 ;
        RECT 121.960 172.700 122.330 175.880 ;
        RECT 122.750 172.700 123.120 175.880 ;
        RECT 105.575 170.740 106.750 171.855 ;
        RECT 110.490 170.745 110.860 171.860 ;
        RECT 103.570 154.325 104.630 155.325 ;
        RECT 103.600 154.295 104.600 154.325 ;
        RECT 82.845 153.455 83.885 153.950 ;
        RECT 86.085 153.475 86.545 153.705 ;
        RECT 88.245 153.455 89.285 153.950 ;
        RECT 90.945 153.455 91.985 153.950 ;
        RECT 94.185 153.475 94.645 153.705 ;
        RECT 96.885 153.475 97.345 153.705 ;
        RECT 83.105 153.305 83.335 153.315 ;
        RECT 83.895 153.305 84.125 153.315 ;
        RECT 85.805 153.305 86.035 153.315 ;
        RECT 86.595 153.305 86.825 153.315 ;
        RECT 88.505 153.305 88.735 153.315 ;
        RECT 89.295 153.305 89.525 153.315 ;
        RECT 91.205 153.305 91.435 153.315 ;
        RECT 91.995 153.305 92.225 153.315 ;
        RECT 93.905 153.305 94.135 153.315 ;
        RECT 94.695 153.305 94.925 153.315 ;
        RECT 96.605 153.305 96.835 153.315 ;
        RECT 97.395 153.305 97.625 153.315 ;
        RECT 82.360 152.675 83.405 153.305 ;
        RECT 83.825 152.675 84.195 153.305 ;
        RECT 83.105 152.665 83.335 152.675 ;
        RECT 83.895 152.665 84.125 152.675 ;
        RECT 83.385 152.275 83.845 152.505 ;
        RECT 85.735 150.125 86.105 153.305 ;
        RECT 86.525 150.125 86.895 153.305 ;
        RECT 87.760 152.675 88.805 153.305 ;
        RECT 89.225 152.675 89.595 153.305 ;
        RECT 90.460 152.675 91.505 153.305 ;
        RECT 91.925 152.675 92.295 153.305 ;
        RECT 88.505 152.665 88.735 152.675 ;
        RECT 89.295 152.665 89.525 152.675 ;
        RECT 91.205 152.665 91.435 152.675 ;
        RECT 91.995 152.665 92.225 152.675 ;
        RECT 88.785 152.275 89.245 152.505 ;
        RECT 91.485 152.275 91.945 152.505 ;
        RECT 93.835 150.125 94.205 153.305 ;
        RECT 94.625 150.125 94.995 153.305 ;
        RECT 96.535 150.125 96.905 153.305 ;
        RECT 97.325 150.125 97.695 153.305 ;
        RECT 80.135 148.170 81.335 149.285 ;
        RECT 85.065 148.170 85.435 149.285 ;
        RECT 80.180 148.140 81.295 148.170 ;
        RECT 85.805 146.815 86.035 150.125 ;
        RECT 86.595 146.815 86.825 150.125 ;
        RECT 87.195 148.170 87.565 149.285 ;
        RECT 93.165 148.170 93.535 149.285 ;
        RECT 93.905 146.815 94.135 150.125 ;
        RECT 94.695 146.815 94.925 150.125 ;
        RECT 95.295 148.170 95.665 149.285 ;
        RECT 95.865 148.170 96.235 149.285 ;
        RECT 96.605 146.815 96.835 150.125 ;
        RECT 97.395 146.815 97.625 150.125 ;
        RECT 97.995 148.170 98.365 149.285 ;
        RECT 99.365 148.140 100.480 153.855 ;
        RECT 105.605 149.285 106.720 170.740 ;
        RECT 111.230 169.390 111.460 172.700 ;
        RECT 112.020 169.390 112.250 172.700 ;
        RECT 112.620 170.745 112.990 171.860 ;
        RECT 118.590 170.745 118.960 171.860 ;
        RECT 119.330 169.390 119.560 172.700 ;
        RECT 120.120 169.390 120.350 172.700 ;
        RECT 120.720 170.745 121.090 171.860 ;
        RECT 121.290 170.745 121.660 171.860 ;
        RECT 122.030 169.390 122.260 172.700 ;
        RECT 122.820 169.390 123.050 172.700 ;
        RECT 123.420 170.745 123.790 171.860 ;
        RECT 124.785 170.745 125.960 171.860 ;
        RECT 111.510 169.200 111.970 169.230 ;
        RECT 119.610 169.200 120.070 169.230 ;
        RECT 122.310 169.200 122.770 169.230 ;
        RECT 111.250 168.800 112.250 169.200 ;
        RECT 119.350 168.800 120.350 169.200 ;
        RECT 122.050 168.800 123.050 169.200 ;
        RECT 124.815 167.770 125.930 170.745 ;
        RECT 113.425 167.025 114.425 167.055 ;
        RECT 117.100 167.025 118.100 167.055 ;
        RECT 111.250 166.575 112.250 167.025 ;
        RECT 111.510 166.565 111.970 166.575 ;
        RECT 110.490 163.970 110.860 165.075 ;
        RECT 111.230 161.350 111.460 166.360 ;
        RECT 112.020 161.350 112.250 166.360 ;
        RECT 113.425 165.995 115.350 167.025 ;
        RECT 112.620 165.025 112.990 165.075 ;
        RECT 112.620 163.970 113.725 165.025 ;
        RECT 108.810 157.565 109.270 157.795 ;
        RECT 108.530 157.350 108.760 157.360 ;
        RECT 109.320 157.350 109.550 157.360 ;
        RECT 107.785 156.370 108.830 157.350 ;
        RECT 109.250 156.370 109.620 157.350 ;
        RECT 111.160 156.370 111.530 161.350 ;
        RECT 111.950 156.370 112.320 161.350 ;
        RECT 112.725 159.275 113.725 163.970 ;
        RECT 114.350 160.925 115.350 165.995 ;
        RECT 116.150 165.995 118.100 167.025 ;
        RECT 119.350 166.575 120.350 167.025 ;
        RECT 122.050 166.575 123.050 167.025 ;
        RECT 119.610 166.565 120.070 166.575 ;
        RECT 122.310 166.565 122.770 166.575 ;
        RECT 116.150 161.670 117.150 165.995 ;
        RECT 118.590 165.025 118.960 165.075 ;
        RECT 117.875 163.970 118.960 165.025 ;
        RECT 114.350 159.925 117.180 160.925 ;
        RECT 117.875 159.275 118.875 163.970 ;
        RECT 119.330 161.350 119.560 166.360 ;
        RECT 120.120 161.350 120.350 166.360 ;
        RECT 120.720 163.970 121.090 165.075 ;
        RECT 121.290 163.970 121.660 165.075 ;
        RECT 122.030 161.350 122.260 166.360 ;
        RECT 122.820 161.350 123.050 166.360 ;
        RECT 125.130 165.115 125.580 167.425 ;
        RECT 123.420 163.970 123.790 165.075 ;
        RECT 112.725 158.275 118.875 159.275 ;
        RECT 114.210 157.565 114.670 157.795 ;
        RECT 116.910 157.565 117.370 157.795 ;
        RECT 113.930 157.350 114.160 157.360 ;
        RECT 114.720 157.350 114.950 157.360 ;
        RECT 116.630 157.350 116.860 157.360 ;
        RECT 117.420 157.350 117.650 157.360 ;
        RECT 113.185 156.370 114.230 157.350 ;
        RECT 114.650 156.370 115.020 157.350 ;
        RECT 115.885 156.370 116.930 157.350 ;
        RECT 117.350 156.370 117.720 157.350 ;
        RECT 119.260 156.370 119.630 161.350 ;
        RECT 120.050 156.370 120.420 161.350 ;
        RECT 121.960 156.370 122.330 161.350 ;
        RECT 122.750 156.370 123.120 161.350 ;
        RECT 108.530 156.360 108.760 156.370 ;
        RECT 109.320 156.360 109.550 156.370 ;
        RECT 111.230 156.360 111.460 156.370 ;
        RECT 112.020 156.360 112.250 156.370 ;
        RECT 113.930 156.360 114.160 156.370 ;
        RECT 114.720 156.360 114.950 156.370 ;
        RECT 116.630 156.360 116.860 156.370 ;
        RECT 117.420 156.360 117.650 156.370 ;
        RECT 119.330 156.360 119.560 156.370 ;
        RECT 120.120 156.360 120.350 156.370 ;
        RECT 122.030 156.360 122.260 156.370 ;
        RECT 122.820 156.360 123.050 156.370 ;
        RECT 108.275 155.700 109.310 156.175 ;
        RECT 111.510 155.925 111.970 156.155 ;
        RECT 113.675 155.700 114.710 156.175 ;
        RECT 116.375 155.700 117.410 156.175 ;
        RECT 119.610 155.925 120.070 156.155 ;
        RECT 122.310 155.925 122.770 156.155 ;
        RECT 125.130 154.205 125.580 156.515 ;
        RECT 129.025 155.325 130.025 176.900 ;
        RECT 131.030 171.855 132.145 193.315 ;
        RECT 136.655 191.965 136.885 195.275 ;
        RECT 137.445 191.965 137.675 195.275 ;
        RECT 138.045 193.320 138.415 194.435 ;
        RECT 144.015 193.320 144.385 194.435 ;
        RECT 144.755 191.965 144.985 195.275 ;
        RECT 145.545 191.965 145.775 195.275 ;
        RECT 146.145 193.320 146.515 194.435 ;
        RECT 146.715 193.320 147.085 194.435 ;
        RECT 147.455 191.965 147.685 195.275 ;
        RECT 148.245 191.965 148.475 195.275 ;
        RECT 148.845 193.320 149.215 194.435 ;
        RECT 136.935 191.775 137.395 191.805 ;
        RECT 145.035 191.775 145.495 191.805 ;
        RECT 147.735 191.775 148.195 191.805 ;
        RECT 136.675 191.375 137.675 191.775 ;
        RECT 144.775 191.375 145.775 191.775 ;
        RECT 147.475 191.375 148.475 191.775 ;
        RECT 138.850 189.600 139.850 189.630 ;
        RECT 142.525 189.600 143.525 189.630 ;
        RECT 136.675 189.150 137.675 189.600 ;
        RECT 136.935 189.140 137.395 189.150 ;
        RECT 135.915 186.545 136.285 187.650 ;
        RECT 136.655 183.925 136.885 188.935 ;
        RECT 137.445 183.925 137.675 188.935 ;
        RECT 138.850 188.570 140.775 189.600 ;
        RECT 138.045 187.600 138.415 187.650 ;
        RECT 138.045 186.545 139.150 187.600 ;
        RECT 134.235 180.140 134.695 180.370 ;
        RECT 133.955 179.925 134.185 179.935 ;
        RECT 134.745 179.925 134.975 179.935 ;
        RECT 133.210 178.945 134.255 179.925 ;
        RECT 134.675 178.945 135.045 179.925 ;
        RECT 136.585 178.945 136.955 183.925 ;
        RECT 137.375 178.945 137.745 183.925 ;
        RECT 138.150 181.850 139.150 186.545 ;
        RECT 139.775 183.500 140.775 188.570 ;
        RECT 141.575 188.570 143.525 189.600 ;
        RECT 144.775 189.150 145.775 189.600 ;
        RECT 147.475 189.150 148.475 189.600 ;
        RECT 145.035 189.140 145.495 189.150 ;
        RECT 147.735 189.140 148.195 189.150 ;
        RECT 141.575 184.245 142.575 188.570 ;
        RECT 144.015 187.600 144.385 187.650 ;
        RECT 143.300 186.545 144.385 187.600 ;
        RECT 139.775 182.500 142.605 183.500 ;
        RECT 143.300 181.850 144.300 186.545 ;
        RECT 144.755 183.925 144.985 188.935 ;
        RECT 145.545 183.925 145.775 188.935 ;
        RECT 146.145 186.545 146.515 187.650 ;
        RECT 146.715 186.545 147.085 187.650 ;
        RECT 147.455 183.925 147.685 188.935 ;
        RECT 148.245 183.925 148.475 188.935 ;
        RECT 148.845 186.545 149.215 187.650 ;
        RECT 138.150 180.850 144.300 181.850 ;
        RECT 139.635 180.140 140.095 180.370 ;
        RECT 142.335 180.140 142.795 180.370 ;
        RECT 139.355 179.925 139.585 179.935 ;
        RECT 140.145 179.925 140.375 179.935 ;
        RECT 142.055 179.925 142.285 179.935 ;
        RECT 142.845 179.925 143.075 179.935 ;
        RECT 138.610 178.945 139.655 179.925 ;
        RECT 140.075 178.945 140.445 179.925 ;
        RECT 141.310 178.945 142.355 179.925 ;
        RECT 142.775 178.945 143.145 179.925 ;
        RECT 144.685 178.945 145.055 183.925 ;
        RECT 145.475 178.945 145.845 183.925 ;
        RECT 147.385 178.945 147.755 183.925 ;
        RECT 148.175 178.945 148.545 183.925 ;
        RECT 133.955 178.935 134.185 178.945 ;
        RECT 134.745 178.935 134.975 178.945 ;
        RECT 136.655 178.935 136.885 178.945 ;
        RECT 137.445 178.935 137.675 178.945 ;
        RECT 139.355 178.935 139.585 178.945 ;
        RECT 140.145 178.935 140.375 178.945 ;
        RECT 142.055 178.935 142.285 178.945 ;
        RECT 142.845 178.935 143.075 178.945 ;
        RECT 144.755 178.935 144.985 178.945 ;
        RECT 145.545 178.935 145.775 178.945 ;
        RECT 147.455 178.935 147.685 178.945 ;
        RECT 148.245 178.935 148.475 178.945 ;
        RECT 133.700 178.275 134.735 178.750 ;
        RECT 136.935 178.500 137.395 178.730 ;
        RECT 139.100 178.275 140.135 178.750 ;
        RECT 141.800 178.275 142.835 178.750 ;
        RECT 145.035 178.500 145.495 178.730 ;
        RECT 147.735 178.500 148.195 178.730 ;
        RECT 133.695 176.030 134.735 176.525 ;
        RECT 136.935 176.050 137.395 176.280 ;
        RECT 139.095 176.030 140.135 176.525 ;
        RECT 141.795 176.030 142.835 176.525 ;
        RECT 145.035 176.050 145.495 176.280 ;
        RECT 147.735 176.050 148.195 176.280 ;
        RECT 133.955 175.880 134.185 175.890 ;
        RECT 134.745 175.880 134.975 175.890 ;
        RECT 136.655 175.880 136.885 175.890 ;
        RECT 137.445 175.880 137.675 175.890 ;
        RECT 139.355 175.880 139.585 175.890 ;
        RECT 140.145 175.880 140.375 175.890 ;
        RECT 142.055 175.880 142.285 175.890 ;
        RECT 142.845 175.880 143.075 175.890 ;
        RECT 144.755 175.880 144.985 175.890 ;
        RECT 145.545 175.880 145.775 175.890 ;
        RECT 147.455 175.880 147.685 175.890 ;
        RECT 148.245 175.880 148.475 175.890 ;
        RECT 133.210 175.250 134.255 175.880 ;
        RECT 134.675 175.250 135.045 175.880 ;
        RECT 133.955 175.240 134.185 175.250 ;
        RECT 134.745 175.240 134.975 175.250 ;
        RECT 134.235 174.850 134.695 175.080 ;
        RECT 136.585 172.700 136.955 175.880 ;
        RECT 137.375 172.700 137.745 175.880 ;
        RECT 138.610 175.250 139.655 175.880 ;
        RECT 140.075 175.250 140.445 175.880 ;
        RECT 141.310 175.250 142.355 175.880 ;
        RECT 142.775 175.250 143.145 175.880 ;
        RECT 139.355 175.240 139.585 175.250 ;
        RECT 140.145 175.240 140.375 175.250 ;
        RECT 142.055 175.240 142.285 175.250 ;
        RECT 142.845 175.240 143.075 175.250 ;
        RECT 139.635 174.850 140.095 175.080 ;
        RECT 142.335 174.850 142.795 175.080 ;
        RECT 144.685 172.700 145.055 175.880 ;
        RECT 145.475 172.700 145.845 175.880 ;
        RECT 147.385 172.700 147.755 175.880 ;
        RECT 148.175 172.700 148.545 175.880 ;
        RECT 131.000 170.740 132.175 171.855 ;
        RECT 135.915 170.745 136.285 171.860 ;
        RECT 128.995 154.325 130.055 155.325 ;
        RECT 129.025 154.295 130.025 154.325 ;
        RECT 108.270 153.455 109.310 153.950 ;
        RECT 111.510 153.475 111.970 153.705 ;
        RECT 113.670 153.455 114.710 153.950 ;
        RECT 116.370 153.455 117.410 153.950 ;
        RECT 119.610 153.475 120.070 153.705 ;
        RECT 122.310 153.475 122.770 153.705 ;
        RECT 108.530 153.305 108.760 153.315 ;
        RECT 109.320 153.305 109.550 153.315 ;
        RECT 111.230 153.305 111.460 153.315 ;
        RECT 112.020 153.305 112.250 153.315 ;
        RECT 113.930 153.305 114.160 153.315 ;
        RECT 114.720 153.305 114.950 153.315 ;
        RECT 116.630 153.305 116.860 153.315 ;
        RECT 117.420 153.305 117.650 153.315 ;
        RECT 119.330 153.305 119.560 153.315 ;
        RECT 120.120 153.305 120.350 153.315 ;
        RECT 122.030 153.305 122.260 153.315 ;
        RECT 122.820 153.305 123.050 153.315 ;
        RECT 107.785 152.675 108.830 153.305 ;
        RECT 109.250 152.675 109.620 153.305 ;
        RECT 108.530 152.665 108.760 152.675 ;
        RECT 109.320 152.665 109.550 152.675 ;
        RECT 108.810 152.275 109.270 152.505 ;
        RECT 111.160 150.125 111.530 153.305 ;
        RECT 111.950 150.125 112.320 153.305 ;
        RECT 113.185 152.675 114.230 153.305 ;
        RECT 114.650 152.675 115.020 153.305 ;
        RECT 115.885 152.675 116.930 153.305 ;
        RECT 117.350 152.675 117.720 153.305 ;
        RECT 113.930 152.665 114.160 152.675 ;
        RECT 114.720 152.665 114.950 152.675 ;
        RECT 116.630 152.665 116.860 152.675 ;
        RECT 117.420 152.665 117.650 152.675 ;
        RECT 114.210 152.275 114.670 152.505 ;
        RECT 116.910 152.275 117.370 152.505 ;
        RECT 119.260 150.125 119.630 153.305 ;
        RECT 120.050 150.125 120.420 153.305 ;
        RECT 121.960 150.125 122.330 153.305 ;
        RECT 122.750 150.125 123.120 153.305 ;
        RECT 105.560 148.170 106.760 149.285 ;
        RECT 110.490 148.170 110.860 149.285 ;
        RECT 105.605 148.140 106.720 148.170 ;
        RECT 111.230 146.815 111.460 150.125 ;
        RECT 112.020 146.815 112.250 150.125 ;
        RECT 112.620 148.170 112.990 149.285 ;
        RECT 118.590 148.170 118.960 149.285 ;
        RECT 119.330 146.815 119.560 150.125 ;
        RECT 120.120 146.815 120.350 150.125 ;
        RECT 120.720 148.170 121.090 149.285 ;
        RECT 121.290 148.170 121.660 149.285 ;
        RECT 122.030 146.815 122.260 150.125 ;
        RECT 122.820 146.815 123.050 150.125 ;
        RECT 123.420 148.170 123.790 149.285 ;
        RECT 124.790 148.140 125.905 153.855 ;
        RECT 131.030 149.285 132.145 170.740 ;
        RECT 136.655 169.390 136.885 172.700 ;
        RECT 137.445 169.390 137.675 172.700 ;
        RECT 138.045 170.745 138.415 171.860 ;
        RECT 144.015 170.745 144.385 171.860 ;
        RECT 144.755 169.390 144.985 172.700 ;
        RECT 145.545 169.390 145.775 172.700 ;
        RECT 146.145 170.745 146.515 171.860 ;
        RECT 146.715 170.745 147.085 171.860 ;
        RECT 147.455 169.390 147.685 172.700 ;
        RECT 148.245 169.390 148.475 172.700 ;
        RECT 148.845 170.745 149.215 171.860 ;
        RECT 150.210 170.745 151.385 171.860 ;
        RECT 136.935 169.200 137.395 169.230 ;
        RECT 145.035 169.200 145.495 169.230 ;
        RECT 147.735 169.200 148.195 169.230 ;
        RECT 136.675 168.800 137.675 169.200 ;
        RECT 144.775 168.800 145.775 169.200 ;
        RECT 147.475 168.800 148.475 169.200 ;
        RECT 150.240 167.770 151.355 170.745 ;
        RECT 138.850 167.025 139.850 167.055 ;
        RECT 142.525 167.025 143.525 167.055 ;
        RECT 136.675 166.575 137.675 167.025 ;
        RECT 136.935 166.565 137.395 166.575 ;
        RECT 135.915 163.970 136.285 165.075 ;
        RECT 136.655 161.350 136.885 166.360 ;
        RECT 137.445 161.350 137.675 166.360 ;
        RECT 138.850 165.995 140.775 167.025 ;
        RECT 138.045 165.025 138.415 165.075 ;
        RECT 138.045 163.970 139.150 165.025 ;
        RECT 134.235 157.565 134.695 157.795 ;
        RECT 133.955 157.350 134.185 157.360 ;
        RECT 134.745 157.350 134.975 157.360 ;
        RECT 133.210 156.370 134.255 157.350 ;
        RECT 134.675 156.370 135.045 157.350 ;
        RECT 136.585 156.370 136.955 161.350 ;
        RECT 137.375 156.370 137.745 161.350 ;
        RECT 138.150 159.275 139.150 163.970 ;
        RECT 139.775 160.925 140.775 165.995 ;
        RECT 141.575 165.995 143.525 167.025 ;
        RECT 144.775 166.575 145.775 167.025 ;
        RECT 147.475 166.575 148.475 167.025 ;
        RECT 145.035 166.565 145.495 166.575 ;
        RECT 147.735 166.565 148.195 166.575 ;
        RECT 141.575 161.670 142.575 165.995 ;
        RECT 144.015 165.025 144.385 165.075 ;
        RECT 143.300 163.970 144.385 165.025 ;
        RECT 139.775 159.925 142.605 160.925 ;
        RECT 143.300 159.275 144.300 163.970 ;
        RECT 144.755 161.350 144.985 166.360 ;
        RECT 145.545 161.350 145.775 166.360 ;
        RECT 146.145 163.970 146.515 165.075 ;
        RECT 146.715 163.970 147.085 165.075 ;
        RECT 147.455 161.350 147.685 166.360 ;
        RECT 148.245 161.350 148.475 166.360 ;
        RECT 150.555 165.115 151.005 167.425 ;
        RECT 148.845 163.970 149.215 165.075 ;
        RECT 138.150 158.275 144.300 159.275 ;
        RECT 139.635 157.565 140.095 157.795 ;
        RECT 142.335 157.565 142.795 157.795 ;
        RECT 139.355 157.350 139.585 157.360 ;
        RECT 140.145 157.350 140.375 157.360 ;
        RECT 142.055 157.350 142.285 157.360 ;
        RECT 142.845 157.350 143.075 157.360 ;
        RECT 138.610 156.370 139.655 157.350 ;
        RECT 140.075 156.370 140.445 157.350 ;
        RECT 141.310 156.370 142.355 157.350 ;
        RECT 142.775 156.370 143.145 157.350 ;
        RECT 144.685 156.370 145.055 161.350 ;
        RECT 145.475 156.370 145.845 161.350 ;
        RECT 147.385 156.370 147.755 161.350 ;
        RECT 148.175 156.370 148.545 161.350 ;
        RECT 133.955 156.360 134.185 156.370 ;
        RECT 134.745 156.360 134.975 156.370 ;
        RECT 136.655 156.360 136.885 156.370 ;
        RECT 137.445 156.360 137.675 156.370 ;
        RECT 139.355 156.360 139.585 156.370 ;
        RECT 140.145 156.360 140.375 156.370 ;
        RECT 142.055 156.360 142.285 156.370 ;
        RECT 142.845 156.360 143.075 156.370 ;
        RECT 144.755 156.360 144.985 156.370 ;
        RECT 145.545 156.360 145.775 156.370 ;
        RECT 147.455 156.360 147.685 156.370 ;
        RECT 148.245 156.360 148.475 156.370 ;
        RECT 133.700 155.700 134.735 156.175 ;
        RECT 136.935 155.925 137.395 156.155 ;
        RECT 139.100 155.700 140.135 156.175 ;
        RECT 141.800 155.700 142.835 156.175 ;
        RECT 145.035 155.925 145.495 156.155 ;
        RECT 147.735 155.925 148.195 156.155 ;
        RECT 150.555 154.205 151.005 156.515 ;
        RECT 133.695 153.455 134.735 153.950 ;
        RECT 136.935 153.475 137.395 153.705 ;
        RECT 139.095 153.455 140.135 153.950 ;
        RECT 141.795 153.455 142.835 153.950 ;
        RECT 145.035 153.475 145.495 153.705 ;
        RECT 147.735 153.475 148.195 153.705 ;
        RECT 133.955 153.305 134.185 153.315 ;
        RECT 134.745 153.305 134.975 153.315 ;
        RECT 136.655 153.305 136.885 153.315 ;
        RECT 137.445 153.305 137.675 153.315 ;
        RECT 139.355 153.305 139.585 153.315 ;
        RECT 140.145 153.305 140.375 153.315 ;
        RECT 142.055 153.305 142.285 153.315 ;
        RECT 142.845 153.305 143.075 153.315 ;
        RECT 144.755 153.305 144.985 153.315 ;
        RECT 145.545 153.305 145.775 153.315 ;
        RECT 147.455 153.305 147.685 153.315 ;
        RECT 148.245 153.305 148.475 153.315 ;
        RECT 133.210 152.675 134.255 153.305 ;
        RECT 134.675 152.675 135.045 153.305 ;
        RECT 133.955 152.665 134.185 152.675 ;
        RECT 134.745 152.665 134.975 152.675 ;
        RECT 134.235 152.275 134.695 152.505 ;
        RECT 136.585 150.125 136.955 153.305 ;
        RECT 137.375 150.125 137.745 153.305 ;
        RECT 138.610 152.675 139.655 153.305 ;
        RECT 140.075 152.675 140.445 153.305 ;
        RECT 141.310 152.675 142.355 153.305 ;
        RECT 142.775 152.675 143.145 153.305 ;
        RECT 139.355 152.665 139.585 152.675 ;
        RECT 140.145 152.665 140.375 152.675 ;
        RECT 142.055 152.665 142.285 152.675 ;
        RECT 142.845 152.665 143.075 152.675 ;
        RECT 139.635 152.275 140.095 152.505 ;
        RECT 142.335 152.275 142.795 152.505 ;
        RECT 144.685 150.125 145.055 153.305 ;
        RECT 145.475 150.125 145.845 153.305 ;
        RECT 147.385 150.125 147.755 153.305 ;
        RECT 148.175 150.125 148.545 153.305 ;
        RECT 130.985 148.170 132.185 149.285 ;
        RECT 135.915 148.170 136.285 149.285 ;
        RECT 131.030 148.140 132.145 148.170 ;
        RECT 136.655 146.815 136.885 150.125 ;
        RECT 137.445 146.815 137.675 150.125 ;
        RECT 138.045 148.170 138.415 149.285 ;
        RECT 144.015 148.170 144.385 149.285 ;
        RECT 144.755 146.815 144.985 150.125 ;
        RECT 145.545 146.815 145.775 150.125 ;
        RECT 146.145 148.170 146.515 149.285 ;
        RECT 146.715 148.170 147.085 149.285 ;
        RECT 147.455 146.815 147.685 150.125 ;
        RECT 148.245 146.815 148.475 150.125 ;
        RECT 148.845 148.170 149.215 149.285 ;
        RECT 150.215 148.140 151.330 153.855 ;
        RECT 9.810 146.625 10.270 146.655 ;
        RECT 17.910 146.625 18.370 146.655 ;
        RECT 20.610 146.625 21.070 146.655 ;
        RECT 35.235 146.625 35.695 146.655 ;
        RECT 43.335 146.625 43.795 146.655 ;
        RECT 46.035 146.625 46.495 146.655 ;
        RECT 60.660 146.625 61.120 146.655 ;
        RECT 68.760 146.625 69.220 146.655 ;
        RECT 71.460 146.625 71.920 146.655 ;
        RECT 86.085 146.625 86.545 146.655 ;
        RECT 94.185 146.625 94.645 146.655 ;
        RECT 96.885 146.625 97.345 146.655 ;
        RECT 111.510 146.625 111.970 146.655 ;
        RECT 119.610 146.625 120.070 146.655 ;
        RECT 122.310 146.625 122.770 146.655 ;
        RECT 136.935 146.625 137.395 146.655 ;
        RECT 145.035 146.625 145.495 146.655 ;
        RECT 147.735 146.625 148.195 146.655 ;
        RECT 9.550 146.225 10.550 146.625 ;
        RECT 17.650 146.225 18.650 146.625 ;
        RECT 20.350 146.225 21.350 146.625 ;
        RECT 34.975 146.225 35.975 146.625 ;
        RECT 43.075 146.225 44.075 146.625 ;
        RECT 45.775 146.225 46.775 146.625 ;
        RECT 60.400 146.225 61.400 146.625 ;
        RECT 68.500 146.225 69.500 146.625 ;
        RECT 71.200 146.225 72.200 146.625 ;
        RECT 85.825 146.225 86.825 146.625 ;
        RECT 93.925 146.225 94.925 146.625 ;
        RECT 96.625 146.225 97.625 146.625 ;
        RECT 111.250 146.225 112.250 146.625 ;
        RECT 119.350 146.225 120.350 146.625 ;
        RECT 122.050 146.225 123.050 146.625 ;
        RECT 136.675 146.225 137.675 146.625 ;
        RECT 144.775 146.225 145.775 146.625 ;
        RECT 147.475 146.225 148.475 146.625 ;
        RECT 7.500 141.550 153.425 142.550 ;
        RECT 11.725 140.175 12.725 140.205 ;
        RECT 15.400 140.175 16.400 140.205 ;
        RECT 37.150 140.175 38.150 140.205 ;
        RECT 40.825 140.175 41.825 140.205 ;
        RECT 9.550 139.725 10.550 140.175 ;
        RECT 9.810 139.715 10.270 139.725 ;
        RECT 8.790 137.120 9.160 138.225 ;
        RECT 9.530 134.500 9.760 139.510 ;
        RECT 10.320 134.500 10.550 139.510 ;
        RECT 11.725 139.145 13.650 140.175 ;
        RECT 10.920 138.175 11.290 138.225 ;
        RECT 10.920 137.120 12.025 138.175 ;
        RECT 7.110 130.715 7.570 130.945 ;
        RECT 6.830 130.500 7.060 130.510 ;
        RECT 7.620 130.500 7.850 130.510 ;
        RECT 6.085 129.520 7.130 130.500 ;
        RECT 7.550 129.520 7.920 130.500 ;
        RECT 9.460 129.520 9.830 134.500 ;
        RECT 10.250 129.520 10.620 134.500 ;
        RECT 11.025 132.425 12.025 137.120 ;
        RECT 12.650 134.075 13.650 139.145 ;
        RECT 14.450 139.145 16.400 140.175 ;
        RECT 17.650 139.725 18.650 140.175 ;
        RECT 20.350 139.725 21.350 140.175 ;
        RECT 27.270 139.975 28.270 140.125 ;
        RECT 17.910 139.715 18.370 139.725 ;
        RECT 20.610 139.715 21.070 139.725 ;
        RECT 23.805 139.715 24.265 139.945 ;
        RECT 26.505 139.715 26.965 139.945 ;
        RECT 27.120 139.525 28.270 139.975 ;
        RECT 29.205 139.715 29.665 139.945 ;
        RECT 34.975 139.725 35.975 140.175 ;
        RECT 35.235 139.715 35.695 139.725 ;
        RECT 14.450 134.820 15.450 139.145 ;
        RECT 16.890 138.175 17.260 138.225 ;
        RECT 16.175 137.120 17.260 138.175 ;
        RECT 12.650 133.075 15.480 134.075 ;
        RECT 16.175 132.425 17.175 137.120 ;
        RECT 17.630 134.500 17.860 139.510 ;
        RECT 18.420 134.500 18.650 139.510 ;
        RECT 19.020 137.120 19.390 138.225 ;
        RECT 19.590 137.120 19.960 138.225 ;
        RECT 20.330 134.500 20.560 139.510 ;
        RECT 21.120 134.500 21.350 139.510 ;
        RECT 23.525 138.510 23.755 139.510 ;
        RECT 24.295 138.495 26.475 139.525 ;
        RECT 26.970 139.500 28.270 139.525 ;
        RECT 28.925 139.500 29.155 139.510 ;
        RECT 29.715 139.500 29.945 139.510 ;
        RECT 26.970 138.975 29.225 139.500 ;
        RECT 26.970 138.570 27.890 138.975 ;
        RECT 27.015 138.510 27.245 138.570 ;
        RECT 28.180 138.520 29.225 138.975 ;
        RECT 29.645 138.520 30.015 139.500 ;
        RECT 28.925 138.510 29.155 138.520 ;
        RECT 29.715 138.510 29.945 138.520 ;
        RECT 21.720 137.120 22.090 138.225 ;
        RECT 23.520 135.625 24.520 138.355 ;
        RECT 26.245 135.625 27.245 138.325 ;
        RECT 28.670 137.850 29.705 138.325 ;
        RECT 34.215 137.120 34.585 138.225 ;
        RECT 28.665 135.605 29.705 136.100 ;
        RECT 23.205 134.800 23.850 135.480 ;
        RECT 24.245 134.800 26.525 135.480 ;
        RECT 27.015 135.405 27.245 135.465 ;
        RECT 28.925 135.455 29.155 135.465 ;
        RECT 29.715 135.455 29.945 135.465 ;
        RECT 26.970 135.250 27.890 135.405 ;
        RECT 28.180 135.250 29.225 135.455 ;
        RECT 26.970 134.825 29.225 135.250 ;
        RECT 29.645 134.825 30.015 135.455 ;
        RECT 27.015 134.815 28.270 134.825 ;
        RECT 28.925 134.815 29.155 134.825 ;
        RECT 29.715 134.815 29.945 134.825 ;
        RECT 27.020 134.800 28.270 134.815 ;
        RECT 11.025 131.425 17.175 132.425 ;
        RECT 12.510 130.715 12.970 130.945 ;
        RECT 15.210 130.715 15.670 130.945 ;
        RECT 12.230 130.500 12.460 130.510 ;
        RECT 13.020 130.500 13.250 130.510 ;
        RECT 14.930 130.500 15.160 130.510 ;
        RECT 15.720 130.500 15.950 130.510 ;
        RECT 11.485 129.520 12.530 130.500 ;
        RECT 12.950 129.520 13.320 130.500 ;
        RECT 14.185 129.520 15.230 130.500 ;
        RECT 15.650 129.520 16.020 130.500 ;
        RECT 17.560 129.520 17.930 134.500 ;
        RECT 18.350 129.520 18.720 134.500 ;
        RECT 20.260 129.520 20.630 134.500 ;
        RECT 21.050 129.520 21.420 134.500 ;
        RECT 23.805 134.425 24.265 134.655 ;
        RECT 26.505 134.425 26.965 134.655 ;
        RECT 27.115 134.250 28.270 134.800 ;
        RECT 29.205 134.425 29.665 134.655 ;
        RECT 34.955 134.500 35.185 139.510 ;
        RECT 35.745 134.500 35.975 139.510 ;
        RECT 37.150 139.145 39.075 140.175 ;
        RECT 36.345 138.175 36.715 138.225 ;
        RECT 36.345 137.120 37.450 138.175 ;
        RECT 27.115 134.200 28.175 134.250 ;
        RECT 6.830 129.510 7.060 129.520 ;
        RECT 7.620 129.510 7.850 129.520 ;
        RECT 9.530 129.510 9.760 129.520 ;
        RECT 10.320 129.510 10.550 129.520 ;
        RECT 12.230 129.510 12.460 129.520 ;
        RECT 13.020 129.510 13.250 129.520 ;
        RECT 14.930 129.510 15.160 129.520 ;
        RECT 15.720 129.510 15.950 129.520 ;
        RECT 17.630 129.510 17.860 129.520 ;
        RECT 18.420 129.510 18.650 129.520 ;
        RECT 20.330 129.510 20.560 129.520 ;
        RECT 21.120 129.510 21.350 129.520 ;
        RECT 6.575 128.850 7.610 129.325 ;
        RECT 9.810 129.075 10.270 129.305 ;
        RECT 11.975 128.850 13.010 129.325 ;
        RECT 14.675 128.850 15.710 129.325 ;
        RECT 17.910 129.075 18.370 129.305 ;
        RECT 20.610 129.075 21.070 129.305 ;
        RECT 3.950 128.475 4.950 128.530 ;
        RECT 24.820 128.510 25.925 133.180 ;
        RECT 32.535 130.715 32.995 130.945 ;
        RECT 32.255 130.500 32.485 130.510 ;
        RECT 33.045 130.500 33.275 130.510 ;
        RECT 31.510 129.520 32.555 130.500 ;
        RECT 32.975 129.520 33.345 130.500 ;
        RECT 34.885 129.520 35.255 134.500 ;
        RECT 35.675 129.520 36.045 134.500 ;
        RECT 36.450 132.425 37.450 137.120 ;
        RECT 38.075 134.075 39.075 139.145 ;
        RECT 39.875 139.145 41.825 140.175 ;
        RECT 43.075 139.725 44.075 140.175 ;
        RECT 45.775 139.725 46.775 140.175 ;
        RECT 43.335 139.715 43.795 139.725 ;
        RECT 46.035 139.715 46.495 139.725 ;
        RECT 39.875 134.820 40.875 139.145 ;
        RECT 42.315 138.175 42.685 138.225 ;
        RECT 41.600 137.120 42.685 138.175 ;
        RECT 38.075 133.075 40.905 134.075 ;
        RECT 41.600 132.425 42.600 137.120 ;
        RECT 43.055 134.500 43.285 139.510 ;
        RECT 43.845 134.500 44.075 139.510 ;
        RECT 44.445 137.120 44.815 138.225 ;
        RECT 45.015 137.120 45.385 138.225 ;
        RECT 45.755 134.500 45.985 139.510 ;
        RECT 46.545 134.500 46.775 139.510 ;
        RECT 47.145 137.120 47.515 138.225 ;
        RECT 36.450 131.425 42.600 132.425 ;
        RECT 37.935 130.715 38.395 130.945 ;
        RECT 40.635 130.715 41.095 130.945 ;
        RECT 37.655 130.500 37.885 130.510 ;
        RECT 38.445 130.500 38.675 130.510 ;
        RECT 40.355 130.500 40.585 130.510 ;
        RECT 41.145 130.500 41.375 130.510 ;
        RECT 36.910 129.520 37.955 130.500 ;
        RECT 38.375 129.520 38.745 130.500 ;
        RECT 39.610 129.520 40.655 130.500 ;
        RECT 41.075 129.520 41.445 130.500 ;
        RECT 42.985 129.520 43.355 134.500 ;
        RECT 43.775 129.520 44.145 134.500 ;
        RECT 45.685 129.520 46.055 134.500 ;
        RECT 46.475 129.520 46.845 134.500 ;
        RECT 32.255 129.510 32.485 129.520 ;
        RECT 33.045 129.510 33.275 129.520 ;
        RECT 34.955 129.510 35.185 129.520 ;
        RECT 35.745 129.510 35.975 129.520 ;
        RECT 37.655 129.510 37.885 129.520 ;
        RECT 38.445 129.510 38.675 129.520 ;
        RECT 40.355 129.510 40.585 129.520 ;
        RECT 41.145 129.510 41.375 129.520 ;
        RECT 43.055 129.510 43.285 129.520 ;
        RECT 43.845 129.510 44.075 129.520 ;
        RECT 45.755 129.510 45.985 129.520 ;
        RECT 46.545 129.510 46.775 129.520 ;
        RECT 32.000 128.850 33.035 129.325 ;
        RECT 35.235 129.075 35.695 129.305 ;
        RECT 37.400 128.850 38.435 129.325 ;
        RECT 40.100 128.850 41.135 129.325 ;
        RECT 43.335 129.075 43.795 129.305 ;
        RECT 46.035 129.075 46.495 129.305 ;
        RECT 29.375 128.510 30.375 128.530 ;
        RECT 3.920 127.475 4.980 128.475 ;
        RECT 3.950 124.250 4.950 127.475 ;
        RECT 24.820 127.405 30.430 128.510 ;
        RECT 50.725 128.475 51.725 141.550 ;
        RECT 62.575 140.175 63.575 140.205 ;
        RECT 66.250 140.175 67.250 140.205 ;
        RECT 88.000 140.175 89.000 140.205 ;
        RECT 91.675 140.175 92.675 140.205 ;
        RECT 60.400 139.725 61.400 140.175 ;
        RECT 60.660 139.715 61.120 139.725 ;
        RECT 59.640 137.120 60.010 138.225 ;
        RECT 60.380 134.500 60.610 139.510 ;
        RECT 61.170 134.500 61.400 139.510 ;
        RECT 62.575 139.145 64.500 140.175 ;
        RECT 61.770 138.175 62.140 138.225 ;
        RECT 61.770 137.120 62.875 138.175 ;
        RECT 57.960 130.715 58.420 130.945 ;
        RECT 57.680 130.500 57.910 130.510 ;
        RECT 58.470 130.500 58.700 130.510 ;
        RECT 56.935 129.520 57.980 130.500 ;
        RECT 58.400 129.520 58.770 130.500 ;
        RECT 60.310 129.520 60.680 134.500 ;
        RECT 61.100 129.520 61.470 134.500 ;
        RECT 61.875 132.425 62.875 137.120 ;
        RECT 63.500 134.075 64.500 139.145 ;
        RECT 65.300 139.145 67.250 140.175 ;
        RECT 68.500 139.725 69.500 140.175 ;
        RECT 71.200 139.725 72.200 140.175 ;
        RECT 78.120 139.975 79.120 140.125 ;
        RECT 68.760 139.715 69.220 139.725 ;
        RECT 71.460 139.715 71.920 139.725 ;
        RECT 74.655 139.715 75.115 139.945 ;
        RECT 77.355 139.715 77.815 139.945 ;
        RECT 77.970 139.525 79.120 139.975 ;
        RECT 80.055 139.715 80.515 139.945 ;
        RECT 85.825 139.725 86.825 140.175 ;
        RECT 86.085 139.715 86.545 139.725 ;
        RECT 65.300 134.820 66.300 139.145 ;
        RECT 67.740 138.175 68.110 138.225 ;
        RECT 67.025 137.120 68.110 138.175 ;
        RECT 63.500 133.075 66.330 134.075 ;
        RECT 67.025 132.425 68.025 137.120 ;
        RECT 68.480 134.500 68.710 139.510 ;
        RECT 69.270 134.500 69.500 139.510 ;
        RECT 69.870 137.120 70.240 138.225 ;
        RECT 70.440 137.120 70.810 138.225 ;
        RECT 71.180 134.500 71.410 139.510 ;
        RECT 71.970 134.500 72.200 139.510 ;
        RECT 74.375 138.510 74.605 139.510 ;
        RECT 75.145 138.495 77.325 139.525 ;
        RECT 77.820 139.500 79.120 139.525 ;
        RECT 79.775 139.500 80.005 139.510 ;
        RECT 80.565 139.500 80.795 139.510 ;
        RECT 77.820 138.975 80.075 139.500 ;
        RECT 77.820 138.570 78.740 138.975 ;
        RECT 77.865 138.510 78.095 138.570 ;
        RECT 79.030 138.520 80.075 138.975 ;
        RECT 80.495 138.520 80.865 139.500 ;
        RECT 79.775 138.510 80.005 138.520 ;
        RECT 80.565 138.510 80.795 138.520 ;
        RECT 72.570 137.120 72.940 138.225 ;
        RECT 74.370 135.625 75.370 138.355 ;
        RECT 77.095 135.625 78.095 138.325 ;
        RECT 79.520 137.850 80.555 138.325 ;
        RECT 85.065 137.120 85.435 138.225 ;
        RECT 79.515 135.605 80.555 136.100 ;
        RECT 74.055 134.800 74.700 135.480 ;
        RECT 75.095 134.800 77.375 135.480 ;
        RECT 77.865 135.405 78.095 135.465 ;
        RECT 79.775 135.455 80.005 135.465 ;
        RECT 80.565 135.455 80.795 135.465 ;
        RECT 77.820 135.250 78.740 135.405 ;
        RECT 79.030 135.250 80.075 135.455 ;
        RECT 77.820 134.825 80.075 135.250 ;
        RECT 80.495 134.825 80.865 135.455 ;
        RECT 77.865 134.815 79.120 134.825 ;
        RECT 79.775 134.815 80.005 134.825 ;
        RECT 80.565 134.815 80.795 134.825 ;
        RECT 77.870 134.800 79.120 134.815 ;
        RECT 61.875 131.425 68.025 132.425 ;
        RECT 63.360 130.715 63.820 130.945 ;
        RECT 66.060 130.715 66.520 130.945 ;
        RECT 63.080 130.500 63.310 130.510 ;
        RECT 63.870 130.500 64.100 130.510 ;
        RECT 65.780 130.500 66.010 130.510 ;
        RECT 66.570 130.500 66.800 130.510 ;
        RECT 62.335 129.520 63.380 130.500 ;
        RECT 63.800 129.520 64.170 130.500 ;
        RECT 65.035 129.520 66.080 130.500 ;
        RECT 66.500 129.520 66.870 130.500 ;
        RECT 68.410 129.520 68.780 134.500 ;
        RECT 69.200 129.520 69.570 134.500 ;
        RECT 71.110 129.520 71.480 134.500 ;
        RECT 71.900 129.520 72.270 134.500 ;
        RECT 74.655 134.425 75.115 134.655 ;
        RECT 77.355 134.425 77.815 134.655 ;
        RECT 77.965 134.250 79.120 134.800 ;
        RECT 80.055 134.425 80.515 134.655 ;
        RECT 85.805 134.500 86.035 139.510 ;
        RECT 86.595 134.500 86.825 139.510 ;
        RECT 88.000 139.145 89.925 140.175 ;
        RECT 87.195 138.175 87.565 138.225 ;
        RECT 87.195 137.120 88.300 138.175 ;
        RECT 77.965 134.200 79.025 134.250 ;
        RECT 57.680 129.510 57.910 129.520 ;
        RECT 58.470 129.510 58.700 129.520 ;
        RECT 60.380 129.510 60.610 129.520 ;
        RECT 61.170 129.510 61.400 129.520 ;
        RECT 63.080 129.510 63.310 129.520 ;
        RECT 63.870 129.510 64.100 129.520 ;
        RECT 65.780 129.510 66.010 129.520 ;
        RECT 66.570 129.510 66.800 129.520 ;
        RECT 68.480 129.510 68.710 129.520 ;
        RECT 69.270 129.510 69.500 129.520 ;
        RECT 71.180 129.510 71.410 129.520 ;
        RECT 71.970 129.510 72.200 129.520 ;
        RECT 57.425 128.850 58.460 129.325 ;
        RECT 60.660 129.075 61.120 129.305 ;
        RECT 62.825 128.850 63.860 129.325 ;
        RECT 65.525 128.850 66.560 129.325 ;
        RECT 68.760 129.075 69.220 129.305 ;
        RECT 71.460 129.075 71.920 129.305 ;
        RECT 54.800 128.475 55.800 128.530 ;
        RECT 75.670 128.510 76.775 133.180 ;
        RECT 83.385 130.715 83.845 130.945 ;
        RECT 83.105 130.500 83.335 130.510 ;
        RECT 83.895 130.500 84.125 130.510 ;
        RECT 82.360 129.520 83.405 130.500 ;
        RECT 83.825 129.520 84.195 130.500 ;
        RECT 85.735 129.520 86.105 134.500 ;
        RECT 86.525 129.520 86.895 134.500 ;
        RECT 87.300 132.425 88.300 137.120 ;
        RECT 88.925 134.075 89.925 139.145 ;
        RECT 90.725 139.145 92.675 140.175 ;
        RECT 93.925 139.725 94.925 140.175 ;
        RECT 96.625 139.725 97.625 140.175 ;
        RECT 94.185 139.715 94.645 139.725 ;
        RECT 96.885 139.715 97.345 139.725 ;
        RECT 90.725 134.820 91.725 139.145 ;
        RECT 93.165 138.175 93.535 138.225 ;
        RECT 92.450 137.120 93.535 138.175 ;
        RECT 88.925 133.075 91.755 134.075 ;
        RECT 92.450 132.425 93.450 137.120 ;
        RECT 93.905 134.500 94.135 139.510 ;
        RECT 94.695 134.500 94.925 139.510 ;
        RECT 95.295 137.120 95.665 138.225 ;
        RECT 95.865 137.120 96.235 138.225 ;
        RECT 96.605 134.500 96.835 139.510 ;
        RECT 97.395 134.500 97.625 139.510 ;
        RECT 97.995 137.120 98.365 138.225 ;
        RECT 87.300 131.425 93.450 132.425 ;
        RECT 88.785 130.715 89.245 130.945 ;
        RECT 91.485 130.715 91.945 130.945 ;
        RECT 88.505 130.500 88.735 130.510 ;
        RECT 89.295 130.500 89.525 130.510 ;
        RECT 91.205 130.500 91.435 130.510 ;
        RECT 91.995 130.500 92.225 130.510 ;
        RECT 87.760 129.520 88.805 130.500 ;
        RECT 89.225 129.520 89.595 130.500 ;
        RECT 90.460 129.520 91.505 130.500 ;
        RECT 91.925 129.520 92.295 130.500 ;
        RECT 93.835 129.520 94.205 134.500 ;
        RECT 94.625 129.520 94.995 134.500 ;
        RECT 96.535 129.520 96.905 134.500 ;
        RECT 97.325 129.520 97.695 134.500 ;
        RECT 83.105 129.510 83.335 129.520 ;
        RECT 83.895 129.510 84.125 129.520 ;
        RECT 85.805 129.510 86.035 129.520 ;
        RECT 86.595 129.510 86.825 129.520 ;
        RECT 88.505 129.510 88.735 129.520 ;
        RECT 89.295 129.510 89.525 129.520 ;
        RECT 91.205 129.510 91.435 129.520 ;
        RECT 91.995 129.510 92.225 129.520 ;
        RECT 93.905 129.510 94.135 129.520 ;
        RECT 94.695 129.510 94.925 129.520 ;
        RECT 96.605 129.510 96.835 129.520 ;
        RECT 97.395 129.510 97.625 129.520 ;
        RECT 82.850 128.850 83.885 129.325 ;
        RECT 86.085 129.075 86.545 129.305 ;
        RECT 88.250 128.850 89.285 129.325 ;
        RECT 90.950 128.850 91.985 129.325 ;
        RECT 94.185 129.075 94.645 129.305 ;
        RECT 96.885 129.075 97.345 129.305 ;
        RECT 80.225 128.510 81.225 128.530 ;
        RECT 50.695 127.475 51.755 128.475 ;
        RECT 54.770 127.475 55.830 128.475 ;
        RECT 6.570 126.605 7.610 127.100 ;
        RECT 9.810 126.625 10.270 126.855 ;
        RECT 11.970 126.605 13.010 127.100 ;
        RECT 14.670 126.605 15.710 127.100 ;
        RECT 17.910 126.625 18.370 126.855 ;
        RECT 20.610 126.625 21.070 126.855 ;
        RECT 6.830 126.455 7.060 126.465 ;
        RECT 7.620 126.455 7.850 126.465 ;
        RECT 9.530 126.455 9.760 126.465 ;
        RECT 10.320 126.455 10.550 126.465 ;
        RECT 12.230 126.455 12.460 126.465 ;
        RECT 13.020 126.455 13.250 126.465 ;
        RECT 14.930 126.455 15.160 126.465 ;
        RECT 15.720 126.455 15.950 126.465 ;
        RECT 17.630 126.455 17.860 126.465 ;
        RECT 18.420 126.455 18.650 126.465 ;
        RECT 20.330 126.455 20.560 126.465 ;
        RECT 21.120 126.455 21.350 126.465 ;
        RECT 6.085 125.825 7.130 126.455 ;
        RECT 7.550 125.825 7.920 126.455 ;
        RECT 6.830 125.815 7.060 125.825 ;
        RECT 7.620 125.815 7.850 125.825 ;
        RECT 7.110 125.425 7.570 125.655 ;
        RECT 1.900 123.250 4.950 124.250 ;
        RECT 9.460 123.275 9.830 126.455 ;
        RECT 10.250 123.275 10.620 126.455 ;
        RECT 11.485 125.825 12.530 126.455 ;
        RECT 12.950 125.825 13.320 126.455 ;
        RECT 14.185 125.825 15.230 126.455 ;
        RECT 15.650 125.825 16.020 126.455 ;
        RECT 12.230 125.815 12.460 125.825 ;
        RECT 13.020 125.815 13.250 125.825 ;
        RECT 14.930 125.815 15.160 125.825 ;
        RECT 15.720 125.815 15.950 125.825 ;
        RECT 12.510 125.425 12.970 125.655 ;
        RECT 15.210 125.425 15.670 125.655 ;
        RECT 17.560 123.275 17.930 126.455 ;
        RECT 18.350 123.275 18.720 126.455 ;
        RECT 20.260 123.275 20.630 126.455 ;
        RECT 21.050 123.275 21.420 126.455 ;
        RECT 29.375 124.250 30.375 127.405 ;
        RECT 31.995 126.605 33.035 127.100 ;
        RECT 35.235 126.625 35.695 126.855 ;
        RECT 37.395 126.605 38.435 127.100 ;
        RECT 40.095 126.605 41.135 127.100 ;
        RECT 43.335 126.625 43.795 126.855 ;
        RECT 46.035 126.625 46.495 126.855 ;
        RECT 32.255 126.455 32.485 126.465 ;
        RECT 33.045 126.455 33.275 126.465 ;
        RECT 34.955 126.455 35.185 126.465 ;
        RECT 35.745 126.455 35.975 126.465 ;
        RECT 37.655 126.455 37.885 126.465 ;
        RECT 38.445 126.455 38.675 126.465 ;
        RECT 40.355 126.455 40.585 126.465 ;
        RECT 41.145 126.455 41.375 126.465 ;
        RECT 43.055 126.455 43.285 126.465 ;
        RECT 43.845 126.455 44.075 126.465 ;
        RECT 45.755 126.455 45.985 126.465 ;
        RECT 46.545 126.455 46.775 126.465 ;
        RECT 31.510 125.825 32.555 126.455 ;
        RECT 32.975 125.825 33.345 126.455 ;
        RECT 32.255 125.815 32.485 125.825 ;
        RECT 33.045 125.815 33.275 125.825 ;
        RECT 32.535 125.425 32.995 125.655 ;
        RECT 1.900 105.900 2.900 123.250 ;
        RECT 3.905 122.430 5.020 122.485 ;
        RECT 3.875 121.315 5.050 122.430 ;
        RECT 8.790 121.320 9.160 122.435 ;
        RECT 1.870 104.900 2.930 105.900 ;
        RECT 1.900 83.325 2.900 104.900 ;
        RECT 3.905 99.855 5.020 121.315 ;
        RECT 9.530 119.965 9.760 123.275 ;
        RECT 10.320 119.965 10.550 123.275 ;
        RECT 10.920 121.320 11.290 122.435 ;
        RECT 16.890 121.320 17.260 122.435 ;
        RECT 17.630 119.965 17.860 123.275 ;
        RECT 18.420 119.965 18.650 123.275 ;
        RECT 19.020 121.320 19.390 122.435 ;
        RECT 19.590 121.320 19.960 122.435 ;
        RECT 20.330 119.965 20.560 123.275 ;
        RECT 21.120 119.965 21.350 123.275 ;
        RECT 27.325 123.250 30.375 124.250 ;
        RECT 34.885 123.275 35.255 126.455 ;
        RECT 35.675 123.275 36.045 126.455 ;
        RECT 36.910 125.825 37.955 126.455 ;
        RECT 38.375 125.825 38.745 126.455 ;
        RECT 39.610 125.825 40.655 126.455 ;
        RECT 41.075 125.825 41.445 126.455 ;
        RECT 37.655 125.815 37.885 125.825 ;
        RECT 38.445 125.815 38.675 125.825 ;
        RECT 40.355 125.815 40.585 125.825 ;
        RECT 41.145 125.815 41.375 125.825 ;
        RECT 37.935 125.425 38.395 125.655 ;
        RECT 40.635 125.425 41.095 125.655 ;
        RECT 42.985 123.275 43.355 126.455 ;
        RECT 43.775 123.275 44.145 126.455 ;
        RECT 45.685 123.275 46.055 126.455 ;
        RECT 46.475 123.275 46.845 126.455 ;
        RECT 54.800 124.250 55.800 127.475 ;
        RECT 75.670 127.405 81.280 128.510 ;
        RECT 101.575 128.475 102.575 141.550 ;
        RECT 113.425 140.175 114.425 140.205 ;
        RECT 117.100 140.175 118.100 140.205 ;
        RECT 138.850 140.175 139.850 140.205 ;
        RECT 142.525 140.175 143.525 140.205 ;
        RECT 111.250 139.725 112.250 140.175 ;
        RECT 111.510 139.715 111.970 139.725 ;
        RECT 110.490 137.120 110.860 138.225 ;
        RECT 111.230 134.500 111.460 139.510 ;
        RECT 112.020 134.500 112.250 139.510 ;
        RECT 113.425 139.145 115.350 140.175 ;
        RECT 112.620 138.175 112.990 138.225 ;
        RECT 112.620 137.120 113.725 138.175 ;
        RECT 108.810 130.715 109.270 130.945 ;
        RECT 108.530 130.500 108.760 130.510 ;
        RECT 109.320 130.500 109.550 130.510 ;
        RECT 107.785 129.520 108.830 130.500 ;
        RECT 109.250 129.520 109.620 130.500 ;
        RECT 111.160 129.520 111.530 134.500 ;
        RECT 111.950 129.520 112.320 134.500 ;
        RECT 112.725 132.425 113.725 137.120 ;
        RECT 114.350 134.075 115.350 139.145 ;
        RECT 116.150 139.145 118.100 140.175 ;
        RECT 119.350 139.725 120.350 140.175 ;
        RECT 122.050 139.725 123.050 140.175 ;
        RECT 128.970 139.975 129.970 140.125 ;
        RECT 119.610 139.715 120.070 139.725 ;
        RECT 122.310 139.715 122.770 139.725 ;
        RECT 125.505 139.715 125.965 139.945 ;
        RECT 128.205 139.715 128.665 139.945 ;
        RECT 128.820 139.525 129.970 139.975 ;
        RECT 130.905 139.715 131.365 139.945 ;
        RECT 136.675 139.725 137.675 140.175 ;
        RECT 136.935 139.715 137.395 139.725 ;
        RECT 116.150 134.820 117.150 139.145 ;
        RECT 118.590 138.175 118.960 138.225 ;
        RECT 117.875 137.120 118.960 138.175 ;
        RECT 114.350 133.075 117.180 134.075 ;
        RECT 117.875 132.425 118.875 137.120 ;
        RECT 119.330 134.500 119.560 139.510 ;
        RECT 120.120 134.500 120.350 139.510 ;
        RECT 120.720 137.120 121.090 138.225 ;
        RECT 121.290 137.120 121.660 138.225 ;
        RECT 122.030 134.500 122.260 139.510 ;
        RECT 122.820 134.500 123.050 139.510 ;
        RECT 125.225 138.510 125.455 139.510 ;
        RECT 125.995 138.495 128.175 139.525 ;
        RECT 128.670 139.500 129.970 139.525 ;
        RECT 130.625 139.500 130.855 139.510 ;
        RECT 131.415 139.500 131.645 139.510 ;
        RECT 128.670 138.975 130.925 139.500 ;
        RECT 128.670 138.570 129.590 138.975 ;
        RECT 128.715 138.510 128.945 138.570 ;
        RECT 129.880 138.520 130.925 138.975 ;
        RECT 131.345 138.520 131.715 139.500 ;
        RECT 130.625 138.510 130.855 138.520 ;
        RECT 131.415 138.510 131.645 138.520 ;
        RECT 123.420 137.120 123.790 138.225 ;
        RECT 125.220 135.625 126.220 138.355 ;
        RECT 127.945 135.625 128.945 138.325 ;
        RECT 130.370 137.850 131.405 138.325 ;
        RECT 135.915 137.120 136.285 138.225 ;
        RECT 130.365 135.605 131.405 136.100 ;
        RECT 124.905 134.800 125.550 135.480 ;
        RECT 125.945 134.800 128.225 135.480 ;
        RECT 128.715 135.405 128.945 135.465 ;
        RECT 130.625 135.455 130.855 135.465 ;
        RECT 131.415 135.455 131.645 135.465 ;
        RECT 128.670 135.250 129.590 135.405 ;
        RECT 129.880 135.250 130.925 135.455 ;
        RECT 128.670 134.825 130.925 135.250 ;
        RECT 131.345 134.825 131.715 135.455 ;
        RECT 128.715 134.815 129.970 134.825 ;
        RECT 130.625 134.815 130.855 134.825 ;
        RECT 131.415 134.815 131.645 134.825 ;
        RECT 128.720 134.800 129.970 134.815 ;
        RECT 112.725 131.425 118.875 132.425 ;
        RECT 114.210 130.715 114.670 130.945 ;
        RECT 116.910 130.715 117.370 130.945 ;
        RECT 113.930 130.500 114.160 130.510 ;
        RECT 114.720 130.500 114.950 130.510 ;
        RECT 116.630 130.500 116.860 130.510 ;
        RECT 117.420 130.500 117.650 130.510 ;
        RECT 113.185 129.520 114.230 130.500 ;
        RECT 114.650 129.520 115.020 130.500 ;
        RECT 115.885 129.520 116.930 130.500 ;
        RECT 117.350 129.520 117.720 130.500 ;
        RECT 119.260 129.520 119.630 134.500 ;
        RECT 120.050 129.520 120.420 134.500 ;
        RECT 121.960 129.520 122.330 134.500 ;
        RECT 122.750 129.520 123.120 134.500 ;
        RECT 125.505 134.425 125.965 134.655 ;
        RECT 128.205 134.425 128.665 134.655 ;
        RECT 128.815 134.250 129.970 134.800 ;
        RECT 130.905 134.425 131.365 134.655 ;
        RECT 136.655 134.500 136.885 139.510 ;
        RECT 137.445 134.500 137.675 139.510 ;
        RECT 138.850 139.145 140.775 140.175 ;
        RECT 138.045 138.175 138.415 138.225 ;
        RECT 138.045 137.120 139.150 138.175 ;
        RECT 128.815 134.200 129.875 134.250 ;
        RECT 108.530 129.510 108.760 129.520 ;
        RECT 109.320 129.510 109.550 129.520 ;
        RECT 111.230 129.510 111.460 129.520 ;
        RECT 112.020 129.510 112.250 129.520 ;
        RECT 113.930 129.510 114.160 129.520 ;
        RECT 114.720 129.510 114.950 129.520 ;
        RECT 116.630 129.510 116.860 129.520 ;
        RECT 117.420 129.510 117.650 129.520 ;
        RECT 119.330 129.510 119.560 129.520 ;
        RECT 120.120 129.510 120.350 129.520 ;
        RECT 122.030 129.510 122.260 129.520 ;
        RECT 122.820 129.510 123.050 129.520 ;
        RECT 108.275 128.850 109.310 129.325 ;
        RECT 111.510 129.075 111.970 129.305 ;
        RECT 113.675 128.850 114.710 129.325 ;
        RECT 116.375 128.850 117.410 129.325 ;
        RECT 119.610 129.075 120.070 129.305 ;
        RECT 122.310 129.075 122.770 129.305 ;
        RECT 105.650 128.475 106.650 128.530 ;
        RECT 126.520 128.510 127.625 133.180 ;
        RECT 134.235 130.715 134.695 130.945 ;
        RECT 133.955 130.500 134.185 130.510 ;
        RECT 134.745 130.500 134.975 130.510 ;
        RECT 133.210 129.520 134.255 130.500 ;
        RECT 134.675 129.520 135.045 130.500 ;
        RECT 136.585 129.520 136.955 134.500 ;
        RECT 137.375 129.520 137.745 134.500 ;
        RECT 138.150 132.425 139.150 137.120 ;
        RECT 139.775 134.075 140.775 139.145 ;
        RECT 141.575 139.145 143.525 140.175 ;
        RECT 144.775 139.725 145.775 140.175 ;
        RECT 147.475 139.725 148.475 140.175 ;
        RECT 145.035 139.715 145.495 139.725 ;
        RECT 147.735 139.715 148.195 139.725 ;
        RECT 141.575 134.820 142.575 139.145 ;
        RECT 144.015 138.175 144.385 138.225 ;
        RECT 143.300 137.120 144.385 138.175 ;
        RECT 139.775 133.075 142.605 134.075 ;
        RECT 143.300 132.425 144.300 137.120 ;
        RECT 144.755 134.500 144.985 139.510 ;
        RECT 145.545 134.500 145.775 139.510 ;
        RECT 146.145 137.120 146.515 138.225 ;
        RECT 146.715 137.120 147.085 138.225 ;
        RECT 147.455 134.500 147.685 139.510 ;
        RECT 148.245 134.500 148.475 139.510 ;
        RECT 148.845 137.120 149.215 138.225 ;
        RECT 138.150 131.425 144.300 132.425 ;
        RECT 139.635 130.715 140.095 130.945 ;
        RECT 142.335 130.715 142.795 130.945 ;
        RECT 139.355 130.500 139.585 130.510 ;
        RECT 140.145 130.500 140.375 130.510 ;
        RECT 142.055 130.500 142.285 130.510 ;
        RECT 142.845 130.500 143.075 130.510 ;
        RECT 138.610 129.520 139.655 130.500 ;
        RECT 140.075 129.520 140.445 130.500 ;
        RECT 141.310 129.520 142.355 130.500 ;
        RECT 142.775 129.520 143.145 130.500 ;
        RECT 144.685 129.520 145.055 134.500 ;
        RECT 145.475 129.520 145.845 134.500 ;
        RECT 147.385 129.520 147.755 134.500 ;
        RECT 148.175 129.520 148.545 134.500 ;
        RECT 133.955 129.510 134.185 129.520 ;
        RECT 134.745 129.510 134.975 129.520 ;
        RECT 136.655 129.510 136.885 129.520 ;
        RECT 137.445 129.510 137.675 129.520 ;
        RECT 139.355 129.510 139.585 129.520 ;
        RECT 140.145 129.510 140.375 129.520 ;
        RECT 142.055 129.510 142.285 129.520 ;
        RECT 142.845 129.510 143.075 129.520 ;
        RECT 144.755 129.510 144.985 129.520 ;
        RECT 145.545 129.510 145.775 129.520 ;
        RECT 147.455 129.510 147.685 129.520 ;
        RECT 148.245 129.510 148.475 129.520 ;
        RECT 133.700 128.850 134.735 129.325 ;
        RECT 136.935 129.075 137.395 129.305 ;
        RECT 139.100 128.850 140.135 129.325 ;
        RECT 141.800 128.850 142.835 129.325 ;
        RECT 145.035 129.075 145.495 129.305 ;
        RECT 147.735 129.075 148.195 129.305 ;
        RECT 131.075 128.510 132.075 128.530 ;
        RECT 101.545 127.475 102.605 128.475 ;
        RECT 105.620 127.475 106.680 128.475 ;
        RECT 57.420 126.605 58.460 127.100 ;
        RECT 60.660 126.625 61.120 126.855 ;
        RECT 62.820 126.605 63.860 127.100 ;
        RECT 65.520 126.605 66.560 127.100 ;
        RECT 68.760 126.625 69.220 126.855 ;
        RECT 71.460 126.625 71.920 126.855 ;
        RECT 57.680 126.455 57.910 126.465 ;
        RECT 58.470 126.455 58.700 126.465 ;
        RECT 60.380 126.455 60.610 126.465 ;
        RECT 61.170 126.455 61.400 126.465 ;
        RECT 63.080 126.455 63.310 126.465 ;
        RECT 63.870 126.455 64.100 126.465 ;
        RECT 65.780 126.455 66.010 126.465 ;
        RECT 66.570 126.455 66.800 126.465 ;
        RECT 68.480 126.455 68.710 126.465 ;
        RECT 69.270 126.455 69.500 126.465 ;
        RECT 71.180 126.455 71.410 126.465 ;
        RECT 71.970 126.455 72.200 126.465 ;
        RECT 56.935 125.825 57.980 126.455 ;
        RECT 58.400 125.825 58.770 126.455 ;
        RECT 57.680 125.815 57.910 125.825 ;
        RECT 58.470 125.815 58.700 125.825 ;
        RECT 57.960 125.425 58.420 125.655 ;
        RECT 21.720 121.320 22.090 122.435 ;
        RECT 9.810 119.775 10.270 119.805 ;
        RECT 17.910 119.775 18.370 119.805 ;
        RECT 20.610 119.775 21.070 119.805 ;
        RECT 9.550 119.375 10.550 119.775 ;
        RECT 17.650 119.375 18.650 119.775 ;
        RECT 20.350 119.375 21.350 119.775 ;
        RECT 11.725 117.600 12.725 117.630 ;
        RECT 15.400 117.600 16.400 117.630 ;
        RECT 9.550 117.150 10.550 117.600 ;
        RECT 9.810 117.140 10.270 117.150 ;
        RECT 8.790 114.545 9.160 115.650 ;
        RECT 9.530 111.925 9.760 116.935 ;
        RECT 10.320 111.925 10.550 116.935 ;
        RECT 11.725 116.570 13.650 117.600 ;
        RECT 10.920 115.600 11.290 115.650 ;
        RECT 10.920 114.545 12.025 115.600 ;
        RECT 7.110 108.140 7.570 108.370 ;
        RECT 6.830 107.925 7.060 107.935 ;
        RECT 7.620 107.925 7.850 107.935 ;
        RECT 6.085 106.945 7.130 107.925 ;
        RECT 7.550 106.945 7.920 107.925 ;
        RECT 9.460 106.945 9.830 111.925 ;
        RECT 10.250 106.945 10.620 111.925 ;
        RECT 11.025 109.850 12.025 114.545 ;
        RECT 12.650 111.500 13.650 116.570 ;
        RECT 14.450 116.570 16.400 117.600 ;
        RECT 17.650 117.150 18.650 117.600 ;
        RECT 20.350 117.150 21.350 117.600 ;
        RECT 17.910 117.140 18.370 117.150 ;
        RECT 20.610 117.140 21.070 117.150 ;
        RECT 14.450 112.245 15.450 116.570 ;
        RECT 16.890 115.600 17.260 115.650 ;
        RECT 16.175 114.545 17.260 115.600 ;
        RECT 12.650 110.500 15.480 111.500 ;
        RECT 16.175 109.850 17.175 114.545 ;
        RECT 17.630 111.925 17.860 116.935 ;
        RECT 18.420 111.925 18.650 116.935 ;
        RECT 19.020 114.545 19.390 115.650 ;
        RECT 19.590 114.545 19.960 115.650 ;
        RECT 20.330 111.925 20.560 116.935 ;
        RECT 21.120 111.925 21.350 116.935 ;
        RECT 21.720 114.545 22.090 115.650 ;
        RECT 11.025 108.850 17.175 109.850 ;
        RECT 12.510 108.140 12.970 108.370 ;
        RECT 15.210 108.140 15.670 108.370 ;
        RECT 12.230 107.925 12.460 107.935 ;
        RECT 13.020 107.925 13.250 107.935 ;
        RECT 14.930 107.925 15.160 107.935 ;
        RECT 15.720 107.925 15.950 107.935 ;
        RECT 11.485 106.945 12.530 107.925 ;
        RECT 12.950 106.945 13.320 107.925 ;
        RECT 14.185 106.945 15.230 107.925 ;
        RECT 15.650 106.945 16.020 107.925 ;
        RECT 17.560 106.945 17.930 111.925 ;
        RECT 18.350 106.945 18.720 111.925 ;
        RECT 20.260 106.945 20.630 111.925 ;
        RECT 21.050 106.945 21.420 111.925 ;
        RECT 6.830 106.935 7.060 106.945 ;
        RECT 7.620 106.935 7.850 106.945 ;
        RECT 9.530 106.935 9.760 106.945 ;
        RECT 10.320 106.935 10.550 106.945 ;
        RECT 12.230 106.935 12.460 106.945 ;
        RECT 13.020 106.935 13.250 106.945 ;
        RECT 14.930 106.935 15.160 106.945 ;
        RECT 15.720 106.935 15.950 106.945 ;
        RECT 17.630 106.935 17.860 106.945 ;
        RECT 18.420 106.935 18.650 106.945 ;
        RECT 20.330 106.935 20.560 106.945 ;
        RECT 21.120 106.935 21.350 106.945 ;
        RECT 6.575 106.275 7.610 106.750 ;
        RECT 9.810 106.500 10.270 106.730 ;
        RECT 11.975 106.275 13.010 106.750 ;
        RECT 14.675 106.275 15.710 106.750 ;
        RECT 17.910 106.500 18.370 106.730 ;
        RECT 20.610 106.500 21.070 106.730 ;
        RECT 27.325 105.900 28.325 123.250 ;
        RECT 29.330 122.430 30.445 122.485 ;
        RECT 29.300 121.315 30.475 122.430 ;
        RECT 34.215 121.320 34.585 122.435 ;
        RECT 27.295 104.900 28.355 105.900 ;
        RECT 6.570 104.030 7.610 104.525 ;
        RECT 9.810 104.050 10.270 104.280 ;
        RECT 11.970 104.030 13.010 104.525 ;
        RECT 14.670 104.030 15.710 104.525 ;
        RECT 17.910 104.050 18.370 104.280 ;
        RECT 20.610 104.050 21.070 104.280 ;
        RECT 6.830 103.880 7.060 103.890 ;
        RECT 7.620 103.880 7.850 103.890 ;
        RECT 9.530 103.880 9.760 103.890 ;
        RECT 10.320 103.880 10.550 103.890 ;
        RECT 12.230 103.880 12.460 103.890 ;
        RECT 13.020 103.880 13.250 103.890 ;
        RECT 14.930 103.880 15.160 103.890 ;
        RECT 15.720 103.880 15.950 103.890 ;
        RECT 17.630 103.880 17.860 103.890 ;
        RECT 18.420 103.880 18.650 103.890 ;
        RECT 20.330 103.880 20.560 103.890 ;
        RECT 21.120 103.880 21.350 103.890 ;
        RECT 6.085 103.250 7.130 103.880 ;
        RECT 7.550 103.250 7.920 103.880 ;
        RECT 6.830 103.240 7.060 103.250 ;
        RECT 7.620 103.240 7.850 103.250 ;
        RECT 7.110 102.850 7.570 103.080 ;
        RECT 9.460 100.700 9.830 103.880 ;
        RECT 10.250 100.700 10.620 103.880 ;
        RECT 11.485 103.250 12.530 103.880 ;
        RECT 12.950 103.250 13.320 103.880 ;
        RECT 14.185 103.250 15.230 103.880 ;
        RECT 15.650 103.250 16.020 103.880 ;
        RECT 12.230 103.240 12.460 103.250 ;
        RECT 13.020 103.240 13.250 103.250 ;
        RECT 14.930 103.240 15.160 103.250 ;
        RECT 15.720 103.240 15.950 103.250 ;
        RECT 12.510 102.850 12.970 103.080 ;
        RECT 15.210 102.850 15.670 103.080 ;
        RECT 17.560 100.700 17.930 103.880 ;
        RECT 18.350 100.700 18.720 103.880 ;
        RECT 20.260 100.700 20.630 103.880 ;
        RECT 21.050 100.700 21.420 103.880 ;
        RECT 3.875 98.740 5.050 99.855 ;
        RECT 8.790 98.745 9.160 99.860 ;
        RECT 1.870 82.325 2.930 83.325 ;
        RECT 1.900 82.295 2.900 82.325 ;
        RECT 3.905 77.285 5.020 98.740 ;
        RECT 9.530 97.390 9.760 100.700 ;
        RECT 10.320 97.390 10.550 100.700 ;
        RECT 10.920 98.745 11.290 99.860 ;
        RECT 16.890 98.745 17.260 99.860 ;
        RECT 17.630 97.390 17.860 100.700 ;
        RECT 18.420 97.390 18.650 100.700 ;
        RECT 19.020 98.745 19.390 99.860 ;
        RECT 19.590 98.745 19.960 99.860 ;
        RECT 20.330 97.390 20.560 100.700 ;
        RECT 21.120 97.390 21.350 100.700 ;
        RECT 21.720 98.745 22.090 99.860 ;
        RECT 23.085 98.745 24.260 99.860 ;
        RECT 9.810 97.200 10.270 97.230 ;
        RECT 17.910 97.200 18.370 97.230 ;
        RECT 20.610 97.200 21.070 97.230 ;
        RECT 9.550 96.800 10.550 97.200 ;
        RECT 17.650 96.800 18.650 97.200 ;
        RECT 20.350 96.800 21.350 97.200 ;
        RECT 23.115 95.770 24.230 98.745 ;
        RECT 11.725 95.025 12.725 95.055 ;
        RECT 15.400 95.025 16.400 95.055 ;
        RECT 9.550 94.575 10.550 95.025 ;
        RECT 9.810 94.565 10.270 94.575 ;
        RECT 8.790 91.970 9.160 93.075 ;
        RECT 9.530 89.350 9.760 94.360 ;
        RECT 10.320 89.350 10.550 94.360 ;
        RECT 11.725 93.995 13.650 95.025 ;
        RECT 10.920 93.025 11.290 93.075 ;
        RECT 10.920 91.970 12.025 93.025 ;
        RECT 7.110 85.565 7.570 85.795 ;
        RECT 6.830 85.350 7.060 85.360 ;
        RECT 7.620 85.350 7.850 85.360 ;
        RECT 6.085 84.370 7.130 85.350 ;
        RECT 7.550 84.370 7.920 85.350 ;
        RECT 9.460 84.370 9.830 89.350 ;
        RECT 10.250 84.370 10.620 89.350 ;
        RECT 11.025 87.275 12.025 91.970 ;
        RECT 12.650 88.925 13.650 93.995 ;
        RECT 14.450 93.995 16.400 95.025 ;
        RECT 17.650 94.575 18.650 95.025 ;
        RECT 20.350 94.575 21.350 95.025 ;
        RECT 17.910 94.565 18.370 94.575 ;
        RECT 20.610 94.565 21.070 94.575 ;
        RECT 14.450 89.670 15.450 93.995 ;
        RECT 16.890 93.025 17.260 93.075 ;
        RECT 16.175 91.970 17.260 93.025 ;
        RECT 12.650 87.925 15.480 88.925 ;
        RECT 16.175 87.275 17.175 91.970 ;
        RECT 17.630 89.350 17.860 94.360 ;
        RECT 18.420 89.350 18.650 94.360 ;
        RECT 19.020 91.970 19.390 93.075 ;
        RECT 19.590 91.970 19.960 93.075 ;
        RECT 20.330 89.350 20.560 94.360 ;
        RECT 21.120 89.350 21.350 94.360 ;
        RECT 23.430 93.115 23.880 95.425 ;
        RECT 21.720 91.970 22.090 93.075 ;
        RECT 11.025 86.275 17.175 87.275 ;
        RECT 12.510 85.565 12.970 85.795 ;
        RECT 15.210 85.565 15.670 85.795 ;
        RECT 12.230 85.350 12.460 85.360 ;
        RECT 13.020 85.350 13.250 85.360 ;
        RECT 14.930 85.350 15.160 85.360 ;
        RECT 15.720 85.350 15.950 85.360 ;
        RECT 11.485 84.370 12.530 85.350 ;
        RECT 12.950 84.370 13.320 85.350 ;
        RECT 14.185 84.370 15.230 85.350 ;
        RECT 15.650 84.370 16.020 85.350 ;
        RECT 17.560 84.370 17.930 89.350 ;
        RECT 18.350 84.370 18.720 89.350 ;
        RECT 20.260 84.370 20.630 89.350 ;
        RECT 21.050 84.370 21.420 89.350 ;
        RECT 6.830 84.360 7.060 84.370 ;
        RECT 7.620 84.360 7.850 84.370 ;
        RECT 9.530 84.360 9.760 84.370 ;
        RECT 10.320 84.360 10.550 84.370 ;
        RECT 12.230 84.360 12.460 84.370 ;
        RECT 13.020 84.360 13.250 84.370 ;
        RECT 14.930 84.360 15.160 84.370 ;
        RECT 15.720 84.360 15.950 84.370 ;
        RECT 17.630 84.360 17.860 84.370 ;
        RECT 18.420 84.360 18.650 84.370 ;
        RECT 20.330 84.360 20.560 84.370 ;
        RECT 21.120 84.360 21.350 84.370 ;
        RECT 6.575 83.700 7.610 84.175 ;
        RECT 9.810 83.925 10.270 84.155 ;
        RECT 11.975 83.700 13.010 84.175 ;
        RECT 14.675 83.700 15.710 84.175 ;
        RECT 17.910 83.925 18.370 84.155 ;
        RECT 20.610 83.925 21.070 84.155 ;
        RECT 23.430 82.205 23.880 84.515 ;
        RECT 27.325 83.325 28.325 104.900 ;
        RECT 29.330 99.855 30.445 121.315 ;
        RECT 34.955 119.965 35.185 123.275 ;
        RECT 35.745 119.965 35.975 123.275 ;
        RECT 36.345 121.320 36.715 122.435 ;
        RECT 42.315 121.320 42.685 122.435 ;
        RECT 43.055 119.965 43.285 123.275 ;
        RECT 43.845 119.965 44.075 123.275 ;
        RECT 44.445 121.320 44.815 122.435 ;
        RECT 45.015 121.320 45.385 122.435 ;
        RECT 45.755 119.965 45.985 123.275 ;
        RECT 46.545 119.965 46.775 123.275 ;
        RECT 52.750 123.250 55.800 124.250 ;
        RECT 60.310 123.275 60.680 126.455 ;
        RECT 61.100 123.275 61.470 126.455 ;
        RECT 62.335 125.825 63.380 126.455 ;
        RECT 63.800 125.825 64.170 126.455 ;
        RECT 65.035 125.825 66.080 126.455 ;
        RECT 66.500 125.825 66.870 126.455 ;
        RECT 63.080 125.815 63.310 125.825 ;
        RECT 63.870 125.815 64.100 125.825 ;
        RECT 65.780 125.815 66.010 125.825 ;
        RECT 66.570 125.815 66.800 125.825 ;
        RECT 63.360 125.425 63.820 125.655 ;
        RECT 66.060 125.425 66.520 125.655 ;
        RECT 68.410 123.275 68.780 126.455 ;
        RECT 69.200 123.275 69.570 126.455 ;
        RECT 71.110 123.275 71.480 126.455 ;
        RECT 71.900 123.275 72.270 126.455 ;
        RECT 80.225 124.250 81.225 127.405 ;
        RECT 82.845 126.605 83.885 127.100 ;
        RECT 86.085 126.625 86.545 126.855 ;
        RECT 88.245 126.605 89.285 127.100 ;
        RECT 90.945 126.605 91.985 127.100 ;
        RECT 94.185 126.625 94.645 126.855 ;
        RECT 96.885 126.625 97.345 126.855 ;
        RECT 83.105 126.455 83.335 126.465 ;
        RECT 83.895 126.455 84.125 126.465 ;
        RECT 85.805 126.455 86.035 126.465 ;
        RECT 86.595 126.455 86.825 126.465 ;
        RECT 88.505 126.455 88.735 126.465 ;
        RECT 89.295 126.455 89.525 126.465 ;
        RECT 91.205 126.455 91.435 126.465 ;
        RECT 91.995 126.455 92.225 126.465 ;
        RECT 93.905 126.455 94.135 126.465 ;
        RECT 94.695 126.455 94.925 126.465 ;
        RECT 96.605 126.455 96.835 126.465 ;
        RECT 97.395 126.455 97.625 126.465 ;
        RECT 82.360 125.825 83.405 126.455 ;
        RECT 83.825 125.825 84.195 126.455 ;
        RECT 83.105 125.815 83.335 125.825 ;
        RECT 83.895 125.815 84.125 125.825 ;
        RECT 83.385 125.425 83.845 125.655 ;
        RECT 47.145 121.320 47.515 122.435 ;
        RECT 35.235 119.775 35.695 119.805 ;
        RECT 43.335 119.775 43.795 119.805 ;
        RECT 46.035 119.775 46.495 119.805 ;
        RECT 34.975 119.375 35.975 119.775 ;
        RECT 43.075 119.375 44.075 119.775 ;
        RECT 45.775 119.375 46.775 119.775 ;
        RECT 37.150 117.600 38.150 117.630 ;
        RECT 40.825 117.600 41.825 117.630 ;
        RECT 34.975 117.150 35.975 117.600 ;
        RECT 35.235 117.140 35.695 117.150 ;
        RECT 34.215 114.545 34.585 115.650 ;
        RECT 34.955 111.925 35.185 116.935 ;
        RECT 35.745 111.925 35.975 116.935 ;
        RECT 37.150 116.570 39.075 117.600 ;
        RECT 36.345 115.600 36.715 115.650 ;
        RECT 36.345 114.545 37.450 115.600 ;
        RECT 32.535 108.140 32.995 108.370 ;
        RECT 32.255 107.925 32.485 107.935 ;
        RECT 33.045 107.925 33.275 107.935 ;
        RECT 31.510 106.945 32.555 107.925 ;
        RECT 32.975 106.945 33.345 107.925 ;
        RECT 34.885 106.945 35.255 111.925 ;
        RECT 35.675 106.945 36.045 111.925 ;
        RECT 36.450 109.850 37.450 114.545 ;
        RECT 38.075 111.500 39.075 116.570 ;
        RECT 39.875 116.570 41.825 117.600 ;
        RECT 43.075 117.150 44.075 117.600 ;
        RECT 45.775 117.150 46.775 117.600 ;
        RECT 43.335 117.140 43.795 117.150 ;
        RECT 46.035 117.140 46.495 117.150 ;
        RECT 39.875 112.245 40.875 116.570 ;
        RECT 42.315 115.600 42.685 115.650 ;
        RECT 41.600 114.545 42.685 115.600 ;
        RECT 38.075 110.500 40.905 111.500 ;
        RECT 41.600 109.850 42.600 114.545 ;
        RECT 43.055 111.925 43.285 116.935 ;
        RECT 43.845 111.925 44.075 116.935 ;
        RECT 44.445 114.545 44.815 115.650 ;
        RECT 45.015 114.545 45.385 115.650 ;
        RECT 45.755 111.925 45.985 116.935 ;
        RECT 46.545 111.925 46.775 116.935 ;
        RECT 47.145 114.545 47.515 115.650 ;
        RECT 36.450 108.850 42.600 109.850 ;
        RECT 37.935 108.140 38.395 108.370 ;
        RECT 40.635 108.140 41.095 108.370 ;
        RECT 37.655 107.925 37.885 107.935 ;
        RECT 38.445 107.925 38.675 107.935 ;
        RECT 40.355 107.925 40.585 107.935 ;
        RECT 41.145 107.925 41.375 107.935 ;
        RECT 36.910 106.945 37.955 107.925 ;
        RECT 38.375 106.945 38.745 107.925 ;
        RECT 39.610 106.945 40.655 107.925 ;
        RECT 41.075 106.945 41.445 107.925 ;
        RECT 42.985 106.945 43.355 111.925 ;
        RECT 43.775 106.945 44.145 111.925 ;
        RECT 45.685 106.945 46.055 111.925 ;
        RECT 46.475 106.945 46.845 111.925 ;
        RECT 32.255 106.935 32.485 106.945 ;
        RECT 33.045 106.935 33.275 106.945 ;
        RECT 34.955 106.935 35.185 106.945 ;
        RECT 35.745 106.935 35.975 106.945 ;
        RECT 37.655 106.935 37.885 106.945 ;
        RECT 38.445 106.935 38.675 106.945 ;
        RECT 40.355 106.935 40.585 106.945 ;
        RECT 41.145 106.935 41.375 106.945 ;
        RECT 43.055 106.935 43.285 106.945 ;
        RECT 43.845 106.935 44.075 106.945 ;
        RECT 45.755 106.935 45.985 106.945 ;
        RECT 46.545 106.935 46.775 106.945 ;
        RECT 32.000 106.275 33.035 106.750 ;
        RECT 35.235 106.500 35.695 106.730 ;
        RECT 37.400 106.275 38.435 106.750 ;
        RECT 40.100 106.275 41.135 106.750 ;
        RECT 43.335 106.500 43.795 106.730 ;
        RECT 46.035 106.500 46.495 106.730 ;
        RECT 52.750 105.900 53.750 123.250 ;
        RECT 54.755 122.430 55.870 122.485 ;
        RECT 54.725 121.315 55.900 122.430 ;
        RECT 59.640 121.320 60.010 122.435 ;
        RECT 52.720 104.900 53.780 105.900 ;
        RECT 31.995 104.030 33.035 104.525 ;
        RECT 35.235 104.050 35.695 104.280 ;
        RECT 37.395 104.030 38.435 104.525 ;
        RECT 40.095 104.030 41.135 104.525 ;
        RECT 43.335 104.050 43.795 104.280 ;
        RECT 46.035 104.050 46.495 104.280 ;
        RECT 32.255 103.880 32.485 103.890 ;
        RECT 33.045 103.880 33.275 103.890 ;
        RECT 34.955 103.880 35.185 103.890 ;
        RECT 35.745 103.880 35.975 103.890 ;
        RECT 37.655 103.880 37.885 103.890 ;
        RECT 38.445 103.880 38.675 103.890 ;
        RECT 40.355 103.880 40.585 103.890 ;
        RECT 41.145 103.880 41.375 103.890 ;
        RECT 43.055 103.880 43.285 103.890 ;
        RECT 43.845 103.880 44.075 103.890 ;
        RECT 45.755 103.880 45.985 103.890 ;
        RECT 46.545 103.880 46.775 103.890 ;
        RECT 31.510 103.250 32.555 103.880 ;
        RECT 32.975 103.250 33.345 103.880 ;
        RECT 32.255 103.240 32.485 103.250 ;
        RECT 33.045 103.240 33.275 103.250 ;
        RECT 32.535 102.850 32.995 103.080 ;
        RECT 34.885 100.700 35.255 103.880 ;
        RECT 35.675 100.700 36.045 103.880 ;
        RECT 36.910 103.250 37.955 103.880 ;
        RECT 38.375 103.250 38.745 103.880 ;
        RECT 39.610 103.250 40.655 103.880 ;
        RECT 41.075 103.250 41.445 103.880 ;
        RECT 37.655 103.240 37.885 103.250 ;
        RECT 38.445 103.240 38.675 103.250 ;
        RECT 40.355 103.240 40.585 103.250 ;
        RECT 41.145 103.240 41.375 103.250 ;
        RECT 37.935 102.850 38.395 103.080 ;
        RECT 40.635 102.850 41.095 103.080 ;
        RECT 42.985 100.700 43.355 103.880 ;
        RECT 43.775 100.700 44.145 103.880 ;
        RECT 45.685 100.700 46.055 103.880 ;
        RECT 46.475 100.700 46.845 103.880 ;
        RECT 29.300 98.740 30.475 99.855 ;
        RECT 34.215 98.745 34.585 99.860 ;
        RECT 27.295 82.325 28.355 83.325 ;
        RECT 27.325 82.295 28.325 82.325 ;
        RECT 6.570 81.455 7.610 81.950 ;
        RECT 9.810 81.475 10.270 81.705 ;
        RECT 11.970 81.455 13.010 81.950 ;
        RECT 14.670 81.455 15.710 81.950 ;
        RECT 17.910 81.475 18.370 81.705 ;
        RECT 20.610 81.475 21.070 81.705 ;
        RECT 6.830 81.305 7.060 81.315 ;
        RECT 7.620 81.305 7.850 81.315 ;
        RECT 9.530 81.305 9.760 81.315 ;
        RECT 10.320 81.305 10.550 81.315 ;
        RECT 12.230 81.305 12.460 81.315 ;
        RECT 13.020 81.305 13.250 81.315 ;
        RECT 14.930 81.305 15.160 81.315 ;
        RECT 15.720 81.305 15.950 81.315 ;
        RECT 17.630 81.305 17.860 81.315 ;
        RECT 18.420 81.305 18.650 81.315 ;
        RECT 20.330 81.305 20.560 81.315 ;
        RECT 21.120 81.305 21.350 81.315 ;
        RECT 6.085 80.675 7.130 81.305 ;
        RECT 7.550 80.675 7.920 81.305 ;
        RECT 6.830 80.665 7.060 80.675 ;
        RECT 7.620 80.665 7.850 80.675 ;
        RECT 7.110 80.275 7.570 80.505 ;
        RECT 9.460 78.125 9.830 81.305 ;
        RECT 10.250 78.125 10.620 81.305 ;
        RECT 11.485 80.675 12.530 81.305 ;
        RECT 12.950 80.675 13.320 81.305 ;
        RECT 14.185 80.675 15.230 81.305 ;
        RECT 15.650 80.675 16.020 81.305 ;
        RECT 12.230 80.665 12.460 80.675 ;
        RECT 13.020 80.665 13.250 80.675 ;
        RECT 14.930 80.665 15.160 80.675 ;
        RECT 15.720 80.665 15.950 80.675 ;
        RECT 12.510 80.275 12.970 80.505 ;
        RECT 15.210 80.275 15.670 80.505 ;
        RECT 17.560 78.125 17.930 81.305 ;
        RECT 18.350 78.125 18.720 81.305 ;
        RECT 20.260 78.125 20.630 81.305 ;
        RECT 21.050 78.125 21.420 81.305 ;
        RECT 3.860 76.170 5.060 77.285 ;
        RECT 8.790 76.170 9.160 77.285 ;
        RECT 3.905 76.140 5.020 76.170 ;
        RECT 9.530 74.815 9.760 78.125 ;
        RECT 10.320 74.815 10.550 78.125 ;
        RECT 10.920 76.170 11.290 77.285 ;
        RECT 16.890 76.170 17.260 77.285 ;
        RECT 17.630 74.815 17.860 78.125 ;
        RECT 18.420 74.815 18.650 78.125 ;
        RECT 19.020 76.170 19.390 77.285 ;
        RECT 19.590 76.170 19.960 77.285 ;
        RECT 20.330 74.815 20.560 78.125 ;
        RECT 21.120 74.815 21.350 78.125 ;
        RECT 21.720 76.170 22.090 77.285 ;
        RECT 23.090 76.140 24.205 81.855 ;
        RECT 29.330 77.285 30.445 98.740 ;
        RECT 34.955 97.390 35.185 100.700 ;
        RECT 35.745 97.390 35.975 100.700 ;
        RECT 36.345 98.745 36.715 99.860 ;
        RECT 42.315 98.745 42.685 99.860 ;
        RECT 43.055 97.390 43.285 100.700 ;
        RECT 43.845 97.390 44.075 100.700 ;
        RECT 44.445 98.745 44.815 99.860 ;
        RECT 45.015 98.745 45.385 99.860 ;
        RECT 45.755 97.390 45.985 100.700 ;
        RECT 46.545 97.390 46.775 100.700 ;
        RECT 47.145 98.745 47.515 99.860 ;
        RECT 48.510 98.745 49.685 99.860 ;
        RECT 35.235 97.200 35.695 97.230 ;
        RECT 43.335 97.200 43.795 97.230 ;
        RECT 46.035 97.200 46.495 97.230 ;
        RECT 34.975 96.800 35.975 97.200 ;
        RECT 43.075 96.800 44.075 97.200 ;
        RECT 45.775 96.800 46.775 97.200 ;
        RECT 48.540 95.770 49.655 98.745 ;
        RECT 37.150 95.025 38.150 95.055 ;
        RECT 40.825 95.025 41.825 95.055 ;
        RECT 34.975 94.575 35.975 95.025 ;
        RECT 35.235 94.565 35.695 94.575 ;
        RECT 34.215 91.970 34.585 93.075 ;
        RECT 34.955 89.350 35.185 94.360 ;
        RECT 35.745 89.350 35.975 94.360 ;
        RECT 37.150 93.995 39.075 95.025 ;
        RECT 36.345 93.025 36.715 93.075 ;
        RECT 36.345 91.970 37.450 93.025 ;
        RECT 32.535 85.565 32.995 85.795 ;
        RECT 32.255 85.350 32.485 85.360 ;
        RECT 33.045 85.350 33.275 85.360 ;
        RECT 31.510 84.370 32.555 85.350 ;
        RECT 32.975 84.370 33.345 85.350 ;
        RECT 34.885 84.370 35.255 89.350 ;
        RECT 35.675 84.370 36.045 89.350 ;
        RECT 36.450 87.275 37.450 91.970 ;
        RECT 38.075 88.925 39.075 93.995 ;
        RECT 39.875 93.995 41.825 95.025 ;
        RECT 43.075 94.575 44.075 95.025 ;
        RECT 45.775 94.575 46.775 95.025 ;
        RECT 43.335 94.565 43.795 94.575 ;
        RECT 46.035 94.565 46.495 94.575 ;
        RECT 39.875 89.670 40.875 93.995 ;
        RECT 42.315 93.025 42.685 93.075 ;
        RECT 41.600 91.970 42.685 93.025 ;
        RECT 38.075 87.925 40.905 88.925 ;
        RECT 41.600 87.275 42.600 91.970 ;
        RECT 43.055 89.350 43.285 94.360 ;
        RECT 43.845 89.350 44.075 94.360 ;
        RECT 44.445 91.970 44.815 93.075 ;
        RECT 45.015 91.970 45.385 93.075 ;
        RECT 45.755 89.350 45.985 94.360 ;
        RECT 46.545 89.350 46.775 94.360 ;
        RECT 48.855 93.115 49.305 95.425 ;
        RECT 47.145 91.970 47.515 93.075 ;
        RECT 36.450 86.275 42.600 87.275 ;
        RECT 37.935 85.565 38.395 85.795 ;
        RECT 40.635 85.565 41.095 85.795 ;
        RECT 37.655 85.350 37.885 85.360 ;
        RECT 38.445 85.350 38.675 85.360 ;
        RECT 40.355 85.350 40.585 85.360 ;
        RECT 41.145 85.350 41.375 85.360 ;
        RECT 36.910 84.370 37.955 85.350 ;
        RECT 38.375 84.370 38.745 85.350 ;
        RECT 39.610 84.370 40.655 85.350 ;
        RECT 41.075 84.370 41.445 85.350 ;
        RECT 42.985 84.370 43.355 89.350 ;
        RECT 43.775 84.370 44.145 89.350 ;
        RECT 45.685 84.370 46.055 89.350 ;
        RECT 46.475 84.370 46.845 89.350 ;
        RECT 32.255 84.360 32.485 84.370 ;
        RECT 33.045 84.360 33.275 84.370 ;
        RECT 34.955 84.360 35.185 84.370 ;
        RECT 35.745 84.360 35.975 84.370 ;
        RECT 37.655 84.360 37.885 84.370 ;
        RECT 38.445 84.360 38.675 84.370 ;
        RECT 40.355 84.360 40.585 84.370 ;
        RECT 41.145 84.360 41.375 84.370 ;
        RECT 43.055 84.360 43.285 84.370 ;
        RECT 43.845 84.360 44.075 84.370 ;
        RECT 45.755 84.360 45.985 84.370 ;
        RECT 46.545 84.360 46.775 84.370 ;
        RECT 32.000 83.700 33.035 84.175 ;
        RECT 35.235 83.925 35.695 84.155 ;
        RECT 37.400 83.700 38.435 84.175 ;
        RECT 40.100 83.700 41.135 84.175 ;
        RECT 43.335 83.925 43.795 84.155 ;
        RECT 46.035 83.925 46.495 84.155 ;
        RECT 48.855 82.205 49.305 84.515 ;
        RECT 52.750 83.325 53.750 104.900 ;
        RECT 54.755 99.855 55.870 121.315 ;
        RECT 60.380 119.965 60.610 123.275 ;
        RECT 61.170 119.965 61.400 123.275 ;
        RECT 61.770 121.320 62.140 122.435 ;
        RECT 67.740 121.320 68.110 122.435 ;
        RECT 68.480 119.965 68.710 123.275 ;
        RECT 69.270 119.965 69.500 123.275 ;
        RECT 69.870 121.320 70.240 122.435 ;
        RECT 70.440 121.320 70.810 122.435 ;
        RECT 71.180 119.965 71.410 123.275 ;
        RECT 71.970 119.965 72.200 123.275 ;
        RECT 78.175 123.250 81.225 124.250 ;
        RECT 85.735 123.275 86.105 126.455 ;
        RECT 86.525 123.275 86.895 126.455 ;
        RECT 87.760 125.825 88.805 126.455 ;
        RECT 89.225 125.825 89.595 126.455 ;
        RECT 90.460 125.825 91.505 126.455 ;
        RECT 91.925 125.825 92.295 126.455 ;
        RECT 88.505 125.815 88.735 125.825 ;
        RECT 89.295 125.815 89.525 125.825 ;
        RECT 91.205 125.815 91.435 125.825 ;
        RECT 91.995 125.815 92.225 125.825 ;
        RECT 88.785 125.425 89.245 125.655 ;
        RECT 91.485 125.425 91.945 125.655 ;
        RECT 93.835 123.275 94.205 126.455 ;
        RECT 94.625 123.275 94.995 126.455 ;
        RECT 96.535 123.275 96.905 126.455 ;
        RECT 97.325 123.275 97.695 126.455 ;
        RECT 105.650 124.250 106.650 127.475 ;
        RECT 126.520 127.405 132.130 128.510 ;
        RECT 152.425 128.475 153.425 141.550 ;
        RECT 152.395 127.475 153.455 128.475 ;
        RECT 108.270 126.605 109.310 127.100 ;
        RECT 111.510 126.625 111.970 126.855 ;
        RECT 113.670 126.605 114.710 127.100 ;
        RECT 116.370 126.605 117.410 127.100 ;
        RECT 119.610 126.625 120.070 126.855 ;
        RECT 122.310 126.625 122.770 126.855 ;
        RECT 108.530 126.455 108.760 126.465 ;
        RECT 109.320 126.455 109.550 126.465 ;
        RECT 111.230 126.455 111.460 126.465 ;
        RECT 112.020 126.455 112.250 126.465 ;
        RECT 113.930 126.455 114.160 126.465 ;
        RECT 114.720 126.455 114.950 126.465 ;
        RECT 116.630 126.455 116.860 126.465 ;
        RECT 117.420 126.455 117.650 126.465 ;
        RECT 119.330 126.455 119.560 126.465 ;
        RECT 120.120 126.455 120.350 126.465 ;
        RECT 122.030 126.455 122.260 126.465 ;
        RECT 122.820 126.455 123.050 126.465 ;
        RECT 107.785 125.825 108.830 126.455 ;
        RECT 109.250 125.825 109.620 126.455 ;
        RECT 108.530 125.815 108.760 125.825 ;
        RECT 109.320 125.815 109.550 125.825 ;
        RECT 108.810 125.425 109.270 125.655 ;
        RECT 72.570 121.320 72.940 122.435 ;
        RECT 60.660 119.775 61.120 119.805 ;
        RECT 68.760 119.775 69.220 119.805 ;
        RECT 71.460 119.775 71.920 119.805 ;
        RECT 60.400 119.375 61.400 119.775 ;
        RECT 68.500 119.375 69.500 119.775 ;
        RECT 71.200 119.375 72.200 119.775 ;
        RECT 62.575 117.600 63.575 117.630 ;
        RECT 66.250 117.600 67.250 117.630 ;
        RECT 60.400 117.150 61.400 117.600 ;
        RECT 60.660 117.140 61.120 117.150 ;
        RECT 59.640 114.545 60.010 115.650 ;
        RECT 60.380 111.925 60.610 116.935 ;
        RECT 61.170 111.925 61.400 116.935 ;
        RECT 62.575 116.570 64.500 117.600 ;
        RECT 61.770 115.600 62.140 115.650 ;
        RECT 61.770 114.545 62.875 115.600 ;
        RECT 57.960 108.140 58.420 108.370 ;
        RECT 57.680 107.925 57.910 107.935 ;
        RECT 58.470 107.925 58.700 107.935 ;
        RECT 56.935 106.945 57.980 107.925 ;
        RECT 58.400 106.945 58.770 107.925 ;
        RECT 60.310 106.945 60.680 111.925 ;
        RECT 61.100 106.945 61.470 111.925 ;
        RECT 61.875 109.850 62.875 114.545 ;
        RECT 63.500 111.500 64.500 116.570 ;
        RECT 65.300 116.570 67.250 117.600 ;
        RECT 68.500 117.150 69.500 117.600 ;
        RECT 71.200 117.150 72.200 117.600 ;
        RECT 68.760 117.140 69.220 117.150 ;
        RECT 71.460 117.140 71.920 117.150 ;
        RECT 65.300 112.245 66.300 116.570 ;
        RECT 67.740 115.600 68.110 115.650 ;
        RECT 67.025 114.545 68.110 115.600 ;
        RECT 63.500 110.500 66.330 111.500 ;
        RECT 67.025 109.850 68.025 114.545 ;
        RECT 68.480 111.925 68.710 116.935 ;
        RECT 69.270 111.925 69.500 116.935 ;
        RECT 69.870 114.545 70.240 115.650 ;
        RECT 70.440 114.545 70.810 115.650 ;
        RECT 71.180 111.925 71.410 116.935 ;
        RECT 71.970 111.925 72.200 116.935 ;
        RECT 72.570 114.545 72.940 115.650 ;
        RECT 61.875 108.850 68.025 109.850 ;
        RECT 63.360 108.140 63.820 108.370 ;
        RECT 66.060 108.140 66.520 108.370 ;
        RECT 63.080 107.925 63.310 107.935 ;
        RECT 63.870 107.925 64.100 107.935 ;
        RECT 65.780 107.925 66.010 107.935 ;
        RECT 66.570 107.925 66.800 107.935 ;
        RECT 62.335 106.945 63.380 107.925 ;
        RECT 63.800 106.945 64.170 107.925 ;
        RECT 65.035 106.945 66.080 107.925 ;
        RECT 66.500 106.945 66.870 107.925 ;
        RECT 68.410 106.945 68.780 111.925 ;
        RECT 69.200 106.945 69.570 111.925 ;
        RECT 71.110 106.945 71.480 111.925 ;
        RECT 71.900 106.945 72.270 111.925 ;
        RECT 57.680 106.935 57.910 106.945 ;
        RECT 58.470 106.935 58.700 106.945 ;
        RECT 60.380 106.935 60.610 106.945 ;
        RECT 61.170 106.935 61.400 106.945 ;
        RECT 63.080 106.935 63.310 106.945 ;
        RECT 63.870 106.935 64.100 106.945 ;
        RECT 65.780 106.935 66.010 106.945 ;
        RECT 66.570 106.935 66.800 106.945 ;
        RECT 68.480 106.935 68.710 106.945 ;
        RECT 69.270 106.935 69.500 106.945 ;
        RECT 71.180 106.935 71.410 106.945 ;
        RECT 71.970 106.935 72.200 106.945 ;
        RECT 57.425 106.275 58.460 106.750 ;
        RECT 60.660 106.500 61.120 106.730 ;
        RECT 62.825 106.275 63.860 106.750 ;
        RECT 65.525 106.275 66.560 106.750 ;
        RECT 68.760 106.500 69.220 106.730 ;
        RECT 71.460 106.500 71.920 106.730 ;
        RECT 78.175 105.900 79.175 123.250 ;
        RECT 80.180 122.430 81.295 122.485 ;
        RECT 80.150 121.315 81.325 122.430 ;
        RECT 85.065 121.320 85.435 122.435 ;
        RECT 78.145 104.900 79.205 105.900 ;
        RECT 57.420 104.030 58.460 104.525 ;
        RECT 60.660 104.050 61.120 104.280 ;
        RECT 62.820 104.030 63.860 104.525 ;
        RECT 65.520 104.030 66.560 104.525 ;
        RECT 68.760 104.050 69.220 104.280 ;
        RECT 71.460 104.050 71.920 104.280 ;
        RECT 57.680 103.880 57.910 103.890 ;
        RECT 58.470 103.880 58.700 103.890 ;
        RECT 60.380 103.880 60.610 103.890 ;
        RECT 61.170 103.880 61.400 103.890 ;
        RECT 63.080 103.880 63.310 103.890 ;
        RECT 63.870 103.880 64.100 103.890 ;
        RECT 65.780 103.880 66.010 103.890 ;
        RECT 66.570 103.880 66.800 103.890 ;
        RECT 68.480 103.880 68.710 103.890 ;
        RECT 69.270 103.880 69.500 103.890 ;
        RECT 71.180 103.880 71.410 103.890 ;
        RECT 71.970 103.880 72.200 103.890 ;
        RECT 56.935 103.250 57.980 103.880 ;
        RECT 58.400 103.250 58.770 103.880 ;
        RECT 57.680 103.240 57.910 103.250 ;
        RECT 58.470 103.240 58.700 103.250 ;
        RECT 57.960 102.850 58.420 103.080 ;
        RECT 60.310 100.700 60.680 103.880 ;
        RECT 61.100 100.700 61.470 103.880 ;
        RECT 62.335 103.250 63.380 103.880 ;
        RECT 63.800 103.250 64.170 103.880 ;
        RECT 65.035 103.250 66.080 103.880 ;
        RECT 66.500 103.250 66.870 103.880 ;
        RECT 63.080 103.240 63.310 103.250 ;
        RECT 63.870 103.240 64.100 103.250 ;
        RECT 65.780 103.240 66.010 103.250 ;
        RECT 66.570 103.240 66.800 103.250 ;
        RECT 63.360 102.850 63.820 103.080 ;
        RECT 66.060 102.850 66.520 103.080 ;
        RECT 68.410 100.700 68.780 103.880 ;
        RECT 69.200 100.700 69.570 103.880 ;
        RECT 71.110 100.700 71.480 103.880 ;
        RECT 71.900 100.700 72.270 103.880 ;
        RECT 54.725 98.740 55.900 99.855 ;
        RECT 59.640 98.745 60.010 99.860 ;
        RECT 52.720 82.325 53.780 83.325 ;
        RECT 52.750 82.295 53.750 82.325 ;
        RECT 31.995 81.455 33.035 81.950 ;
        RECT 35.235 81.475 35.695 81.705 ;
        RECT 37.395 81.455 38.435 81.950 ;
        RECT 40.095 81.455 41.135 81.950 ;
        RECT 43.335 81.475 43.795 81.705 ;
        RECT 46.035 81.475 46.495 81.705 ;
        RECT 32.255 81.305 32.485 81.315 ;
        RECT 33.045 81.305 33.275 81.315 ;
        RECT 34.955 81.305 35.185 81.315 ;
        RECT 35.745 81.305 35.975 81.315 ;
        RECT 37.655 81.305 37.885 81.315 ;
        RECT 38.445 81.305 38.675 81.315 ;
        RECT 40.355 81.305 40.585 81.315 ;
        RECT 41.145 81.305 41.375 81.315 ;
        RECT 43.055 81.305 43.285 81.315 ;
        RECT 43.845 81.305 44.075 81.315 ;
        RECT 45.755 81.305 45.985 81.315 ;
        RECT 46.545 81.305 46.775 81.315 ;
        RECT 31.510 80.675 32.555 81.305 ;
        RECT 32.975 80.675 33.345 81.305 ;
        RECT 32.255 80.665 32.485 80.675 ;
        RECT 33.045 80.665 33.275 80.675 ;
        RECT 32.535 80.275 32.995 80.505 ;
        RECT 34.885 78.125 35.255 81.305 ;
        RECT 35.675 78.125 36.045 81.305 ;
        RECT 36.910 80.675 37.955 81.305 ;
        RECT 38.375 80.675 38.745 81.305 ;
        RECT 39.610 80.675 40.655 81.305 ;
        RECT 41.075 80.675 41.445 81.305 ;
        RECT 37.655 80.665 37.885 80.675 ;
        RECT 38.445 80.665 38.675 80.675 ;
        RECT 40.355 80.665 40.585 80.675 ;
        RECT 41.145 80.665 41.375 80.675 ;
        RECT 37.935 80.275 38.395 80.505 ;
        RECT 40.635 80.275 41.095 80.505 ;
        RECT 42.985 78.125 43.355 81.305 ;
        RECT 43.775 78.125 44.145 81.305 ;
        RECT 45.685 78.125 46.055 81.305 ;
        RECT 46.475 78.125 46.845 81.305 ;
        RECT 29.285 76.170 30.485 77.285 ;
        RECT 34.215 76.170 34.585 77.285 ;
        RECT 29.330 76.140 30.445 76.170 ;
        RECT 34.955 74.815 35.185 78.125 ;
        RECT 35.745 74.815 35.975 78.125 ;
        RECT 36.345 76.170 36.715 77.285 ;
        RECT 42.315 76.170 42.685 77.285 ;
        RECT 43.055 74.815 43.285 78.125 ;
        RECT 43.845 74.815 44.075 78.125 ;
        RECT 44.445 76.170 44.815 77.285 ;
        RECT 45.015 76.170 45.385 77.285 ;
        RECT 45.755 74.815 45.985 78.125 ;
        RECT 46.545 74.815 46.775 78.125 ;
        RECT 47.145 76.170 47.515 77.285 ;
        RECT 48.515 76.140 49.630 81.855 ;
        RECT 54.755 77.285 55.870 98.740 ;
        RECT 60.380 97.390 60.610 100.700 ;
        RECT 61.170 97.390 61.400 100.700 ;
        RECT 61.770 98.745 62.140 99.860 ;
        RECT 67.740 98.745 68.110 99.860 ;
        RECT 68.480 97.390 68.710 100.700 ;
        RECT 69.270 97.390 69.500 100.700 ;
        RECT 69.870 98.745 70.240 99.860 ;
        RECT 70.440 98.745 70.810 99.860 ;
        RECT 71.180 97.390 71.410 100.700 ;
        RECT 71.970 97.390 72.200 100.700 ;
        RECT 72.570 98.745 72.940 99.860 ;
        RECT 73.935 98.745 75.110 99.860 ;
        RECT 60.660 97.200 61.120 97.230 ;
        RECT 68.760 97.200 69.220 97.230 ;
        RECT 71.460 97.200 71.920 97.230 ;
        RECT 60.400 96.800 61.400 97.200 ;
        RECT 68.500 96.800 69.500 97.200 ;
        RECT 71.200 96.800 72.200 97.200 ;
        RECT 73.965 95.770 75.080 98.745 ;
        RECT 62.575 95.025 63.575 95.055 ;
        RECT 66.250 95.025 67.250 95.055 ;
        RECT 60.400 94.575 61.400 95.025 ;
        RECT 60.660 94.565 61.120 94.575 ;
        RECT 59.640 91.970 60.010 93.075 ;
        RECT 60.380 89.350 60.610 94.360 ;
        RECT 61.170 89.350 61.400 94.360 ;
        RECT 62.575 93.995 64.500 95.025 ;
        RECT 61.770 93.025 62.140 93.075 ;
        RECT 61.770 91.970 62.875 93.025 ;
        RECT 57.960 85.565 58.420 85.795 ;
        RECT 57.680 85.350 57.910 85.360 ;
        RECT 58.470 85.350 58.700 85.360 ;
        RECT 56.935 84.370 57.980 85.350 ;
        RECT 58.400 84.370 58.770 85.350 ;
        RECT 60.310 84.370 60.680 89.350 ;
        RECT 61.100 84.370 61.470 89.350 ;
        RECT 61.875 87.275 62.875 91.970 ;
        RECT 63.500 88.925 64.500 93.995 ;
        RECT 65.300 93.995 67.250 95.025 ;
        RECT 68.500 94.575 69.500 95.025 ;
        RECT 71.200 94.575 72.200 95.025 ;
        RECT 68.760 94.565 69.220 94.575 ;
        RECT 71.460 94.565 71.920 94.575 ;
        RECT 65.300 89.670 66.300 93.995 ;
        RECT 67.740 93.025 68.110 93.075 ;
        RECT 67.025 91.970 68.110 93.025 ;
        RECT 63.500 87.925 66.330 88.925 ;
        RECT 67.025 87.275 68.025 91.970 ;
        RECT 68.480 89.350 68.710 94.360 ;
        RECT 69.270 89.350 69.500 94.360 ;
        RECT 69.870 91.970 70.240 93.075 ;
        RECT 70.440 91.970 70.810 93.075 ;
        RECT 71.180 89.350 71.410 94.360 ;
        RECT 71.970 89.350 72.200 94.360 ;
        RECT 74.280 93.115 74.730 95.425 ;
        RECT 72.570 91.970 72.940 93.075 ;
        RECT 61.875 86.275 68.025 87.275 ;
        RECT 63.360 85.565 63.820 85.795 ;
        RECT 66.060 85.565 66.520 85.795 ;
        RECT 63.080 85.350 63.310 85.360 ;
        RECT 63.870 85.350 64.100 85.360 ;
        RECT 65.780 85.350 66.010 85.360 ;
        RECT 66.570 85.350 66.800 85.360 ;
        RECT 62.335 84.370 63.380 85.350 ;
        RECT 63.800 84.370 64.170 85.350 ;
        RECT 65.035 84.370 66.080 85.350 ;
        RECT 66.500 84.370 66.870 85.350 ;
        RECT 68.410 84.370 68.780 89.350 ;
        RECT 69.200 84.370 69.570 89.350 ;
        RECT 71.110 84.370 71.480 89.350 ;
        RECT 71.900 84.370 72.270 89.350 ;
        RECT 57.680 84.360 57.910 84.370 ;
        RECT 58.470 84.360 58.700 84.370 ;
        RECT 60.380 84.360 60.610 84.370 ;
        RECT 61.170 84.360 61.400 84.370 ;
        RECT 63.080 84.360 63.310 84.370 ;
        RECT 63.870 84.360 64.100 84.370 ;
        RECT 65.780 84.360 66.010 84.370 ;
        RECT 66.570 84.360 66.800 84.370 ;
        RECT 68.480 84.360 68.710 84.370 ;
        RECT 69.270 84.360 69.500 84.370 ;
        RECT 71.180 84.360 71.410 84.370 ;
        RECT 71.970 84.360 72.200 84.370 ;
        RECT 57.425 83.700 58.460 84.175 ;
        RECT 60.660 83.925 61.120 84.155 ;
        RECT 62.825 83.700 63.860 84.175 ;
        RECT 65.525 83.700 66.560 84.175 ;
        RECT 68.760 83.925 69.220 84.155 ;
        RECT 71.460 83.925 71.920 84.155 ;
        RECT 74.280 82.205 74.730 84.515 ;
        RECT 78.175 83.325 79.175 104.900 ;
        RECT 80.180 99.855 81.295 121.315 ;
        RECT 85.805 119.965 86.035 123.275 ;
        RECT 86.595 119.965 86.825 123.275 ;
        RECT 87.195 121.320 87.565 122.435 ;
        RECT 93.165 121.320 93.535 122.435 ;
        RECT 93.905 119.965 94.135 123.275 ;
        RECT 94.695 119.965 94.925 123.275 ;
        RECT 95.295 121.320 95.665 122.435 ;
        RECT 95.865 121.320 96.235 122.435 ;
        RECT 96.605 119.965 96.835 123.275 ;
        RECT 97.395 119.965 97.625 123.275 ;
        RECT 103.600 123.250 106.650 124.250 ;
        RECT 111.160 123.275 111.530 126.455 ;
        RECT 111.950 123.275 112.320 126.455 ;
        RECT 113.185 125.825 114.230 126.455 ;
        RECT 114.650 125.825 115.020 126.455 ;
        RECT 115.885 125.825 116.930 126.455 ;
        RECT 117.350 125.825 117.720 126.455 ;
        RECT 113.930 125.815 114.160 125.825 ;
        RECT 114.720 125.815 114.950 125.825 ;
        RECT 116.630 125.815 116.860 125.825 ;
        RECT 117.420 125.815 117.650 125.825 ;
        RECT 114.210 125.425 114.670 125.655 ;
        RECT 116.910 125.425 117.370 125.655 ;
        RECT 119.260 123.275 119.630 126.455 ;
        RECT 120.050 123.275 120.420 126.455 ;
        RECT 121.960 123.275 122.330 126.455 ;
        RECT 122.750 123.275 123.120 126.455 ;
        RECT 131.075 124.250 132.075 127.405 ;
        RECT 133.695 126.605 134.735 127.100 ;
        RECT 136.935 126.625 137.395 126.855 ;
        RECT 139.095 126.605 140.135 127.100 ;
        RECT 141.795 126.605 142.835 127.100 ;
        RECT 145.035 126.625 145.495 126.855 ;
        RECT 147.735 126.625 148.195 126.855 ;
        RECT 133.955 126.455 134.185 126.465 ;
        RECT 134.745 126.455 134.975 126.465 ;
        RECT 136.655 126.455 136.885 126.465 ;
        RECT 137.445 126.455 137.675 126.465 ;
        RECT 139.355 126.455 139.585 126.465 ;
        RECT 140.145 126.455 140.375 126.465 ;
        RECT 142.055 126.455 142.285 126.465 ;
        RECT 142.845 126.455 143.075 126.465 ;
        RECT 144.755 126.455 144.985 126.465 ;
        RECT 145.545 126.455 145.775 126.465 ;
        RECT 147.455 126.455 147.685 126.465 ;
        RECT 148.245 126.455 148.475 126.465 ;
        RECT 133.210 125.825 134.255 126.455 ;
        RECT 134.675 125.825 135.045 126.455 ;
        RECT 133.955 125.815 134.185 125.825 ;
        RECT 134.745 125.815 134.975 125.825 ;
        RECT 134.235 125.425 134.695 125.655 ;
        RECT 97.995 121.320 98.365 122.435 ;
        RECT 86.085 119.775 86.545 119.805 ;
        RECT 94.185 119.775 94.645 119.805 ;
        RECT 96.885 119.775 97.345 119.805 ;
        RECT 85.825 119.375 86.825 119.775 ;
        RECT 93.925 119.375 94.925 119.775 ;
        RECT 96.625 119.375 97.625 119.775 ;
        RECT 88.000 117.600 89.000 117.630 ;
        RECT 91.675 117.600 92.675 117.630 ;
        RECT 85.825 117.150 86.825 117.600 ;
        RECT 86.085 117.140 86.545 117.150 ;
        RECT 85.065 114.545 85.435 115.650 ;
        RECT 85.805 111.925 86.035 116.935 ;
        RECT 86.595 111.925 86.825 116.935 ;
        RECT 88.000 116.570 89.925 117.600 ;
        RECT 87.195 115.600 87.565 115.650 ;
        RECT 87.195 114.545 88.300 115.600 ;
        RECT 83.385 108.140 83.845 108.370 ;
        RECT 83.105 107.925 83.335 107.935 ;
        RECT 83.895 107.925 84.125 107.935 ;
        RECT 82.360 106.945 83.405 107.925 ;
        RECT 83.825 106.945 84.195 107.925 ;
        RECT 85.735 106.945 86.105 111.925 ;
        RECT 86.525 106.945 86.895 111.925 ;
        RECT 87.300 109.850 88.300 114.545 ;
        RECT 88.925 111.500 89.925 116.570 ;
        RECT 90.725 116.570 92.675 117.600 ;
        RECT 93.925 117.150 94.925 117.600 ;
        RECT 96.625 117.150 97.625 117.600 ;
        RECT 94.185 117.140 94.645 117.150 ;
        RECT 96.885 117.140 97.345 117.150 ;
        RECT 90.725 112.245 91.725 116.570 ;
        RECT 93.165 115.600 93.535 115.650 ;
        RECT 92.450 114.545 93.535 115.600 ;
        RECT 88.925 110.500 91.755 111.500 ;
        RECT 92.450 109.850 93.450 114.545 ;
        RECT 93.905 111.925 94.135 116.935 ;
        RECT 94.695 111.925 94.925 116.935 ;
        RECT 95.295 114.545 95.665 115.650 ;
        RECT 95.865 114.545 96.235 115.650 ;
        RECT 96.605 111.925 96.835 116.935 ;
        RECT 97.395 111.925 97.625 116.935 ;
        RECT 97.995 114.545 98.365 115.650 ;
        RECT 87.300 108.850 93.450 109.850 ;
        RECT 88.785 108.140 89.245 108.370 ;
        RECT 91.485 108.140 91.945 108.370 ;
        RECT 88.505 107.925 88.735 107.935 ;
        RECT 89.295 107.925 89.525 107.935 ;
        RECT 91.205 107.925 91.435 107.935 ;
        RECT 91.995 107.925 92.225 107.935 ;
        RECT 87.760 106.945 88.805 107.925 ;
        RECT 89.225 106.945 89.595 107.925 ;
        RECT 90.460 106.945 91.505 107.925 ;
        RECT 91.925 106.945 92.295 107.925 ;
        RECT 93.835 106.945 94.205 111.925 ;
        RECT 94.625 106.945 94.995 111.925 ;
        RECT 96.535 106.945 96.905 111.925 ;
        RECT 97.325 106.945 97.695 111.925 ;
        RECT 83.105 106.935 83.335 106.945 ;
        RECT 83.895 106.935 84.125 106.945 ;
        RECT 85.805 106.935 86.035 106.945 ;
        RECT 86.595 106.935 86.825 106.945 ;
        RECT 88.505 106.935 88.735 106.945 ;
        RECT 89.295 106.935 89.525 106.945 ;
        RECT 91.205 106.935 91.435 106.945 ;
        RECT 91.995 106.935 92.225 106.945 ;
        RECT 93.905 106.935 94.135 106.945 ;
        RECT 94.695 106.935 94.925 106.945 ;
        RECT 96.605 106.935 96.835 106.945 ;
        RECT 97.395 106.935 97.625 106.945 ;
        RECT 82.850 106.275 83.885 106.750 ;
        RECT 86.085 106.500 86.545 106.730 ;
        RECT 88.250 106.275 89.285 106.750 ;
        RECT 90.950 106.275 91.985 106.750 ;
        RECT 94.185 106.500 94.645 106.730 ;
        RECT 96.885 106.500 97.345 106.730 ;
        RECT 103.600 105.900 104.600 123.250 ;
        RECT 105.605 122.430 106.720 122.485 ;
        RECT 105.575 121.315 106.750 122.430 ;
        RECT 110.490 121.320 110.860 122.435 ;
        RECT 103.570 104.900 104.630 105.900 ;
        RECT 82.845 104.030 83.885 104.525 ;
        RECT 86.085 104.050 86.545 104.280 ;
        RECT 88.245 104.030 89.285 104.525 ;
        RECT 90.945 104.030 91.985 104.525 ;
        RECT 94.185 104.050 94.645 104.280 ;
        RECT 96.885 104.050 97.345 104.280 ;
        RECT 83.105 103.880 83.335 103.890 ;
        RECT 83.895 103.880 84.125 103.890 ;
        RECT 85.805 103.880 86.035 103.890 ;
        RECT 86.595 103.880 86.825 103.890 ;
        RECT 88.505 103.880 88.735 103.890 ;
        RECT 89.295 103.880 89.525 103.890 ;
        RECT 91.205 103.880 91.435 103.890 ;
        RECT 91.995 103.880 92.225 103.890 ;
        RECT 93.905 103.880 94.135 103.890 ;
        RECT 94.695 103.880 94.925 103.890 ;
        RECT 96.605 103.880 96.835 103.890 ;
        RECT 97.395 103.880 97.625 103.890 ;
        RECT 82.360 103.250 83.405 103.880 ;
        RECT 83.825 103.250 84.195 103.880 ;
        RECT 83.105 103.240 83.335 103.250 ;
        RECT 83.895 103.240 84.125 103.250 ;
        RECT 83.385 102.850 83.845 103.080 ;
        RECT 85.735 100.700 86.105 103.880 ;
        RECT 86.525 100.700 86.895 103.880 ;
        RECT 87.760 103.250 88.805 103.880 ;
        RECT 89.225 103.250 89.595 103.880 ;
        RECT 90.460 103.250 91.505 103.880 ;
        RECT 91.925 103.250 92.295 103.880 ;
        RECT 88.505 103.240 88.735 103.250 ;
        RECT 89.295 103.240 89.525 103.250 ;
        RECT 91.205 103.240 91.435 103.250 ;
        RECT 91.995 103.240 92.225 103.250 ;
        RECT 88.785 102.850 89.245 103.080 ;
        RECT 91.485 102.850 91.945 103.080 ;
        RECT 93.835 100.700 94.205 103.880 ;
        RECT 94.625 100.700 94.995 103.880 ;
        RECT 96.535 100.700 96.905 103.880 ;
        RECT 97.325 100.700 97.695 103.880 ;
        RECT 80.150 98.740 81.325 99.855 ;
        RECT 85.065 98.745 85.435 99.860 ;
        RECT 78.145 82.325 79.205 83.325 ;
        RECT 78.175 82.295 79.175 82.325 ;
        RECT 57.420 81.455 58.460 81.950 ;
        RECT 60.660 81.475 61.120 81.705 ;
        RECT 62.820 81.455 63.860 81.950 ;
        RECT 65.520 81.455 66.560 81.950 ;
        RECT 68.760 81.475 69.220 81.705 ;
        RECT 71.460 81.475 71.920 81.705 ;
        RECT 57.680 81.305 57.910 81.315 ;
        RECT 58.470 81.305 58.700 81.315 ;
        RECT 60.380 81.305 60.610 81.315 ;
        RECT 61.170 81.305 61.400 81.315 ;
        RECT 63.080 81.305 63.310 81.315 ;
        RECT 63.870 81.305 64.100 81.315 ;
        RECT 65.780 81.305 66.010 81.315 ;
        RECT 66.570 81.305 66.800 81.315 ;
        RECT 68.480 81.305 68.710 81.315 ;
        RECT 69.270 81.305 69.500 81.315 ;
        RECT 71.180 81.305 71.410 81.315 ;
        RECT 71.970 81.305 72.200 81.315 ;
        RECT 56.935 80.675 57.980 81.305 ;
        RECT 58.400 80.675 58.770 81.305 ;
        RECT 57.680 80.665 57.910 80.675 ;
        RECT 58.470 80.665 58.700 80.675 ;
        RECT 57.960 80.275 58.420 80.505 ;
        RECT 60.310 78.125 60.680 81.305 ;
        RECT 61.100 78.125 61.470 81.305 ;
        RECT 62.335 80.675 63.380 81.305 ;
        RECT 63.800 80.675 64.170 81.305 ;
        RECT 65.035 80.675 66.080 81.305 ;
        RECT 66.500 80.675 66.870 81.305 ;
        RECT 63.080 80.665 63.310 80.675 ;
        RECT 63.870 80.665 64.100 80.675 ;
        RECT 65.780 80.665 66.010 80.675 ;
        RECT 66.570 80.665 66.800 80.675 ;
        RECT 63.360 80.275 63.820 80.505 ;
        RECT 66.060 80.275 66.520 80.505 ;
        RECT 68.410 78.125 68.780 81.305 ;
        RECT 69.200 78.125 69.570 81.305 ;
        RECT 71.110 78.125 71.480 81.305 ;
        RECT 71.900 78.125 72.270 81.305 ;
        RECT 54.710 76.170 55.910 77.285 ;
        RECT 59.640 76.170 60.010 77.285 ;
        RECT 54.755 76.140 55.870 76.170 ;
        RECT 60.380 74.815 60.610 78.125 ;
        RECT 61.170 74.815 61.400 78.125 ;
        RECT 61.770 76.170 62.140 77.285 ;
        RECT 67.740 76.170 68.110 77.285 ;
        RECT 68.480 74.815 68.710 78.125 ;
        RECT 69.270 74.815 69.500 78.125 ;
        RECT 69.870 76.170 70.240 77.285 ;
        RECT 70.440 76.170 70.810 77.285 ;
        RECT 71.180 74.815 71.410 78.125 ;
        RECT 71.970 74.815 72.200 78.125 ;
        RECT 72.570 76.170 72.940 77.285 ;
        RECT 73.940 76.140 75.055 81.855 ;
        RECT 80.180 77.285 81.295 98.740 ;
        RECT 85.805 97.390 86.035 100.700 ;
        RECT 86.595 97.390 86.825 100.700 ;
        RECT 87.195 98.745 87.565 99.860 ;
        RECT 93.165 98.745 93.535 99.860 ;
        RECT 93.905 97.390 94.135 100.700 ;
        RECT 94.695 97.390 94.925 100.700 ;
        RECT 95.295 98.745 95.665 99.860 ;
        RECT 95.865 98.745 96.235 99.860 ;
        RECT 96.605 97.390 96.835 100.700 ;
        RECT 97.395 97.390 97.625 100.700 ;
        RECT 97.995 98.745 98.365 99.860 ;
        RECT 99.360 98.745 100.535 99.860 ;
        RECT 86.085 97.200 86.545 97.230 ;
        RECT 94.185 97.200 94.645 97.230 ;
        RECT 96.885 97.200 97.345 97.230 ;
        RECT 85.825 96.800 86.825 97.200 ;
        RECT 93.925 96.800 94.925 97.200 ;
        RECT 96.625 96.800 97.625 97.200 ;
        RECT 99.390 95.770 100.505 98.745 ;
        RECT 88.000 95.025 89.000 95.055 ;
        RECT 91.675 95.025 92.675 95.055 ;
        RECT 85.825 94.575 86.825 95.025 ;
        RECT 86.085 94.565 86.545 94.575 ;
        RECT 85.065 91.970 85.435 93.075 ;
        RECT 85.805 89.350 86.035 94.360 ;
        RECT 86.595 89.350 86.825 94.360 ;
        RECT 88.000 93.995 89.925 95.025 ;
        RECT 87.195 93.025 87.565 93.075 ;
        RECT 87.195 91.970 88.300 93.025 ;
        RECT 83.385 85.565 83.845 85.795 ;
        RECT 83.105 85.350 83.335 85.360 ;
        RECT 83.895 85.350 84.125 85.360 ;
        RECT 82.360 84.370 83.405 85.350 ;
        RECT 83.825 84.370 84.195 85.350 ;
        RECT 85.735 84.370 86.105 89.350 ;
        RECT 86.525 84.370 86.895 89.350 ;
        RECT 87.300 87.275 88.300 91.970 ;
        RECT 88.925 88.925 89.925 93.995 ;
        RECT 90.725 93.995 92.675 95.025 ;
        RECT 93.925 94.575 94.925 95.025 ;
        RECT 96.625 94.575 97.625 95.025 ;
        RECT 94.185 94.565 94.645 94.575 ;
        RECT 96.885 94.565 97.345 94.575 ;
        RECT 90.725 89.670 91.725 93.995 ;
        RECT 93.165 93.025 93.535 93.075 ;
        RECT 92.450 91.970 93.535 93.025 ;
        RECT 88.925 87.925 91.755 88.925 ;
        RECT 92.450 87.275 93.450 91.970 ;
        RECT 93.905 89.350 94.135 94.360 ;
        RECT 94.695 89.350 94.925 94.360 ;
        RECT 95.295 91.970 95.665 93.075 ;
        RECT 95.865 91.970 96.235 93.075 ;
        RECT 96.605 89.350 96.835 94.360 ;
        RECT 97.395 89.350 97.625 94.360 ;
        RECT 99.705 93.115 100.155 95.425 ;
        RECT 97.995 91.970 98.365 93.075 ;
        RECT 87.300 86.275 93.450 87.275 ;
        RECT 88.785 85.565 89.245 85.795 ;
        RECT 91.485 85.565 91.945 85.795 ;
        RECT 88.505 85.350 88.735 85.360 ;
        RECT 89.295 85.350 89.525 85.360 ;
        RECT 91.205 85.350 91.435 85.360 ;
        RECT 91.995 85.350 92.225 85.360 ;
        RECT 87.760 84.370 88.805 85.350 ;
        RECT 89.225 84.370 89.595 85.350 ;
        RECT 90.460 84.370 91.505 85.350 ;
        RECT 91.925 84.370 92.295 85.350 ;
        RECT 93.835 84.370 94.205 89.350 ;
        RECT 94.625 84.370 94.995 89.350 ;
        RECT 96.535 84.370 96.905 89.350 ;
        RECT 97.325 84.370 97.695 89.350 ;
        RECT 83.105 84.360 83.335 84.370 ;
        RECT 83.895 84.360 84.125 84.370 ;
        RECT 85.805 84.360 86.035 84.370 ;
        RECT 86.595 84.360 86.825 84.370 ;
        RECT 88.505 84.360 88.735 84.370 ;
        RECT 89.295 84.360 89.525 84.370 ;
        RECT 91.205 84.360 91.435 84.370 ;
        RECT 91.995 84.360 92.225 84.370 ;
        RECT 93.905 84.360 94.135 84.370 ;
        RECT 94.695 84.360 94.925 84.370 ;
        RECT 96.605 84.360 96.835 84.370 ;
        RECT 97.395 84.360 97.625 84.370 ;
        RECT 82.850 83.700 83.885 84.175 ;
        RECT 86.085 83.925 86.545 84.155 ;
        RECT 88.250 83.700 89.285 84.175 ;
        RECT 90.950 83.700 91.985 84.175 ;
        RECT 94.185 83.925 94.645 84.155 ;
        RECT 96.885 83.925 97.345 84.155 ;
        RECT 99.705 82.205 100.155 84.515 ;
        RECT 103.600 83.325 104.600 104.900 ;
        RECT 105.605 99.855 106.720 121.315 ;
        RECT 111.230 119.965 111.460 123.275 ;
        RECT 112.020 119.965 112.250 123.275 ;
        RECT 112.620 121.320 112.990 122.435 ;
        RECT 118.590 121.320 118.960 122.435 ;
        RECT 119.330 119.965 119.560 123.275 ;
        RECT 120.120 119.965 120.350 123.275 ;
        RECT 120.720 121.320 121.090 122.435 ;
        RECT 121.290 121.320 121.660 122.435 ;
        RECT 122.030 119.965 122.260 123.275 ;
        RECT 122.820 119.965 123.050 123.275 ;
        RECT 129.025 123.250 132.075 124.250 ;
        RECT 136.585 123.275 136.955 126.455 ;
        RECT 137.375 123.275 137.745 126.455 ;
        RECT 138.610 125.825 139.655 126.455 ;
        RECT 140.075 125.825 140.445 126.455 ;
        RECT 141.310 125.825 142.355 126.455 ;
        RECT 142.775 125.825 143.145 126.455 ;
        RECT 139.355 125.815 139.585 125.825 ;
        RECT 140.145 125.815 140.375 125.825 ;
        RECT 142.055 125.815 142.285 125.825 ;
        RECT 142.845 125.815 143.075 125.825 ;
        RECT 139.635 125.425 140.095 125.655 ;
        RECT 142.335 125.425 142.795 125.655 ;
        RECT 144.685 123.275 145.055 126.455 ;
        RECT 145.475 123.275 145.845 126.455 ;
        RECT 147.385 123.275 147.755 126.455 ;
        RECT 148.175 123.275 148.545 126.455 ;
        RECT 123.420 121.320 123.790 122.435 ;
        RECT 111.510 119.775 111.970 119.805 ;
        RECT 119.610 119.775 120.070 119.805 ;
        RECT 122.310 119.775 122.770 119.805 ;
        RECT 111.250 119.375 112.250 119.775 ;
        RECT 119.350 119.375 120.350 119.775 ;
        RECT 122.050 119.375 123.050 119.775 ;
        RECT 113.425 117.600 114.425 117.630 ;
        RECT 117.100 117.600 118.100 117.630 ;
        RECT 111.250 117.150 112.250 117.600 ;
        RECT 111.510 117.140 111.970 117.150 ;
        RECT 110.490 114.545 110.860 115.650 ;
        RECT 111.230 111.925 111.460 116.935 ;
        RECT 112.020 111.925 112.250 116.935 ;
        RECT 113.425 116.570 115.350 117.600 ;
        RECT 112.620 115.600 112.990 115.650 ;
        RECT 112.620 114.545 113.725 115.600 ;
        RECT 108.810 108.140 109.270 108.370 ;
        RECT 108.530 107.925 108.760 107.935 ;
        RECT 109.320 107.925 109.550 107.935 ;
        RECT 107.785 106.945 108.830 107.925 ;
        RECT 109.250 106.945 109.620 107.925 ;
        RECT 111.160 106.945 111.530 111.925 ;
        RECT 111.950 106.945 112.320 111.925 ;
        RECT 112.725 109.850 113.725 114.545 ;
        RECT 114.350 111.500 115.350 116.570 ;
        RECT 116.150 116.570 118.100 117.600 ;
        RECT 119.350 117.150 120.350 117.600 ;
        RECT 122.050 117.150 123.050 117.600 ;
        RECT 119.610 117.140 120.070 117.150 ;
        RECT 122.310 117.140 122.770 117.150 ;
        RECT 116.150 112.245 117.150 116.570 ;
        RECT 118.590 115.600 118.960 115.650 ;
        RECT 117.875 114.545 118.960 115.600 ;
        RECT 114.350 110.500 117.180 111.500 ;
        RECT 117.875 109.850 118.875 114.545 ;
        RECT 119.330 111.925 119.560 116.935 ;
        RECT 120.120 111.925 120.350 116.935 ;
        RECT 120.720 114.545 121.090 115.650 ;
        RECT 121.290 114.545 121.660 115.650 ;
        RECT 122.030 111.925 122.260 116.935 ;
        RECT 122.820 111.925 123.050 116.935 ;
        RECT 123.420 114.545 123.790 115.650 ;
        RECT 112.725 108.850 118.875 109.850 ;
        RECT 114.210 108.140 114.670 108.370 ;
        RECT 116.910 108.140 117.370 108.370 ;
        RECT 113.930 107.925 114.160 107.935 ;
        RECT 114.720 107.925 114.950 107.935 ;
        RECT 116.630 107.925 116.860 107.935 ;
        RECT 117.420 107.925 117.650 107.935 ;
        RECT 113.185 106.945 114.230 107.925 ;
        RECT 114.650 106.945 115.020 107.925 ;
        RECT 115.885 106.945 116.930 107.925 ;
        RECT 117.350 106.945 117.720 107.925 ;
        RECT 119.260 106.945 119.630 111.925 ;
        RECT 120.050 106.945 120.420 111.925 ;
        RECT 121.960 106.945 122.330 111.925 ;
        RECT 122.750 106.945 123.120 111.925 ;
        RECT 108.530 106.935 108.760 106.945 ;
        RECT 109.320 106.935 109.550 106.945 ;
        RECT 111.230 106.935 111.460 106.945 ;
        RECT 112.020 106.935 112.250 106.945 ;
        RECT 113.930 106.935 114.160 106.945 ;
        RECT 114.720 106.935 114.950 106.945 ;
        RECT 116.630 106.935 116.860 106.945 ;
        RECT 117.420 106.935 117.650 106.945 ;
        RECT 119.330 106.935 119.560 106.945 ;
        RECT 120.120 106.935 120.350 106.945 ;
        RECT 122.030 106.935 122.260 106.945 ;
        RECT 122.820 106.935 123.050 106.945 ;
        RECT 108.275 106.275 109.310 106.750 ;
        RECT 111.510 106.500 111.970 106.730 ;
        RECT 113.675 106.275 114.710 106.750 ;
        RECT 116.375 106.275 117.410 106.750 ;
        RECT 119.610 106.500 120.070 106.730 ;
        RECT 122.310 106.500 122.770 106.730 ;
        RECT 129.025 105.900 130.025 123.250 ;
        RECT 131.030 122.430 132.145 122.485 ;
        RECT 131.000 121.315 132.175 122.430 ;
        RECT 135.915 121.320 136.285 122.435 ;
        RECT 128.995 104.900 130.055 105.900 ;
        RECT 108.270 104.030 109.310 104.525 ;
        RECT 111.510 104.050 111.970 104.280 ;
        RECT 113.670 104.030 114.710 104.525 ;
        RECT 116.370 104.030 117.410 104.525 ;
        RECT 119.610 104.050 120.070 104.280 ;
        RECT 122.310 104.050 122.770 104.280 ;
        RECT 108.530 103.880 108.760 103.890 ;
        RECT 109.320 103.880 109.550 103.890 ;
        RECT 111.230 103.880 111.460 103.890 ;
        RECT 112.020 103.880 112.250 103.890 ;
        RECT 113.930 103.880 114.160 103.890 ;
        RECT 114.720 103.880 114.950 103.890 ;
        RECT 116.630 103.880 116.860 103.890 ;
        RECT 117.420 103.880 117.650 103.890 ;
        RECT 119.330 103.880 119.560 103.890 ;
        RECT 120.120 103.880 120.350 103.890 ;
        RECT 122.030 103.880 122.260 103.890 ;
        RECT 122.820 103.880 123.050 103.890 ;
        RECT 107.785 103.250 108.830 103.880 ;
        RECT 109.250 103.250 109.620 103.880 ;
        RECT 108.530 103.240 108.760 103.250 ;
        RECT 109.320 103.240 109.550 103.250 ;
        RECT 108.810 102.850 109.270 103.080 ;
        RECT 111.160 100.700 111.530 103.880 ;
        RECT 111.950 100.700 112.320 103.880 ;
        RECT 113.185 103.250 114.230 103.880 ;
        RECT 114.650 103.250 115.020 103.880 ;
        RECT 115.885 103.250 116.930 103.880 ;
        RECT 117.350 103.250 117.720 103.880 ;
        RECT 113.930 103.240 114.160 103.250 ;
        RECT 114.720 103.240 114.950 103.250 ;
        RECT 116.630 103.240 116.860 103.250 ;
        RECT 117.420 103.240 117.650 103.250 ;
        RECT 114.210 102.850 114.670 103.080 ;
        RECT 116.910 102.850 117.370 103.080 ;
        RECT 119.260 100.700 119.630 103.880 ;
        RECT 120.050 100.700 120.420 103.880 ;
        RECT 121.960 100.700 122.330 103.880 ;
        RECT 122.750 100.700 123.120 103.880 ;
        RECT 105.575 98.740 106.750 99.855 ;
        RECT 110.490 98.745 110.860 99.860 ;
        RECT 103.570 82.325 104.630 83.325 ;
        RECT 103.600 82.295 104.600 82.325 ;
        RECT 82.845 81.455 83.885 81.950 ;
        RECT 86.085 81.475 86.545 81.705 ;
        RECT 88.245 81.455 89.285 81.950 ;
        RECT 90.945 81.455 91.985 81.950 ;
        RECT 94.185 81.475 94.645 81.705 ;
        RECT 96.885 81.475 97.345 81.705 ;
        RECT 83.105 81.305 83.335 81.315 ;
        RECT 83.895 81.305 84.125 81.315 ;
        RECT 85.805 81.305 86.035 81.315 ;
        RECT 86.595 81.305 86.825 81.315 ;
        RECT 88.505 81.305 88.735 81.315 ;
        RECT 89.295 81.305 89.525 81.315 ;
        RECT 91.205 81.305 91.435 81.315 ;
        RECT 91.995 81.305 92.225 81.315 ;
        RECT 93.905 81.305 94.135 81.315 ;
        RECT 94.695 81.305 94.925 81.315 ;
        RECT 96.605 81.305 96.835 81.315 ;
        RECT 97.395 81.305 97.625 81.315 ;
        RECT 82.360 80.675 83.405 81.305 ;
        RECT 83.825 80.675 84.195 81.305 ;
        RECT 83.105 80.665 83.335 80.675 ;
        RECT 83.895 80.665 84.125 80.675 ;
        RECT 83.385 80.275 83.845 80.505 ;
        RECT 85.735 78.125 86.105 81.305 ;
        RECT 86.525 78.125 86.895 81.305 ;
        RECT 87.760 80.675 88.805 81.305 ;
        RECT 89.225 80.675 89.595 81.305 ;
        RECT 90.460 80.675 91.505 81.305 ;
        RECT 91.925 80.675 92.295 81.305 ;
        RECT 88.505 80.665 88.735 80.675 ;
        RECT 89.295 80.665 89.525 80.675 ;
        RECT 91.205 80.665 91.435 80.675 ;
        RECT 91.995 80.665 92.225 80.675 ;
        RECT 88.785 80.275 89.245 80.505 ;
        RECT 91.485 80.275 91.945 80.505 ;
        RECT 93.835 78.125 94.205 81.305 ;
        RECT 94.625 78.125 94.995 81.305 ;
        RECT 96.535 78.125 96.905 81.305 ;
        RECT 97.325 78.125 97.695 81.305 ;
        RECT 80.135 76.170 81.335 77.285 ;
        RECT 85.065 76.170 85.435 77.285 ;
        RECT 80.180 76.140 81.295 76.170 ;
        RECT 85.805 74.815 86.035 78.125 ;
        RECT 86.595 74.815 86.825 78.125 ;
        RECT 87.195 76.170 87.565 77.285 ;
        RECT 93.165 76.170 93.535 77.285 ;
        RECT 93.905 74.815 94.135 78.125 ;
        RECT 94.695 74.815 94.925 78.125 ;
        RECT 95.295 76.170 95.665 77.285 ;
        RECT 95.865 76.170 96.235 77.285 ;
        RECT 96.605 74.815 96.835 78.125 ;
        RECT 97.395 74.815 97.625 78.125 ;
        RECT 97.995 76.170 98.365 77.285 ;
        RECT 99.365 76.140 100.480 81.855 ;
        RECT 105.605 77.285 106.720 98.740 ;
        RECT 111.230 97.390 111.460 100.700 ;
        RECT 112.020 97.390 112.250 100.700 ;
        RECT 112.620 98.745 112.990 99.860 ;
        RECT 118.590 98.745 118.960 99.860 ;
        RECT 119.330 97.390 119.560 100.700 ;
        RECT 120.120 97.390 120.350 100.700 ;
        RECT 120.720 98.745 121.090 99.860 ;
        RECT 121.290 98.745 121.660 99.860 ;
        RECT 122.030 97.390 122.260 100.700 ;
        RECT 122.820 97.390 123.050 100.700 ;
        RECT 123.420 98.745 123.790 99.860 ;
        RECT 124.785 98.745 125.960 99.860 ;
        RECT 111.510 97.200 111.970 97.230 ;
        RECT 119.610 97.200 120.070 97.230 ;
        RECT 122.310 97.200 122.770 97.230 ;
        RECT 111.250 96.800 112.250 97.200 ;
        RECT 119.350 96.800 120.350 97.200 ;
        RECT 122.050 96.800 123.050 97.200 ;
        RECT 124.815 95.770 125.930 98.745 ;
        RECT 113.425 95.025 114.425 95.055 ;
        RECT 117.100 95.025 118.100 95.055 ;
        RECT 111.250 94.575 112.250 95.025 ;
        RECT 111.510 94.565 111.970 94.575 ;
        RECT 110.490 91.970 110.860 93.075 ;
        RECT 111.230 89.350 111.460 94.360 ;
        RECT 112.020 89.350 112.250 94.360 ;
        RECT 113.425 93.995 115.350 95.025 ;
        RECT 112.620 93.025 112.990 93.075 ;
        RECT 112.620 91.970 113.725 93.025 ;
        RECT 108.810 85.565 109.270 85.795 ;
        RECT 108.530 85.350 108.760 85.360 ;
        RECT 109.320 85.350 109.550 85.360 ;
        RECT 107.785 84.370 108.830 85.350 ;
        RECT 109.250 84.370 109.620 85.350 ;
        RECT 111.160 84.370 111.530 89.350 ;
        RECT 111.950 84.370 112.320 89.350 ;
        RECT 112.725 87.275 113.725 91.970 ;
        RECT 114.350 88.925 115.350 93.995 ;
        RECT 116.150 93.995 118.100 95.025 ;
        RECT 119.350 94.575 120.350 95.025 ;
        RECT 122.050 94.575 123.050 95.025 ;
        RECT 119.610 94.565 120.070 94.575 ;
        RECT 122.310 94.565 122.770 94.575 ;
        RECT 116.150 89.670 117.150 93.995 ;
        RECT 118.590 93.025 118.960 93.075 ;
        RECT 117.875 91.970 118.960 93.025 ;
        RECT 114.350 87.925 117.180 88.925 ;
        RECT 117.875 87.275 118.875 91.970 ;
        RECT 119.330 89.350 119.560 94.360 ;
        RECT 120.120 89.350 120.350 94.360 ;
        RECT 120.720 91.970 121.090 93.075 ;
        RECT 121.290 91.970 121.660 93.075 ;
        RECT 122.030 89.350 122.260 94.360 ;
        RECT 122.820 89.350 123.050 94.360 ;
        RECT 125.130 93.115 125.580 95.425 ;
        RECT 123.420 91.970 123.790 93.075 ;
        RECT 112.725 86.275 118.875 87.275 ;
        RECT 114.210 85.565 114.670 85.795 ;
        RECT 116.910 85.565 117.370 85.795 ;
        RECT 113.930 85.350 114.160 85.360 ;
        RECT 114.720 85.350 114.950 85.360 ;
        RECT 116.630 85.350 116.860 85.360 ;
        RECT 117.420 85.350 117.650 85.360 ;
        RECT 113.185 84.370 114.230 85.350 ;
        RECT 114.650 84.370 115.020 85.350 ;
        RECT 115.885 84.370 116.930 85.350 ;
        RECT 117.350 84.370 117.720 85.350 ;
        RECT 119.260 84.370 119.630 89.350 ;
        RECT 120.050 84.370 120.420 89.350 ;
        RECT 121.960 84.370 122.330 89.350 ;
        RECT 122.750 84.370 123.120 89.350 ;
        RECT 108.530 84.360 108.760 84.370 ;
        RECT 109.320 84.360 109.550 84.370 ;
        RECT 111.230 84.360 111.460 84.370 ;
        RECT 112.020 84.360 112.250 84.370 ;
        RECT 113.930 84.360 114.160 84.370 ;
        RECT 114.720 84.360 114.950 84.370 ;
        RECT 116.630 84.360 116.860 84.370 ;
        RECT 117.420 84.360 117.650 84.370 ;
        RECT 119.330 84.360 119.560 84.370 ;
        RECT 120.120 84.360 120.350 84.370 ;
        RECT 122.030 84.360 122.260 84.370 ;
        RECT 122.820 84.360 123.050 84.370 ;
        RECT 108.275 83.700 109.310 84.175 ;
        RECT 111.510 83.925 111.970 84.155 ;
        RECT 113.675 83.700 114.710 84.175 ;
        RECT 116.375 83.700 117.410 84.175 ;
        RECT 119.610 83.925 120.070 84.155 ;
        RECT 122.310 83.925 122.770 84.155 ;
        RECT 125.130 82.205 125.580 84.515 ;
        RECT 129.025 83.325 130.025 104.900 ;
        RECT 131.030 99.855 132.145 121.315 ;
        RECT 136.655 119.965 136.885 123.275 ;
        RECT 137.445 119.965 137.675 123.275 ;
        RECT 138.045 121.320 138.415 122.435 ;
        RECT 144.015 121.320 144.385 122.435 ;
        RECT 144.755 119.965 144.985 123.275 ;
        RECT 145.545 119.965 145.775 123.275 ;
        RECT 146.145 121.320 146.515 122.435 ;
        RECT 146.715 121.320 147.085 122.435 ;
        RECT 147.455 119.965 147.685 123.275 ;
        RECT 148.245 119.965 148.475 123.275 ;
        RECT 148.845 121.320 149.215 122.435 ;
        RECT 136.935 119.775 137.395 119.805 ;
        RECT 145.035 119.775 145.495 119.805 ;
        RECT 147.735 119.775 148.195 119.805 ;
        RECT 136.675 119.375 137.675 119.775 ;
        RECT 144.775 119.375 145.775 119.775 ;
        RECT 147.475 119.375 148.475 119.775 ;
        RECT 138.850 117.600 139.850 117.630 ;
        RECT 142.525 117.600 143.525 117.630 ;
        RECT 136.675 117.150 137.675 117.600 ;
        RECT 136.935 117.140 137.395 117.150 ;
        RECT 135.915 114.545 136.285 115.650 ;
        RECT 136.655 111.925 136.885 116.935 ;
        RECT 137.445 111.925 137.675 116.935 ;
        RECT 138.850 116.570 140.775 117.600 ;
        RECT 138.045 115.600 138.415 115.650 ;
        RECT 138.045 114.545 139.150 115.600 ;
        RECT 134.235 108.140 134.695 108.370 ;
        RECT 133.955 107.925 134.185 107.935 ;
        RECT 134.745 107.925 134.975 107.935 ;
        RECT 133.210 106.945 134.255 107.925 ;
        RECT 134.675 106.945 135.045 107.925 ;
        RECT 136.585 106.945 136.955 111.925 ;
        RECT 137.375 106.945 137.745 111.925 ;
        RECT 138.150 109.850 139.150 114.545 ;
        RECT 139.775 111.500 140.775 116.570 ;
        RECT 141.575 116.570 143.525 117.600 ;
        RECT 144.775 117.150 145.775 117.600 ;
        RECT 147.475 117.150 148.475 117.600 ;
        RECT 145.035 117.140 145.495 117.150 ;
        RECT 147.735 117.140 148.195 117.150 ;
        RECT 141.575 112.245 142.575 116.570 ;
        RECT 144.015 115.600 144.385 115.650 ;
        RECT 143.300 114.545 144.385 115.600 ;
        RECT 139.775 110.500 142.605 111.500 ;
        RECT 143.300 109.850 144.300 114.545 ;
        RECT 144.755 111.925 144.985 116.935 ;
        RECT 145.545 111.925 145.775 116.935 ;
        RECT 146.145 114.545 146.515 115.650 ;
        RECT 146.715 114.545 147.085 115.650 ;
        RECT 147.455 111.925 147.685 116.935 ;
        RECT 148.245 111.925 148.475 116.935 ;
        RECT 148.845 114.545 149.215 115.650 ;
        RECT 138.150 108.850 144.300 109.850 ;
        RECT 139.635 108.140 140.095 108.370 ;
        RECT 142.335 108.140 142.795 108.370 ;
        RECT 139.355 107.925 139.585 107.935 ;
        RECT 140.145 107.925 140.375 107.935 ;
        RECT 142.055 107.925 142.285 107.935 ;
        RECT 142.845 107.925 143.075 107.935 ;
        RECT 138.610 106.945 139.655 107.925 ;
        RECT 140.075 106.945 140.445 107.925 ;
        RECT 141.310 106.945 142.355 107.925 ;
        RECT 142.775 106.945 143.145 107.925 ;
        RECT 144.685 106.945 145.055 111.925 ;
        RECT 145.475 106.945 145.845 111.925 ;
        RECT 147.385 106.945 147.755 111.925 ;
        RECT 148.175 106.945 148.545 111.925 ;
        RECT 133.955 106.935 134.185 106.945 ;
        RECT 134.745 106.935 134.975 106.945 ;
        RECT 136.655 106.935 136.885 106.945 ;
        RECT 137.445 106.935 137.675 106.945 ;
        RECT 139.355 106.935 139.585 106.945 ;
        RECT 140.145 106.935 140.375 106.945 ;
        RECT 142.055 106.935 142.285 106.945 ;
        RECT 142.845 106.935 143.075 106.945 ;
        RECT 144.755 106.935 144.985 106.945 ;
        RECT 145.545 106.935 145.775 106.945 ;
        RECT 147.455 106.935 147.685 106.945 ;
        RECT 148.245 106.935 148.475 106.945 ;
        RECT 133.700 106.275 134.735 106.750 ;
        RECT 136.935 106.500 137.395 106.730 ;
        RECT 139.100 106.275 140.135 106.750 ;
        RECT 141.800 106.275 142.835 106.750 ;
        RECT 145.035 106.500 145.495 106.730 ;
        RECT 147.735 106.500 148.195 106.730 ;
        RECT 133.695 104.030 134.735 104.525 ;
        RECT 136.935 104.050 137.395 104.280 ;
        RECT 139.095 104.030 140.135 104.525 ;
        RECT 141.795 104.030 142.835 104.525 ;
        RECT 145.035 104.050 145.495 104.280 ;
        RECT 147.735 104.050 148.195 104.280 ;
        RECT 133.955 103.880 134.185 103.890 ;
        RECT 134.745 103.880 134.975 103.890 ;
        RECT 136.655 103.880 136.885 103.890 ;
        RECT 137.445 103.880 137.675 103.890 ;
        RECT 139.355 103.880 139.585 103.890 ;
        RECT 140.145 103.880 140.375 103.890 ;
        RECT 142.055 103.880 142.285 103.890 ;
        RECT 142.845 103.880 143.075 103.890 ;
        RECT 144.755 103.880 144.985 103.890 ;
        RECT 145.545 103.880 145.775 103.890 ;
        RECT 147.455 103.880 147.685 103.890 ;
        RECT 148.245 103.880 148.475 103.890 ;
        RECT 133.210 103.250 134.255 103.880 ;
        RECT 134.675 103.250 135.045 103.880 ;
        RECT 133.955 103.240 134.185 103.250 ;
        RECT 134.745 103.240 134.975 103.250 ;
        RECT 134.235 102.850 134.695 103.080 ;
        RECT 136.585 100.700 136.955 103.880 ;
        RECT 137.375 100.700 137.745 103.880 ;
        RECT 138.610 103.250 139.655 103.880 ;
        RECT 140.075 103.250 140.445 103.880 ;
        RECT 141.310 103.250 142.355 103.880 ;
        RECT 142.775 103.250 143.145 103.880 ;
        RECT 139.355 103.240 139.585 103.250 ;
        RECT 140.145 103.240 140.375 103.250 ;
        RECT 142.055 103.240 142.285 103.250 ;
        RECT 142.845 103.240 143.075 103.250 ;
        RECT 139.635 102.850 140.095 103.080 ;
        RECT 142.335 102.850 142.795 103.080 ;
        RECT 144.685 100.700 145.055 103.880 ;
        RECT 145.475 100.700 145.845 103.880 ;
        RECT 147.385 100.700 147.755 103.880 ;
        RECT 148.175 100.700 148.545 103.880 ;
        RECT 131.000 98.740 132.175 99.855 ;
        RECT 135.915 98.745 136.285 99.860 ;
        RECT 128.995 82.325 130.055 83.325 ;
        RECT 129.025 82.295 130.025 82.325 ;
        RECT 108.270 81.455 109.310 81.950 ;
        RECT 111.510 81.475 111.970 81.705 ;
        RECT 113.670 81.455 114.710 81.950 ;
        RECT 116.370 81.455 117.410 81.950 ;
        RECT 119.610 81.475 120.070 81.705 ;
        RECT 122.310 81.475 122.770 81.705 ;
        RECT 108.530 81.305 108.760 81.315 ;
        RECT 109.320 81.305 109.550 81.315 ;
        RECT 111.230 81.305 111.460 81.315 ;
        RECT 112.020 81.305 112.250 81.315 ;
        RECT 113.930 81.305 114.160 81.315 ;
        RECT 114.720 81.305 114.950 81.315 ;
        RECT 116.630 81.305 116.860 81.315 ;
        RECT 117.420 81.305 117.650 81.315 ;
        RECT 119.330 81.305 119.560 81.315 ;
        RECT 120.120 81.305 120.350 81.315 ;
        RECT 122.030 81.305 122.260 81.315 ;
        RECT 122.820 81.305 123.050 81.315 ;
        RECT 107.785 80.675 108.830 81.305 ;
        RECT 109.250 80.675 109.620 81.305 ;
        RECT 108.530 80.665 108.760 80.675 ;
        RECT 109.320 80.665 109.550 80.675 ;
        RECT 108.810 80.275 109.270 80.505 ;
        RECT 111.160 78.125 111.530 81.305 ;
        RECT 111.950 78.125 112.320 81.305 ;
        RECT 113.185 80.675 114.230 81.305 ;
        RECT 114.650 80.675 115.020 81.305 ;
        RECT 115.885 80.675 116.930 81.305 ;
        RECT 117.350 80.675 117.720 81.305 ;
        RECT 113.930 80.665 114.160 80.675 ;
        RECT 114.720 80.665 114.950 80.675 ;
        RECT 116.630 80.665 116.860 80.675 ;
        RECT 117.420 80.665 117.650 80.675 ;
        RECT 114.210 80.275 114.670 80.505 ;
        RECT 116.910 80.275 117.370 80.505 ;
        RECT 119.260 78.125 119.630 81.305 ;
        RECT 120.050 78.125 120.420 81.305 ;
        RECT 121.960 78.125 122.330 81.305 ;
        RECT 122.750 78.125 123.120 81.305 ;
        RECT 105.560 76.170 106.760 77.285 ;
        RECT 110.490 76.170 110.860 77.285 ;
        RECT 105.605 76.140 106.720 76.170 ;
        RECT 111.230 74.815 111.460 78.125 ;
        RECT 112.020 74.815 112.250 78.125 ;
        RECT 112.620 76.170 112.990 77.285 ;
        RECT 118.590 76.170 118.960 77.285 ;
        RECT 119.330 74.815 119.560 78.125 ;
        RECT 120.120 74.815 120.350 78.125 ;
        RECT 120.720 76.170 121.090 77.285 ;
        RECT 121.290 76.170 121.660 77.285 ;
        RECT 122.030 74.815 122.260 78.125 ;
        RECT 122.820 74.815 123.050 78.125 ;
        RECT 123.420 76.170 123.790 77.285 ;
        RECT 124.790 76.140 125.905 81.855 ;
        RECT 131.030 77.285 132.145 98.740 ;
        RECT 136.655 97.390 136.885 100.700 ;
        RECT 137.445 97.390 137.675 100.700 ;
        RECT 138.045 98.745 138.415 99.860 ;
        RECT 144.015 98.745 144.385 99.860 ;
        RECT 144.755 97.390 144.985 100.700 ;
        RECT 145.545 97.390 145.775 100.700 ;
        RECT 146.145 98.745 146.515 99.860 ;
        RECT 146.715 98.745 147.085 99.860 ;
        RECT 147.455 97.390 147.685 100.700 ;
        RECT 148.245 97.390 148.475 100.700 ;
        RECT 148.845 98.745 149.215 99.860 ;
        RECT 150.210 98.745 151.385 99.860 ;
        RECT 136.935 97.200 137.395 97.230 ;
        RECT 145.035 97.200 145.495 97.230 ;
        RECT 147.735 97.200 148.195 97.230 ;
        RECT 136.675 96.800 137.675 97.200 ;
        RECT 144.775 96.800 145.775 97.200 ;
        RECT 147.475 96.800 148.475 97.200 ;
        RECT 150.240 95.770 151.355 98.745 ;
        RECT 138.850 95.025 139.850 95.055 ;
        RECT 142.525 95.025 143.525 95.055 ;
        RECT 136.675 94.575 137.675 95.025 ;
        RECT 136.935 94.565 137.395 94.575 ;
        RECT 135.915 91.970 136.285 93.075 ;
        RECT 136.655 89.350 136.885 94.360 ;
        RECT 137.445 89.350 137.675 94.360 ;
        RECT 138.850 93.995 140.775 95.025 ;
        RECT 138.045 93.025 138.415 93.075 ;
        RECT 138.045 91.970 139.150 93.025 ;
        RECT 134.235 85.565 134.695 85.795 ;
        RECT 133.955 85.350 134.185 85.360 ;
        RECT 134.745 85.350 134.975 85.360 ;
        RECT 133.210 84.370 134.255 85.350 ;
        RECT 134.675 84.370 135.045 85.350 ;
        RECT 136.585 84.370 136.955 89.350 ;
        RECT 137.375 84.370 137.745 89.350 ;
        RECT 138.150 87.275 139.150 91.970 ;
        RECT 139.775 88.925 140.775 93.995 ;
        RECT 141.575 93.995 143.525 95.025 ;
        RECT 144.775 94.575 145.775 95.025 ;
        RECT 147.475 94.575 148.475 95.025 ;
        RECT 145.035 94.565 145.495 94.575 ;
        RECT 147.735 94.565 148.195 94.575 ;
        RECT 141.575 89.670 142.575 93.995 ;
        RECT 144.015 93.025 144.385 93.075 ;
        RECT 143.300 91.970 144.385 93.025 ;
        RECT 139.775 87.925 142.605 88.925 ;
        RECT 143.300 87.275 144.300 91.970 ;
        RECT 144.755 89.350 144.985 94.360 ;
        RECT 145.545 89.350 145.775 94.360 ;
        RECT 146.145 91.970 146.515 93.075 ;
        RECT 146.715 91.970 147.085 93.075 ;
        RECT 147.455 89.350 147.685 94.360 ;
        RECT 148.245 89.350 148.475 94.360 ;
        RECT 150.555 93.115 151.005 95.425 ;
        RECT 148.845 91.970 149.215 93.075 ;
        RECT 138.150 86.275 144.300 87.275 ;
        RECT 139.635 85.565 140.095 85.795 ;
        RECT 142.335 85.565 142.795 85.795 ;
        RECT 139.355 85.350 139.585 85.360 ;
        RECT 140.145 85.350 140.375 85.360 ;
        RECT 142.055 85.350 142.285 85.360 ;
        RECT 142.845 85.350 143.075 85.360 ;
        RECT 138.610 84.370 139.655 85.350 ;
        RECT 140.075 84.370 140.445 85.350 ;
        RECT 141.310 84.370 142.355 85.350 ;
        RECT 142.775 84.370 143.145 85.350 ;
        RECT 144.685 84.370 145.055 89.350 ;
        RECT 145.475 84.370 145.845 89.350 ;
        RECT 147.385 84.370 147.755 89.350 ;
        RECT 148.175 84.370 148.545 89.350 ;
        RECT 133.955 84.360 134.185 84.370 ;
        RECT 134.745 84.360 134.975 84.370 ;
        RECT 136.655 84.360 136.885 84.370 ;
        RECT 137.445 84.360 137.675 84.370 ;
        RECT 139.355 84.360 139.585 84.370 ;
        RECT 140.145 84.360 140.375 84.370 ;
        RECT 142.055 84.360 142.285 84.370 ;
        RECT 142.845 84.360 143.075 84.370 ;
        RECT 144.755 84.360 144.985 84.370 ;
        RECT 145.545 84.360 145.775 84.370 ;
        RECT 147.455 84.360 147.685 84.370 ;
        RECT 148.245 84.360 148.475 84.370 ;
        RECT 133.700 83.700 134.735 84.175 ;
        RECT 136.935 83.925 137.395 84.155 ;
        RECT 139.100 83.700 140.135 84.175 ;
        RECT 141.800 83.700 142.835 84.175 ;
        RECT 145.035 83.925 145.495 84.155 ;
        RECT 147.735 83.925 148.195 84.155 ;
        RECT 150.555 82.205 151.005 84.515 ;
        RECT 133.695 81.455 134.735 81.950 ;
        RECT 136.935 81.475 137.395 81.705 ;
        RECT 139.095 81.455 140.135 81.950 ;
        RECT 141.795 81.455 142.835 81.950 ;
        RECT 145.035 81.475 145.495 81.705 ;
        RECT 147.735 81.475 148.195 81.705 ;
        RECT 133.955 81.305 134.185 81.315 ;
        RECT 134.745 81.305 134.975 81.315 ;
        RECT 136.655 81.305 136.885 81.315 ;
        RECT 137.445 81.305 137.675 81.315 ;
        RECT 139.355 81.305 139.585 81.315 ;
        RECT 140.145 81.305 140.375 81.315 ;
        RECT 142.055 81.305 142.285 81.315 ;
        RECT 142.845 81.305 143.075 81.315 ;
        RECT 144.755 81.305 144.985 81.315 ;
        RECT 145.545 81.305 145.775 81.315 ;
        RECT 147.455 81.305 147.685 81.315 ;
        RECT 148.245 81.305 148.475 81.315 ;
        RECT 133.210 80.675 134.255 81.305 ;
        RECT 134.675 80.675 135.045 81.305 ;
        RECT 133.955 80.665 134.185 80.675 ;
        RECT 134.745 80.665 134.975 80.675 ;
        RECT 134.235 80.275 134.695 80.505 ;
        RECT 136.585 78.125 136.955 81.305 ;
        RECT 137.375 78.125 137.745 81.305 ;
        RECT 138.610 80.675 139.655 81.305 ;
        RECT 140.075 80.675 140.445 81.305 ;
        RECT 141.310 80.675 142.355 81.305 ;
        RECT 142.775 80.675 143.145 81.305 ;
        RECT 139.355 80.665 139.585 80.675 ;
        RECT 140.145 80.665 140.375 80.675 ;
        RECT 142.055 80.665 142.285 80.675 ;
        RECT 142.845 80.665 143.075 80.675 ;
        RECT 139.635 80.275 140.095 80.505 ;
        RECT 142.335 80.275 142.795 80.505 ;
        RECT 144.685 78.125 145.055 81.305 ;
        RECT 145.475 78.125 145.845 81.305 ;
        RECT 147.385 78.125 147.755 81.305 ;
        RECT 148.175 78.125 148.545 81.305 ;
        RECT 130.985 76.170 132.185 77.285 ;
        RECT 135.915 76.170 136.285 77.285 ;
        RECT 131.030 76.140 132.145 76.170 ;
        RECT 136.655 74.815 136.885 78.125 ;
        RECT 137.445 74.815 137.675 78.125 ;
        RECT 138.045 76.170 138.415 77.285 ;
        RECT 144.015 76.170 144.385 77.285 ;
        RECT 144.755 74.815 144.985 78.125 ;
        RECT 145.545 74.815 145.775 78.125 ;
        RECT 146.145 76.170 146.515 77.285 ;
        RECT 146.715 76.170 147.085 77.285 ;
        RECT 147.455 74.815 147.685 78.125 ;
        RECT 148.245 74.815 148.475 78.125 ;
        RECT 148.845 76.170 149.215 77.285 ;
        RECT 150.215 76.140 151.330 81.855 ;
        RECT 9.810 74.625 10.270 74.655 ;
        RECT 17.910 74.625 18.370 74.655 ;
        RECT 20.610 74.625 21.070 74.655 ;
        RECT 35.235 74.625 35.695 74.655 ;
        RECT 43.335 74.625 43.795 74.655 ;
        RECT 46.035 74.625 46.495 74.655 ;
        RECT 60.660 74.625 61.120 74.655 ;
        RECT 68.760 74.625 69.220 74.655 ;
        RECT 71.460 74.625 71.920 74.655 ;
        RECT 86.085 74.625 86.545 74.655 ;
        RECT 94.185 74.625 94.645 74.655 ;
        RECT 96.885 74.625 97.345 74.655 ;
        RECT 111.510 74.625 111.970 74.655 ;
        RECT 119.610 74.625 120.070 74.655 ;
        RECT 122.310 74.625 122.770 74.655 ;
        RECT 136.935 74.625 137.395 74.655 ;
        RECT 145.035 74.625 145.495 74.655 ;
        RECT 147.735 74.625 148.195 74.655 ;
        RECT 9.550 74.225 10.550 74.625 ;
        RECT 17.650 74.225 18.650 74.625 ;
        RECT 20.350 74.225 21.350 74.625 ;
        RECT 34.975 74.225 35.975 74.625 ;
        RECT 43.075 74.225 44.075 74.625 ;
        RECT 45.775 74.225 46.775 74.625 ;
        RECT 60.400 74.225 61.400 74.625 ;
        RECT 68.500 74.225 69.500 74.625 ;
        RECT 71.200 74.225 72.200 74.625 ;
        RECT 85.825 74.225 86.825 74.625 ;
        RECT 93.925 74.225 94.925 74.625 ;
        RECT 96.625 74.225 97.625 74.625 ;
        RECT 111.250 74.225 112.250 74.625 ;
        RECT 119.350 74.225 120.350 74.625 ;
        RECT 122.050 74.225 123.050 74.625 ;
        RECT 136.675 74.225 137.675 74.625 ;
        RECT 144.775 74.225 145.775 74.625 ;
        RECT 147.475 74.225 148.475 74.625 ;
        RECT 7.500 69.550 153.425 70.550 ;
        RECT 11.725 68.175 12.725 68.205 ;
        RECT 15.400 68.175 16.400 68.205 ;
        RECT 37.150 68.175 38.150 68.205 ;
        RECT 40.825 68.175 41.825 68.205 ;
        RECT 9.550 67.725 10.550 68.175 ;
        RECT 9.810 67.715 10.270 67.725 ;
        RECT 8.790 65.120 9.160 66.225 ;
        RECT 9.530 62.500 9.760 67.510 ;
        RECT 10.320 62.500 10.550 67.510 ;
        RECT 11.725 67.145 13.650 68.175 ;
        RECT 10.920 66.175 11.290 66.225 ;
        RECT 10.920 65.120 12.025 66.175 ;
        RECT 7.110 58.715 7.570 58.945 ;
        RECT 6.830 58.500 7.060 58.510 ;
        RECT 7.620 58.500 7.850 58.510 ;
        RECT 6.085 57.520 7.130 58.500 ;
        RECT 7.550 57.520 7.920 58.500 ;
        RECT 9.460 57.520 9.830 62.500 ;
        RECT 10.250 57.520 10.620 62.500 ;
        RECT 11.025 60.425 12.025 65.120 ;
        RECT 12.650 62.075 13.650 67.145 ;
        RECT 14.450 67.145 16.400 68.175 ;
        RECT 17.650 67.725 18.650 68.175 ;
        RECT 20.350 67.725 21.350 68.175 ;
        RECT 27.270 67.975 28.270 68.125 ;
        RECT 17.910 67.715 18.370 67.725 ;
        RECT 20.610 67.715 21.070 67.725 ;
        RECT 23.805 67.715 24.265 67.945 ;
        RECT 26.505 67.715 26.965 67.945 ;
        RECT 27.120 67.525 28.270 67.975 ;
        RECT 29.205 67.715 29.665 67.945 ;
        RECT 34.975 67.725 35.975 68.175 ;
        RECT 35.235 67.715 35.695 67.725 ;
        RECT 14.450 62.820 15.450 67.145 ;
        RECT 16.890 66.175 17.260 66.225 ;
        RECT 16.175 65.120 17.260 66.175 ;
        RECT 12.650 61.075 15.480 62.075 ;
        RECT 16.175 60.425 17.175 65.120 ;
        RECT 17.630 62.500 17.860 67.510 ;
        RECT 18.420 62.500 18.650 67.510 ;
        RECT 19.020 65.120 19.390 66.225 ;
        RECT 19.590 65.120 19.960 66.225 ;
        RECT 20.330 62.500 20.560 67.510 ;
        RECT 21.120 62.500 21.350 67.510 ;
        RECT 23.525 66.510 23.755 67.510 ;
        RECT 24.295 66.495 26.475 67.525 ;
        RECT 26.970 67.500 28.270 67.525 ;
        RECT 28.925 67.500 29.155 67.510 ;
        RECT 29.715 67.500 29.945 67.510 ;
        RECT 26.970 66.975 29.225 67.500 ;
        RECT 26.970 66.570 27.890 66.975 ;
        RECT 27.015 66.510 27.245 66.570 ;
        RECT 28.180 66.520 29.225 66.975 ;
        RECT 29.645 66.520 30.015 67.500 ;
        RECT 28.925 66.510 29.155 66.520 ;
        RECT 29.715 66.510 29.945 66.520 ;
        RECT 21.720 65.120 22.090 66.225 ;
        RECT 23.520 63.625 24.520 66.355 ;
        RECT 26.245 63.625 27.245 66.325 ;
        RECT 28.670 65.850 29.705 66.325 ;
        RECT 34.215 65.120 34.585 66.225 ;
        RECT 28.665 63.605 29.705 64.100 ;
        RECT 23.205 62.800 23.850 63.480 ;
        RECT 24.245 62.800 26.525 63.480 ;
        RECT 27.015 63.405 27.245 63.465 ;
        RECT 28.925 63.455 29.155 63.465 ;
        RECT 29.715 63.455 29.945 63.465 ;
        RECT 26.970 63.250 27.890 63.405 ;
        RECT 28.180 63.250 29.225 63.455 ;
        RECT 26.970 62.825 29.225 63.250 ;
        RECT 29.645 62.825 30.015 63.455 ;
        RECT 27.015 62.815 28.270 62.825 ;
        RECT 28.925 62.815 29.155 62.825 ;
        RECT 29.715 62.815 29.945 62.825 ;
        RECT 27.020 62.800 28.270 62.815 ;
        RECT 11.025 59.425 17.175 60.425 ;
        RECT 12.510 58.715 12.970 58.945 ;
        RECT 15.210 58.715 15.670 58.945 ;
        RECT 12.230 58.500 12.460 58.510 ;
        RECT 13.020 58.500 13.250 58.510 ;
        RECT 14.930 58.500 15.160 58.510 ;
        RECT 15.720 58.500 15.950 58.510 ;
        RECT 11.485 57.520 12.530 58.500 ;
        RECT 12.950 57.520 13.320 58.500 ;
        RECT 14.185 57.520 15.230 58.500 ;
        RECT 15.650 57.520 16.020 58.500 ;
        RECT 17.560 57.520 17.930 62.500 ;
        RECT 18.350 57.520 18.720 62.500 ;
        RECT 20.260 57.520 20.630 62.500 ;
        RECT 21.050 57.520 21.420 62.500 ;
        RECT 23.805 62.425 24.265 62.655 ;
        RECT 26.505 62.425 26.965 62.655 ;
        RECT 27.115 62.250 28.270 62.800 ;
        RECT 29.205 62.425 29.665 62.655 ;
        RECT 34.955 62.500 35.185 67.510 ;
        RECT 35.745 62.500 35.975 67.510 ;
        RECT 37.150 67.145 39.075 68.175 ;
        RECT 36.345 66.175 36.715 66.225 ;
        RECT 36.345 65.120 37.450 66.175 ;
        RECT 27.115 62.200 28.175 62.250 ;
        RECT 6.830 57.510 7.060 57.520 ;
        RECT 7.620 57.510 7.850 57.520 ;
        RECT 9.530 57.510 9.760 57.520 ;
        RECT 10.320 57.510 10.550 57.520 ;
        RECT 12.230 57.510 12.460 57.520 ;
        RECT 13.020 57.510 13.250 57.520 ;
        RECT 14.930 57.510 15.160 57.520 ;
        RECT 15.720 57.510 15.950 57.520 ;
        RECT 17.630 57.510 17.860 57.520 ;
        RECT 18.420 57.510 18.650 57.520 ;
        RECT 20.330 57.510 20.560 57.520 ;
        RECT 21.120 57.510 21.350 57.520 ;
        RECT 6.575 56.850 7.610 57.325 ;
        RECT 9.810 57.075 10.270 57.305 ;
        RECT 11.975 56.850 13.010 57.325 ;
        RECT 14.675 56.850 15.710 57.325 ;
        RECT 17.910 57.075 18.370 57.305 ;
        RECT 20.610 57.075 21.070 57.305 ;
        RECT 3.950 56.475 4.950 56.530 ;
        RECT 24.820 56.510 25.925 61.180 ;
        RECT 32.535 58.715 32.995 58.945 ;
        RECT 32.255 58.500 32.485 58.510 ;
        RECT 33.045 58.500 33.275 58.510 ;
        RECT 31.510 57.520 32.555 58.500 ;
        RECT 32.975 57.520 33.345 58.500 ;
        RECT 34.885 57.520 35.255 62.500 ;
        RECT 35.675 57.520 36.045 62.500 ;
        RECT 36.450 60.425 37.450 65.120 ;
        RECT 38.075 62.075 39.075 67.145 ;
        RECT 39.875 67.145 41.825 68.175 ;
        RECT 43.075 67.725 44.075 68.175 ;
        RECT 45.775 67.725 46.775 68.175 ;
        RECT 43.335 67.715 43.795 67.725 ;
        RECT 46.035 67.715 46.495 67.725 ;
        RECT 39.875 62.820 40.875 67.145 ;
        RECT 42.315 66.175 42.685 66.225 ;
        RECT 41.600 65.120 42.685 66.175 ;
        RECT 38.075 61.075 40.905 62.075 ;
        RECT 41.600 60.425 42.600 65.120 ;
        RECT 43.055 62.500 43.285 67.510 ;
        RECT 43.845 62.500 44.075 67.510 ;
        RECT 44.445 65.120 44.815 66.225 ;
        RECT 45.015 65.120 45.385 66.225 ;
        RECT 45.755 62.500 45.985 67.510 ;
        RECT 46.545 62.500 46.775 67.510 ;
        RECT 47.145 65.120 47.515 66.225 ;
        RECT 36.450 59.425 42.600 60.425 ;
        RECT 37.935 58.715 38.395 58.945 ;
        RECT 40.635 58.715 41.095 58.945 ;
        RECT 37.655 58.500 37.885 58.510 ;
        RECT 38.445 58.500 38.675 58.510 ;
        RECT 40.355 58.500 40.585 58.510 ;
        RECT 41.145 58.500 41.375 58.510 ;
        RECT 36.910 57.520 37.955 58.500 ;
        RECT 38.375 57.520 38.745 58.500 ;
        RECT 39.610 57.520 40.655 58.500 ;
        RECT 41.075 57.520 41.445 58.500 ;
        RECT 42.985 57.520 43.355 62.500 ;
        RECT 43.775 57.520 44.145 62.500 ;
        RECT 45.685 57.520 46.055 62.500 ;
        RECT 46.475 57.520 46.845 62.500 ;
        RECT 32.255 57.510 32.485 57.520 ;
        RECT 33.045 57.510 33.275 57.520 ;
        RECT 34.955 57.510 35.185 57.520 ;
        RECT 35.745 57.510 35.975 57.520 ;
        RECT 37.655 57.510 37.885 57.520 ;
        RECT 38.445 57.510 38.675 57.520 ;
        RECT 40.355 57.510 40.585 57.520 ;
        RECT 41.145 57.510 41.375 57.520 ;
        RECT 43.055 57.510 43.285 57.520 ;
        RECT 43.845 57.510 44.075 57.520 ;
        RECT 45.755 57.510 45.985 57.520 ;
        RECT 46.545 57.510 46.775 57.520 ;
        RECT 32.000 56.850 33.035 57.325 ;
        RECT 35.235 57.075 35.695 57.305 ;
        RECT 37.400 56.850 38.435 57.325 ;
        RECT 40.100 56.850 41.135 57.325 ;
        RECT 43.335 57.075 43.795 57.305 ;
        RECT 46.035 57.075 46.495 57.305 ;
        RECT 29.375 56.510 30.375 56.530 ;
        RECT 3.920 55.475 4.980 56.475 ;
        RECT 3.950 52.250 4.950 55.475 ;
        RECT 24.820 55.405 30.430 56.510 ;
        RECT 50.725 56.475 51.725 69.550 ;
        RECT 62.575 68.175 63.575 68.205 ;
        RECT 66.250 68.175 67.250 68.205 ;
        RECT 88.000 68.175 89.000 68.205 ;
        RECT 91.675 68.175 92.675 68.205 ;
        RECT 60.400 67.725 61.400 68.175 ;
        RECT 60.660 67.715 61.120 67.725 ;
        RECT 59.640 65.120 60.010 66.225 ;
        RECT 60.380 62.500 60.610 67.510 ;
        RECT 61.170 62.500 61.400 67.510 ;
        RECT 62.575 67.145 64.500 68.175 ;
        RECT 61.770 66.175 62.140 66.225 ;
        RECT 61.770 65.120 62.875 66.175 ;
        RECT 57.960 58.715 58.420 58.945 ;
        RECT 57.680 58.500 57.910 58.510 ;
        RECT 58.470 58.500 58.700 58.510 ;
        RECT 56.935 57.520 57.980 58.500 ;
        RECT 58.400 57.520 58.770 58.500 ;
        RECT 60.310 57.520 60.680 62.500 ;
        RECT 61.100 57.520 61.470 62.500 ;
        RECT 61.875 60.425 62.875 65.120 ;
        RECT 63.500 62.075 64.500 67.145 ;
        RECT 65.300 67.145 67.250 68.175 ;
        RECT 68.500 67.725 69.500 68.175 ;
        RECT 71.200 67.725 72.200 68.175 ;
        RECT 78.120 67.975 79.120 68.125 ;
        RECT 68.760 67.715 69.220 67.725 ;
        RECT 71.460 67.715 71.920 67.725 ;
        RECT 74.655 67.715 75.115 67.945 ;
        RECT 77.355 67.715 77.815 67.945 ;
        RECT 77.970 67.525 79.120 67.975 ;
        RECT 80.055 67.715 80.515 67.945 ;
        RECT 85.825 67.725 86.825 68.175 ;
        RECT 86.085 67.715 86.545 67.725 ;
        RECT 65.300 62.820 66.300 67.145 ;
        RECT 67.740 66.175 68.110 66.225 ;
        RECT 67.025 65.120 68.110 66.175 ;
        RECT 63.500 61.075 66.330 62.075 ;
        RECT 67.025 60.425 68.025 65.120 ;
        RECT 68.480 62.500 68.710 67.510 ;
        RECT 69.270 62.500 69.500 67.510 ;
        RECT 69.870 65.120 70.240 66.225 ;
        RECT 70.440 65.120 70.810 66.225 ;
        RECT 71.180 62.500 71.410 67.510 ;
        RECT 71.970 62.500 72.200 67.510 ;
        RECT 74.375 66.510 74.605 67.510 ;
        RECT 75.145 66.495 77.325 67.525 ;
        RECT 77.820 67.500 79.120 67.525 ;
        RECT 79.775 67.500 80.005 67.510 ;
        RECT 80.565 67.500 80.795 67.510 ;
        RECT 77.820 66.975 80.075 67.500 ;
        RECT 77.820 66.570 78.740 66.975 ;
        RECT 77.865 66.510 78.095 66.570 ;
        RECT 79.030 66.520 80.075 66.975 ;
        RECT 80.495 66.520 80.865 67.500 ;
        RECT 79.775 66.510 80.005 66.520 ;
        RECT 80.565 66.510 80.795 66.520 ;
        RECT 72.570 65.120 72.940 66.225 ;
        RECT 74.370 63.625 75.370 66.355 ;
        RECT 77.095 63.625 78.095 66.325 ;
        RECT 79.520 65.850 80.555 66.325 ;
        RECT 85.065 65.120 85.435 66.225 ;
        RECT 79.515 63.605 80.555 64.100 ;
        RECT 74.055 62.800 74.700 63.480 ;
        RECT 75.095 62.800 77.375 63.480 ;
        RECT 77.865 63.405 78.095 63.465 ;
        RECT 79.775 63.455 80.005 63.465 ;
        RECT 80.565 63.455 80.795 63.465 ;
        RECT 77.820 63.250 78.740 63.405 ;
        RECT 79.030 63.250 80.075 63.455 ;
        RECT 77.820 62.825 80.075 63.250 ;
        RECT 80.495 62.825 80.865 63.455 ;
        RECT 77.865 62.815 79.120 62.825 ;
        RECT 79.775 62.815 80.005 62.825 ;
        RECT 80.565 62.815 80.795 62.825 ;
        RECT 77.870 62.800 79.120 62.815 ;
        RECT 61.875 59.425 68.025 60.425 ;
        RECT 63.360 58.715 63.820 58.945 ;
        RECT 66.060 58.715 66.520 58.945 ;
        RECT 63.080 58.500 63.310 58.510 ;
        RECT 63.870 58.500 64.100 58.510 ;
        RECT 65.780 58.500 66.010 58.510 ;
        RECT 66.570 58.500 66.800 58.510 ;
        RECT 62.335 57.520 63.380 58.500 ;
        RECT 63.800 57.520 64.170 58.500 ;
        RECT 65.035 57.520 66.080 58.500 ;
        RECT 66.500 57.520 66.870 58.500 ;
        RECT 68.410 57.520 68.780 62.500 ;
        RECT 69.200 57.520 69.570 62.500 ;
        RECT 71.110 57.520 71.480 62.500 ;
        RECT 71.900 57.520 72.270 62.500 ;
        RECT 74.655 62.425 75.115 62.655 ;
        RECT 77.355 62.425 77.815 62.655 ;
        RECT 77.965 62.250 79.120 62.800 ;
        RECT 80.055 62.425 80.515 62.655 ;
        RECT 85.805 62.500 86.035 67.510 ;
        RECT 86.595 62.500 86.825 67.510 ;
        RECT 88.000 67.145 89.925 68.175 ;
        RECT 87.195 66.175 87.565 66.225 ;
        RECT 87.195 65.120 88.300 66.175 ;
        RECT 77.965 62.200 79.025 62.250 ;
        RECT 57.680 57.510 57.910 57.520 ;
        RECT 58.470 57.510 58.700 57.520 ;
        RECT 60.380 57.510 60.610 57.520 ;
        RECT 61.170 57.510 61.400 57.520 ;
        RECT 63.080 57.510 63.310 57.520 ;
        RECT 63.870 57.510 64.100 57.520 ;
        RECT 65.780 57.510 66.010 57.520 ;
        RECT 66.570 57.510 66.800 57.520 ;
        RECT 68.480 57.510 68.710 57.520 ;
        RECT 69.270 57.510 69.500 57.520 ;
        RECT 71.180 57.510 71.410 57.520 ;
        RECT 71.970 57.510 72.200 57.520 ;
        RECT 57.425 56.850 58.460 57.325 ;
        RECT 60.660 57.075 61.120 57.305 ;
        RECT 62.825 56.850 63.860 57.325 ;
        RECT 65.525 56.850 66.560 57.325 ;
        RECT 68.760 57.075 69.220 57.305 ;
        RECT 71.460 57.075 71.920 57.305 ;
        RECT 54.800 56.475 55.800 56.530 ;
        RECT 75.670 56.510 76.775 61.180 ;
        RECT 83.385 58.715 83.845 58.945 ;
        RECT 83.105 58.500 83.335 58.510 ;
        RECT 83.895 58.500 84.125 58.510 ;
        RECT 82.360 57.520 83.405 58.500 ;
        RECT 83.825 57.520 84.195 58.500 ;
        RECT 85.735 57.520 86.105 62.500 ;
        RECT 86.525 57.520 86.895 62.500 ;
        RECT 87.300 60.425 88.300 65.120 ;
        RECT 88.925 62.075 89.925 67.145 ;
        RECT 90.725 67.145 92.675 68.175 ;
        RECT 93.925 67.725 94.925 68.175 ;
        RECT 96.625 67.725 97.625 68.175 ;
        RECT 94.185 67.715 94.645 67.725 ;
        RECT 96.885 67.715 97.345 67.725 ;
        RECT 90.725 62.820 91.725 67.145 ;
        RECT 93.165 66.175 93.535 66.225 ;
        RECT 92.450 65.120 93.535 66.175 ;
        RECT 88.925 61.075 91.755 62.075 ;
        RECT 92.450 60.425 93.450 65.120 ;
        RECT 93.905 62.500 94.135 67.510 ;
        RECT 94.695 62.500 94.925 67.510 ;
        RECT 95.295 65.120 95.665 66.225 ;
        RECT 95.865 65.120 96.235 66.225 ;
        RECT 96.605 62.500 96.835 67.510 ;
        RECT 97.395 62.500 97.625 67.510 ;
        RECT 97.995 65.120 98.365 66.225 ;
        RECT 87.300 59.425 93.450 60.425 ;
        RECT 88.785 58.715 89.245 58.945 ;
        RECT 91.485 58.715 91.945 58.945 ;
        RECT 88.505 58.500 88.735 58.510 ;
        RECT 89.295 58.500 89.525 58.510 ;
        RECT 91.205 58.500 91.435 58.510 ;
        RECT 91.995 58.500 92.225 58.510 ;
        RECT 87.760 57.520 88.805 58.500 ;
        RECT 89.225 57.520 89.595 58.500 ;
        RECT 90.460 57.520 91.505 58.500 ;
        RECT 91.925 57.520 92.295 58.500 ;
        RECT 93.835 57.520 94.205 62.500 ;
        RECT 94.625 57.520 94.995 62.500 ;
        RECT 96.535 57.520 96.905 62.500 ;
        RECT 97.325 57.520 97.695 62.500 ;
        RECT 83.105 57.510 83.335 57.520 ;
        RECT 83.895 57.510 84.125 57.520 ;
        RECT 85.805 57.510 86.035 57.520 ;
        RECT 86.595 57.510 86.825 57.520 ;
        RECT 88.505 57.510 88.735 57.520 ;
        RECT 89.295 57.510 89.525 57.520 ;
        RECT 91.205 57.510 91.435 57.520 ;
        RECT 91.995 57.510 92.225 57.520 ;
        RECT 93.905 57.510 94.135 57.520 ;
        RECT 94.695 57.510 94.925 57.520 ;
        RECT 96.605 57.510 96.835 57.520 ;
        RECT 97.395 57.510 97.625 57.520 ;
        RECT 82.850 56.850 83.885 57.325 ;
        RECT 86.085 57.075 86.545 57.305 ;
        RECT 88.250 56.850 89.285 57.325 ;
        RECT 90.950 56.850 91.985 57.325 ;
        RECT 94.185 57.075 94.645 57.305 ;
        RECT 96.885 57.075 97.345 57.305 ;
        RECT 80.225 56.510 81.225 56.530 ;
        RECT 50.695 55.475 51.755 56.475 ;
        RECT 54.770 55.475 55.830 56.475 ;
        RECT 6.570 54.605 7.610 55.100 ;
        RECT 9.810 54.625 10.270 54.855 ;
        RECT 11.970 54.605 13.010 55.100 ;
        RECT 14.670 54.605 15.710 55.100 ;
        RECT 17.910 54.625 18.370 54.855 ;
        RECT 20.610 54.625 21.070 54.855 ;
        RECT 6.830 54.455 7.060 54.465 ;
        RECT 7.620 54.455 7.850 54.465 ;
        RECT 9.530 54.455 9.760 54.465 ;
        RECT 10.320 54.455 10.550 54.465 ;
        RECT 12.230 54.455 12.460 54.465 ;
        RECT 13.020 54.455 13.250 54.465 ;
        RECT 14.930 54.455 15.160 54.465 ;
        RECT 15.720 54.455 15.950 54.465 ;
        RECT 17.630 54.455 17.860 54.465 ;
        RECT 18.420 54.455 18.650 54.465 ;
        RECT 20.330 54.455 20.560 54.465 ;
        RECT 21.120 54.455 21.350 54.465 ;
        RECT 6.085 53.825 7.130 54.455 ;
        RECT 7.550 53.825 7.920 54.455 ;
        RECT 6.830 53.815 7.060 53.825 ;
        RECT 7.620 53.815 7.850 53.825 ;
        RECT 7.110 53.425 7.570 53.655 ;
        RECT 1.900 51.250 4.950 52.250 ;
        RECT 9.460 51.275 9.830 54.455 ;
        RECT 10.250 51.275 10.620 54.455 ;
        RECT 11.485 53.825 12.530 54.455 ;
        RECT 12.950 53.825 13.320 54.455 ;
        RECT 14.185 53.825 15.230 54.455 ;
        RECT 15.650 53.825 16.020 54.455 ;
        RECT 12.230 53.815 12.460 53.825 ;
        RECT 13.020 53.815 13.250 53.825 ;
        RECT 14.930 53.815 15.160 53.825 ;
        RECT 15.720 53.815 15.950 53.825 ;
        RECT 12.510 53.425 12.970 53.655 ;
        RECT 15.210 53.425 15.670 53.655 ;
        RECT 17.560 51.275 17.930 54.455 ;
        RECT 18.350 51.275 18.720 54.455 ;
        RECT 20.260 51.275 20.630 54.455 ;
        RECT 21.050 51.275 21.420 54.455 ;
        RECT 29.375 52.250 30.375 55.405 ;
        RECT 31.995 54.605 33.035 55.100 ;
        RECT 35.235 54.625 35.695 54.855 ;
        RECT 37.395 54.605 38.435 55.100 ;
        RECT 40.095 54.605 41.135 55.100 ;
        RECT 43.335 54.625 43.795 54.855 ;
        RECT 46.035 54.625 46.495 54.855 ;
        RECT 32.255 54.455 32.485 54.465 ;
        RECT 33.045 54.455 33.275 54.465 ;
        RECT 34.955 54.455 35.185 54.465 ;
        RECT 35.745 54.455 35.975 54.465 ;
        RECT 37.655 54.455 37.885 54.465 ;
        RECT 38.445 54.455 38.675 54.465 ;
        RECT 40.355 54.455 40.585 54.465 ;
        RECT 41.145 54.455 41.375 54.465 ;
        RECT 43.055 54.455 43.285 54.465 ;
        RECT 43.845 54.455 44.075 54.465 ;
        RECT 45.755 54.455 45.985 54.465 ;
        RECT 46.545 54.455 46.775 54.465 ;
        RECT 31.510 53.825 32.555 54.455 ;
        RECT 32.975 53.825 33.345 54.455 ;
        RECT 32.255 53.815 32.485 53.825 ;
        RECT 33.045 53.815 33.275 53.825 ;
        RECT 32.535 53.425 32.995 53.655 ;
        RECT 1.900 33.900 2.900 51.250 ;
        RECT 3.905 50.430 5.020 50.485 ;
        RECT 3.875 49.315 5.050 50.430 ;
        RECT 8.790 49.320 9.160 50.435 ;
        RECT 1.870 32.900 2.930 33.900 ;
        RECT 1.900 11.325 2.900 32.900 ;
        RECT 3.905 27.855 5.020 49.315 ;
        RECT 9.530 47.965 9.760 51.275 ;
        RECT 10.320 47.965 10.550 51.275 ;
        RECT 10.920 49.320 11.290 50.435 ;
        RECT 16.890 49.320 17.260 50.435 ;
        RECT 17.630 47.965 17.860 51.275 ;
        RECT 18.420 47.965 18.650 51.275 ;
        RECT 19.020 49.320 19.390 50.435 ;
        RECT 19.590 49.320 19.960 50.435 ;
        RECT 20.330 47.965 20.560 51.275 ;
        RECT 21.120 47.965 21.350 51.275 ;
        RECT 27.325 51.250 30.375 52.250 ;
        RECT 34.885 51.275 35.255 54.455 ;
        RECT 35.675 51.275 36.045 54.455 ;
        RECT 36.910 53.825 37.955 54.455 ;
        RECT 38.375 53.825 38.745 54.455 ;
        RECT 39.610 53.825 40.655 54.455 ;
        RECT 41.075 53.825 41.445 54.455 ;
        RECT 37.655 53.815 37.885 53.825 ;
        RECT 38.445 53.815 38.675 53.825 ;
        RECT 40.355 53.815 40.585 53.825 ;
        RECT 41.145 53.815 41.375 53.825 ;
        RECT 37.935 53.425 38.395 53.655 ;
        RECT 40.635 53.425 41.095 53.655 ;
        RECT 42.985 51.275 43.355 54.455 ;
        RECT 43.775 51.275 44.145 54.455 ;
        RECT 45.685 51.275 46.055 54.455 ;
        RECT 46.475 51.275 46.845 54.455 ;
        RECT 54.800 52.250 55.800 55.475 ;
        RECT 75.670 55.405 81.280 56.510 ;
        RECT 101.575 56.475 102.575 69.550 ;
        RECT 113.425 68.175 114.425 68.205 ;
        RECT 117.100 68.175 118.100 68.205 ;
        RECT 138.850 68.175 139.850 68.205 ;
        RECT 142.525 68.175 143.525 68.205 ;
        RECT 111.250 67.725 112.250 68.175 ;
        RECT 111.510 67.715 111.970 67.725 ;
        RECT 110.490 65.120 110.860 66.225 ;
        RECT 111.230 62.500 111.460 67.510 ;
        RECT 112.020 62.500 112.250 67.510 ;
        RECT 113.425 67.145 115.350 68.175 ;
        RECT 112.620 66.175 112.990 66.225 ;
        RECT 112.620 65.120 113.725 66.175 ;
        RECT 108.810 58.715 109.270 58.945 ;
        RECT 108.530 58.500 108.760 58.510 ;
        RECT 109.320 58.500 109.550 58.510 ;
        RECT 107.785 57.520 108.830 58.500 ;
        RECT 109.250 57.520 109.620 58.500 ;
        RECT 111.160 57.520 111.530 62.500 ;
        RECT 111.950 57.520 112.320 62.500 ;
        RECT 112.725 60.425 113.725 65.120 ;
        RECT 114.350 62.075 115.350 67.145 ;
        RECT 116.150 67.145 118.100 68.175 ;
        RECT 119.350 67.725 120.350 68.175 ;
        RECT 122.050 67.725 123.050 68.175 ;
        RECT 128.970 67.975 129.970 68.125 ;
        RECT 119.610 67.715 120.070 67.725 ;
        RECT 122.310 67.715 122.770 67.725 ;
        RECT 125.505 67.715 125.965 67.945 ;
        RECT 128.205 67.715 128.665 67.945 ;
        RECT 128.820 67.525 129.970 67.975 ;
        RECT 130.905 67.715 131.365 67.945 ;
        RECT 136.675 67.725 137.675 68.175 ;
        RECT 136.935 67.715 137.395 67.725 ;
        RECT 116.150 62.820 117.150 67.145 ;
        RECT 118.590 66.175 118.960 66.225 ;
        RECT 117.875 65.120 118.960 66.175 ;
        RECT 114.350 61.075 117.180 62.075 ;
        RECT 117.875 60.425 118.875 65.120 ;
        RECT 119.330 62.500 119.560 67.510 ;
        RECT 120.120 62.500 120.350 67.510 ;
        RECT 120.720 65.120 121.090 66.225 ;
        RECT 121.290 65.120 121.660 66.225 ;
        RECT 122.030 62.500 122.260 67.510 ;
        RECT 122.820 62.500 123.050 67.510 ;
        RECT 125.225 66.510 125.455 67.510 ;
        RECT 125.995 66.495 128.175 67.525 ;
        RECT 128.670 67.500 129.970 67.525 ;
        RECT 130.625 67.500 130.855 67.510 ;
        RECT 131.415 67.500 131.645 67.510 ;
        RECT 128.670 66.975 130.925 67.500 ;
        RECT 128.670 66.570 129.590 66.975 ;
        RECT 128.715 66.510 128.945 66.570 ;
        RECT 129.880 66.520 130.925 66.975 ;
        RECT 131.345 66.520 131.715 67.500 ;
        RECT 130.625 66.510 130.855 66.520 ;
        RECT 131.415 66.510 131.645 66.520 ;
        RECT 123.420 65.120 123.790 66.225 ;
        RECT 125.220 63.625 126.220 66.355 ;
        RECT 127.945 63.625 128.945 66.325 ;
        RECT 130.370 65.850 131.405 66.325 ;
        RECT 135.915 65.120 136.285 66.225 ;
        RECT 130.365 63.605 131.405 64.100 ;
        RECT 124.905 62.800 125.550 63.480 ;
        RECT 125.945 62.800 128.225 63.480 ;
        RECT 128.715 63.405 128.945 63.465 ;
        RECT 130.625 63.455 130.855 63.465 ;
        RECT 131.415 63.455 131.645 63.465 ;
        RECT 128.670 63.250 129.590 63.405 ;
        RECT 129.880 63.250 130.925 63.455 ;
        RECT 128.670 62.825 130.925 63.250 ;
        RECT 131.345 62.825 131.715 63.455 ;
        RECT 128.715 62.815 129.970 62.825 ;
        RECT 130.625 62.815 130.855 62.825 ;
        RECT 131.415 62.815 131.645 62.825 ;
        RECT 128.720 62.800 129.970 62.815 ;
        RECT 112.725 59.425 118.875 60.425 ;
        RECT 114.210 58.715 114.670 58.945 ;
        RECT 116.910 58.715 117.370 58.945 ;
        RECT 113.930 58.500 114.160 58.510 ;
        RECT 114.720 58.500 114.950 58.510 ;
        RECT 116.630 58.500 116.860 58.510 ;
        RECT 117.420 58.500 117.650 58.510 ;
        RECT 113.185 57.520 114.230 58.500 ;
        RECT 114.650 57.520 115.020 58.500 ;
        RECT 115.885 57.520 116.930 58.500 ;
        RECT 117.350 57.520 117.720 58.500 ;
        RECT 119.260 57.520 119.630 62.500 ;
        RECT 120.050 57.520 120.420 62.500 ;
        RECT 121.960 57.520 122.330 62.500 ;
        RECT 122.750 57.520 123.120 62.500 ;
        RECT 125.505 62.425 125.965 62.655 ;
        RECT 128.205 62.425 128.665 62.655 ;
        RECT 128.815 62.250 129.970 62.800 ;
        RECT 130.905 62.425 131.365 62.655 ;
        RECT 136.655 62.500 136.885 67.510 ;
        RECT 137.445 62.500 137.675 67.510 ;
        RECT 138.850 67.145 140.775 68.175 ;
        RECT 138.045 66.175 138.415 66.225 ;
        RECT 138.045 65.120 139.150 66.175 ;
        RECT 128.815 62.200 129.875 62.250 ;
        RECT 108.530 57.510 108.760 57.520 ;
        RECT 109.320 57.510 109.550 57.520 ;
        RECT 111.230 57.510 111.460 57.520 ;
        RECT 112.020 57.510 112.250 57.520 ;
        RECT 113.930 57.510 114.160 57.520 ;
        RECT 114.720 57.510 114.950 57.520 ;
        RECT 116.630 57.510 116.860 57.520 ;
        RECT 117.420 57.510 117.650 57.520 ;
        RECT 119.330 57.510 119.560 57.520 ;
        RECT 120.120 57.510 120.350 57.520 ;
        RECT 122.030 57.510 122.260 57.520 ;
        RECT 122.820 57.510 123.050 57.520 ;
        RECT 108.275 56.850 109.310 57.325 ;
        RECT 111.510 57.075 111.970 57.305 ;
        RECT 113.675 56.850 114.710 57.325 ;
        RECT 116.375 56.850 117.410 57.325 ;
        RECT 119.610 57.075 120.070 57.305 ;
        RECT 122.310 57.075 122.770 57.305 ;
        RECT 105.650 56.475 106.650 56.530 ;
        RECT 126.520 56.510 127.625 61.180 ;
        RECT 134.235 58.715 134.695 58.945 ;
        RECT 133.955 58.500 134.185 58.510 ;
        RECT 134.745 58.500 134.975 58.510 ;
        RECT 133.210 57.520 134.255 58.500 ;
        RECT 134.675 57.520 135.045 58.500 ;
        RECT 136.585 57.520 136.955 62.500 ;
        RECT 137.375 57.520 137.745 62.500 ;
        RECT 138.150 60.425 139.150 65.120 ;
        RECT 139.775 62.075 140.775 67.145 ;
        RECT 141.575 67.145 143.525 68.175 ;
        RECT 144.775 67.725 145.775 68.175 ;
        RECT 147.475 67.725 148.475 68.175 ;
        RECT 145.035 67.715 145.495 67.725 ;
        RECT 147.735 67.715 148.195 67.725 ;
        RECT 141.575 62.820 142.575 67.145 ;
        RECT 144.015 66.175 144.385 66.225 ;
        RECT 143.300 65.120 144.385 66.175 ;
        RECT 139.775 61.075 142.605 62.075 ;
        RECT 143.300 60.425 144.300 65.120 ;
        RECT 144.755 62.500 144.985 67.510 ;
        RECT 145.545 62.500 145.775 67.510 ;
        RECT 146.145 65.120 146.515 66.225 ;
        RECT 146.715 65.120 147.085 66.225 ;
        RECT 147.455 62.500 147.685 67.510 ;
        RECT 148.245 62.500 148.475 67.510 ;
        RECT 148.845 65.120 149.215 66.225 ;
        RECT 138.150 59.425 144.300 60.425 ;
        RECT 139.635 58.715 140.095 58.945 ;
        RECT 142.335 58.715 142.795 58.945 ;
        RECT 139.355 58.500 139.585 58.510 ;
        RECT 140.145 58.500 140.375 58.510 ;
        RECT 142.055 58.500 142.285 58.510 ;
        RECT 142.845 58.500 143.075 58.510 ;
        RECT 138.610 57.520 139.655 58.500 ;
        RECT 140.075 57.520 140.445 58.500 ;
        RECT 141.310 57.520 142.355 58.500 ;
        RECT 142.775 57.520 143.145 58.500 ;
        RECT 144.685 57.520 145.055 62.500 ;
        RECT 145.475 57.520 145.845 62.500 ;
        RECT 147.385 57.520 147.755 62.500 ;
        RECT 148.175 57.520 148.545 62.500 ;
        RECT 133.955 57.510 134.185 57.520 ;
        RECT 134.745 57.510 134.975 57.520 ;
        RECT 136.655 57.510 136.885 57.520 ;
        RECT 137.445 57.510 137.675 57.520 ;
        RECT 139.355 57.510 139.585 57.520 ;
        RECT 140.145 57.510 140.375 57.520 ;
        RECT 142.055 57.510 142.285 57.520 ;
        RECT 142.845 57.510 143.075 57.520 ;
        RECT 144.755 57.510 144.985 57.520 ;
        RECT 145.545 57.510 145.775 57.520 ;
        RECT 147.455 57.510 147.685 57.520 ;
        RECT 148.245 57.510 148.475 57.520 ;
        RECT 133.700 56.850 134.735 57.325 ;
        RECT 136.935 57.075 137.395 57.305 ;
        RECT 139.100 56.850 140.135 57.325 ;
        RECT 141.800 56.850 142.835 57.325 ;
        RECT 145.035 57.075 145.495 57.305 ;
        RECT 147.735 57.075 148.195 57.305 ;
        RECT 131.075 56.510 132.075 56.530 ;
        RECT 101.545 55.475 102.605 56.475 ;
        RECT 105.620 55.475 106.680 56.475 ;
        RECT 57.420 54.605 58.460 55.100 ;
        RECT 60.660 54.625 61.120 54.855 ;
        RECT 62.820 54.605 63.860 55.100 ;
        RECT 65.520 54.605 66.560 55.100 ;
        RECT 68.760 54.625 69.220 54.855 ;
        RECT 71.460 54.625 71.920 54.855 ;
        RECT 57.680 54.455 57.910 54.465 ;
        RECT 58.470 54.455 58.700 54.465 ;
        RECT 60.380 54.455 60.610 54.465 ;
        RECT 61.170 54.455 61.400 54.465 ;
        RECT 63.080 54.455 63.310 54.465 ;
        RECT 63.870 54.455 64.100 54.465 ;
        RECT 65.780 54.455 66.010 54.465 ;
        RECT 66.570 54.455 66.800 54.465 ;
        RECT 68.480 54.455 68.710 54.465 ;
        RECT 69.270 54.455 69.500 54.465 ;
        RECT 71.180 54.455 71.410 54.465 ;
        RECT 71.970 54.455 72.200 54.465 ;
        RECT 56.935 53.825 57.980 54.455 ;
        RECT 58.400 53.825 58.770 54.455 ;
        RECT 57.680 53.815 57.910 53.825 ;
        RECT 58.470 53.815 58.700 53.825 ;
        RECT 57.960 53.425 58.420 53.655 ;
        RECT 21.720 49.320 22.090 50.435 ;
        RECT 9.810 47.775 10.270 47.805 ;
        RECT 17.910 47.775 18.370 47.805 ;
        RECT 20.610 47.775 21.070 47.805 ;
        RECT 9.550 47.375 10.550 47.775 ;
        RECT 17.650 47.375 18.650 47.775 ;
        RECT 20.350 47.375 21.350 47.775 ;
        RECT 11.725 45.600 12.725 45.630 ;
        RECT 15.400 45.600 16.400 45.630 ;
        RECT 9.550 45.150 10.550 45.600 ;
        RECT 9.810 45.140 10.270 45.150 ;
        RECT 8.790 42.545 9.160 43.650 ;
        RECT 9.530 39.925 9.760 44.935 ;
        RECT 10.320 39.925 10.550 44.935 ;
        RECT 11.725 44.570 13.650 45.600 ;
        RECT 10.920 43.600 11.290 43.650 ;
        RECT 10.920 42.545 12.025 43.600 ;
        RECT 7.110 36.140 7.570 36.370 ;
        RECT 6.830 35.925 7.060 35.935 ;
        RECT 7.620 35.925 7.850 35.935 ;
        RECT 6.085 34.945 7.130 35.925 ;
        RECT 7.550 34.945 7.920 35.925 ;
        RECT 9.460 34.945 9.830 39.925 ;
        RECT 10.250 34.945 10.620 39.925 ;
        RECT 11.025 37.850 12.025 42.545 ;
        RECT 12.650 39.500 13.650 44.570 ;
        RECT 14.450 44.570 16.400 45.600 ;
        RECT 17.650 45.150 18.650 45.600 ;
        RECT 20.350 45.150 21.350 45.600 ;
        RECT 17.910 45.140 18.370 45.150 ;
        RECT 20.610 45.140 21.070 45.150 ;
        RECT 14.450 40.245 15.450 44.570 ;
        RECT 16.890 43.600 17.260 43.650 ;
        RECT 16.175 42.545 17.260 43.600 ;
        RECT 12.650 38.500 15.480 39.500 ;
        RECT 16.175 37.850 17.175 42.545 ;
        RECT 17.630 39.925 17.860 44.935 ;
        RECT 18.420 39.925 18.650 44.935 ;
        RECT 19.020 42.545 19.390 43.650 ;
        RECT 19.590 42.545 19.960 43.650 ;
        RECT 20.330 39.925 20.560 44.935 ;
        RECT 21.120 39.925 21.350 44.935 ;
        RECT 21.720 42.545 22.090 43.650 ;
        RECT 11.025 36.850 17.175 37.850 ;
        RECT 12.510 36.140 12.970 36.370 ;
        RECT 15.210 36.140 15.670 36.370 ;
        RECT 12.230 35.925 12.460 35.935 ;
        RECT 13.020 35.925 13.250 35.935 ;
        RECT 14.930 35.925 15.160 35.935 ;
        RECT 15.720 35.925 15.950 35.935 ;
        RECT 11.485 34.945 12.530 35.925 ;
        RECT 12.950 34.945 13.320 35.925 ;
        RECT 14.185 34.945 15.230 35.925 ;
        RECT 15.650 34.945 16.020 35.925 ;
        RECT 17.560 34.945 17.930 39.925 ;
        RECT 18.350 34.945 18.720 39.925 ;
        RECT 20.260 34.945 20.630 39.925 ;
        RECT 21.050 34.945 21.420 39.925 ;
        RECT 6.830 34.935 7.060 34.945 ;
        RECT 7.620 34.935 7.850 34.945 ;
        RECT 9.530 34.935 9.760 34.945 ;
        RECT 10.320 34.935 10.550 34.945 ;
        RECT 12.230 34.935 12.460 34.945 ;
        RECT 13.020 34.935 13.250 34.945 ;
        RECT 14.930 34.935 15.160 34.945 ;
        RECT 15.720 34.935 15.950 34.945 ;
        RECT 17.630 34.935 17.860 34.945 ;
        RECT 18.420 34.935 18.650 34.945 ;
        RECT 20.330 34.935 20.560 34.945 ;
        RECT 21.120 34.935 21.350 34.945 ;
        RECT 6.575 34.275 7.610 34.750 ;
        RECT 9.810 34.500 10.270 34.730 ;
        RECT 11.975 34.275 13.010 34.750 ;
        RECT 14.675 34.275 15.710 34.750 ;
        RECT 17.910 34.500 18.370 34.730 ;
        RECT 20.610 34.500 21.070 34.730 ;
        RECT 27.325 33.900 28.325 51.250 ;
        RECT 29.330 50.430 30.445 50.485 ;
        RECT 29.300 49.315 30.475 50.430 ;
        RECT 34.215 49.320 34.585 50.435 ;
        RECT 27.295 32.900 28.355 33.900 ;
        RECT 6.570 32.030 7.610 32.525 ;
        RECT 9.810 32.050 10.270 32.280 ;
        RECT 11.970 32.030 13.010 32.525 ;
        RECT 14.670 32.030 15.710 32.525 ;
        RECT 17.910 32.050 18.370 32.280 ;
        RECT 20.610 32.050 21.070 32.280 ;
        RECT 6.830 31.880 7.060 31.890 ;
        RECT 7.620 31.880 7.850 31.890 ;
        RECT 9.530 31.880 9.760 31.890 ;
        RECT 10.320 31.880 10.550 31.890 ;
        RECT 12.230 31.880 12.460 31.890 ;
        RECT 13.020 31.880 13.250 31.890 ;
        RECT 14.930 31.880 15.160 31.890 ;
        RECT 15.720 31.880 15.950 31.890 ;
        RECT 17.630 31.880 17.860 31.890 ;
        RECT 18.420 31.880 18.650 31.890 ;
        RECT 20.330 31.880 20.560 31.890 ;
        RECT 21.120 31.880 21.350 31.890 ;
        RECT 6.085 31.250 7.130 31.880 ;
        RECT 7.550 31.250 7.920 31.880 ;
        RECT 6.830 31.240 7.060 31.250 ;
        RECT 7.620 31.240 7.850 31.250 ;
        RECT 7.110 30.850 7.570 31.080 ;
        RECT 9.460 28.700 9.830 31.880 ;
        RECT 10.250 28.700 10.620 31.880 ;
        RECT 11.485 31.250 12.530 31.880 ;
        RECT 12.950 31.250 13.320 31.880 ;
        RECT 14.185 31.250 15.230 31.880 ;
        RECT 15.650 31.250 16.020 31.880 ;
        RECT 12.230 31.240 12.460 31.250 ;
        RECT 13.020 31.240 13.250 31.250 ;
        RECT 14.930 31.240 15.160 31.250 ;
        RECT 15.720 31.240 15.950 31.250 ;
        RECT 12.510 30.850 12.970 31.080 ;
        RECT 15.210 30.850 15.670 31.080 ;
        RECT 17.560 28.700 17.930 31.880 ;
        RECT 18.350 28.700 18.720 31.880 ;
        RECT 20.260 28.700 20.630 31.880 ;
        RECT 21.050 28.700 21.420 31.880 ;
        RECT 3.875 26.740 5.050 27.855 ;
        RECT 8.790 26.745 9.160 27.860 ;
        RECT 1.870 10.325 2.930 11.325 ;
        RECT 1.900 10.295 2.900 10.325 ;
        RECT 3.905 5.285 5.020 26.740 ;
        RECT 9.530 25.390 9.760 28.700 ;
        RECT 10.320 25.390 10.550 28.700 ;
        RECT 10.920 26.745 11.290 27.860 ;
        RECT 16.890 26.745 17.260 27.860 ;
        RECT 17.630 25.390 17.860 28.700 ;
        RECT 18.420 25.390 18.650 28.700 ;
        RECT 19.020 26.745 19.390 27.860 ;
        RECT 19.590 26.745 19.960 27.860 ;
        RECT 20.330 25.390 20.560 28.700 ;
        RECT 21.120 25.390 21.350 28.700 ;
        RECT 21.720 26.745 22.090 27.860 ;
        RECT 23.085 26.745 24.260 27.860 ;
        RECT 9.810 25.200 10.270 25.230 ;
        RECT 17.910 25.200 18.370 25.230 ;
        RECT 20.610 25.200 21.070 25.230 ;
        RECT 9.550 24.800 10.550 25.200 ;
        RECT 17.650 24.800 18.650 25.200 ;
        RECT 20.350 24.800 21.350 25.200 ;
        RECT 23.115 23.770 24.230 26.745 ;
        RECT 11.725 23.025 12.725 23.055 ;
        RECT 15.400 23.025 16.400 23.055 ;
        RECT 9.550 22.575 10.550 23.025 ;
        RECT 9.810 22.565 10.270 22.575 ;
        RECT 8.790 19.970 9.160 21.075 ;
        RECT 9.530 17.350 9.760 22.360 ;
        RECT 10.320 17.350 10.550 22.360 ;
        RECT 11.725 21.995 13.650 23.025 ;
        RECT 10.920 21.025 11.290 21.075 ;
        RECT 10.920 19.970 12.025 21.025 ;
        RECT 7.110 13.565 7.570 13.795 ;
        RECT 6.830 13.350 7.060 13.360 ;
        RECT 7.620 13.350 7.850 13.360 ;
        RECT 6.085 12.370 7.130 13.350 ;
        RECT 7.550 12.370 7.920 13.350 ;
        RECT 9.460 12.370 9.830 17.350 ;
        RECT 10.250 12.370 10.620 17.350 ;
        RECT 11.025 15.275 12.025 19.970 ;
        RECT 12.650 16.925 13.650 21.995 ;
        RECT 14.450 21.995 16.400 23.025 ;
        RECT 17.650 22.575 18.650 23.025 ;
        RECT 20.350 22.575 21.350 23.025 ;
        RECT 17.910 22.565 18.370 22.575 ;
        RECT 20.610 22.565 21.070 22.575 ;
        RECT 14.450 17.670 15.450 21.995 ;
        RECT 16.890 21.025 17.260 21.075 ;
        RECT 16.175 19.970 17.260 21.025 ;
        RECT 12.650 15.925 15.480 16.925 ;
        RECT 16.175 15.275 17.175 19.970 ;
        RECT 17.630 17.350 17.860 22.360 ;
        RECT 18.420 17.350 18.650 22.360 ;
        RECT 19.020 19.970 19.390 21.075 ;
        RECT 19.590 19.970 19.960 21.075 ;
        RECT 20.330 17.350 20.560 22.360 ;
        RECT 21.120 17.350 21.350 22.360 ;
        RECT 23.430 21.115 23.880 23.425 ;
        RECT 21.720 19.970 22.090 21.075 ;
        RECT 11.025 14.275 17.175 15.275 ;
        RECT 12.510 13.565 12.970 13.795 ;
        RECT 15.210 13.565 15.670 13.795 ;
        RECT 12.230 13.350 12.460 13.360 ;
        RECT 13.020 13.350 13.250 13.360 ;
        RECT 14.930 13.350 15.160 13.360 ;
        RECT 15.720 13.350 15.950 13.360 ;
        RECT 11.485 12.370 12.530 13.350 ;
        RECT 12.950 12.370 13.320 13.350 ;
        RECT 14.185 12.370 15.230 13.350 ;
        RECT 15.650 12.370 16.020 13.350 ;
        RECT 17.560 12.370 17.930 17.350 ;
        RECT 18.350 12.370 18.720 17.350 ;
        RECT 20.260 12.370 20.630 17.350 ;
        RECT 21.050 12.370 21.420 17.350 ;
        RECT 6.830 12.360 7.060 12.370 ;
        RECT 7.620 12.360 7.850 12.370 ;
        RECT 9.530 12.360 9.760 12.370 ;
        RECT 10.320 12.360 10.550 12.370 ;
        RECT 12.230 12.360 12.460 12.370 ;
        RECT 13.020 12.360 13.250 12.370 ;
        RECT 14.930 12.360 15.160 12.370 ;
        RECT 15.720 12.360 15.950 12.370 ;
        RECT 17.630 12.360 17.860 12.370 ;
        RECT 18.420 12.360 18.650 12.370 ;
        RECT 20.330 12.360 20.560 12.370 ;
        RECT 21.120 12.360 21.350 12.370 ;
        RECT 6.575 11.700 7.610 12.175 ;
        RECT 9.810 11.925 10.270 12.155 ;
        RECT 11.975 11.700 13.010 12.175 ;
        RECT 14.675 11.700 15.710 12.175 ;
        RECT 17.910 11.925 18.370 12.155 ;
        RECT 20.610 11.925 21.070 12.155 ;
        RECT 23.430 10.205 23.880 12.515 ;
        RECT 27.325 11.325 28.325 32.900 ;
        RECT 29.330 27.855 30.445 49.315 ;
        RECT 34.955 47.965 35.185 51.275 ;
        RECT 35.745 47.965 35.975 51.275 ;
        RECT 36.345 49.320 36.715 50.435 ;
        RECT 42.315 49.320 42.685 50.435 ;
        RECT 43.055 47.965 43.285 51.275 ;
        RECT 43.845 47.965 44.075 51.275 ;
        RECT 44.445 49.320 44.815 50.435 ;
        RECT 45.015 49.320 45.385 50.435 ;
        RECT 45.755 47.965 45.985 51.275 ;
        RECT 46.545 47.965 46.775 51.275 ;
        RECT 52.750 51.250 55.800 52.250 ;
        RECT 60.310 51.275 60.680 54.455 ;
        RECT 61.100 51.275 61.470 54.455 ;
        RECT 62.335 53.825 63.380 54.455 ;
        RECT 63.800 53.825 64.170 54.455 ;
        RECT 65.035 53.825 66.080 54.455 ;
        RECT 66.500 53.825 66.870 54.455 ;
        RECT 63.080 53.815 63.310 53.825 ;
        RECT 63.870 53.815 64.100 53.825 ;
        RECT 65.780 53.815 66.010 53.825 ;
        RECT 66.570 53.815 66.800 53.825 ;
        RECT 63.360 53.425 63.820 53.655 ;
        RECT 66.060 53.425 66.520 53.655 ;
        RECT 68.410 51.275 68.780 54.455 ;
        RECT 69.200 51.275 69.570 54.455 ;
        RECT 71.110 51.275 71.480 54.455 ;
        RECT 71.900 51.275 72.270 54.455 ;
        RECT 80.225 52.250 81.225 55.405 ;
        RECT 82.845 54.605 83.885 55.100 ;
        RECT 86.085 54.625 86.545 54.855 ;
        RECT 88.245 54.605 89.285 55.100 ;
        RECT 90.945 54.605 91.985 55.100 ;
        RECT 94.185 54.625 94.645 54.855 ;
        RECT 96.885 54.625 97.345 54.855 ;
        RECT 83.105 54.455 83.335 54.465 ;
        RECT 83.895 54.455 84.125 54.465 ;
        RECT 85.805 54.455 86.035 54.465 ;
        RECT 86.595 54.455 86.825 54.465 ;
        RECT 88.505 54.455 88.735 54.465 ;
        RECT 89.295 54.455 89.525 54.465 ;
        RECT 91.205 54.455 91.435 54.465 ;
        RECT 91.995 54.455 92.225 54.465 ;
        RECT 93.905 54.455 94.135 54.465 ;
        RECT 94.695 54.455 94.925 54.465 ;
        RECT 96.605 54.455 96.835 54.465 ;
        RECT 97.395 54.455 97.625 54.465 ;
        RECT 82.360 53.825 83.405 54.455 ;
        RECT 83.825 53.825 84.195 54.455 ;
        RECT 83.105 53.815 83.335 53.825 ;
        RECT 83.895 53.815 84.125 53.825 ;
        RECT 83.385 53.425 83.845 53.655 ;
        RECT 47.145 49.320 47.515 50.435 ;
        RECT 35.235 47.775 35.695 47.805 ;
        RECT 43.335 47.775 43.795 47.805 ;
        RECT 46.035 47.775 46.495 47.805 ;
        RECT 34.975 47.375 35.975 47.775 ;
        RECT 43.075 47.375 44.075 47.775 ;
        RECT 45.775 47.375 46.775 47.775 ;
        RECT 37.150 45.600 38.150 45.630 ;
        RECT 40.825 45.600 41.825 45.630 ;
        RECT 34.975 45.150 35.975 45.600 ;
        RECT 35.235 45.140 35.695 45.150 ;
        RECT 34.215 42.545 34.585 43.650 ;
        RECT 34.955 39.925 35.185 44.935 ;
        RECT 35.745 39.925 35.975 44.935 ;
        RECT 37.150 44.570 39.075 45.600 ;
        RECT 36.345 43.600 36.715 43.650 ;
        RECT 36.345 42.545 37.450 43.600 ;
        RECT 32.535 36.140 32.995 36.370 ;
        RECT 32.255 35.925 32.485 35.935 ;
        RECT 33.045 35.925 33.275 35.935 ;
        RECT 31.510 34.945 32.555 35.925 ;
        RECT 32.975 34.945 33.345 35.925 ;
        RECT 34.885 34.945 35.255 39.925 ;
        RECT 35.675 34.945 36.045 39.925 ;
        RECT 36.450 37.850 37.450 42.545 ;
        RECT 38.075 39.500 39.075 44.570 ;
        RECT 39.875 44.570 41.825 45.600 ;
        RECT 43.075 45.150 44.075 45.600 ;
        RECT 45.775 45.150 46.775 45.600 ;
        RECT 43.335 45.140 43.795 45.150 ;
        RECT 46.035 45.140 46.495 45.150 ;
        RECT 39.875 40.245 40.875 44.570 ;
        RECT 42.315 43.600 42.685 43.650 ;
        RECT 41.600 42.545 42.685 43.600 ;
        RECT 38.075 38.500 40.905 39.500 ;
        RECT 41.600 37.850 42.600 42.545 ;
        RECT 43.055 39.925 43.285 44.935 ;
        RECT 43.845 39.925 44.075 44.935 ;
        RECT 44.445 42.545 44.815 43.650 ;
        RECT 45.015 42.545 45.385 43.650 ;
        RECT 45.755 39.925 45.985 44.935 ;
        RECT 46.545 39.925 46.775 44.935 ;
        RECT 47.145 42.545 47.515 43.650 ;
        RECT 36.450 36.850 42.600 37.850 ;
        RECT 37.935 36.140 38.395 36.370 ;
        RECT 40.635 36.140 41.095 36.370 ;
        RECT 37.655 35.925 37.885 35.935 ;
        RECT 38.445 35.925 38.675 35.935 ;
        RECT 40.355 35.925 40.585 35.935 ;
        RECT 41.145 35.925 41.375 35.935 ;
        RECT 36.910 34.945 37.955 35.925 ;
        RECT 38.375 34.945 38.745 35.925 ;
        RECT 39.610 34.945 40.655 35.925 ;
        RECT 41.075 34.945 41.445 35.925 ;
        RECT 42.985 34.945 43.355 39.925 ;
        RECT 43.775 34.945 44.145 39.925 ;
        RECT 45.685 34.945 46.055 39.925 ;
        RECT 46.475 34.945 46.845 39.925 ;
        RECT 32.255 34.935 32.485 34.945 ;
        RECT 33.045 34.935 33.275 34.945 ;
        RECT 34.955 34.935 35.185 34.945 ;
        RECT 35.745 34.935 35.975 34.945 ;
        RECT 37.655 34.935 37.885 34.945 ;
        RECT 38.445 34.935 38.675 34.945 ;
        RECT 40.355 34.935 40.585 34.945 ;
        RECT 41.145 34.935 41.375 34.945 ;
        RECT 43.055 34.935 43.285 34.945 ;
        RECT 43.845 34.935 44.075 34.945 ;
        RECT 45.755 34.935 45.985 34.945 ;
        RECT 46.545 34.935 46.775 34.945 ;
        RECT 32.000 34.275 33.035 34.750 ;
        RECT 35.235 34.500 35.695 34.730 ;
        RECT 37.400 34.275 38.435 34.750 ;
        RECT 40.100 34.275 41.135 34.750 ;
        RECT 43.335 34.500 43.795 34.730 ;
        RECT 46.035 34.500 46.495 34.730 ;
        RECT 52.750 33.900 53.750 51.250 ;
        RECT 54.755 50.430 55.870 50.485 ;
        RECT 54.725 49.315 55.900 50.430 ;
        RECT 59.640 49.320 60.010 50.435 ;
        RECT 52.720 32.900 53.780 33.900 ;
        RECT 31.995 32.030 33.035 32.525 ;
        RECT 35.235 32.050 35.695 32.280 ;
        RECT 37.395 32.030 38.435 32.525 ;
        RECT 40.095 32.030 41.135 32.525 ;
        RECT 43.335 32.050 43.795 32.280 ;
        RECT 46.035 32.050 46.495 32.280 ;
        RECT 32.255 31.880 32.485 31.890 ;
        RECT 33.045 31.880 33.275 31.890 ;
        RECT 34.955 31.880 35.185 31.890 ;
        RECT 35.745 31.880 35.975 31.890 ;
        RECT 37.655 31.880 37.885 31.890 ;
        RECT 38.445 31.880 38.675 31.890 ;
        RECT 40.355 31.880 40.585 31.890 ;
        RECT 41.145 31.880 41.375 31.890 ;
        RECT 43.055 31.880 43.285 31.890 ;
        RECT 43.845 31.880 44.075 31.890 ;
        RECT 45.755 31.880 45.985 31.890 ;
        RECT 46.545 31.880 46.775 31.890 ;
        RECT 31.510 31.250 32.555 31.880 ;
        RECT 32.975 31.250 33.345 31.880 ;
        RECT 32.255 31.240 32.485 31.250 ;
        RECT 33.045 31.240 33.275 31.250 ;
        RECT 32.535 30.850 32.995 31.080 ;
        RECT 34.885 28.700 35.255 31.880 ;
        RECT 35.675 28.700 36.045 31.880 ;
        RECT 36.910 31.250 37.955 31.880 ;
        RECT 38.375 31.250 38.745 31.880 ;
        RECT 39.610 31.250 40.655 31.880 ;
        RECT 41.075 31.250 41.445 31.880 ;
        RECT 37.655 31.240 37.885 31.250 ;
        RECT 38.445 31.240 38.675 31.250 ;
        RECT 40.355 31.240 40.585 31.250 ;
        RECT 41.145 31.240 41.375 31.250 ;
        RECT 37.935 30.850 38.395 31.080 ;
        RECT 40.635 30.850 41.095 31.080 ;
        RECT 42.985 28.700 43.355 31.880 ;
        RECT 43.775 28.700 44.145 31.880 ;
        RECT 45.685 28.700 46.055 31.880 ;
        RECT 46.475 28.700 46.845 31.880 ;
        RECT 29.300 26.740 30.475 27.855 ;
        RECT 34.215 26.745 34.585 27.860 ;
        RECT 27.295 10.325 28.355 11.325 ;
        RECT 27.325 10.295 28.325 10.325 ;
        RECT 6.570 9.455 7.610 9.950 ;
        RECT 9.810 9.475 10.270 9.705 ;
        RECT 11.970 9.455 13.010 9.950 ;
        RECT 14.670 9.455 15.710 9.950 ;
        RECT 17.910 9.475 18.370 9.705 ;
        RECT 20.610 9.475 21.070 9.705 ;
        RECT 6.830 9.305 7.060 9.315 ;
        RECT 7.620 9.305 7.850 9.315 ;
        RECT 9.530 9.305 9.760 9.315 ;
        RECT 10.320 9.305 10.550 9.315 ;
        RECT 12.230 9.305 12.460 9.315 ;
        RECT 13.020 9.305 13.250 9.315 ;
        RECT 14.930 9.305 15.160 9.315 ;
        RECT 15.720 9.305 15.950 9.315 ;
        RECT 17.630 9.305 17.860 9.315 ;
        RECT 18.420 9.305 18.650 9.315 ;
        RECT 20.330 9.305 20.560 9.315 ;
        RECT 21.120 9.305 21.350 9.315 ;
        RECT 6.085 8.675 7.130 9.305 ;
        RECT 7.550 8.675 7.920 9.305 ;
        RECT 6.830 8.665 7.060 8.675 ;
        RECT 7.620 8.665 7.850 8.675 ;
        RECT 7.110 8.275 7.570 8.505 ;
        RECT 9.460 6.125 9.830 9.305 ;
        RECT 10.250 6.125 10.620 9.305 ;
        RECT 11.485 8.675 12.530 9.305 ;
        RECT 12.950 8.675 13.320 9.305 ;
        RECT 14.185 8.675 15.230 9.305 ;
        RECT 15.650 8.675 16.020 9.305 ;
        RECT 12.230 8.665 12.460 8.675 ;
        RECT 13.020 8.665 13.250 8.675 ;
        RECT 14.930 8.665 15.160 8.675 ;
        RECT 15.720 8.665 15.950 8.675 ;
        RECT 12.510 8.275 12.970 8.505 ;
        RECT 15.210 8.275 15.670 8.505 ;
        RECT 17.560 6.125 17.930 9.305 ;
        RECT 18.350 6.125 18.720 9.305 ;
        RECT 20.260 6.125 20.630 9.305 ;
        RECT 21.050 6.125 21.420 9.305 ;
        RECT 3.860 4.170 5.060 5.285 ;
        RECT 8.790 4.170 9.160 5.285 ;
        RECT 3.905 4.140 5.020 4.170 ;
        RECT 9.530 2.815 9.760 6.125 ;
        RECT 10.320 2.815 10.550 6.125 ;
        RECT 10.920 4.170 11.290 5.285 ;
        RECT 16.890 4.170 17.260 5.285 ;
        RECT 17.630 2.815 17.860 6.125 ;
        RECT 18.420 2.815 18.650 6.125 ;
        RECT 19.020 4.170 19.390 5.285 ;
        RECT 19.590 4.170 19.960 5.285 ;
        RECT 20.330 2.815 20.560 6.125 ;
        RECT 21.120 2.815 21.350 6.125 ;
        RECT 21.720 4.170 22.090 5.285 ;
        RECT 23.090 4.140 24.205 9.855 ;
        RECT 29.330 5.285 30.445 26.740 ;
        RECT 34.955 25.390 35.185 28.700 ;
        RECT 35.745 25.390 35.975 28.700 ;
        RECT 36.345 26.745 36.715 27.860 ;
        RECT 42.315 26.745 42.685 27.860 ;
        RECT 43.055 25.390 43.285 28.700 ;
        RECT 43.845 25.390 44.075 28.700 ;
        RECT 44.445 26.745 44.815 27.860 ;
        RECT 45.015 26.745 45.385 27.860 ;
        RECT 45.755 25.390 45.985 28.700 ;
        RECT 46.545 25.390 46.775 28.700 ;
        RECT 47.145 26.745 47.515 27.860 ;
        RECT 48.510 26.745 49.685 27.860 ;
        RECT 35.235 25.200 35.695 25.230 ;
        RECT 43.335 25.200 43.795 25.230 ;
        RECT 46.035 25.200 46.495 25.230 ;
        RECT 34.975 24.800 35.975 25.200 ;
        RECT 43.075 24.800 44.075 25.200 ;
        RECT 45.775 24.800 46.775 25.200 ;
        RECT 48.540 23.770 49.655 26.745 ;
        RECT 37.150 23.025 38.150 23.055 ;
        RECT 40.825 23.025 41.825 23.055 ;
        RECT 34.975 22.575 35.975 23.025 ;
        RECT 35.235 22.565 35.695 22.575 ;
        RECT 34.215 19.970 34.585 21.075 ;
        RECT 34.955 17.350 35.185 22.360 ;
        RECT 35.745 17.350 35.975 22.360 ;
        RECT 37.150 21.995 39.075 23.025 ;
        RECT 36.345 21.025 36.715 21.075 ;
        RECT 36.345 19.970 37.450 21.025 ;
        RECT 32.535 13.565 32.995 13.795 ;
        RECT 32.255 13.350 32.485 13.360 ;
        RECT 33.045 13.350 33.275 13.360 ;
        RECT 31.510 12.370 32.555 13.350 ;
        RECT 32.975 12.370 33.345 13.350 ;
        RECT 34.885 12.370 35.255 17.350 ;
        RECT 35.675 12.370 36.045 17.350 ;
        RECT 36.450 15.275 37.450 19.970 ;
        RECT 38.075 16.925 39.075 21.995 ;
        RECT 39.875 21.995 41.825 23.025 ;
        RECT 43.075 22.575 44.075 23.025 ;
        RECT 45.775 22.575 46.775 23.025 ;
        RECT 43.335 22.565 43.795 22.575 ;
        RECT 46.035 22.565 46.495 22.575 ;
        RECT 39.875 17.670 40.875 21.995 ;
        RECT 42.315 21.025 42.685 21.075 ;
        RECT 41.600 19.970 42.685 21.025 ;
        RECT 38.075 15.925 40.905 16.925 ;
        RECT 41.600 15.275 42.600 19.970 ;
        RECT 43.055 17.350 43.285 22.360 ;
        RECT 43.845 17.350 44.075 22.360 ;
        RECT 44.445 19.970 44.815 21.075 ;
        RECT 45.015 19.970 45.385 21.075 ;
        RECT 45.755 17.350 45.985 22.360 ;
        RECT 46.545 17.350 46.775 22.360 ;
        RECT 48.855 21.115 49.305 23.425 ;
        RECT 47.145 19.970 47.515 21.075 ;
        RECT 36.450 14.275 42.600 15.275 ;
        RECT 37.935 13.565 38.395 13.795 ;
        RECT 40.635 13.565 41.095 13.795 ;
        RECT 37.655 13.350 37.885 13.360 ;
        RECT 38.445 13.350 38.675 13.360 ;
        RECT 40.355 13.350 40.585 13.360 ;
        RECT 41.145 13.350 41.375 13.360 ;
        RECT 36.910 12.370 37.955 13.350 ;
        RECT 38.375 12.370 38.745 13.350 ;
        RECT 39.610 12.370 40.655 13.350 ;
        RECT 41.075 12.370 41.445 13.350 ;
        RECT 42.985 12.370 43.355 17.350 ;
        RECT 43.775 12.370 44.145 17.350 ;
        RECT 45.685 12.370 46.055 17.350 ;
        RECT 46.475 12.370 46.845 17.350 ;
        RECT 32.255 12.360 32.485 12.370 ;
        RECT 33.045 12.360 33.275 12.370 ;
        RECT 34.955 12.360 35.185 12.370 ;
        RECT 35.745 12.360 35.975 12.370 ;
        RECT 37.655 12.360 37.885 12.370 ;
        RECT 38.445 12.360 38.675 12.370 ;
        RECT 40.355 12.360 40.585 12.370 ;
        RECT 41.145 12.360 41.375 12.370 ;
        RECT 43.055 12.360 43.285 12.370 ;
        RECT 43.845 12.360 44.075 12.370 ;
        RECT 45.755 12.360 45.985 12.370 ;
        RECT 46.545 12.360 46.775 12.370 ;
        RECT 32.000 11.700 33.035 12.175 ;
        RECT 35.235 11.925 35.695 12.155 ;
        RECT 37.400 11.700 38.435 12.175 ;
        RECT 40.100 11.700 41.135 12.175 ;
        RECT 43.335 11.925 43.795 12.155 ;
        RECT 46.035 11.925 46.495 12.155 ;
        RECT 48.855 10.205 49.305 12.515 ;
        RECT 52.750 11.325 53.750 32.900 ;
        RECT 54.755 27.855 55.870 49.315 ;
        RECT 60.380 47.965 60.610 51.275 ;
        RECT 61.170 47.965 61.400 51.275 ;
        RECT 61.770 49.320 62.140 50.435 ;
        RECT 67.740 49.320 68.110 50.435 ;
        RECT 68.480 47.965 68.710 51.275 ;
        RECT 69.270 47.965 69.500 51.275 ;
        RECT 69.870 49.320 70.240 50.435 ;
        RECT 70.440 49.320 70.810 50.435 ;
        RECT 71.180 47.965 71.410 51.275 ;
        RECT 71.970 47.965 72.200 51.275 ;
        RECT 78.175 51.250 81.225 52.250 ;
        RECT 85.735 51.275 86.105 54.455 ;
        RECT 86.525 51.275 86.895 54.455 ;
        RECT 87.760 53.825 88.805 54.455 ;
        RECT 89.225 53.825 89.595 54.455 ;
        RECT 90.460 53.825 91.505 54.455 ;
        RECT 91.925 53.825 92.295 54.455 ;
        RECT 88.505 53.815 88.735 53.825 ;
        RECT 89.295 53.815 89.525 53.825 ;
        RECT 91.205 53.815 91.435 53.825 ;
        RECT 91.995 53.815 92.225 53.825 ;
        RECT 88.785 53.425 89.245 53.655 ;
        RECT 91.485 53.425 91.945 53.655 ;
        RECT 93.835 51.275 94.205 54.455 ;
        RECT 94.625 51.275 94.995 54.455 ;
        RECT 96.535 51.275 96.905 54.455 ;
        RECT 97.325 51.275 97.695 54.455 ;
        RECT 105.650 52.250 106.650 55.475 ;
        RECT 126.520 55.405 132.130 56.510 ;
        RECT 152.425 56.475 153.425 69.550 ;
        RECT 152.395 55.475 153.455 56.475 ;
        RECT 108.270 54.605 109.310 55.100 ;
        RECT 111.510 54.625 111.970 54.855 ;
        RECT 113.670 54.605 114.710 55.100 ;
        RECT 116.370 54.605 117.410 55.100 ;
        RECT 119.610 54.625 120.070 54.855 ;
        RECT 122.310 54.625 122.770 54.855 ;
        RECT 108.530 54.455 108.760 54.465 ;
        RECT 109.320 54.455 109.550 54.465 ;
        RECT 111.230 54.455 111.460 54.465 ;
        RECT 112.020 54.455 112.250 54.465 ;
        RECT 113.930 54.455 114.160 54.465 ;
        RECT 114.720 54.455 114.950 54.465 ;
        RECT 116.630 54.455 116.860 54.465 ;
        RECT 117.420 54.455 117.650 54.465 ;
        RECT 119.330 54.455 119.560 54.465 ;
        RECT 120.120 54.455 120.350 54.465 ;
        RECT 122.030 54.455 122.260 54.465 ;
        RECT 122.820 54.455 123.050 54.465 ;
        RECT 107.785 53.825 108.830 54.455 ;
        RECT 109.250 53.825 109.620 54.455 ;
        RECT 108.530 53.815 108.760 53.825 ;
        RECT 109.320 53.815 109.550 53.825 ;
        RECT 108.810 53.425 109.270 53.655 ;
        RECT 72.570 49.320 72.940 50.435 ;
        RECT 60.660 47.775 61.120 47.805 ;
        RECT 68.760 47.775 69.220 47.805 ;
        RECT 71.460 47.775 71.920 47.805 ;
        RECT 60.400 47.375 61.400 47.775 ;
        RECT 68.500 47.375 69.500 47.775 ;
        RECT 71.200 47.375 72.200 47.775 ;
        RECT 62.575 45.600 63.575 45.630 ;
        RECT 66.250 45.600 67.250 45.630 ;
        RECT 60.400 45.150 61.400 45.600 ;
        RECT 60.660 45.140 61.120 45.150 ;
        RECT 59.640 42.545 60.010 43.650 ;
        RECT 60.380 39.925 60.610 44.935 ;
        RECT 61.170 39.925 61.400 44.935 ;
        RECT 62.575 44.570 64.500 45.600 ;
        RECT 61.770 43.600 62.140 43.650 ;
        RECT 61.770 42.545 62.875 43.600 ;
        RECT 57.960 36.140 58.420 36.370 ;
        RECT 57.680 35.925 57.910 35.935 ;
        RECT 58.470 35.925 58.700 35.935 ;
        RECT 56.935 34.945 57.980 35.925 ;
        RECT 58.400 34.945 58.770 35.925 ;
        RECT 60.310 34.945 60.680 39.925 ;
        RECT 61.100 34.945 61.470 39.925 ;
        RECT 61.875 37.850 62.875 42.545 ;
        RECT 63.500 39.500 64.500 44.570 ;
        RECT 65.300 44.570 67.250 45.600 ;
        RECT 68.500 45.150 69.500 45.600 ;
        RECT 71.200 45.150 72.200 45.600 ;
        RECT 68.760 45.140 69.220 45.150 ;
        RECT 71.460 45.140 71.920 45.150 ;
        RECT 65.300 40.245 66.300 44.570 ;
        RECT 67.740 43.600 68.110 43.650 ;
        RECT 67.025 42.545 68.110 43.600 ;
        RECT 63.500 38.500 66.330 39.500 ;
        RECT 67.025 37.850 68.025 42.545 ;
        RECT 68.480 39.925 68.710 44.935 ;
        RECT 69.270 39.925 69.500 44.935 ;
        RECT 69.870 42.545 70.240 43.650 ;
        RECT 70.440 42.545 70.810 43.650 ;
        RECT 71.180 39.925 71.410 44.935 ;
        RECT 71.970 39.925 72.200 44.935 ;
        RECT 72.570 42.545 72.940 43.650 ;
        RECT 61.875 36.850 68.025 37.850 ;
        RECT 63.360 36.140 63.820 36.370 ;
        RECT 66.060 36.140 66.520 36.370 ;
        RECT 63.080 35.925 63.310 35.935 ;
        RECT 63.870 35.925 64.100 35.935 ;
        RECT 65.780 35.925 66.010 35.935 ;
        RECT 66.570 35.925 66.800 35.935 ;
        RECT 62.335 34.945 63.380 35.925 ;
        RECT 63.800 34.945 64.170 35.925 ;
        RECT 65.035 34.945 66.080 35.925 ;
        RECT 66.500 34.945 66.870 35.925 ;
        RECT 68.410 34.945 68.780 39.925 ;
        RECT 69.200 34.945 69.570 39.925 ;
        RECT 71.110 34.945 71.480 39.925 ;
        RECT 71.900 34.945 72.270 39.925 ;
        RECT 57.680 34.935 57.910 34.945 ;
        RECT 58.470 34.935 58.700 34.945 ;
        RECT 60.380 34.935 60.610 34.945 ;
        RECT 61.170 34.935 61.400 34.945 ;
        RECT 63.080 34.935 63.310 34.945 ;
        RECT 63.870 34.935 64.100 34.945 ;
        RECT 65.780 34.935 66.010 34.945 ;
        RECT 66.570 34.935 66.800 34.945 ;
        RECT 68.480 34.935 68.710 34.945 ;
        RECT 69.270 34.935 69.500 34.945 ;
        RECT 71.180 34.935 71.410 34.945 ;
        RECT 71.970 34.935 72.200 34.945 ;
        RECT 57.425 34.275 58.460 34.750 ;
        RECT 60.660 34.500 61.120 34.730 ;
        RECT 62.825 34.275 63.860 34.750 ;
        RECT 65.525 34.275 66.560 34.750 ;
        RECT 68.760 34.500 69.220 34.730 ;
        RECT 71.460 34.500 71.920 34.730 ;
        RECT 78.175 33.900 79.175 51.250 ;
        RECT 80.180 50.430 81.295 50.485 ;
        RECT 80.150 49.315 81.325 50.430 ;
        RECT 85.065 49.320 85.435 50.435 ;
        RECT 78.145 32.900 79.205 33.900 ;
        RECT 57.420 32.030 58.460 32.525 ;
        RECT 60.660 32.050 61.120 32.280 ;
        RECT 62.820 32.030 63.860 32.525 ;
        RECT 65.520 32.030 66.560 32.525 ;
        RECT 68.760 32.050 69.220 32.280 ;
        RECT 71.460 32.050 71.920 32.280 ;
        RECT 57.680 31.880 57.910 31.890 ;
        RECT 58.470 31.880 58.700 31.890 ;
        RECT 60.380 31.880 60.610 31.890 ;
        RECT 61.170 31.880 61.400 31.890 ;
        RECT 63.080 31.880 63.310 31.890 ;
        RECT 63.870 31.880 64.100 31.890 ;
        RECT 65.780 31.880 66.010 31.890 ;
        RECT 66.570 31.880 66.800 31.890 ;
        RECT 68.480 31.880 68.710 31.890 ;
        RECT 69.270 31.880 69.500 31.890 ;
        RECT 71.180 31.880 71.410 31.890 ;
        RECT 71.970 31.880 72.200 31.890 ;
        RECT 56.935 31.250 57.980 31.880 ;
        RECT 58.400 31.250 58.770 31.880 ;
        RECT 57.680 31.240 57.910 31.250 ;
        RECT 58.470 31.240 58.700 31.250 ;
        RECT 57.960 30.850 58.420 31.080 ;
        RECT 60.310 28.700 60.680 31.880 ;
        RECT 61.100 28.700 61.470 31.880 ;
        RECT 62.335 31.250 63.380 31.880 ;
        RECT 63.800 31.250 64.170 31.880 ;
        RECT 65.035 31.250 66.080 31.880 ;
        RECT 66.500 31.250 66.870 31.880 ;
        RECT 63.080 31.240 63.310 31.250 ;
        RECT 63.870 31.240 64.100 31.250 ;
        RECT 65.780 31.240 66.010 31.250 ;
        RECT 66.570 31.240 66.800 31.250 ;
        RECT 63.360 30.850 63.820 31.080 ;
        RECT 66.060 30.850 66.520 31.080 ;
        RECT 68.410 28.700 68.780 31.880 ;
        RECT 69.200 28.700 69.570 31.880 ;
        RECT 71.110 28.700 71.480 31.880 ;
        RECT 71.900 28.700 72.270 31.880 ;
        RECT 54.725 26.740 55.900 27.855 ;
        RECT 59.640 26.745 60.010 27.860 ;
        RECT 52.720 10.325 53.780 11.325 ;
        RECT 52.750 10.295 53.750 10.325 ;
        RECT 31.995 9.455 33.035 9.950 ;
        RECT 35.235 9.475 35.695 9.705 ;
        RECT 37.395 9.455 38.435 9.950 ;
        RECT 40.095 9.455 41.135 9.950 ;
        RECT 43.335 9.475 43.795 9.705 ;
        RECT 46.035 9.475 46.495 9.705 ;
        RECT 32.255 9.305 32.485 9.315 ;
        RECT 33.045 9.305 33.275 9.315 ;
        RECT 34.955 9.305 35.185 9.315 ;
        RECT 35.745 9.305 35.975 9.315 ;
        RECT 37.655 9.305 37.885 9.315 ;
        RECT 38.445 9.305 38.675 9.315 ;
        RECT 40.355 9.305 40.585 9.315 ;
        RECT 41.145 9.305 41.375 9.315 ;
        RECT 43.055 9.305 43.285 9.315 ;
        RECT 43.845 9.305 44.075 9.315 ;
        RECT 45.755 9.305 45.985 9.315 ;
        RECT 46.545 9.305 46.775 9.315 ;
        RECT 31.510 8.675 32.555 9.305 ;
        RECT 32.975 8.675 33.345 9.305 ;
        RECT 32.255 8.665 32.485 8.675 ;
        RECT 33.045 8.665 33.275 8.675 ;
        RECT 32.535 8.275 32.995 8.505 ;
        RECT 34.885 6.125 35.255 9.305 ;
        RECT 35.675 6.125 36.045 9.305 ;
        RECT 36.910 8.675 37.955 9.305 ;
        RECT 38.375 8.675 38.745 9.305 ;
        RECT 39.610 8.675 40.655 9.305 ;
        RECT 41.075 8.675 41.445 9.305 ;
        RECT 37.655 8.665 37.885 8.675 ;
        RECT 38.445 8.665 38.675 8.675 ;
        RECT 40.355 8.665 40.585 8.675 ;
        RECT 41.145 8.665 41.375 8.675 ;
        RECT 37.935 8.275 38.395 8.505 ;
        RECT 40.635 8.275 41.095 8.505 ;
        RECT 42.985 6.125 43.355 9.305 ;
        RECT 43.775 6.125 44.145 9.305 ;
        RECT 45.685 6.125 46.055 9.305 ;
        RECT 46.475 6.125 46.845 9.305 ;
        RECT 29.285 4.170 30.485 5.285 ;
        RECT 34.215 4.170 34.585 5.285 ;
        RECT 29.330 4.140 30.445 4.170 ;
        RECT 34.955 2.815 35.185 6.125 ;
        RECT 35.745 2.815 35.975 6.125 ;
        RECT 36.345 4.170 36.715 5.285 ;
        RECT 42.315 4.170 42.685 5.285 ;
        RECT 43.055 2.815 43.285 6.125 ;
        RECT 43.845 2.815 44.075 6.125 ;
        RECT 44.445 4.170 44.815 5.285 ;
        RECT 45.015 4.170 45.385 5.285 ;
        RECT 45.755 2.815 45.985 6.125 ;
        RECT 46.545 2.815 46.775 6.125 ;
        RECT 47.145 4.170 47.515 5.285 ;
        RECT 48.515 4.140 49.630 9.855 ;
        RECT 54.755 5.285 55.870 26.740 ;
        RECT 60.380 25.390 60.610 28.700 ;
        RECT 61.170 25.390 61.400 28.700 ;
        RECT 61.770 26.745 62.140 27.860 ;
        RECT 67.740 26.745 68.110 27.860 ;
        RECT 68.480 25.390 68.710 28.700 ;
        RECT 69.270 25.390 69.500 28.700 ;
        RECT 69.870 26.745 70.240 27.860 ;
        RECT 70.440 26.745 70.810 27.860 ;
        RECT 71.180 25.390 71.410 28.700 ;
        RECT 71.970 25.390 72.200 28.700 ;
        RECT 72.570 26.745 72.940 27.860 ;
        RECT 73.935 26.745 75.110 27.860 ;
        RECT 60.660 25.200 61.120 25.230 ;
        RECT 68.760 25.200 69.220 25.230 ;
        RECT 71.460 25.200 71.920 25.230 ;
        RECT 60.400 24.800 61.400 25.200 ;
        RECT 68.500 24.800 69.500 25.200 ;
        RECT 71.200 24.800 72.200 25.200 ;
        RECT 73.965 23.770 75.080 26.745 ;
        RECT 62.575 23.025 63.575 23.055 ;
        RECT 66.250 23.025 67.250 23.055 ;
        RECT 60.400 22.575 61.400 23.025 ;
        RECT 60.660 22.565 61.120 22.575 ;
        RECT 59.640 19.970 60.010 21.075 ;
        RECT 60.380 17.350 60.610 22.360 ;
        RECT 61.170 17.350 61.400 22.360 ;
        RECT 62.575 21.995 64.500 23.025 ;
        RECT 61.770 21.025 62.140 21.075 ;
        RECT 61.770 19.970 62.875 21.025 ;
        RECT 57.960 13.565 58.420 13.795 ;
        RECT 57.680 13.350 57.910 13.360 ;
        RECT 58.470 13.350 58.700 13.360 ;
        RECT 56.935 12.370 57.980 13.350 ;
        RECT 58.400 12.370 58.770 13.350 ;
        RECT 60.310 12.370 60.680 17.350 ;
        RECT 61.100 12.370 61.470 17.350 ;
        RECT 61.875 15.275 62.875 19.970 ;
        RECT 63.500 16.925 64.500 21.995 ;
        RECT 65.300 21.995 67.250 23.025 ;
        RECT 68.500 22.575 69.500 23.025 ;
        RECT 71.200 22.575 72.200 23.025 ;
        RECT 68.760 22.565 69.220 22.575 ;
        RECT 71.460 22.565 71.920 22.575 ;
        RECT 65.300 17.670 66.300 21.995 ;
        RECT 67.740 21.025 68.110 21.075 ;
        RECT 67.025 19.970 68.110 21.025 ;
        RECT 63.500 15.925 66.330 16.925 ;
        RECT 67.025 15.275 68.025 19.970 ;
        RECT 68.480 17.350 68.710 22.360 ;
        RECT 69.270 17.350 69.500 22.360 ;
        RECT 69.870 19.970 70.240 21.075 ;
        RECT 70.440 19.970 70.810 21.075 ;
        RECT 71.180 17.350 71.410 22.360 ;
        RECT 71.970 17.350 72.200 22.360 ;
        RECT 74.280 21.115 74.730 23.425 ;
        RECT 72.570 19.970 72.940 21.075 ;
        RECT 61.875 14.275 68.025 15.275 ;
        RECT 63.360 13.565 63.820 13.795 ;
        RECT 66.060 13.565 66.520 13.795 ;
        RECT 63.080 13.350 63.310 13.360 ;
        RECT 63.870 13.350 64.100 13.360 ;
        RECT 65.780 13.350 66.010 13.360 ;
        RECT 66.570 13.350 66.800 13.360 ;
        RECT 62.335 12.370 63.380 13.350 ;
        RECT 63.800 12.370 64.170 13.350 ;
        RECT 65.035 12.370 66.080 13.350 ;
        RECT 66.500 12.370 66.870 13.350 ;
        RECT 68.410 12.370 68.780 17.350 ;
        RECT 69.200 12.370 69.570 17.350 ;
        RECT 71.110 12.370 71.480 17.350 ;
        RECT 71.900 12.370 72.270 17.350 ;
        RECT 57.680 12.360 57.910 12.370 ;
        RECT 58.470 12.360 58.700 12.370 ;
        RECT 60.380 12.360 60.610 12.370 ;
        RECT 61.170 12.360 61.400 12.370 ;
        RECT 63.080 12.360 63.310 12.370 ;
        RECT 63.870 12.360 64.100 12.370 ;
        RECT 65.780 12.360 66.010 12.370 ;
        RECT 66.570 12.360 66.800 12.370 ;
        RECT 68.480 12.360 68.710 12.370 ;
        RECT 69.270 12.360 69.500 12.370 ;
        RECT 71.180 12.360 71.410 12.370 ;
        RECT 71.970 12.360 72.200 12.370 ;
        RECT 57.425 11.700 58.460 12.175 ;
        RECT 60.660 11.925 61.120 12.155 ;
        RECT 62.825 11.700 63.860 12.175 ;
        RECT 65.525 11.700 66.560 12.175 ;
        RECT 68.760 11.925 69.220 12.155 ;
        RECT 71.460 11.925 71.920 12.155 ;
        RECT 74.280 10.205 74.730 12.515 ;
        RECT 78.175 11.325 79.175 32.900 ;
        RECT 80.180 27.855 81.295 49.315 ;
        RECT 85.805 47.965 86.035 51.275 ;
        RECT 86.595 47.965 86.825 51.275 ;
        RECT 87.195 49.320 87.565 50.435 ;
        RECT 93.165 49.320 93.535 50.435 ;
        RECT 93.905 47.965 94.135 51.275 ;
        RECT 94.695 47.965 94.925 51.275 ;
        RECT 95.295 49.320 95.665 50.435 ;
        RECT 95.865 49.320 96.235 50.435 ;
        RECT 96.605 47.965 96.835 51.275 ;
        RECT 97.395 47.965 97.625 51.275 ;
        RECT 103.600 51.250 106.650 52.250 ;
        RECT 111.160 51.275 111.530 54.455 ;
        RECT 111.950 51.275 112.320 54.455 ;
        RECT 113.185 53.825 114.230 54.455 ;
        RECT 114.650 53.825 115.020 54.455 ;
        RECT 115.885 53.825 116.930 54.455 ;
        RECT 117.350 53.825 117.720 54.455 ;
        RECT 113.930 53.815 114.160 53.825 ;
        RECT 114.720 53.815 114.950 53.825 ;
        RECT 116.630 53.815 116.860 53.825 ;
        RECT 117.420 53.815 117.650 53.825 ;
        RECT 114.210 53.425 114.670 53.655 ;
        RECT 116.910 53.425 117.370 53.655 ;
        RECT 119.260 51.275 119.630 54.455 ;
        RECT 120.050 51.275 120.420 54.455 ;
        RECT 121.960 51.275 122.330 54.455 ;
        RECT 122.750 51.275 123.120 54.455 ;
        RECT 131.075 52.250 132.075 55.405 ;
        RECT 133.695 54.605 134.735 55.100 ;
        RECT 136.935 54.625 137.395 54.855 ;
        RECT 139.095 54.605 140.135 55.100 ;
        RECT 141.795 54.605 142.835 55.100 ;
        RECT 145.035 54.625 145.495 54.855 ;
        RECT 147.735 54.625 148.195 54.855 ;
        RECT 133.955 54.455 134.185 54.465 ;
        RECT 134.745 54.455 134.975 54.465 ;
        RECT 136.655 54.455 136.885 54.465 ;
        RECT 137.445 54.455 137.675 54.465 ;
        RECT 139.355 54.455 139.585 54.465 ;
        RECT 140.145 54.455 140.375 54.465 ;
        RECT 142.055 54.455 142.285 54.465 ;
        RECT 142.845 54.455 143.075 54.465 ;
        RECT 144.755 54.455 144.985 54.465 ;
        RECT 145.545 54.455 145.775 54.465 ;
        RECT 147.455 54.455 147.685 54.465 ;
        RECT 148.245 54.455 148.475 54.465 ;
        RECT 133.210 53.825 134.255 54.455 ;
        RECT 134.675 53.825 135.045 54.455 ;
        RECT 133.955 53.815 134.185 53.825 ;
        RECT 134.745 53.815 134.975 53.825 ;
        RECT 134.235 53.425 134.695 53.655 ;
        RECT 97.995 49.320 98.365 50.435 ;
        RECT 86.085 47.775 86.545 47.805 ;
        RECT 94.185 47.775 94.645 47.805 ;
        RECT 96.885 47.775 97.345 47.805 ;
        RECT 85.825 47.375 86.825 47.775 ;
        RECT 93.925 47.375 94.925 47.775 ;
        RECT 96.625 47.375 97.625 47.775 ;
        RECT 88.000 45.600 89.000 45.630 ;
        RECT 91.675 45.600 92.675 45.630 ;
        RECT 85.825 45.150 86.825 45.600 ;
        RECT 86.085 45.140 86.545 45.150 ;
        RECT 85.065 42.545 85.435 43.650 ;
        RECT 85.805 39.925 86.035 44.935 ;
        RECT 86.595 39.925 86.825 44.935 ;
        RECT 88.000 44.570 89.925 45.600 ;
        RECT 87.195 43.600 87.565 43.650 ;
        RECT 87.195 42.545 88.300 43.600 ;
        RECT 83.385 36.140 83.845 36.370 ;
        RECT 83.105 35.925 83.335 35.935 ;
        RECT 83.895 35.925 84.125 35.935 ;
        RECT 82.360 34.945 83.405 35.925 ;
        RECT 83.825 34.945 84.195 35.925 ;
        RECT 85.735 34.945 86.105 39.925 ;
        RECT 86.525 34.945 86.895 39.925 ;
        RECT 87.300 37.850 88.300 42.545 ;
        RECT 88.925 39.500 89.925 44.570 ;
        RECT 90.725 44.570 92.675 45.600 ;
        RECT 93.925 45.150 94.925 45.600 ;
        RECT 96.625 45.150 97.625 45.600 ;
        RECT 94.185 45.140 94.645 45.150 ;
        RECT 96.885 45.140 97.345 45.150 ;
        RECT 90.725 40.245 91.725 44.570 ;
        RECT 93.165 43.600 93.535 43.650 ;
        RECT 92.450 42.545 93.535 43.600 ;
        RECT 88.925 38.500 91.755 39.500 ;
        RECT 92.450 37.850 93.450 42.545 ;
        RECT 93.905 39.925 94.135 44.935 ;
        RECT 94.695 39.925 94.925 44.935 ;
        RECT 95.295 42.545 95.665 43.650 ;
        RECT 95.865 42.545 96.235 43.650 ;
        RECT 96.605 39.925 96.835 44.935 ;
        RECT 97.395 39.925 97.625 44.935 ;
        RECT 97.995 42.545 98.365 43.650 ;
        RECT 87.300 36.850 93.450 37.850 ;
        RECT 88.785 36.140 89.245 36.370 ;
        RECT 91.485 36.140 91.945 36.370 ;
        RECT 88.505 35.925 88.735 35.935 ;
        RECT 89.295 35.925 89.525 35.935 ;
        RECT 91.205 35.925 91.435 35.935 ;
        RECT 91.995 35.925 92.225 35.935 ;
        RECT 87.760 34.945 88.805 35.925 ;
        RECT 89.225 34.945 89.595 35.925 ;
        RECT 90.460 34.945 91.505 35.925 ;
        RECT 91.925 34.945 92.295 35.925 ;
        RECT 93.835 34.945 94.205 39.925 ;
        RECT 94.625 34.945 94.995 39.925 ;
        RECT 96.535 34.945 96.905 39.925 ;
        RECT 97.325 34.945 97.695 39.925 ;
        RECT 83.105 34.935 83.335 34.945 ;
        RECT 83.895 34.935 84.125 34.945 ;
        RECT 85.805 34.935 86.035 34.945 ;
        RECT 86.595 34.935 86.825 34.945 ;
        RECT 88.505 34.935 88.735 34.945 ;
        RECT 89.295 34.935 89.525 34.945 ;
        RECT 91.205 34.935 91.435 34.945 ;
        RECT 91.995 34.935 92.225 34.945 ;
        RECT 93.905 34.935 94.135 34.945 ;
        RECT 94.695 34.935 94.925 34.945 ;
        RECT 96.605 34.935 96.835 34.945 ;
        RECT 97.395 34.935 97.625 34.945 ;
        RECT 82.850 34.275 83.885 34.750 ;
        RECT 86.085 34.500 86.545 34.730 ;
        RECT 88.250 34.275 89.285 34.750 ;
        RECT 90.950 34.275 91.985 34.750 ;
        RECT 94.185 34.500 94.645 34.730 ;
        RECT 96.885 34.500 97.345 34.730 ;
        RECT 103.600 33.900 104.600 51.250 ;
        RECT 105.605 50.430 106.720 50.485 ;
        RECT 105.575 49.315 106.750 50.430 ;
        RECT 110.490 49.320 110.860 50.435 ;
        RECT 103.570 32.900 104.630 33.900 ;
        RECT 82.845 32.030 83.885 32.525 ;
        RECT 86.085 32.050 86.545 32.280 ;
        RECT 88.245 32.030 89.285 32.525 ;
        RECT 90.945 32.030 91.985 32.525 ;
        RECT 94.185 32.050 94.645 32.280 ;
        RECT 96.885 32.050 97.345 32.280 ;
        RECT 83.105 31.880 83.335 31.890 ;
        RECT 83.895 31.880 84.125 31.890 ;
        RECT 85.805 31.880 86.035 31.890 ;
        RECT 86.595 31.880 86.825 31.890 ;
        RECT 88.505 31.880 88.735 31.890 ;
        RECT 89.295 31.880 89.525 31.890 ;
        RECT 91.205 31.880 91.435 31.890 ;
        RECT 91.995 31.880 92.225 31.890 ;
        RECT 93.905 31.880 94.135 31.890 ;
        RECT 94.695 31.880 94.925 31.890 ;
        RECT 96.605 31.880 96.835 31.890 ;
        RECT 97.395 31.880 97.625 31.890 ;
        RECT 82.360 31.250 83.405 31.880 ;
        RECT 83.825 31.250 84.195 31.880 ;
        RECT 83.105 31.240 83.335 31.250 ;
        RECT 83.895 31.240 84.125 31.250 ;
        RECT 83.385 30.850 83.845 31.080 ;
        RECT 85.735 28.700 86.105 31.880 ;
        RECT 86.525 28.700 86.895 31.880 ;
        RECT 87.760 31.250 88.805 31.880 ;
        RECT 89.225 31.250 89.595 31.880 ;
        RECT 90.460 31.250 91.505 31.880 ;
        RECT 91.925 31.250 92.295 31.880 ;
        RECT 88.505 31.240 88.735 31.250 ;
        RECT 89.295 31.240 89.525 31.250 ;
        RECT 91.205 31.240 91.435 31.250 ;
        RECT 91.995 31.240 92.225 31.250 ;
        RECT 88.785 30.850 89.245 31.080 ;
        RECT 91.485 30.850 91.945 31.080 ;
        RECT 93.835 28.700 94.205 31.880 ;
        RECT 94.625 28.700 94.995 31.880 ;
        RECT 96.535 28.700 96.905 31.880 ;
        RECT 97.325 28.700 97.695 31.880 ;
        RECT 80.150 26.740 81.325 27.855 ;
        RECT 85.065 26.745 85.435 27.860 ;
        RECT 78.145 10.325 79.205 11.325 ;
        RECT 78.175 10.295 79.175 10.325 ;
        RECT 57.420 9.455 58.460 9.950 ;
        RECT 60.660 9.475 61.120 9.705 ;
        RECT 62.820 9.455 63.860 9.950 ;
        RECT 65.520 9.455 66.560 9.950 ;
        RECT 68.760 9.475 69.220 9.705 ;
        RECT 71.460 9.475 71.920 9.705 ;
        RECT 57.680 9.305 57.910 9.315 ;
        RECT 58.470 9.305 58.700 9.315 ;
        RECT 60.380 9.305 60.610 9.315 ;
        RECT 61.170 9.305 61.400 9.315 ;
        RECT 63.080 9.305 63.310 9.315 ;
        RECT 63.870 9.305 64.100 9.315 ;
        RECT 65.780 9.305 66.010 9.315 ;
        RECT 66.570 9.305 66.800 9.315 ;
        RECT 68.480 9.305 68.710 9.315 ;
        RECT 69.270 9.305 69.500 9.315 ;
        RECT 71.180 9.305 71.410 9.315 ;
        RECT 71.970 9.305 72.200 9.315 ;
        RECT 56.935 8.675 57.980 9.305 ;
        RECT 58.400 8.675 58.770 9.305 ;
        RECT 57.680 8.665 57.910 8.675 ;
        RECT 58.470 8.665 58.700 8.675 ;
        RECT 57.960 8.275 58.420 8.505 ;
        RECT 60.310 6.125 60.680 9.305 ;
        RECT 61.100 6.125 61.470 9.305 ;
        RECT 62.335 8.675 63.380 9.305 ;
        RECT 63.800 8.675 64.170 9.305 ;
        RECT 65.035 8.675 66.080 9.305 ;
        RECT 66.500 8.675 66.870 9.305 ;
        RECT 63.080 8.665 63.310 8.675 ;
        RECT 63.870 8.665 64.100 8.675 ;
        RECT 65.780 8.665 66.010 8.675 ;
        RECT 66.570 8.665 66.800 8.675 ;
        RECT 63.360 8.275 63.820 8.505 ;
        RECT 66.060 8.275 66.520 8.505 ;
        RECT 68.410 6.125 68.780 9.305 ;
        RECT 69.200 6.125 69.570 9.305 ;
        RECT 71.110 6.125 71.480 9.305 ;
        RECT 71.900 6.125 72.270 9.305 ;
        RECT 54.710 4.170 55.910 5.285 ;
        RECT 59.640 4.170 60.010 5.285 ;
        RECT 54.755 4.140 55.870 4.170 ;
        RECT 60.380 2.815 60.610 6.125 ;
        RECT 61.170 2.815 61.400 6.125 ;
        RECT 61.770 4.170 62.140 5.285 ;
        RECT 67.740 4.170 68.110 5.285 ;
        RECT 68.480 2.815 68.710 6.125 ;
        RECT 69.270 2.815 69.500 6.125 ;
        RECT 69.870 4.170 70.240 5.285 ;
        RECT 70.440 4.170 70.810 5.285 ;
        RECT 71.180 2.815 71.410 6.125 ;
        RECT 71.970 2.815 72.200 6.125 ;
        RECT 72.570 4.170 72.940 5.285 ;
        RECT 73.940 4.140 75.055 9.855 ;
        RECT 80.180 5.285 81.295 26.740 ;
        RECT 85.805 25.390 86.035 28.700 ;
        RECT 86.595 25.390 86.825 28.700 ;
        RECT 87.195 26.745 87.565 27.860 ;
        RECT 93.165 26.745 93.535 27.860 ;
        RECT 93.905 25.390 94.135 28.700 ;
        RECT 94.695 25.390 94.925 28.700 ;
        RECT 95.295 26.745 95.665 27.860 ;
        RECT 95.865 26.745 96.235 27.860 ;
        RECT 96.605 25.390 96.835 28.700 ;
        RECT 97.395 25.390 97.625 28.700 ;
        RECT 97.995 26.745 98.365 27.860 ;
        RECT 99.360 26.745 100.535 27.860 ;
        RECT 86.085 25.200 86.545 25.230 ;
        RECT 94.185 25.200 94.645 25.230 ;
        RECT 96.885 25.200 97.345 25.230 ;
        RECT 85.825 24.800 86.825 25.200 ;
        RECT 93.925 24.800 94.925 25.200 ;
        RECT 96.625 24.800 97.625 25.200 ;
        RECT 99.390 23.770 100.505 26.745 ;
        RECT 88.000 23.025 89.000 23.055 ;
        RECT 91.675 23.025 92.675 23.055 ;
        RECT 85.825 22.575 86.825 23.025 ;
        RECT 86.085 22.565 86.545 22.575 ;
        RECT 85.065 19.970 85.435 21.075 ;
        RECT 85.805 17.350 86.035 22.360 ;
        RECT 86.595 17.350 86.825 22.360 ;
        RECT 88.000 21.995 89.925 23.025 ;
        RECT 87.195 21.025 87.565 21.075 ;
        RECT 87.195 19.970 88.300 21.025 ;
        RECT 83.385 13.565 83.845 13.795 ;
        RECT 83.105 13.350 83.335 13.360 ;
        RECT 83.895 13.350 84.125 13.360 ;
        RECT 82.360 12.370 83.405 13.350 ;
        RECT 83.825 12.370 84.195 13.350 ;
        RECT 85.735 12.370 86.105 17.350 ;
        RECT 86.525 12.370 86.895 17.350 ;
        RECT 87.300 15.275 88.300 19.970 ;
        RECT 88.925 16.925 89.925 21.995 ;
        RECT 90.725 21.995 92.675 23.025 ;
        RECT 93.925 22.575 94.925 23.025 ;
        RECT 96.625 22.575 97.625 23.025 ;
        RECT 94.185 22.565 94.645 22.575 ;
        RECT 96.885 22.565 97.345 22.575 ;
        RECT 90.725 17.670 91.725 21.995 ;
        RECT 93.165 21.025 93.535 21.075 ;
        RECT 92.450 19.970 93.535 21.025 ;
        RECT 88.925 15.925 91.755 16.925 ;
        RECT 92.450 15.275 93.450 19.970 ;
        RECT 93.905 17.350 94.135 22.360 ;
        RECT 94.695 17.350 94.925 22.360 ;
        RECT 95.295 19.970 95.665 21.075 ;
        RECT 95.865 19.970 96.235 21.075 ;
        RECT 96.605 17.350 96.835 22.360 ;
        RECT 97.395 17.350 97.625 22.360 ;
        RECT 99.705 21.115 100.155 23.425 ;
        RECT 97.995 19.970 98.365 21.075 ;
        RECT 87.300 14.275 93.450 15.275 ;
        RECT 88.785 13.565 89.245 13.795 ;
        RECT 91.485 13.565 91.945 13.795 ;
        RECT 88.505 13.350 88.735 13.360 ;
        RECT 89.295 13.350 89.525 13.360 ;
        RECT 91.205 13.350 91.435 13.360 ;
        RECT 91.995 13.350 92.225 13.360 ;
        RECT 87.760 12.370 88.805 13.350 ;
        RECT 89.225 12.370 89.595 13.350 ;
        RECT 90.460 12.370 91.505 13.350 ;
        RECT 91.925 12.370 92.295 13.350 ;
        RECT 93.835 12.370 94.205 17.350 ;
        RECT 94.625 12.370 94.995 17.350 ;
        RECT 96.535 12.370 96.905 17.350 ;
        RECT 97.325 12.370 97.695 17.350 ;
        RECT 83.105 12.360 83.335 12.370 ;
        RECT 83.895 12.360 84.125 12.370 ;
        RECT 85.805 12.360 86.035 12.370 ;
        RECT 86.595 12.360 86.825 12.370 ;
        RECT 88.505 12.360 88.735 12.370 ;
        RECT 89.295 12.360 89.525 12.370 ;
        RECT 91.205 12.360 91.435 12.370 ;
        RECT 91.995 12.360 92.225 12.370 ;
        RECT 93.905 12.360 94.135 12.370 ;
        RECT 94.695 12.360 94.925 12.370 ;
        RECT 96.605 12.360 96.835 12.370 ;
        RECT 97.395 12.360 97.625 12.370 ;
        RECT 82.850 11.700 83.885 12.175 ;
        RECT 86.085 11.925 86.545 12.155 ;
        RECT 88.250 11.700 89.285 12.175 ;
        RECT 90.950 11.700 91.985 12.175 ;
        RECT 94.185 11.925 94.645 12.155 ;
        RECT 96.885 11.925 97.345 12.155 ;
        RECT 99.705 10.205 100.155 12.515 ;
        RECT 103.600 11.325 104.600 32.900 ;
        RECT 105.605 27.855 106.720 49.315 ;
        RECT 111.230 47.965 111.460 51.275 ;
        RECT 112.020 47.965 112.250 51.275 ;
        RECT 112.620 49.320 112.990 50.435 ;
        RECT 118.590 49.320 118.960 50.435 ;
        RECT 119.330 47.965 119.560 51.275 ;
        RECT 120.120 47.965 120.350 51.275 ;
        RECT 120.720 49.320 121.090 50.435 ;
        RECT 121.290 49.320 121.660 50.435 ;
        RECT 122.030 47.965 122.260 51.275 ;
        RECT 122.820 47.965 123.050 51.275 ;
        RECT 129.025 51.250 132.075 52.250 ;
        RECT 136.585 51.275 136.955 54.455 ;
        RECT 137.375 51.275 137.745 54.455 ;
        RECT 138.610 53.825 139.655 54.455 ;
        RECT 140.075 53.825 140.445 54.455 ;
        RECT 141.310 53.825 142.355 54.455 ;
        RECT 142.775 53.825 143.145 54.455 ;
        RECT 139.355 53.815 139.585 53.825 ;
        RECT 140.145 53.815 140.375 53.825 ;
        RECT 142.055 53.815 142.285 53.825 ;
        RECT 142.845 53.815 143.075 53.825 ;
        RECT 139.635 53.425 140.095 53.655 ;
        RECT 142.335 53.425 142.795 53.655 ;
        RECT 144.685 51.275 145.055 54.455 ;
        RECT 145.475 51.275 145.845 54.455 ;
        RECT 147.385 51.275 147.755 54.455 ;
        RECT 148.175 51.275 148.545 54.455 ;
        RECT 123.420 49.320 123.790 50.435 ;
        RECT 111.510 47.775 111.970 47.805 ;
        RECT 119.610 47.775 120.070 47.805 ;
        RECT 122.310 47.775 122.770 47.805 ;
        RECT 111.250 47.375 112.250 47.775 ;
        RECT 119.350 47.375 120.350 47.775 ;
        RECT 122.050 47.375 123.050 47.775 ;
        RECT 113.425 45.600 114.425 45.630 ;
        RECT 117.100 45.600 118.100 45.630 ;
        RECT 111.250 45.150 112.250 45.600 ;
        RECT 111.510 45.140 111.970 45.150 ;
        RECT 110.490 42.545 110.860 43.650 ;
        RECT 111.230 39.925 111.460 44.935 ;
        RECT 112.020 39.925 112.250 44.935 ;
        RECT 113.425 44.570 115.350 45.600 ;
        RECT 112.620 43.600 112.990 43.650 ;
        RECT 112.620 42.545 113.725 43.600 ;
        RECT 108.810 36.140 109.270 36.370 ;
        RECT 108.530 35.925 108.760 35.935 ;
        RECT 109.320 35.925 109.550 35.935 ;
        RECT 107.785 34.945 108.830 35.925 ;
        RECT 109.250 34.945 109.620 35.925 ;
        RECT 111.160 34.945 111.530 39.925 ;
        RECT 111.950 34.945 112.320 39.925 ;
        RECT 112.725 37.850 113.725 42.545 ;
        RECT 114.350 39.500 115.350 44.570 ;
        RECT 116.150 44.570 118.100 45.600 ;
        RECT 119.350 45.150 120.350 45.600 ;
        RECT 122.050 45.150 123.050 45.600 ;
        RECT 119.610 45.140 120.070 45.150 ;
        RECT 122.310 45.140 122.770 45.150 ;
        RECT 116.150 40.245 117.150 44.570 ;
        RECT 118.590 43.600 118.960 43.650 ;
        RECT 117.875 42.545 118.960 43.600 ;
        RECT 114.350 38.500 117.180 39.500 ;
        RECT 117.875 37.850 118.875 42.545 ;
        RECT 119.330 39.925 119.560 44.935 ;
        RECT 120.120 39.925 120.350 44.935 ;
        RECT 120.720 42.545 121.090 43.650 ;
        RECT 121.290 42.545 121.660 43.650 ;
        RECT 122.030 39.925 122.260 44.935 ;
        RECT 122.820 39.925 123.050 44.935 ;
        RECT 123.420 42.545 123.790 43.650 ;
        RECT 112.725 36.850 118.875 37.850 ;
        RECT 114.210 36.140 114.670 36.370 ;
        RECT 116.910 36.140 117.370 36.370 ;
        RECT 113.930 35.925 114.160 35.935 ;
        RECT 114.720 35.925 114.950 35.935 ;
        RECT 116.630 35.925 116.860 35.935 ;
        RECT 117.420 35.925 117.650 35.935 ;
        RECT 113.185 34.945 114.230 35.925 ;
        RECT 114.650 34.945 115.020 35.925 ;
        RECT 115.885 34.945 116.930 35.925 ;
        RECT 117.350 34.945 117.720 35.925 ;
        RECT 119.260 34.945 119.630 39.925 ;
        RECT 120.050 34.945 120.420 39.925 ;
        RECT 121.960 34.945 122.330 39.925 ;
        RECT 122.750 34.945 123.120 39.925 ;
        RECT 108.530 34.935 108.760 34.945 ;
        RECT 109.320 34.935 109.550 34.945 ;
        RECT 111.230 34.935 111.460 34.945 ;
        RECT 112.020 34.935 112.250 34.945 ;
        RECT 113.930 34.935 114.160 34.945 ;
        RECT 114.720 34.935 114.950 34.945 ;
        RECT 116.630 34.935 116.860 34.945 ;
        RECT 117.420 34.935 117.650 34.945 ;
        RECT 119.330 34.935 119.560 34.945 ;
        RECT 120.120 34.935 120.350 34.945 ;
        RECT 122.030 34.935 122.260 34.945 ;
        RECT 122.820 34.935 123.050 34.945 ;
        RECT 108.275 34.275 109.310 34.750 ;
        RECT 111.510 34.500 111.970 34.730 ;
        RECT 113.675 34.275 114.710 34.750 ;
        RECT 116.375 34.275 117.410 34.750 ;
        RECT 119.610 34.500 120.070 34.730 ;
        RECT 122.310 34.500 122.770 34.730 ;
        RECT 129.025 33.900 130.025 51.250 ;
        RECT 131.030 50.430 132.145 50.485 ;
        RECT 131.000 49.315 132.175 50.430 ;
        RECT 135.915 49.320 136.285 50.435 ;
        RECT 128.995 32.900 130.055 33.900 ;
        RECT 108.270 32.030 109.310 32.525 ;
        RECT 111.510 32.050 111.970 32.280 ;
        RECT 113.670 32.030 114.710 32.525 ;
        RECT 116.370 32.030 117.410 32.525 ;
        RECT 119.610 32.050 120.070 32.280 ;
        RECT 122.310 32.050 122.770 32.280 ;
        RECT 108.530 31.880 108.760 31.890 ;
        RECT 109.320 31.880 109.550 31.890 ;
        RECT 111.230 31.880 111.460 31.890 ;
        RECT 112.020 31.880 112.250 31.890 ;
        RECT 113.930 31.880 114.160 31.890 ;
        RECT 114.720 31.880 114.950 31.890 ;
        RECT 116.630 31.880 116.860 31.890 ;
        RECT 117.420 31.880 117.650 31.890 ;
        RECT 119.330 31.880 119.560 31.890 ;
        RECT 120.120 31.880 120.350 31.890 ;
        RECT 122.030 31.880 122.260 31.890 ;
        RECT 122.820 31.880 123.050 31.890 ;
        RECT 107.785 31.250 108.830 31.880 ;
        RECT 109.250 31.250 109.620 31.880 ;
        RECT 108.530 31.240 108.760 31.250 ;
        RECT 109.320 31.240 109.550 31.250 ;
        RECT 108.810 30.850 109.270 31.080 ;
        RECT 111.160 28.700 111.530 31.880 ;
        RECT 111.950 28.700 112.320 31.880 ;
        RECT 113.185 31.250 114.230 31.880 ;
        RECT 114.650 31.250 115.020 31.880 ;
        RECT 115.885 31.250 116.930 31.880 ;
        RECT 117.350 31.250 117.720 31.880 ;
        RECT 113.930 31.240 114.160 31.250 ;
        RECT 114.720 31.240 114.950 31.250 ;
        RECT 116.630 31.240 116.860 31.250 ;
        RECT 117.420 31.240 117.650 31.250 ;
        RECT 114.210 30.850 114.670 31.080 ;
        RECT 116.910 30.850 117.370 31.080 ;
        RECT 119.260 28.700 119.630 31.880 ;
        RECT 120.050 28.700 120.420 31.880 ;
        RECT 121.960 28.700 122.330 31.880 ;
        RECT 122.750 28.700 123.120 31.880 ;
        RECT 105.575 26.740 106.750 27.855 ;
        RECT 110.490 26.745 110.860 27.860 ;
        RECT 103.570 10.325 104.630 11.325 ;
        RECT 103.600 10.295 104.600 10.325 ;
        RECT 82.845 9.455 83.885 9.950 ;
        RECT 86.085 9.475 86.545 9.705 ;
        RECT 88.245 9.455 89.285 9.950 ;
        RECT 90.945 9.455 91.985 9.950 ;
        RECT 94.185 9.475 94.645 9.705 ;
        RECT 96.885 9.475 97.345 9.705 ;
        RECT 83.105 9.305 83.335 9.315 ;
        RECT 83.895 9.305 84.125 9.315 ;
        RECT 85.805 9.305 86.035 9.315 ;
        RECT 86.595 9.305 86.825 9.315 ;
        RECT 88.505 9.305 88.735 9.315 ;
        RECT 89.295 9.305 89.525 9.315 ;
        RECT 91.205 9.305 91.435 9.315 ;
        RECT 91.995 9.305 92.225 9.315 ;
        RECT 93.905 9.305 94.135 9.315 ;
        RECT 94.695 9.305 94.925 9.315 ;
        RECT 96.605 9.305 96.835 9.315 ;
        RECT 97.395 9.305 97.625 9.315 ;
        RECT 82.360 8.675 83.405 9.305 ;
        RECT 83.825 8.675 84.195 9.305 ;
        RECT 83.105 8.665 83.335 8.675 ;
        RECT 83.895 8.665 84.125 8.675 ;
        RECT 83.385 8.275 83.845 8.505 ;
        RECT 85.735 6.125 86.105 9.305 ;
        RECT 86.525 6.125 86.895 9.305 ;
        RECT 87.760 8.675 88.805 9.305 ;
        RECT 89.225 8.675 89.595 9.305 ;
        RECT 90.460 8.675 91.505 9.305 ;
        RECT 91.925 8.675 92.295 9.305 ;
        RECT 88.505 8.665 88.735 8.675 ;
        RECT 89.295 8.665 89.525 8.675 ;
        RECT 91.205 8.665 91.435 8.675 ;
        RECT 91.995 8.665 92.225 8.675 ;
        RECT 88.785 8.275 89.245 8.505 ;
        RECT 91.485 8.275 91.945 8.505 ;
        RECT 93.835 6.125 94.205 9.305 ;
        RECT 94.625 6.125 94.995 9.305 ;
        RECT 96.535 6.125 96.905 9.305 ;
        RECT 97.325 6.125 97.695 9.305 ;
        RECT 80.135 4.170 81.335 5.285 ;
        RECT 85.065 4.170 85.435 5.285 ;
        RECT 80.180 4.140 81.295 4.170 ;
        RECT 85.805 2.815 86.035 6.125 ;
        RECT 86.595 2.815 86.825 6.125 ;
        RECT 87.195 4.170 87.565 5.285 ;
        RECT 93.165 4.170 93.535 5.285 ;
        RECT 93.905 2.815 94.135 6.125 ;
        RECT 94.695 2.815 94.925 6.125 ;
        RECT 95.295 4.170 95.665 5.285 ;
        RECT 95.865 4.170 96.235 5.285 ;
        RECT 96.605 2.815 96.835 6.125 ;
        RECT 97.395 2.815 97.625 6.125 ;
        RECT 97.995 4.170 98.365 5.285 ;
        RECT 99.365 4.140 100.480 9.855 ;
        RECT 105.605 5.285 106.720 26.740 ;
        RECT 111.230 25.390 111.460 28.700 ;
        RECT 112.020 25.390 112.250 28.700 ;
        RECT 112.620 26.745 112.990 27.860 ;
        RECT 118.590 26.745 118.960 27.860 ;
        RECT 119.330 25.390 119.560 28.700 ;
        RECT 120.120 25.390 120.350 28.700 ;
        RECT 120.720 26.745 121.090 27.860 ;
        RECT 121.290 26.745 121.660 27.860 ;
        RECT 122.030 25.390 122.260 28.700 ;
        RECT 122.820 25.390 123.050 28.700 ;
        RECT 123.420 26.745 123.790 27.860 ;
        RECT 124.785 26.745 125.960 27.860 ;
        RECT 111.510 25.200 111.970 25.230 ;
        RECT 119.610 25.200 120.070 25.230 ;
        RECT 122.310 25.200 122.770 25.230 ;
        RECT 111.250 24.800 112.250 25.200 ;
        RECT 119.350 24.800 120.350 25.200 ;
        RECT 122.050 24.800 123.050 25.200 ;
        RECT 124.815 23.770 125.930 26.745 ;
        RECT 113.425 23.025 114.425 23.055 ;
        RECT 117.100 23.025 118.100 23.055 ;
        RECT 111.250 22.575 112.250 23.025 ;
        RECT 111.510 22.565 111.970 22.575 ;
        RECT 110.490 19.970 110.860 21.075 ;
        RECT 111.230 17.350 111.460 22.360 ;
        RECT 112.020 17.350 112.250 22.360 ;
        RECT 113.425 21.995 115.350 23.025 ;
        RECT 112.620 21.025 112.990 21.075 ;
        RECT 112.620 19.970 113.725 21.025 ;
        RECT 108.810 13.565 109.270 13.795 ;
        RECT 108.530 13.350 108.760 13.360 ;
        RECT 109.320 13.350 109.550 13.360 ;
        RECT 107.785 12.370 108.830 13.350 ;
        RECT 109.250 12.370 109.620 13.350 ;
        RECT 111.160 12.370 111.530 17.350 ;
        RECT 111.950 12.370 112.320 17.350 ;
        RECT 112.725 15.275 113.725 19.970 ;
        RECT 114.350 16.925 115.350 21.995 ;
        RECT 116.150 21.995 118.100 23.025 ;
        RECT 119.350 22.575 120.350 23.025 ;
        RECT 122.050 22.575 123.050 23.025 ;
        RECT 119.610 22.565 120.070 22.575 ;
        RECT 122.310 22.565 122.770 22.575 ;
        RECT 116.150 17.670 117.150 21.995 ;
        RECT 118.590 21.025 118.960 21.075 ;
        RECT 117.875 19.970 118.960 21.025 ;
        RECT 114.350 15.925 117.180 16.925 ;
        RECT 117.875 15.275 118.875 19.970 ;
        RECT 119.330 17.350 119.560 22.360 ;
        RECT 120.120 17.350 120.350 22.360 ;
        RECT 120.720 19.970 121.090 21.075 ;
        RECT 121.290 19.970 121.660 21.075 ;
        RECT 122.030 17.350 122.260 22.360 ;
        RECT 122.820 17.350 123.050 22.360 ;
        RECT 125.130 21.115 125.580 23.425 ;
        RECT 123.420 19.970 123.790 21.075 ;
        RECT 112.725 14.275 118.875 15.275 ;
        RECT 114.210 13.565 114.670 13.795 ;
        RECT 116.910 13.565 117.370 13.795 ;
        RECT 113.930 13.350 114.160 13.360 ;
        RECT 114.720 13.350 114.950 13.360 ;
        RECT 116.630 13.350 116.860 13.360 ;
        RECT 117.420 13.350 117.650 13.360 ;
        RECT 113.185 12.370 114.230 13.350 ;
        RECT 114.650 12.370 115.020 13.350 ;
        RECT 115.885 12.370 116.930 13.350 ;
        RECT 117.350 12.370 117.720 13.350 ;
        RECT 119.260 12.370 119.630 17.350 ;
        RECT 120.050 12.370 120.420 17.350 ;
        RECT 121.960 12.370 122.330 17.350 ;
        RECT 122.750 12.370 123.120 17.350 ;
        RECT 108.530 12.360 108.760 12.370 ;
        RECT 109.320 12.360 109.550 12.370 ;
        RECT 111.230 12.360 111.460 12.370 ;
        RECT 112.020 12.360 112.250 12.370 ;
        RECT 113.930 12.360 114.160 12.370 ;
        RECT 114.720 12.360 114.950 12.370 ;
        RECT 116.630 12.360 116.860 12.370 ;
        RECT 117.420 12.360 117.650 12.370 ;
        RECT 119.330 12.360 119.560 12.370 ;
        RECT 120.120 12.360 120.350 12.370 ;
        RECT 122.030 12.360 122.260 12.370 ;
        RECT 122.820 12.360 123.050 12.370 ;
        RECT 108.275 11.700 109.310 12.175 ;
        RECT 111.510 11.925 111.970 12.155 ;
        RECT 113.675 11.700 114.710 12.175 ;
        RECT 116.375 11.700 117.410 12.175 ;
        RECT 119.610 11.925 120.070 12.155 ;
        RECT 122.310 11.925 122.770 12.155 ;
        RECT 125.130 10.205 125.580 12.515 ;
        RECT 129.025 11.325 130.025 32.900 ;
        RECT 131.030 27.855 132.145 49.315 ;
        RECT 136.655 47.965 136.885 51.275 ;
        RECT 137.445 47.965 137.675 51.275 ;
        RECT 138.045 49.320 138.415 50.435 ;
        RECT 144.015 49.320 144.385 50.435 ;
        RECT 144.755 47.965 144.985 51.275 ;
        RECT 145.545 47.965 145.775 51.275 ;
        RECT 146.145 49.320 146.515 50.435 ;
        RECT 146.715 49.320 147.085 50.435 ;
        RECT 147.455 47.965 147.685 51.275 ;
        RECT 148.245 47.965 148.475 51.275 ;
        RECT 148.845 49.320 149.215 50.435 ;
        RECT 136.935 47.775 137.395 47.805 ;
        RECT 145.035 47.775 145.495 47.805 ;
        RECT 147.735 47.775 148.195 47.805 ;
        RECT 136.675 47.375 137.675 47.775 ;
        RECT 144.775 47.375 145.775 47.775 ;
        RECT 147.475 47.375 148.475 47.775 ;
        RECT 138.850 45.600 139.850 45.630 ;
        RECT 142.525 45.600 143.525 45.630 ;
        RECT 136.675 45.150 137.675 45.600 ;
        RECT 136.935 45.140 137.395 45.150 ;
        RECT 135.915 42.545 136.285 43.650 ;
        RECT 136.655 39.925 136.885 44.935 ;
        RECT 137.445 39.925 137.675 44.935 ;
        RECT 138.850 44.570 140.775 45.600 ;
        RECT 138.045 43.600 138.415 43.650 ;
        RECT 138.045 42.545 139.150 43.600 ;
        RECT 134.235 36.140 134.695 36.370 ;
        RECT 133.955 35.925 134.185 35.935 ;
        RECT 134.745 35.925 134.975 35.935 ;
        RECT 133.210 34.945 134.255 35.925 ;
        RECT 134.675 34.945 135.045 35.925 ;
        RECT 136.585 34.945 136.955 39.925 ;
        RECT 137.375 34.945 137.745 39.925 ;
        RECT 138.150 37.850 139.150 42.545 ;
        RECT 139.775 39.500 140.775 44.570 ;
        RECT 141.575 44.570 143.525 45.600 ;
        RECT 144.775 45.150 145.775 45.600 ;
        RECT 147.475 45.150 148.475 45.600 ;
        RECT 145.035 45.140 145.495 45.150 ;
        RECT 147.735 45.140 148.195 45.150 ;
        RECT 141.575 40.245 142.575 44.570 ;
        RECT 144.015 43.600 144.385 43.650 ;
        RECT 143.300 42.545 144.385 43.600 ;
        RECT 139.775 38.500 142.605 39.500 ;
        RECT 143.300 37.850 144.300 42.545 ;
        RECT 144.755 39.925 144.985 44.935 ;
        RECT 145.545 39.925 145.775 44.935 ;
        RECT 146.145 42.545 146.515 43.650 ;
        RECT 146.715 42.545 147.085 43.650 ;
        RECT 147.455 39.925 147.685 44.935 ;
        RECT 148.245 39.925 148.475 44.935 ;
        RECT 148.845 42.545 149.215 43.650 ;
        RECT 138.150 36.850 144.300 37.850 ;
        RECT 139.635 36.140 140.095 36.370 ;
        RECT 142.335 36.140 142.795 36.370 ;
        RECT 139.355 35.925 139.585 35.935 ;
        RECT 140.145 35.925 140.375 35.935 ;
        RECT 142.055 35.925 142.285 35.935 ;
        RECT 142.845 35.925 143.075 35.935 ;
        RECT 138.610 34.945 139.655 35.925 ;
        RECT 140.075 34.945 140.445 35.925 ;
        RECT 141.310 34.945 142.355 35.925 ;
        RECT 142.775 34.945 143.145 35.925 ;
        RECT 144.685 34.945 145.055 39.925 ;
        RECT 145.475 34.945 145.845 39.925 ;
        RECT 147.385 34.945 147.755 39.925 ;
        RECT 148.175 34.945 148.545 39.925 ;
        RECT 133.955 34.935 134.185 34.945 ;
        RECT 134.745 34.935 134.975 34.945 ;
        RECT 136.655 34.935 136.885 34.945 ;
        RECT 137.445 34.935 137.675 34.945 ;
        RECT 139.355 34.935 139.585 34.945 ;
        RECT 140.145 34.935 140.375 34.945 ;
        RECT 142.055 34.935 142.285 34.945 ;
        RECT 142.845 34.935 143.075 34.945 ;
        RECT 144.755 34.935 144.985 34.945 ;
        RECT 145.545 34.935 145.775 34.945 ;
        RECT 147.455 34.935 147.685 34.945 ;
        RECT 148.245 34.935 148.475 34.945 ;
        RECT 133.700 34.275 134.735 34.750 ;
        RECT 136.935 34.500 137.395 34.730 ;
        RECT 139.100 34.275 140.135 34.750 ;
        RECT 141.800 34.275 142.835 34.750 ;
        RECT 145.035 34.500 145.495 34.730 ;
        RECT 147.735 34.500 148.195 34.730 ;
        RECT 133.695 32.030 134.735 32.525 ;
        RECT 136.935 32.050 137.395 32.280 ;
        RECT 139.095 32.030 140.135 32.525 ;
        RECT 141.795 32.030 142.835 32.525 ;
        RECT 145.035 32.050 145.495 32.280 ;
        RECT 147.735 32.050 148.195 32.280 ;
        RECT 133.955 31.880 134.185 31.890 ;
        RECT 134.745 31.880 134.975 31.890 ;
        RECT 136.655 31.880 136.885 31.890 ;
        RECT 137.445 31.880 137.675 31.890 ;
        RECT 139.355 31.880 139.585 31.890 ;
        RECT 140.145 31.880 140.375 31.890 ;
        RECT 142.055 31.880 142.285 31.890 ;
        RECT 142.845 31.880 143.075 31.890 ;
        RECT 144.755 31.880 144.985 31.890 ;
        RECT 145.545 31.880 145.775 31.890 ;
        RECT 147.455 31.880 147.685 31.890 ;
        RECT 148.245 31.880 148.475 31.890 ;
        RECT 133.210 31.250 134.255 31.880 ;
        RECT 134.675 31.250 135.045 31.880 ;
        RECT 133.955 31.240 134.185 31.250 ;
        RECT 134.745 31.240 134.975 31.250 ;
        RECT 134.235 30.850 134.695 31.080 ;
        RECT 136.585 28.700 136.955 31.880 ;
        RECT 137.375 28.700 137.745 31.880 ;
        RECT 138.610 31.250 139.655 31.880 ;
        RECT 140.075 31.250 140.445 31.880 ;
        RECT 141.310 31.250 142.355 31.880 ;
        RECT 142.775 31.250 143.145 31.880 ;
        RECT 139.355 31.240 139.585 31.250 ;
        RECT 140.145 31.240 140.375 31.250 ;
        RECT 142.055 31.240 142.285 31.250 ;
        RECT 142.845 31.240 143.075 31.250 ;
        RECT 139.635 30.850 140.095 31.080 ;
        RECT 142.335 30.850 142.795 31.080 ;
        RECT 144.685 28.700 145.055 31.880 ;
        RECT 145.475 28.700 145.845 31.880 ;
        RECT 147.385 28.700 147.755 31.880 ;
        RECT 148.175 28.700 148.545 31.880 ;
        RECT 131.000 26.740 132.175 27.855 ;
        RECT 135.915 26.745 136.285 27.860 ;
        RECT 128.995 10.325 130.055 11.325 ;
        RECT 129.025 10.295 130.025 10.325 ;
        RECT 108.270 9.455 109.310 9.950 ;
        RECT 111.510 9.475 111.970 9.705 ;
        RECT 113.670 9.455 114.710 9.950 ;
        RECT 116.370 9.455 117.410 9.950 ;
        RECT 119.610 9.475 120.070 9.705 ;
        RECT 122.310 9.475 122.770 9.705 ;
        RECT 108.530 9.305 108.760 9.315 ;
        RECT 109.320 9.305 109.550 9.315 ;
        RECT 111.230 9.305 111.460 9.315 ;
        RECT 112.020 9.305 112.250 9.315 ;
        RECT 113.930 9.305 114.160 9.315 ;
        RECT 114.720 9.305 114.950 9.315 ;
        RECT 116.630 9.305 116.860 9.315 ;
        RECT 117.420 9.305 117.650 9.315 ;
        RECT 119.330 9.305 119.560 9.315 ;
        RECT 120.120 9.305 120.350 9.315 ;
        RECT 122.030 9.305 122.260 9.315 ;
        RECT 122.820 9.305 123.050 9.315 ;
        RECT 107.785 8.675 108.830 9.305 ;
        RECT 109.250 8.675 109.620 9.305 ;
        RECT 108.530 8.665 108.760 8.675 ;
        RECT 109.320 8.665 109.550 8.675 ;
        RECT 108.810 8.275 109.270 8.505 ;
        RECT 111.160 6.125 111.530 9.305 ;
        RECT 111.950 6.125 112.320 9.305 ;
        RECT 113.185 8.675 114.230 9.305 ;
        RECT 114.650 8.675 115.020 9.305 ;
        RECT 115.885 8.675 116.930 9.305 ;
        RECT 117.350 8.675 117.720 9.305 ;
        RECT 113.930 8.665 114.160 8.675 ;
        RECT 114.720 8.665 114.950 8.675 ;
        RECT 116.630 8.665 116.860 8.675 ;
        RECT 117.420 8.665 117.650 8.675 ;
        RECT 114.210 8.275 114.670 8.505 ;
        RECT 116.910 8.275 117.370 8.505 ;
        RECT 119.260 6.125 119.630 9.305 ;
        RECT 120.050 6.125 120.420 9.305 ;
        RECT 121.960 6.125 122.330 9.305 ;
        RECT 122.750 6.125 123.120 9.305 ;
        RECT 105.560 4.170 106.760 5.285 ;
        RECT 110.490 4.170 110.860 5.285 ;
        RECT 105.605 4.140 106.720 4.170 ;
        RECT 111.230 2.815 111.460 6.125 ;
        RECT 112.020 2.815 112.250 6.125 ;
        RECT 112.620 4.170 112.990 5.285 ;
        RECT 118.590 4.170 118.960 5.285 ;
        RECT 119.330 2.815 119.560 6.125 ;
        RECT 120.120 2.815 120.350 6.125 ;
        RECT 120.720 4.170 121.090 5.285 ;
        RECT 121.290 4.170 121.660 5.285 ;
        RECT 122.030 2.815 122.260 6.125 ;
        RECT 122.820 2.815 123.050 6.125 ;
        RECT 123.420 4.170 123.790 5.285 ;
        RECT 124.790 4.140 125.905 9.855 ;
        RECT 131.030 5.285 132.145 26.740 ;
        RECT 136.655 25.390 136.885 28.700 ;
        RECT 137.445 25.390 137.675 28.700 ;
        RECT 138.045 26.745 138.415 27.860 ;
        RECT 144.015 26.745 144.385 27.860 ;
        RECT 144.755 25.390 144.985 28.700 ;
        RECT 145.545 25.390 145.775 28.700 ;
        RECT 146.145 26.745 146.515 27.860 ;
        RECT 146.715 26.745 147.085 27.860 ;
        RECT 147.455 25.390 147.685 28.700 ;
        RECT 148.245 25.390 148.475 28.700 ;
        RECT 148.845 26.745 149.215 27.860 ;
        RECT 150.210 26.745 151.385 27.860 ;
        RECT 136.935 25.200 137.395 25.230 ;
        RECT 145.035 25.200 145.495 25.230 ;
        RECT 147.735 25.200 148.195 25.230 ;
        RECT 136.675 24.800 137.675 25.200 ;
        RECT 144.775 24.800 145.775 25.200 ;
        RECT 147.475 24.800 148.475 25.200 ;
        RECT 150.240 23.770 151.355 26.745 ;
        RECT 138.850 23.025 139.850 23.055 ;
        RECT 142.525 23.025 143.525 23.055 ;
        RECT 136.675 22.575 137.675 23.025 ;
        RECT 136.935 22.565 137.395 22.575 ;
        RECT 135.915 19.970 136.285 21.075 ;
        RECT 136.655 17.350 136.885 22.360 ;
        RECT 137.445 17.350 137.675 22.360 ;
        RECT 138.850 21.995 140.775 23.025 ;
        RECT 138.045 21.025 138.415 21.075 ;
        RECT 138.045 19.970 139.150 21.025 ;
        RECT 134.235 13.565 134.695 13.795 ;
        RECT 133.955 13.350 134.185 13.360 ;
        RECT 134.745 13.350 134.975 13.360 ;
        RECT 133.210 12.370 134.255 13.350 ;
        RECT 134.675 12.370 135.045 13.350 ;
        RECT 136.585 12.370 136.955 17.350 ;
        RECT 137.375 12.370 137.745 17.350 ;
        RECT 138.150 15.275 139.150 19.970 ;
        RECT 139.775 16.925 140.775 21.995 ;
        RECT 141.575 21.995 143.525 23.025 ;
        RECT 144.775 22.575 145.775 23.025 ;
        RECT 147.475 22.575 148.475 23.025 ;
        RECT 145.035 22.565 145.495 22.575 ;
        RECT 147.735 22.565 148.195 22.575 ;
        RECT 141.575 17.670 142.575 21.995 ;
        RECT 144.015 21.025 144.385 21.075 ;
        RECT 143.300 19.970 144.385 21.025 ;
        RECT 139.775 15.925 142.605 16.925 ;
        RECT 143.300 15.275 144.300 19.970 ;
        RECT 144.755 17.350 144.985 22.360 ;
        RECT 145.545 17.350 145.775 22.360 ;
        RECT 146.145 19.970 146.515 21.075 ;
        RECT 146.715 19.970 147.085 21.075 ;
        RECT 147.455 17.350 147.685 22.360 ;
        RECT 148.245 17.350 148.475 22.360 ;
        RECT 150.555 21.115 151.005 23.425 ;
        RECT 148.845 19.970 149.215 21.075 ;
        RECT 138.150 14.275 144.300 15.275 ;
        RECT 139.635 13.565 140.095 13.795 ;
        RECT 142.335 13.565 142.795 13.795 ;
        RECT 139.355 13.350 139.585 13.360 ;
        RECT 140.145 13.350 140.375 13.360 ;
        RECT 142.055 13.350 142.285 13.360 ;
        RECT 142.845 13.350 143.075 13.360 ;
        RECT 138.610 12.370 139.655 13.350 ;
        RECT 140.075 12.370 140.445 13.350 ;
        RECT 141.310 12.370 142.355 13.350 ;
        RECT 142.775 12.370 143.145 13.350 ;
        RECT 144.685 12.370 145.055 17.350 ;
        RECT 145.475 12.370 145.845 17.350 ;
        RECT 147.385 12.370 147.755 17.350 ;
        RECT 148.175 12.370 148.545 17.350 ;
        RECT 133.955 12.360 134.185 12.370 ;
        RECT 134.745 12.360 134.975 12.370 ;
        RECT 136.655 12.360 136.885 12.370 ;
        RECT 137.445 12.360 137.675 12.370 ;
        RECT 139.355 12.360 139.585 12.370 ;
        RECT 140.145 12.360 140.375 12.370 ;
        RECT 142.055 12.360 142.285 12.370 ;
        RECT 142.845 12.360 143.075 12.370 ;
        RECT 144.755 12.360 144.985 12.370 ;
        RECT 145.545 12.360 145.775 12.370 ;
        RECT 147.455 12.360 147.685 12.370 ;
        RECT 148.245 12.360 148.475 12.370 ;
        RECT 133.700 11.700 134.735 12.175 ;
        RECT 136.935 11.925 137.395 12.155 ;
        RECT 139.100 11.700 140.135 12.175 ;
        RECT 141.800 11.700 142.835 12.175 ;
        RECT 145.035 11.925 145.495 12.155 ;
        RECT 147.735 11.925 148.195 12.155 ;
        RECT 150.555 10.205 151.005 12.515 ;
        RECT 133.695 9.455 134.735 9.950 ;
        RECT 136.935 9.475 137.395 9.705 ;
        RECT 139.095 9.455 140.135 9.950 ;
        RECT 141.795 9.455 142.835 9.950 ;
        RECT 145.035 9.475 145.495 9.705 ;
        RECT 147.735 9.475 148.195 9.705 ;
        RECT 133.955 9.305 134.185 9.315 ;
        RECT 134.745 9.305 134.975 9.315 ;
        RECT 136.655 9.305 136.885 9.315 ;
        RECT 137.445 9.305 137.675 9.315 ;
        RECT 139.355 9.305 139.585 9.315 ;
        RECT 140.145 9.305 140.375 9.315 ;
        RECT 142.055 9.305 142.285 9.315 ;
        RECT 142.845 9.305 143.075 9.315 ;
        RECT 144.755 9.305 144.985 9.315 ;
        RECT 145.545 9.305 145.775 9.315 ;
        RECT 147.455 9.305 147.685 9.315 ;
        RECT 148.245 9.305 148.475 9.315 ;
        RECT 133.210 8.675 134.255 9.305 ;
        RECT 134.675 8.675 135.045 9.305 ;
        RECT 133.955 8.665 134.185 8.675 ;
        RECT 134.745 8.665 134.975 8.675 ;
        RECT 134.235 8.275 134.695 8.505 ;
        RECT 136.585 6.125 136.955 9.305 ;
        RECT 137.375 6.125 137.745 9.305 ;
        RECT 138.610 8.675 139.655 9.305 ;
        RECT 140.075 8.675 140.445 9.305 ;
        RECT 141.310 8.675 142.355 9.305 ;
        RECT 142.775 8.675 143.145 9.305 ;
        RECT 139.355 8.665 139.585 8.675 ;
        RECT 140.145 8.665 140.375 8.675 ;
        RECT 142.055 8.665 142.285 8.675 ;
        RECT 142.845 8.665 143.075 8.675 ;
        RECT 139.635 8.275 140.095 8.505 ;
        RECT 142.335 8.275 142.795 8.505 ;
        RECT 144.685 6.125 145.055 9.305 ;
        RECT 145.475 6.125 145.845 9.305 ;
        RECT 147.385 6.125 147.755 9.305 ;
        RECT 148.175 6.125 148.545 9.305 ;
        RECT 130.985 4.170 132.185 5.285 ;
        RECT 135.915 4.170 136.285 5.285 ;
        RECT 131.030 4.140 132.145 4.170 ;
        RECT 136.655 2.815 136.885 6.125 ;
        RECT 137.445 2.815 137.675 6.125 ;
        RECT 138.045 4.170 138.415 5.285 ;
        RECT 144.015 4.170 144.385 5.285 ;
        RECT 144.755 2.815 144.985 6.125 ;
        RECT 145.545 2.815 145.775 6.125 ;
        RECT 146.145 4.170 146.515 5.285 ;
        RECT 146.715 4.170 147.085 5.285 ;
        RECT 147.455 2.815 147.685 6.125 ;
        RECT 148.245 2.815 148.475 6.125 ;
        RECT 148.845 4.170 149.215 5.285 ;
        RECT 150.215 4.140 151.330 9.855 ;
        RECT 9.810 2.625 10.270 2.655 ;
        RECT 17.910 2.625 18.370 2.655 ;
        RECT 20.610 2.625 21.070 2.655 ;
        RECT 35.235 2.625 35.695 2.655 ;
        RECT 43.335 2.625 43.795 2.655 ;
        RECT 46.035 2.625 46.495 2.655 ;
        RECT 60.660 2.625 61.120 2.655 ;
        RECT 68.760 2.625 69.220 2.655 ;
        RECT 71.460 2.625 71.920 2.655 ;
        RECT 86.085 2.625 86.545 2.655 ;
        RECT 94.185 2.625 94.645 2.655 ;
        RECT 96.885 2.625 97.345 2.655 ;
        RECT 111.510 2.625 111.970 2.655 ;
        RECT 119.610 2.625 120.070 2.655 ;
        RECT 122.310 2.625 122.770 2.655 ;
        RECT 136.935 2.625 137.395 2.655 ;
        RECT 145.035 2.625 145.495 2.655 ;
        RECT 147.735 2.625 148.195 2.655 ;
        RECT 9.550 2.225 10.550 2.625 ;
        RECT 17.650 2.225 18.650 2.625 ;
        RECT 20.350 2.225 21.350 2.625 ;
        RECT 34.975 2.225 35.975 2.625 ;
        RECT 43.075 2.225 44.075 2.625 ;
        RECT 45.775 2.225 46.775 2.625 ;
        RECT 60.400 2.225 61.400 2.625 ;
        RECT 68.500 2.225 69.500 2.625 ;
        RECT 71.200 2.225 72.200 2.625 ;
        RECT 85.825 2.225 86.825 2.625 ;
        RECT 93.925 2.225 94.925 2.625 ;
        RECT 96.625 2.225 97.625 2.625 ;
        RECT 111.250 2.225 112.250 2.625 ;
        RECT 119.350 2.225 120.350 2.625 ;
        RECT 122.050 2.225 123.050 2.625 ;
        RECT 136.675 2.225 137.675 2.625 ;
        RECT 144.775 2.225 145.775 2.625 ;
        RECT 147.475 2.225 148.475 2.625 ;
      LAYER met2 ;
        RECT 139.800 225.300 140.800 225.345 ;
        RECT 35.170 224.300 36.230 225.300 ;
        RECT 86.020 224.300 87.080 225.300 ;
        RECT 136.870 224.300 140.845 225.300 ;
        RECT 33.170 222.550 34.230 223.550 ;
        RECT 31.170 220.800 32.230 221.800 ;
        RECT 9.745 219.050 10.805 220.050 ;
        RECT 7.730 217.300 8.820 218.300 ;
        RECT 5.800 216.550 6.750 216.570 ;
        RECT 5.745 215.550 6.805 216.550 ;
        RECT 5.800 215.530 6.750 215.550 ;
        RECT 7.775 215.545 8.775 217.300 ;
        RECT 9.775 215.550 10.775 219.050 ;
        RECT 31.200 215.550 32.200 220.800 ;
        RECT 33.200 215.550 34.200 222.550 ;
        RECT 35.200 215.550 36.200 224.300 ;
        RECT 84.020 222.550 85.080 223.550 ;
        RECT 82.020 220.800 83.080 221.800 ;
        RECT 60.595 219.050 61.655 220.050 ;
        RECT 58.580 217.300 59.670 218.300 ;
        RECT 56.650 216.550 57.600 216.570 ;
        RECT 56.595 215.550 57.655 216.550 ;
        RECT 7.800 215.525 8.750 215.545 ;
        RECT 9.800 215.530 10.750 215.550 ;
        RECT 31.225 215.530 32.175 215.550 ;
        RECT 33.225 215.530 34.175 215.550 ;
        RECT 35.225 215.530 36.175 215.550 ;
        RECT 56.650 215.530 57.600 215.550 ;
        RECT 58.625 215.545 59.625 217.300 ;
        RECT 60.625 215.550 61.625 219.050 ;
        RECT 82.050 215.550 83.050 220.800 ;
        RECT 84.050 215.550 85.050 222.550 ;
        RECT 86.050 215.550 87.050 224.300 ;
        RECT 134.900 223.550 135.900 223.595 ;
        RECT 134.870 222.550 135.930 223.550 ;
        RECT 111.445 219.050 112.505 220.050 ;
        RECT 109.430 217.300 110.520 218.300 ;
        RECT 107.500 216.550 108.450 216.570 ;
        RECT 107.445 215.550 108.505 216.550 ;
        RECT 58.650 215.525 59.600 215.545 ;
        RECT 60.650 215.530 61.600 215.550 ;
        RECT 82.075 215.530 83.025 215.550 ;
        RECT 84.075 215.530 85.025 215.550 ;
        RECT 86.075 215.530 87.025 215.550 ;
        RECT 107.500 215.530 108.450 215.550 ;
        RECT 109.475 215.545 110.475 217.300 ;
        RECT 111.475 215.550 112.475 219.050 ;
        RECT 121.425 216.550 122.425 221.845 ;
        RECT 125.075 218.300 126.075 221.845 ;
        RECT 128.775 220.050 129.775 221.845 ;
        RECT 132.900 221.800 133.900 221.845 ;
        RECT 132.870 220.800 133.930 221.800 ;
        RECT 128.745 219.050 129.805 220.050 ;
        RECT 125.045 217.300 126.105 218.300 ;
        RECT 121.395 215.550 122.455 216.550 ;
        RECT 132.900 215.550 133.900 220.800 ;
        RECT 134.900 215.550 135.900 222.550 ;
        RECT 136.900 215.550 137.900 224.300 ;
        RECT 139.800 224.255 140.800 224.300 ;
        RECT 109.500 215.525 110.450 215.545 ;
        RECT 111.500 215.530 112.450 215.550 ;
        RECT 132.925 215.530 133.875 215.550 ;
        RECT 134.925 215.530 135.875 215.550 ;
        RECT 136.925 215.530 137.875 215.550 ;
        RECT 23.545 214.550 24.495 214.570 ;
        RECT 74.395 214.550 75.345 214.570 ;
        RECT 125.245 214.550 126.195 214.570 ;
        RECT 150.550 214.550 151.500 214.570 ;
        RECT 23.525 213.550 151.525 214.550 ;
        RECT 23.545 213.530 24.495 213.550 ;
        RECT 74.395 213.530 75.345 213.550 ;
        RECT 125.245 213.530 126.195 213.550 ;
        RECT 150.550 213.530 151.500 213.550 ;
        RECT 9.575 212.175 10.525 212.195 ;
        RECT 20.375 212.175 21.325 212.195 ;
        RECT 9.550 211.175 12.755 212.175 ;
        RECT 13.530 211.175 14.620 212.175 ;
        RECT 15.370 211.175 18.650 212.175 ;
        RECT 20.350 211.175 21.350 212.175 ;
        RECT 21.795 212.000 32.470 213.000 ;
        RECT 35.000 212.175 35.950 212.195 ;
        RECT 45.800 212.175 46.750 212.195 ;
        RECT 60.425 212.175 61.375 212.195 ;
        RECT 71.225 212.175 72.175 212.195 ;
        RECT 9.575 211.155 10.525 211.175 ;
        RECT 5.995 210.225 7.100 210.270 ;
        RECT 5.965 209.125 12.025 210.225 ;
        RECT 13.575 210.200 14.575 211.175 ;
        RECT 20.375 211.155 21.325 211.175 ;
        RECT 21.795 210.225 22.795 212.000 ;
        RECT 23.520 210.325 24.520 211.220 ;
        RECT 12.650 209.200 14.575 210.200 ;
        RECT 5.965 209.120 11.290 209.125 ;
        RECT 5.995 209.075 7.100 209.120 ;
        RECT 6.050 202.975 7.050 209.075 ;
        RECT 12.650 207.825 13.650 209.200 ;
        RECT 16.175 209.150 22.795 210.225 ;
        RECT 23.490 209.325 24.550 210.325 ;
        RECT 16.175 209.125 22.100 209.150 ;
        RECT 16.890 209.120 19.400 209.125 ;
        RECT 19.590 209.120 22.090 209.125 ;
        RECT 24.870 208.575 25.870 211.525 ;
        RECT 27.145 210.975 29.170 212.000 ;
        RECT 29.645 210.975 30.590 211.500 ;
        RECT 27.145 210.945 28.145 210.975 ;
        RECT 26.245 210.295 27.245 210.340 ;
        RECT 26.215 209.295 27.275 210.295 ;
        RECT 28.665 209.850 29.705 210.325 ;
        RECT 28.665 209.475 29.170 209.850 ;
        RECT 30.015 209.475 30.590 210.975 ;
        RECT 31.470 210.270 32.470 212.000 ;
        RECT 34.975 211.175 38.180 212.175 ;
        RECT 38.955 211.175 40.045 212.175 ;
        RECT 40.795 211.175 44.075 212.175 ;
        RECT 45.775 211.175 46.775 212.175 ;
        RECT 60.400 211.175 63.605 212.175 ;
        RECT 64.380 211.175 65.470 212.175 ;
        RECT 66.220 211.175 69.500 212.175 ;
        RECT 71.200 211.175 72.200 212.175 ;
        RECT 72.645 212.000 83.320 213.000 ;
        RECT 85.850 212.175 86.800 212.195 ;
        RECT 96.650 212.175 97.600 212.195 ;
        RECT 111.275 212.175 112.225 212.195 ;
        RECT 122.075 212.175 123.025 212.195 ;
        RECT 35.000 211.155 35.950 211.175 ;
        RECT 31.420 210.225 32.525 210.270 ;
        RECT 26.245 209.250 27.245 209.295 ;
        RECT 28.170 208.575 29.170 209.475 ;
        RECT 16.175 208.340 17.175 208.385 ;
        RECT 20.370 208.340 21.320 208.360 ;
        RECT 12.630 206.875 13.670 207.825 ;
        RECT 12.650 206.850 13.650 206.875 ;
        RECT 14.405 206.850 15.495 207.850 ;
        RECT 16.175 207.340 21.345 208.340 ;
        RECT 24.870 208.100 29.170 208.575 ;
        RECT 29.550 208.475 30.640 209.475 ;
        RECT 31.390 209.125 37.450 210.225 ;
        RECT 39.000 210.200 40.000 211.175 ;
        RECT 45.800 211.155 46.750 211.175 ;
        RECT 60.425 211.155 61.375 211.175 ;
        RECT 56.845 210.225 57.950 210.270 ;
        RECT 38.075 209.200 40.000 210.200 ;
        RECT 31.390 209.120 36.715 209.125 ;
        RECT 31.420 209.075 32.525 209.120 ;
        RECT 24.870 207.650 29.705 208.100 ;
        RECT 23.020 207.605 29.705 207.650 ;
        RECT 23.020 207.575 29.170 207.605 ;
        RECT 16.175 207.295 17.175 207.340 ;
        RECT 20.370 207.320 21.320 207.340 ;
        RECT 23.020 206.650 25.870 207.575 ;
        RECT 27.145 207.200 28.145 207.230 ;
        RECT 30.015 207.200 30.590 208.475 ;
        RECT 27.145 206.825 29.225 207.200 ;
        RECT 29.645 206.825 30.590 207.200 ;
        RECT 6.050 201.975 7.075 202.975 ;
        RECT 7.550 201.975 8.495 202.500 ;
        RECT 6.570 200.850 7.610 201.325 ;
        RECT 3.950 200.500 4.950 200.505 ;
        RECT 3.920 200.475 4.980 200.500 ;
        RECT 6.570 200.475 7.075 200.850 ;
        RECT 7.920 200.520 8.495 201.975 ;
        RECT 3.875 200.450 7.075 200.475 ;
        RECT 3.875 199.500 7.095 200.450 ;
        RECT 3.875 199.475 7.075 199.500 ;
        RECT 3.950 199.445 4.950 199.475 ;
        RECT 6.570 199.100 7.075 199.475 ;
        RECT 7.500 199.430 8.500 200.520 ;
        RECT 9.460 200.475 9.830 206.500 ;
        RECT 8.825 199.475 9.830 200.475 ;
        RECT 6.570 198.605 7.610 199.100 ;
        RECT 7.920 198.200 8.495 199.430 ;
        RECT 6.075 197.825 7.130 198.200 ;
        RECT 7.550 197.825 8.495 198.200 ;
        RECT 3.905 194.455 5.020 194.460 ;
        RECT 3.875 194.435 5.050 194.455 ;
        RECT 6.075 194.435 7.075 197.825 ;
        RECT 8.830 196.275 9.830 199.475 ;
        RECT 7.630 195.275 9.830 196.275 ;
        RECT 10.250 200.520 10.620 206.500 ;
        RECT 14.450 206.075 15.450 206.105 ;
        RECT 14.450 205.075 17.220 206.075 ;
        RECT 14.450 205.045 15.450 205.075 ;
        RECT 11.475 201.975 12.475 204.425 ;
        RECT 12.950 201.975 13.895 202.500 ;
        RECT 14.175 201.975 15.175 204.425 ;
        RECT 15.650 201.975 16.595 202.500 ;
        RECT 11.970 200.850 13.010 201.325 ;
        RECT 10.250 200.475 11.250 200.520 ;
        RECT 11.970 200.475 12.475 200.850 ;
        RECT 13.320 200.475 13.895 201.975 ;
        RECT 14.670 200.850 15.710 201.325 ;
        RECT 14.670 200.475 15.175 200.850 ;
        RECT 16.020 200.475 16.595 201.975 ;
        RECT 17.560 200.475 17.930 206.500 ;
        RECT 18.350 200.475 18.720 206.500 ;
        RECT 20.260 200.475 20.630 206.500 ;
        RECT 10.250 200.450 12.475 200.475 ;
        RECT 10.250 199.505 12.495 200.450 ;
        RECT 10.250 199.475 12.475 199.505 ;
        RECT 12.855 199.475 15.175 200.475 ;
        RECT 15.600 199.475 17.930 200.475 ;
        RECT 18.305 199.475 19.395 200.475 ;
        RECT 10.250 199.430 11.250 199.475 ;
        RECT 10.250 195.275 10.620 199.430 ;
        RECT 11.970 199.100 12.475 199.475 ;
        RECT 11.970 198.605 13.010 199.100 ;
        RECT 13.320 198.200 13.895 199.475 ;
        RECT 14.670 199.100 15.175 199.475 ;
        RECT 14.670 198.605 15.710 199.100 ;
        RECT 16.020 198.200 16.595 199.475 ;
        RECT 11.475 197.825 12.530 198.200 ;
        RECT 12.950 197.825 13.895 198.200 ;
        RECT 14.175 197.825 15.230 198.200 ;
        RECT 15.650 197.825 16.595 198.200 ;
        RECT 11.475 196.950 12.475 197.825 ;
        RECT 14.175 196.950 15.175 197.825 ;
        RECT 11.475 195.950 15.175 196.950 ;
        RECT 15.750 196.275 16.750 196.320 ;
        RECT 16.930 196.275 17.930 199.475 ;
        RECT 11.475 194.435 12.475 195.950 ;
        RECT 15.750 195.275 17.930 196.275 ;
        RECT 18.350 195.275 18.720 199.475 ;
        RECT 19.625 197.975 20.630 200.475 ;
        RECT 21.050 200.475 21.420 206.500 ;
        RECT 27.145 206.200 29.170 206.825 ;
        RECT 27.145 206.170 28.370 206.200 ;
        RECT 24.820 205.155 25.925 205.200 ;
        RECT 24.775 204.050 25.970 205.155 ;
        RECT 24.790 204.045 25.955 204.050 ;
        RECT 23.425 200.475 24.375 200.500 ;
        RECT 21.050 199.475 26.300 200.475 ;
        RECT 19.605 197.025 20.645 197.975 ;
        RECT 19.625 197.000 20.630 197.025 ;
        RECT 20.260 195.275 20.630 197.000 ;
        RECT 21.050 195.275 21.420 199.475 ;
        RECT 23.425 199.460 24.375 199.475 ;
        RECT 15.750 195.230 16.750 195.275 ;
        RECT 27.370 194.435 28.370 206.170 ;
        RECT 31.475 202.975 32.475 209.075 ;
        RECT 38.075 207.825 39.075 209.200 ;
        RECT 41.600 209.125 62.875 210.225 ;
        RECT 64.425 210.200 65.425 211.175 ;
        RECT 71.225 211.155 72.175 211.175 ;
        RECT 72.645 210.225 73.645 212.000 ;
        RECT 74.370 210.325 75.370 211.220 ;
        RECT 63.500 209.200 65.425 210.200 ;
        RECT 42.315 209.120 44.825 209.125 ;
        RECT 45.015 209.120 62.140 209.125 ;
        RECT 56.845 209.075 57.950 209.120 ;
        RECT 38.055 206.875 39.095 207.825 ;
        RECT 38.075 206.850 39.075 206.875 ;
        RECT 39.830 206.850 40.920 207.850 ;
        RECT 31.475 201.975 32.500 202.975 ;
        RECT 32.975 201.975 33.920 202.500 ;
        RECT 31.995 200.850 33.035 201.325 ;
        RECT 29.375 200.500 30.375 200.505 ;
        RECT 29.345 200.475 30.405 200.500 ;
        RECT 31.995 200.475 32.500 200.850 ;
        RECT 33.345 200.520 33.920 201.975 ;
        RECT 29.300 200.450 32.500 200.475 ;
        RECT 29.300 199.500 32.520 200.450 ;
        RECT 29.300 199.475 32.500 199.500 ;
        RECT 29.375 199.445 30.375 199.475 ;
        RECT 31.995 199.100 32.500 199.475 ;
        RECT 32.925 199.430 33.925 200.520 ;
        RECT 34.885 200.475 35.255 206.500 ;
        RECT 34.250 199.475 35.255 200.475 ;
        RECT 31.995 198.605 33.035 199.100 ;
        RECT 33.345 198.200 33.920 199.430 ;
        RECT 31.500 197.825 32.555 198.200 ;
        RECT 32.975 197.825 33.920 198.200 ;
        RECT 29.330 194.455 30.445 194.460 ;
        RECT 29.300 194.435 30.475 194.455 ;
        RECT 31.500 194.435 32.500 197.825 ;
        RECT 34.255 196.275 35.255 199.475 ;
        RECT 33.055 195.275 35.255 196.275 ;
        RECT 35.675 200.520 36.045 206.500 ;
        RECT 39.875 206.075 40.875 206.105 ;
        RECT 39.875 205.075 42.645 206.075 ;
        RECT 39.875 205.045 40.875 205.075 ;
        RECT 36.900 201.975 37.900 204.425 ;
        RECT 38.375 201.975 39.320 202.500 ;
        RECT 39.600 201.975 40.600 204.425 ;
        RECT 41.075 201.975 42.020 202.500 ;
        RECT 37.395 200.850 38.435 201.325 ;
        RECT 35.675 200.475 36.675 200.520 ;
        RECT 37.395 200.475 37.900 200.850 ;
        RECT 38.745 200.475 39.320 201.975 ;
        RECT 40.095 200.850 41.135 201.325 ;
        RECT 40.095 200.475 40.600 200.850 ;
        RECT 41.445 200.475 42.020 201.975 ;
        RECT 42.985 200.475 43.355 206.500 ;
        RECT 43.775 200.475 44.145 206.500 ;
        RECT 45.685 200.475 46.055 206.500 ;
        RECT 35.675 200.450 37.900 200.475 ;
        RECT 35.675 199.505 37.920 200.450 ;
        RECT 35.675 199.475 37.900 199.505 ;
        RECT 38.280 199.475 40.600 200.475 ;
        RECT 41.025 199.475 43.355 200.475 ;
        RECT 43.730 199.475 44.820 200.475 ;
        RECT 35.675 199.430 36.675 199.475 ;
        RECT 35.675 195.275 36.045 199.430 ;
        RECT 37.395 199.100 37.900 199.475 ;
        RECT 37.395 198.605 38.435 199.100 ;
        RECT 38.745 198.200 39.320 199.475 ;
        RECT 40.095 199.100 40.600 199.475 ;
        RECT 40.095 198.605 41.135 199.100 ;
        RECT 41.445 198.200 42.020 199.475 ;
        RECT 36.900 197.825 37.955 198.200 ;
        RECT 38.375 197.825 39.320 198.200 ;
        RECT 39.600 197.825 40.655 198.200 ;
        RECT 41.075 197.825 42.020 198.200 ;
        RECT 36.900 196.950 37.900 197.825 ;
        RECT 39.600 196.950 40.600 197.825 ;
        RECT 36.900 195.950 40.600 196.950 ;
        RECT 41.175 196.275 42.175 196.320 ;
        RECT 42.355 196.275 43.355 199.475 ;
        RECT 36.900 194.435 37.900 195.950 ;
        RECT 41.175 195.275 43.355 196.275 ;
        RECT 43.775 195.275 44.145 199.475 ;
        RECT 45.050 197.975 46.055 200.475 ;
        RECT 46.475 200.475 46.845 206.500 ;
        RECT 56.900 202.975 57.900 209.075 ;
        RECT 63.500 207.825 64.500 209.200 ;
        RECT 67.025 209.150 73.645 210.225 ;
        RECT 74.340 209.325 75.400 210.325 ;
        RECT 67.025 209.125 72.950 209.150 ;
        RECT 67.740 209.120 70.250 209.125 ;
        RECT 70.440 209.120 72.940 209.125 ;
        RECT 75.720 208.575 76.720 211.525 ;
        RECT 77.995 210.975 80.020 212.000 ;
        RECT 80.495 210.975 81.440 211.500 ;
        RECT 77.995 210.945 78.995 210.975 ;
        RECT 77.095 210.295 78.095 210.340 ;
        RECT 77.065 209.295 78.125 210.295 ;
        RECT 79.515 209.850 80.555 210.325 ;
        RECT 79.515 209.475 80.020 209.850 ;
        RECT 80.865 209.475 81.440 210.975 ;
        RECT 82.320 210.270 83.320 212.000 ;
        RECT 85.825 211.175 89.030 212.175 ;
        RECT 89.805 211.175 90.895 212.175 ;
        RECT 91.645 211.175 94.925 212.175 ;
        RECT 96.625 211.175 97.625 212.175 ;
        RECT 111.250 211.175 114.455 212.175 ;
        RECT 115.230 211.175 116.320 212.175 ;
        RECT 117.070 211.175 120.350 212.175 ;
        RECT 122.050 211.175 123.050 212.175 ;
        RECT 123.495 212.000 134.170 213.000 ;
        RECT 136.700 212.175 137.650 212.195 ;
        RECT 147.500 212.175 148.450 212.195 ;
        RECT 85.850 211.155 86.800 211.175 ;
        RECT 82.270 210.225 83.375 210.270 ;
        RECT 77.095 209.250 78.095 209.295 ;
        RECT 79.020 208.575 80.020 209.475 ;
        RECT 67.025 208.340 68.025 208.385 ;
        RECT 71.220 208.340 72.170 208.360 ;
        RECT 63.480 206.875 64.520 207.825 ;
        RECT 63.500 206.850 64.500 206.875 ;
        RECT 65.255 206.850 66.345 207.850 ;
        RECT 67.025 207.340 72.195 208.340 ;
        RECT 75.720 208.100 80.020 208.575 ;
        RECT 80.400 208.475 81.490 209.475 ;
        RECT 82.240 209.125 88.300 210.225 ;
        RECT 89.850 210.200 90.850 211.175 ;
        RECT 96.650 211.155 97.600 211.175 ;
        RECT 111.275 211.155 112.225 211.175 ;
        RECT 107.695 210.225 108.800 210.270 ;
        RECT 88.925 209.200 90.850 210.200 ;
        RECT 82.240 209.120 87.565 209.125 ;
        RECT 82.270 209.075 83.375 209.120 ;
        RECT 75.720 207.650 80.555 208.100 ;
        RECT 73.870 207.605 80.555 207.650 ;
        RECT 73.870 207.575 80.020 207.605 ;
        RECT 67.025 207.295 68.025 207.340 ;
        RECT 71.220 207.320 72.170 207.340 ;
        RECT 73.870 206.650 76.720 207.575 ;
        RECT 77.995 207.200 78.995 207.230 ;
        RECT 80.865 207.200 81.440 208.475 ;
        RECT 77.995 206.825 80.075 207.200 ;
        RECT 80.495 206.825 81.440 207.200 ;
        RECT 56.900 201.975 57.925 202.975 ;
        RECT 58.400 201.975 59.345 202.500 ;
        RECT 57.420 200.850 58.460 201.325 ;
        RECT 50.725 200.475 51.725 200.505 ;
        RECT 54.800 200.500 55.800 200.505 ;
        RECT 54.770 200.475 55.830 200.500 ;
        RECT 57.420 200.475 57.925 200.850 ;
        RECT 58.770 200.520 59.345 201.975 ;
        RECT 46.475 199.475 51.725 200.475 ;
        RECT 54.725 200.450 57.925 200.475 ;
        RECT 54.725 199.500 57.945 200.450 ;
        RECT 54.725 199.475 57.925 199.500 ;
        RECT 45.030 197.025 46.070 197.975 ;
        RECT 45.050 197.000 46.055 197.025 ;
        RECT 45.685 195.275 46.055 197.000 ;
        RECT 46.475 195.275 46.845 199.475 ;
        RECT 50.725 199.445 51.725 199.475 ;
        RECT 54.800 199.445 55.800 199.475 ;
        RECT 57.420 199.100 57.925 199.475 ;
        RECT 58.350 199.430 59.350 200.520 ;
        RECT 60.310 200.475 60.680 206.500 ;
        RECT 59.675 199.475 60.680 200.475 ;
        RECT 57.420 198.605 58.460 199.100 ;
        RECT 58.770 198.200 59.345 199.430 ;
        RECT 56.925 197.825 57.980 198.200 ;
        RECT 58.400 197.825 59.345 198.200 ;
        RECT 41.175 195.230 42.175 195.275 ;
        RECT 54.755 194.455 55.870 194.460 ;
        RECT 54.725 194.435 55.900 194.455 ;
        RECT 56.925 194.435 57.925 197.825 ;
        RECT 59.680 196.275 60.680 199.475 ;
        RECT 58.480 195.275 60.680 196.275 ;
        RECT 61.100 200.520 61.470 206.500 ;
        RECT 65.300 206.075 66.300 206.105 ;
        RECT 65.300 205.075 68.070 206.075 ;
        RECT 65.300 205.045 66.300 205.075 ;
        RECT 62.325 201.975 63.325 204.425 ;
        RECT 63.800 201.975 64.745 202.500 ;
        RECT 65.025 201.975 66.025 204.425 ;
        RECT 66.500 201.975 67.445 202.500 ;
        RECT 62.820 200.850 63.860 201.325 ;
        RECT 61.100 200.475 62.100 200.520 ;
        RECT 62.820 200.475 63.325 200.850 ;
        RECT 64.170 200.475 64.745 201.975 ;
        RECT 65.520 200.850 66.560 201.325 ;
        RECT 65.520 200.475 66.025 200.850 ;
        RECT 66.870 200.475 67.445 201.975 ;
        RECT 68.410 200.475 68.780 206.500 ;
        RECT 69.200 200.475 69.570 206.500 ;
        RECT 71.110 200.475 71.480 206.500 ;
        RECT 61.100 200.450 63.325 200.475 ;
        RECT 61.100 199.505 63.345 200.450 ;
        RECT 61.100 199.475 63.325 199.505 ;
        RECT 63.705 199.475 66.025 200.475 ;
        RECT 66.450 199.475 68.780 200.475 ;
        RECT 69.155 199.475 70.245 200.475 ;
        RECT 61.100 199.430 62.100 199.475 ;
        RECT 61.100 195.275 61.470 199.430 ;
        RECT 62.820 199.100 63.325 199.475 ;
        RECT 62.820 198.605 63.860 199.100 ;
        RECT 64.170 198.200 64.745 199.475 ;
        RECT 65.520 199.100 66.025 199.475 ;
        RECT 65.520 198.605 66.560 199.100 ;
        RECT 66.870 198.200 67.445 199.475 ;
        RECT 62.325 197.825 63.380 198.200 ;
        RECT 63.800 197.825 64.745 198.200 ;
        RECT 65.025 197.825 66.080 198.200 ;
        RECT 66.500 197.825 67.445 198.200 ;
        RECT 62.325 196.950 63.325 197.825 ;
        RECT 65.025 196.950 66.025 197.825 ;
        RECT 62.325 195.950 66.025 196.950 ;
        RECT 66.600 196.275 67.600 196.320 ;
        RECT 67.780 196.275 68.780 199.475 ;
        RECT 62.325 194.435 63.325 195.950 ;
        RECT 66.600 195.275 68.780 196.275 ;
        RECT 69.200 195.275 69.570 199.475 ;
        RECT 70.475 197.975 71.480 200.475 ;
        RECT 71.900 200.475 72.270 206.500 ;
        RECT 77.995 206.200 80.020 206.825 ;
        RECT 77.995 206.170 79.220 206.200 ;
        RECT 75.670 205.155 76.775 205.200 ;
        RECT 75.625 204.050 76.820 205.155 ;
        RECT 75.640 204.045 76.805 204.050 ;
        RECT 74.275 200.475 75.225 200.500 ;
        RECT 71.900 199.475 77.150 200.475 ;
        RECT 70.455 197.025 71.495 197.975 ;
        RECT 70.475 197.000 71.480 197.025 ;
        RECT 71.110 195.275 71.480 197.000 ;
        RECT 71.900 195.275 72.270 199.475 ;
        RECT 74.275 199.460 75.225 199.475 ;
        RECT 66.600 195.230 67.600 195.275 ;
        RECT 78.220 194.435 79.220 206.170 ;
        RECT 82.325 202.975 83.325 209.075 ;
        RECT 88.925 207.825 89.925 209.200 ;
        RECT 92.450 209.125 113.725 210.225 ;
        RECT 115.275 210.200 116.275 211.175 ;
        RECT 122.075 211.155 123.025 211.175 ;
        RECT 123.495 210.225 124.495 212.000 ;
        RECT 125.220 210.325 126.220 211.220 ;
        RECT 114.350 209.200 116.275 210.200 ;
        RECT 93.165 209.120 95.675 209.125 ;
        RECT 95.865 209.120 112.990 209.125 ;
        RECT 107.695 209.075 108.800 209.120 ;
        RECT 88.905 206.875 89.945 207.825 ;
        RECT 88.925 206.850 89.925 206.875 ;
        RECT 90.680 206.850 91.770 207.850 ;
        RECT 82.325 201.975 83.350 202.975 ;
        RECT 83.825 201.975 84.770 202.500 ;
        RECT 82.845 200.850 83.885 201.325 ;
        RECT 80.225 200.500 81.225 200.505 ;
        RECT 80.195 200.475 81.255 200.500 ;
        RECT 82.845 200.475 83.350 200.850 ;
        RECT 84.195 200.520 84.770 201.975 ;
        RECT 80.150 200.450 83.350 200.475 ;
        RECT 80.150 199.500 83.370 200.450 ;
        RECT 80.150 199.475 83.350 199.500 ;
        RECT 80.225 199.445 81.225 199.475 ;
        RECT 82.845 199.100 83.350 199.475 ;
        RECT 83.775 199.430 84.775 200.520 ;
        RECT 85.735 200.475 86.105 206.500 ;
        RECT 85.100 199.475 86.105 200.475 ;
        RECT 82.845 198.605 83.885 199.100 ;
        RECT 84.195 198.200 84.770 199.430 ;
        RECT 82.350 197.825 83.405 198.200 ;
        RECT 83.825 197.825 84.770 198.200 ;
        RECT 80.180 194.455 81.295 194.460 ;
        RECT 80.150 194.435 81.325 194.455 ;
        RECT 82.350 194.435 83.350 197.825 ;
        RECT 85.105 196.275 86.105 199.475 ;
        RECT 83.905 195.275 86.105 196.275 ;
        RECT 86.525 200.520 86.895 206.500 ;
        RECT 90.725 206.075 91.725 206.105 ;
        RECT 90.725 205.075 93.495 206.075 ;
        RECT 90.725 205.045 91.725 205.075 ;
        RECT 87.750 201.975 88.750 204.425 ;
        RECT 89.225 201.975 90.170 202.500 ;
        RECT 90.450 201.975 91.450 204.425 ;
        RECT 91.925 201.975 92.870 202.500 ;
        RECT 88.245 200.850 89.285 201.325 ;
        RECT 86.525 200.475 87.525 200.520 ;
        RECT 88.245 200.475 88.750 200.850 ;
        RECT 89.595 200.475 90.170 201.975 ;
        RECT 90.945 200.850 91.985 201.325 ;
        RECT 90.945 200.475 91.450 200.850 ;
        RECT 92.295 200.475 92.870 201.975 ;
        RECT 93.835 200.475 94.205 206.500 ;
        RECT 94.625 200.475 94.995 206.500 ;
        RECT 96.535 200.475 96.905 206.500 ;
        RECT 86.525 200.450 88.750 200.475 ;
        RECT 86.525 199.505 88.770 200.450 ;
        RECT 86.525 199.475 88.750 199.505 ;
        RECT 89.130 199.475 91.450 200.475 ;
        RECT 91.875 199.475 94.205 200.475 ;
        RECT 94.580 199.475 95.670 200.475 ;
        RECT 86.525 199.430 87.525 199.475 ;
        RECT 86.525 195.275 86.895 199.430 ;
        RECT 88.245 199.100 88.750 199.475 ;
        RECT 88.245 198.605 89.285 199.100 ;
        RECT 89.595 198.200 90.170 199.475 ;
        RECT 90.945 199.100 91.450 199.475 ;
        RECT 90.945 198.605 91.985 199.100 ;
        RECT 92.295 198.200 92.870 199.475 ;
        RECT 87.750 197.825 88.805 198.200 ;
        RECT 89.225 197.825 90.170 198.200 ;
        RECT 90.450 197.825 91.505 198.200 ;
        RECT 91.925 197.825 92.870 198.200 ;
        RECT 87.750 196.950 88.750 197.825 ;
        RECT 90.450 196.950 91.450 197.825 ;
        RECT 87.750 195.950 91.450 196.950 ;
        RECT 92.025 196.275 93.025 196.320 ;
        RECT 93.205 196.275 94.205 199.475 ;
        RECT 87.750 194.435 88.750 195.950 ;
        RECT 92.025 195.275 94.205 196.275 ;
        RECT 94.625 195.275 94.995 199.475 ;
        RECT 95.900 197.975 96.905 200.475 ;
        RECT 97.325 200.475 97.695 206.500 ;
        RECT 107.750 202.975 108.750 209.075 ;
        RECT 114.350 207.825 115.350 209.200 ;
        RECT 117.875 209.150 124.495 210.225 ;
        RECT 125.190 209.325 126.250 210.325 ;
        RECT 117.875 209.125 123.800 209.150 ;
        RECT 118.590 209.120 121.100 209.125 ;
        RECT 121.290 209.120 123.790 209.125 ;
        RECT 126.570 208.575 127.570 211.525 ;
        RECT 128.845 210.975 130.870 212.000 ;
        RECT 131.345 210.975 132.290 211.500 ;
        RECT 128.845 210.945 129.845 210.975 ;
        RECT 127.945 210.295 128.945 210.340 ;
        RECT 127.915 209.295 128.975 210.295 ;
        RECT 130.365 209.850 131.405 210.325 ;
        RECT 130.365 209.475 130.870 209.850 ;
        RECT 131.715 209.475 132.290 210.975 ;
        RECT 133.170 210.270 134.170 212.000 ;
        RECT 136.675 211.175 139.880 212.175 ;
        RECT 140.655 211.175 141.745 212.175 ;
        RECT 142.495 211.175 145.775 212.175 ;
        RECT 147.475 211.175 148.475 212.175 ;
        RECT 136.700 211.155 137.650 211.175 ;
        RECT 133.120 210.225 134.225 210.270 ;
        RECT 127.945 209.250 128.945 209.295 ;
        RECT 129.870 208.575 130.870 209.475 ;
        RECT 117.875 208.340 118.875 208.385 ;
        RECT 122.070 208.340 123.020 208.360 ;
        RECT 114.330 206.875 115.370 207.825 ;
        RECT 114.350 206.850 115.350 206.875 ;
        RECT 116.105 206.850 117.195 207.850 ;
        RECT 117.875 207.340 123.045 208.340 ;
        RECT 126.570 208.100 130.870 208.575 ;
        RECT 131.250 208.475 132.340 209.475 ;
        RECT 133.090 209.125 139.150 210.225 ;
        RECT 140.700 210.200 141.700 211.175 ;
        RECT 147.500 211.155 148.450 211.175 ;
        RECT 139.775 209.200 141.700 210.200 ;
        RECT 133.090 209.120 138.415 209.125 ;
        RECT 133.120 209.075 134.225 209.120 ;
        RECT 126.570 207.650 131.405 208.100 ;
        RECT 124.720 207.605 131.405 207.650 ;
        RECT 124.720 207.575 130.870 207.605 ;
        RECT 117.875 207.295 118.875 207.340 ;
        RECT 122.070 207.320 123.020 207.340 ;
        RECT 124.720 206.650 127.570 207.575 ;
        RECT 128.845 207.200 129.845 207.230 ;
        RECT 131.715 207.200 132.290 208.475 ;
        RECT 128.845 206.825 130.925 207.200 ;
        RECT 131.345 206.825 132.290 207.200 ;
        RECT 107.750 201.975 108.775 202.975 ;
        RECT 109.250 201.975 110.195 202.500 ;
        RECT 108.270 200.850 109.310 201.325 ;
        RECT 101.575 200.475 102.575 200.505 ;
        RECT 105.650 200.500 106.650 200.505 ;
        RECT 105.620 200.475 106.680 200.500 ;
        RECT 108.270 200.475 108.775 200.850 ;
        RECT 109.620 200.520 110.195 201.975 ;
        RECT 97.325 199.475 102.575 200.475 ;
        RECT 105.575 200.450 108.775 200.475 ;
        RECT 105.575 199.500 108.795 200.450 ;
        RECT 105.575 199.475 108.775 199.500 ;
        RECT 95.880 197.025 96.920 197.975 ;
        RECT 95.900 197.000 96.905 197.025 ;
        RECT 96.535 195.275 96.905 197.000 ;
        RECT 97.325 195.275 97.695 199.475 ;
        RECT 101.575 199.445 102.575 199.475 ;
        RECT 105.650 199.445 106.650 199.475 ;
        RECT 108.270 199.100 108.775 199.475 ;
        RECT 109.200 199.430 110.200 200.520 ;
        RECT 111.160 200.475 111.530 206.500 ;
        RECT 110.525 199.475 111.530 200.475 ;
        RECT 108.270 198.605 109.310 199.100 ;
        RECT 109.620 198.200 110.195 199.430 ;
        RECT 107.775 197.825 108.830 198.200 ;
        RECT 109.250 197.825 110.195 198.200 ;
        RECT 92.025 195.230 93.025 195.275 ;
        RECT 105.605 194.455 106.720 194.460 ;
        RECT 105.575 194.435 106.750 194.455 ;
        RECT 107.775 194.435 108.775 197.825 ;
        RECT 110.530 196.275 111.530 199.475 ;
        RECT 109.330 195.275 111.530 196.275 ;
        RECT 111.950 200.520 112.320 206.500 ;
        RECT 116.150 206.075 117.150 206.105 ;
        RECT 116.150 205.075 118.920 206.075 ;
        RECT 116.150 205.045 117.150 205.075 ;
        RECT 113.175 201.975 114.175 204.425 ;
        RECT 114.650 201.975 115.595 202.500 ;
        RECT 115.875 201.975 116.875 204.425 ;
        RECT 117.350 201.975 118.295 202.500 ;
        RECT 113.670 200.850 114.710 201.325 ;
        RECT 111.950 200.475 112.950 200.520 ;
        RECT 113.670 200.475 114.175 200.850 ;
        RECT 115.020 200.475 115.595 201.975 ;
        RECT 116.370 200.850 117.410 201.325 ;
        RECT 116.370 200.475 116.875 200.850 ;
        RECT 117.720 200.475 118.295 201.975 ;
        RECT 119.260 200.475 119.630 206.500 ;
        RECT 120.050 200.475 120.420 206.500 ;
        RECT 121.960 200.475 122.330 206.500 ;
        RECT 111.950 200.450 114.175 200.475 ;
        RECT 111.950 199.505 114.195 200.450 ;
        RECT 111.950 199.475 114.175 199.505 ;
        RECT 114.555 199.475 116.875 200.475 ;
        RECT 117.300 199.475 119.630 200.475 ;
        RECT 120.005 199.475 121.095 200.475 ;
        RECT 111.950 199.430 112.950 199.475 ;
        RECT 111.950 195.275 112.320 199.430 ;
        RECT 113.670 199.100 114.175 199.475 ;
        RECT 113.670 198.605 114.710 199.100 ;
        RECT 115.020 198.200 115.595 199.475 ;
        RECT 116.370 199.100 116.875 199.475 ;
        RECT 116.370 198.605 117.410 199.100 ;
        RECT 117.720 198.200 118.295 199.475 ;
        RECT 113.175 197.825 114.230 198.200 ;
        RECT 114.650 197.825 115.595 198.200 ;
        RECT 115.875 197.825 116.930 198.200 ;
        RECT 117.350 197.825 118.295 198.200 ;
        RECT 113.175 196.950 114.175 197.825 ;
        RECT 115.875 196.950 116.875 197.825 ;
        RECT 113.175 195.950 116.875 196.950 ;
        RECT 117.450 196.275 118.450 196.320 ;
        RECT 118.630 196.275 119.630 199.475 ;
        RECT 113.175 194.435 114.175 195.950 ;
        RECT 117.450 195.275 119.630 196.275 ;
        RECT 120.050 195.275 120.420 199.475 ;
        RECT 121.325 197.975 122.330 200.475 ;
        RECT 122.750 200.475 123.120 206.500 ;
        RECT 128.845 206.200 130.870 206.825 ;
        RECT 128.845 206.170 130.070 206.200 ;
        RECT 126.520 205.155 127.625 205.200 ;
        RECT 126.475 204.050 127.670 205.155 ;
        RECT 126.490 204.045 127.655 204.050 ;
        RECT 125.125 200.475 126.075 200.500 ;
        RECT 122.750 199.475 128.000 200.475 ;
        RECT 121.305 197.025 122.345 197.975 ;
        RECT 121.325 197.000 122.330 197.025 ;
        RECT 121.960 195.275 122.330 197.000 ;
        RECT 122.750 195.275 123.120 199.475 ;
        RECT 125.125 199.460 126.075 199.475 ;
        RECT 117.450 195.230 118.450 195.275 ;
        RECT 129.070 194.435 130.070 206.170 ;
        RECT 133.175 202.975 134.175 209.075 ;
        RECT 139.775 207.825 140.775 209.200 ;
        RECT 143.300 209.125 149.225 210.225 ;
        RECT 144.015 209.120 146.525 209.125 ;
        RECT 146.715 209.120 149.215 209.125 ;
        RECT 139.755 206.875 140.795 207.825 ;
        RECT 139.775 206.850 140.775 206.875 ;
        RECT 141.530 206.850 142.620 207.850 ;
        RECT 133.175 201.975 134.200 202.975 ;
        RECT 134.675 201.975 135.620 202.500 ;
        RECT 133.695 200.850 134.735 201.325 ;
        RECT 131.075 200.500 132.075 200.505 ;
        RECT 131.045 200.475 132.105 200.500 ;
        RECT 133.695 200.475 134.200 200.850 ;
        RECT 135.045 200.520 135.620 201.975 ;
        RECT 131.000 200.450 134.200 200.475 ;
        RECT 131.000 199.500 134.220 200.450 ;
        RECT 131.000 199.475 134.200 199.500 ;
        RECT 131.075 199.445 132.075 199.475 ;
        RECT 133.695 199.100 134.200 199.475 ;
        RECT 134.625 199.430 135.625 200.520 ;
        RECT 136.585 200.475 136.955 206.500 ;
        RECT 135.950 199.475 136.955 200.475 ;
        RECT 133.695 198.605 134.735 199.100 ;
        RECT 135.045 198.200 135.620 199.430 ;
        RECT 133.200 197.825 134.255 198.200 ;
        RECT 134.675 197.825 135.620 198.200 ;
        RECT 131.030 194.455 132.145 194.460 ;
        RECT 131.000 194.435 132.175 194.455 ;
        RECT 133.200 194.435 134.200 197.825 ;
        RECT 135.955 196.275 136.955 199.475 ;
        RECT 134.755 195.275 136.955 196.275 ;
        RECT 137.375 200.520 137.745 206.500 ;
        RECT 141.575 206.075 142.575 206.105 ;
        RECT 141.575 205.075 144.345 206.075 ;
        RECT 141.575 205.045 142.575 205.075 ;
        RECT 138.600 201.975 139.600 204.425 ;
        RECT 140.075 201.975 141.020 202.500 ;
        RECT 141.300 201.975 142.300 204.425 ;
        RECT 142.775 201.975 143.720 202.500 ;
        RECT 139.095 200.850 140.135 201.325 ;
        RECT 137.375 200.475 138.375 200.520 ;
        RECT 139.095 200.475 139.600 200.850 ;
        RECT 140.445 200.475 141.020 201.975 ;
        RECT 141.795 200.850 142.835 201.325 ;
        RECT 141.795 200.475 142.300 200.850 ;
        RECT 143.145 200.475 143.720 201.975 ;
        RECT 144.685 200.475 145.055 206.500 ;
        RECT 145.475 200.475 145.845 206.500 ;
        RECT 147.385 200.475 147.755 206.500 ;
        RECT 137.375 200.450 139.600 200.475 ;
        RECT 137.375 199.505 139.620 200.450 ;
        RECT 137.375 199.475 139.600 199.505 ;
        RECT 139.980 199.475 142.300 200.475 ;
        RECT 142.725 199.475 145.055 200.475 ;
        RECT 145.430 199.475 146.520 200.475 ;
        RECT 137.375 199.430 138.375 199.475 ;
        RECT 137.375 195.275 137.745 199.430 ;
        RECT 139.095 199.100 139.600 199.475 ;
        RECT 139.095 198.605 140.135 199.100 ;
        RECT 140.445 198.200 141.020 199.475 ;
        RECT 141.795 199.100 142.300 199.475 ;
        RECT 141.795 198.605 142.835 199.100 ;
        RECT 143.145 198.200 143.720 199.475 ;
        RECT 138.600 197.825 139.655 198.200 ;
        RECT 140.075 197.825 141.020 198.200 ;
        RECT 141.300 197.825 142.355 198.200 ;
        RECT 142.775 197.825 143.720 198.200 ;
        RECT 138.600 196.950 139.600 197.825 ;
        RECT 141.300 196.950 142.300 197.825 ;
        RECT 138.600 195.950 142.300 196.950 ;
        RECT 142.875 196.275 143.875 196.320 ;
        RECT 144.055 196.275 145.055 199.475 ;
        RECT 138.600 194.435 139.600 195.950 ;
        RECT 142.875 195.275 145.055 196.275 ;
        RECT 145.475 195.275 145.845 199.475 ;
        RECT 146.750 197.975 147.755 200.475 ;
        RECT 148.175 200.475 148.545 206.500 ;
        RECT 152.425 200.475 153.425 200.505 ;
        RECT 148.175 199.475 153.425 200.475 ;
        RECT 146.730 197.025 147.770 197.975 ;
        RECT 146.750 197.000 147.755 197.025 ;
        RECT 147.385 195.275 147.755 197.000 ;
        RECT 148.175 195.275 148.545 199.475 ;
        RECT 152.425 199.445 153.425 199.475 ;
        RECT 142.875 195.230 143.875 195.275 ;
        RECT 1.850 194.425 14.575 194.435 ;
        RECT 15.350 194.425 19.390 194.435 ;
        RECT 19.590 194.425 40.000 194.435 ;
        RECT 40.775 194.425 44.815 194.435 ;
        RECT 45.015 194.425 65.425 194.435 ;
        RECT 66.200 194.425 70.240 194.435 ;
        RECT 70.440 194.425 90.850 194.435 ;
        RECT 91.625 194.425 95.665 194.435 ;
        RECT 95.865 194.425 116.275 194.435 ;
        RECT 117.050 194.425 121.090 194.435 ;
        RECT 121.290 194.425 141.700 194.435 ;
        RECT 142.475 194.425 146.515 194.435 ;
        RECT 146.715 194.425 149.215 194.435 ;
        RECT 1.850 193.325 149.215 194.425 ;
        RECT 1.850 193.320 19.390 193.325 ;
        RECT 19.590 193.320 44.815 193.325 ;
        RECT 45.015 193.320 70.240 193.325 ;
        RECT 70.440 193.320 95.665 193.325 ;
        RECT 95.865 193.320 121.090 193.325 ;
        RECT 121.290 193.320 146.515 193.325 ;
        RECT 146.715 193.320 149.215 193.325 ;
        RECT 3.905 193.315 6.480 193.320 ;
        RECT 29.330 193.315 31.905 193.320 ;
        RECT 54.755 193.315 57.330 193.320 ;
        RECT 80.180 193.315 82.755 193.320 ;
        RECT 105.605 193.315 108.180 193.320 ;
        RECT 131.030 193.315 133.605 193.320 ;
        RECT 3.905 193.285 5.020 193.315 ;
        RECT 29.330 193.285 30.445 193.315 ;
        RECT 54.755 193.285 55.870 193.315 ;
        RECT 80.180 193.285 81.295 193.315 ;
        RECT 105.605 193.285 106.720 193.315 ;
        RECT 131.030 193.285 132.145 193.315 ;
        RECT 19.370 192.375 21.325 192.395 ;
        RECT 44.795 192.375 46.750 192.395 ;
        RECT 70.220 192.375 72.175 192.395 ;
        RECT 95.645 192.375 97.600 192.395 ;
        RECT 121.070 192.375 123.025 192.395 ;
        RECT 146.495 192.375 148.450 192.395 ;
        RECT 9.550 192.350 10.550 192.375 ;
        RECT 15.750 192.350 16.750 192.375 ;
        RECT 17.650 192.350 18.650 192.375 ;
        RECT 9.530 191.400 10.570 192.350 ;
        RECT 15.730 191.400 16.770 192.350 ;
        RECT 17.630 191.400 18.670 192.350 ;
        RECT 9.550 191.375 10.550 191.400 ;
        RECT 15.750 191.375 16.750 191.400 ;
        RECT 17.650 191.375 18.650 191.400 ;
        RECT 19.365 191.375 21.350 192.375 ;
        RECT 34.975 192.350 35.975 192.375 ;
        RECT 41.175 192.350 42.175 192.375 ;
        RECT 43.075 192.350 44.075 192.375 ;
        RECT 34.955 191.400 35.995 192.350 ;
        RECT 41.155 191.400 42.195 192.350 ;
        RECT 43.055 191.400 44.095 192.350 ;
        RECT 34.975 191.375 35.975 191.400 ;
        RECT 41.175 191.375 42.175 191.400 ;
        RECT 43.075 191.375 44.075 191.400 ;
        RECT 44.790 191.375 46.775 192.375 ;
        RECT 60.400 192.350 61.400 192.375 ;
        RECT 66.600 192.350 67.600 192.375 ;
        RECT 68.500 192.350 69.500 192.375 ;
        RECT 60.380 191.400 61.420 192.350 ;
        RECT 66.580 191.400 67.620 192.350 ;
        RECT 68.480 191.400 69.520 192.350 ;
        RECT 60.400 191.375 61.400 191.400 ;
        RECT 66.600 191.375 67.600 191.400 ;
        RECT 68.500 191.375 69.500 191.400 ;
        RECT 70.215 191.375 72.200 192.375 ;
        RECT 85.825 192.350 86.825 192.375 ;
        RECT 92.025 192.350 93.025 192.375 ;
        RECT 93.925 192.350 94.925 192.375 ;
        RECT 85.805 191.400 86.845 192.350 ;
        RECT 92.005 191.400 93.045 192.350 ;
        RECT 93.905 191.400 94.945 192.350 ;
        RECT 85.825 191.375 86.825 191.400 ;
        RECT 92.025 191.375 93.025 191.400 ;
        RECT 93.925 191.375 94.925 191.400 ;
        RECT 95.640 191.375 97.625 192.375 ;
        RECT 111.250 192.350 112.250 192.375 ;
        RECT 117.450 192.350 118.450 192.375 ;
        RECT 119.350 192.350 120.350 192.375 ;
        RECT 111.230 191.400 112.270 192.350 ;
        RECT 117.430 191.400 118.470 192.350 ;
        RECT 119.330 191.400 120.370 192.350 ;
        RECT 111.250 191.375 112.250 191.400 ;
        RECT 117.450 191.375 118.450 191.400 ;
        RECT 119.350 191.375 120.350 191.400 ;
        RECT 121.065 191.375 123.050 192.375 ;
        RECT 136.675 192.350 137.675 192.375 ;
        RECT 142.875 192.350 143.875 192.375 ;
        RECT 144.775 192.350 145.775 192.375 ;
        RECT 136.655 191.400 137.695 192.350 ;
        RECT 142.855 191.400 143.895 192.350 ;
        RECT 144.755 191.400 145.795 192.350 ;
        RECT 136.675 191.375 137.675 191.400 ;
        RECT 142.875 191.375 143.875 191.400 ;
        RECT 144.775 191.375 145.775 191.400 ;
        RECT 146.490 191.375 148.475 192.375 ;
        RECT 19.370 191.355 21.325 191.375 ;
        RECT 44.795 191.355 46.750 191.375 ;
        RECT 70.220 191.355 72.175 191.375 ;
        RECT 95.645 191.355 97.600 191.375 ;
        RECT 121.070 191.355 123.025 191.375 ;
        RECT 146.495 191.355 148.450 191.375 ;
        RECT 9.575 189.600 10.525 189.620 ;
        RECT 20.375 189.600 21.325 189.620 ;
        RECT 35.000 189.600 35.950 189.620 ;
        RECT 45.800 189.600 46.750 189.620 ;
        RECT 60.425 189.600 61.375 189.620 ;
        RECT 71.225 189.600 72.175 189.620 ;
        RECT 85.850 189.600 86.800 189.620 ;
        RECT 96.650 189.600 97.600 189.620 ;
        RECT 111.275 189.600 112.225 189.620 ;
        RECT 122.075 189.600 123.025 189.620 ;
        RECT 136.700 189.600 137.650 189.620 ;
        RECT 147.500 189.600 148.450 189.620 ;
        RECT 9.550 188.600 12.755 189.600 ;
        RECT 13.530 188.600 14.620 189.600 ;
        RECT 15.370 188.600 18.650 189.600 ;
        RECT 20.350 188.600 21.350 189.600 ;
        RECT 34.975 188.600 38.180 189.600 ;
        RECT 38.955 188.600 40.045 189.600 ;
        RECT 40.795 188.600 44.075 189.600 ;
        RECT 45.775 188.600 46.775 189.600 ;
        RECT 60.400 188.600 63.605 189.600 ;
        RECT 64.380 188.600 65.470 189.600 ;
        RECT 66.220 188.600 69.500 189.600 ;
        RECT 71.200 188.600 72.200 189.600 ;
        RECT 85.825 188.600 89.030 189.600 ;
        RECT 89.805 188.600 90.895 189.600 ;
        RECT 91.645 188.600 94.925 189.600 ;
        RECT 96.625 188.600 97.625 189.600 ;
        RECT 111.250 188.600 114.455 189.600 ;
        RECT 115.230 188.600 116.320 189.600 ;
        RECT 117.070 188.600 120.350 189.600 ;
        RECT 122.050 188.600 123.050 189.600 ;
        RECT 136.675 188.600 139.880 189.600 ;
        RECT 140.655 188.600 141.745 189.600 ;
        RECT 142.495 188.600 145.775 189.600 ;
        RECT 147.475 188.600 148.475 189.600 ;
        RECT 9.575 188.580 10.525 188.600 ;
        RECT 3.925 187.655 4.980 187.675 ;
        RECT 3.575 187.650 6.000 187.655 ;
        RECT 1.850 186.550 12.025 187.650 ;
        RECT 13.575 187.625 14.575 188.600 ;
        RECT 20.375 188.580 21.325 188.600 ;
        RECT 35.000 188.580 35.950 188.600 ;
        RECT 29.350 187.655 30.405 187.675 ;
        RECT 29.000 187.650 31.425 187.655 ;
        RECT 12.650 186.625 14.575 187.625 ;
        RECT 1.850 186.545 11.290 186.550 ;
        RECT 3.925 186.530 4.980 186.545 ;
        RECT 6.050 180.400 7.050 186.545 ;
        RECT 12.650 185.250 13.650 186.625 ;
        RECT 16.175 186.550 37.450 187.650 ;
        RECT 39.000 187.625 40.000 188.600 ;
        RECT 45.800 188.580 46.750 188.600 ;
        RECT 60.425 188.580 61.375 188.600 ;
        RECT 54.775 187.655 55.830 187.675 ;
        RECT 54.425 187.650 56.850 187.655 ;
        RECT 38.075 186.625 40.000 187.625 ;
        RECT 16.890 186.545 19.400 186.550 ;
        RECT 19.590 186.545 36.715 186.550 ;
        RECT 29.350 186.530 30.405 186.545 ;
        RECT 12.630 184.300 13.670 185.250 ;
        RECT 12.650 184.275 13.650 184.300 ;
        RECT 14.405 184.275 15.495 185.275 ;
        RECT 6.050 179.400 7.075 180.400 ;
        RECT 7.550 179.400 8.495 179.925 ;
        RECT 6.570 178.275 7.610 178.750 ;
        RECT 1.900 177.925 2.900 177.930 ;
        RECT 1.870 177.900 2.930 177.925 ;
        RECT 6.570 177.900 7.075 178.275 ;
        RECT 7.920 177.945 8.495 179.400 ;
        RECT 1.850 177.875 7.075 177.900 ;
        RECT 1.850 176.925 7.095 177.875 ;
        RECT 1.850 176.900 7.075 176.925 ;
        RECT 1.900 176.870 2.900 176.900 ;
        RECT 6.570 176.525 7.075 176.900 ;
        RECT 7.500 176.855 8.500 177.945 ;
        RECT 9.460 177.900 9.830 183.925 ;
        RECT 8.825 176.900 9.830 177.900 ;
        RECT 6.570 176.030 7.610 176.525 ;
        RECT 7.920 175.625 8.495 176.855 ;
        RECT 6.075 175.250 7.130 175.625 ;
        RECT 7.550 175.250 8.495 175.625 ;
        RECT 3.905 171.860 5.020 171.885 ;
        RECT 6.075 171.860 7.075 175.250 ;
        RECT 8.830 173.700 9.830 176.900 ;
        RECT 7.630 172.700 9.830 173.700 ;
        RECT 10.250 177.945 10.620 183.925 ;
        RECT 14.450 183.500 15.450 183.530 ;
        RECT 14.450 182.500 17.220 183.500 ;
        RECT 14.450 182.470 15.450 182.500 ;
        RECT 11.475 179.400 12.475 181.850 ;
        RECT 12.950 179.400 13.895 179.925 ;
        RECT 14.175 179.400 15.175 181.850 ;
        RECT 15.650 179.400 16.595 179.925 ;
        RECT 11.970 178.275 13.010 178.750 ;
        RECT 10.250 177.900 11.250 177.945 ;
        RECT 11.970 177.900 12.475 178.275 ;
        RECT 13.320 177.900 13.895 179.400 ;
        RECT 14.670 178.275 15.710 178.750 ;
        RECT 14.670 177.900 15.175 178.275 ;
        RECT 16.020 177.900 16.595 179.400 ;
        RECT 17.560 177.900 17.930 183.925 ;
        RECT 18.350 177.900 18.720 183.925 ;
        RECT 20.260 177.900 20.630 183.925 ;
        RECT 10.250 177.875 12.475 177.900 ;
        RECT 10.250 176.930 12.495 177.875 ;
        RECT 10.250 176.900 12.475 176.930 ;
        RECT 12.855 176.900 15.175 177.900 ;
        RECT 15.600 176.900 17.930 177.900 ;
        RECT 18.305 176.900 19.395 177.900 ;
        RECT 10.250 176.855 11.250 176.900 ;
        RECT 10.250 172.700 10.620 176.855 ;
        RECT 11.970 176.525 12.475 176.900 ;
        RECT 11.970 176.030 13.010 176.525 ;
        RECT 13.320 175.625 13.895 176.900 ;
        RECT 14.670 176.525 15.175 176.900 ;
        RECT 14.670 176.030 15.710 176.525 ;
        RECT 16.020 175.625 16.595 176.900 ;
        RECT 11.475 175.250 12.530 175.625 ;
        RECT 12.950 175.250 13.895 175.625 ;
        RECT 14.175 175.250 15.230 175.625 ;
        RECT 15.650 175.250 16.595 175.625 ;
        RECT 11.475 174.375 12.475 175.250 ;
        RECT 14.175 174.375 15.175 175.250 ;
        RECT 11.475 173.375 15.175 174.375 ;
        RECT 15.750 173.700 16.750 173.745 ;
        RECT 16.930 173.700 17.930 176.900 ;
        RECT 11.475 171.860 12.475 173.375 ;
        RECT 15.750 172.700 17.930 173.700 ;
        RECT 18.350 172.700 18.720 176.900 ;
        RECT 19.625 175.900 20.630 177.900 ;
        RECT 21.050 177.925 21.420 183.925 ;
        RECT 31.475 180.400 32.475 186.545 ;
        RECT 38.075 185.250 39.075 186.625 ;
        RECT 41.600 186.550 62.875 187.650 ;
        RECT 64.425 187.625 65.425 188.600 ;
        RECT 71.225 188.580 72.175 188.600 ;
        RECT 85.850 188.580 86.800 188.600 ;
        RECT 80.200 187.655 81.255 187.675 ;
        RECT 79.850 187.650 82.275 187.655 ;
        RECT 63.500 186.625 65.425 187.625 ;
        RECT 42.315 186.545 44.825 186.550 ;
        RECT 45.015 186.545 62.140 186.550 ;
        RECT 54.775 186.530 55.830 186.545 ;
        RECT 38.055 184.300 39.095 185.250 ;
        RECT 38.075 184.275 39.075 184.300 ;
        RECT 39.830 184.275 40.920 185.275 ;
        RECT 31.475 179.400 32.500 180.400 ;
        RECT 32.975 179.400 33.920 179.925 ;
        RECT 31.995 178.275 33.035 178.750 ;
        RECT 27.325 177.925 28.325 177.930 ;
        RECT 21.050 177.900 22.375 177.925 ;
        RECT 27.295 177.900 28.355 177.925 ;
        RECT 31.995 177.900 32.500 178.275 ;
        RECT 33.345 177.945 33.920 179.400 ;
        RECT 21.050 176.900 26.250 177.900 ;
        RECT 27.275 177.875 32.500 177.900 ;
        RECT 27.275 176.925 32.520 177.875 ;
        RECT 27.275 176.900 32.500 176.925 ;
        RECT 21.050 176.885 22.375 176.900 ;
        RECT 19.605 174.950 20.645 175.900 ;
        RECT 19.625 174.925 20.630 174.950 ;
        RECT 20.260 172.700 20.630 174.925 ;
        RECT 21.050 172.700 21.420 176.885 ;
        RECT 23.155 173.775 24.155 176.900 ;
        RECT 27.325 176.870 28.325 176.900 ;
        RECT 31.995 176.525 32.500 176.900 ;
        RECT 32.925 176.855 33.925 177.945 ;
        RECT 34.885 177.900 35.255 183.925 ;
        RECT 34.250 176.900 35.255 177.900 ;
        RECT 31.995 176.030 33.035 176.525 ;
        RECT 33.345 175.625 33.920 176.855 ;
        RECT 31.500 175.250 32.555 175.625 ;
        RECT 32.975 175.250 33.920 175.625 ;
        RECT 23.135 172.825 24.175 173.775 ;
        RECT 23.155 172.800 24.155 172.825 ;
        RECT 15.750 172.655 16.750 172.700 ;
        RECT 23.115 171.860 24.230 171.890 ;
        RECT 29.330 171.860 30.445 171.885 ;
        RECT 31.500 171.860 32.500 175.250 ;
        RECT 34.255 173.700 35.255 176.900 ;
        RECT 33.055 172.700 35.255 173.700 ;
        RECT 35.675 177.945 36.045 183.925 ;
        RECT 39.875 183.500 40.875 183.530 ;
        RECT 39.875 182.500 42.645 183.500 ;
        RECT 39.875 182.470 40.875 182.500 ;
        RECT 36.900 179.400 37.900 181.850 ;
        RECT 38.375 179.400 39.320 179.925 ;
        RECT 39.600 179.400 40.600 181.850 ;
        RECT 41.075 179.400 42.020 179.925 ;
        RECT 37.395 178.275 38.435 178.750 ;
        RECT 35.675 177.900 36.675 177.945 ;
        RECT 37.395 177.900 37.900 178.275 ;
        RECT 38.745 177.900 39.320 179.400 ;
        RECT 40.095 178.275 41.135 178.750 ;
        RECT 40.095 177.900 40.600 178.275 ;
        RECT 41.445 177.900 42.020 179.400 ;
        RECT 42.985 177.900 43.355 183.925 ;
        RECT 43.775 177.900 44.145 183.925 ;
        RECT 45.685 177.900 46.055 183.925 ;
        RECT 35.675 177.875 37.900 177.900 ;
        RECT 35.675 176.930 37.920 177.875 ;
        RECT 35.675 176.900 37.900 176.930 ;
        RECT 38.280 176.900 40.600 177.900 ;
        RECT 41.025 176.900 43.355 177.900 ;
        RECT 43.730 176.900 44.820 177.900 ;
        RECT 35.675 176.855 36.675 176.900 ;
        RECT 35.675 172.700 36.045 176.855 ;
        RECT 37.395 176.525 37.900 176.900 ;
        RECT 37.395 176.030 38.435 176.525 ;
        RECT 38.745 175.625 39.320 176.900 ;
        RECT 40.095 176.525 40.600 176.900 ;
        RECT 40.095 176.030 41.135 176.525 ;
        RECT 41.445 175.625 42.020 176.900 ;
        RECT 36.900 175.250 37.955 175.625 ;
        RECT 38.375 175.250 39.320 175.625 ;
        RECT 39.600 175.250 40.655 175.625 ;
        RECT 41.075 175.250 42.020 175.625 ;
        RECT 36.900 174.375 37.900 175.250 ;
        RECT 39.600 174.375 40.600 175.250 ;
        RECT 36.900 173.375 40.600 174.375 ;
        RECT 41.175 173.700 42.175 173.745 ;
        RECT 42.355 173.700 43.355 176.900 ;
        RECT 36.900 171.860 37.900 173.375 ;
        RECT 41.175 172.700 43.355 173.700 ;
        RECT 43.775 172.700 44.145 176.900 ;
        RECT 45.050 175.900 46.055 177.900 ;
        RECT 46.475 177.900 46.845 183.925 ;
        RECT 56.900 180.400 57.900 186.545 ;
        RECT 63.500 185.250 64.500 186.625 ;
        RECT 67.025 186.550 88.300 187.650 ;
        RECT 89.850 187.625 90.850 188.600 ;
        RECT 96.650 188.580 97.600 188.600 ;
        RECT 111.275 188.580 112.225 188.600 ;
        RECT 105.625 187.655 106.680 187.675 ;
        RECT 105.275 187.650 107.700 187.655 ;
        RECT 88.925 186.625 90.850 187.625 ;
        RECT 67.740 186.545 70.250 186.550 ;
        RECT 70.440 186.545 87.565 186.550 ;
        RECT 80.200 186.530 81.255 186.545 ;
        RECT 63.480 184.300 64.520 185.250 ;
        RECT 63.500 184.275 64.500 184.300 ;
        RECT 65.255 184.275 66.345 185.275 ;
        RECT 56.900 179.400 57.925 180.400 ;
        RECT 58.400 179.400 59.345 179.925 ;
        RECT 57.420 178.275 58.460 178.750 ;
        RECT 52.750 177.925 53.750 177.930 ;
        RECT 52.720 177.900 53.780 177.925 ;
        RECT 57.420 177.900 57.925 178.275 ;
        RECT 58.770 177.945 59.345 179.400 ;
        RECT 46.475 176.900 51.720 177.900 ;
        RECT 52.700 177.875 57.925 177.900 ;
        RECT 52.700 176.925 57.945 177.875 ;
        RECT 52.700 176.900 57.925 176.925 ;
        RECT 45.030 174.950 46.070 175.900 ;
        RECT 45.050 174.925 46.055 174.950 ;
        RECT 45.685 172.700 46.055 174.925 ;
        RECT 46.475 172.700 46.845 176.900 ;
        RECT 48.580 173.775 49.580 176.900 ;
        RECT 52.750 176.870 53.750 176.900 ;
        RECT 57.420 176.525 57.925 176.900 ;
        RECT 58.350 176.855 59.350 177.945 ;
        RECT 60.310 177.900 60.680 183.925 ;
        RECT 59.675 176.900 60.680 177.900 ;
        RECT 57.420 176.030 58.460 176.525 ;
        RECT 58.770 175.625 59.345 176.855 ;
        RECT 56.925 175.250 57.980 175.625 ;
        RECT 58.400 175.250 59.345 175.625 ;
        RECT 48.560 172.825 49.600 173.775 ;
        RECT 48.580 172.800 49.580 172.825 ;
        RECT 41.175 172.655 42.175 172.700 ;
        RECT 48.540 171.860 49.655 171.890 ;
        RECT 54.755 171.860 55.870 171.885 ;
        RECT 56.925 171.860 57.925 175.250 ;
        RECT 59.680 173.700 60.680 176.900 ;
        RECT 58.480 172.700 60.680 173.700 ;
        RECT 61.100 177.945 61.470 183.925 ;
        RECT 65.300 183.500 66.300 183.530 ;
        RECT 65.300 182.500 68.070 183.500 ;
        RECT 65.300 182.470 66.300 182.500 ;
        RECT 62.325 179.400 63.325 181.850 ;
        RECT 63.800 179.400 64.745 179.925 ;
        RECT 65.025 179.400 66.025 181.850 ;
        RECT 66.500 179.400 67.445 179.925 ;
        RECT 62.820 178.275 63.860 178.750 ;
        RECT 61.100 177.900 62.100 177.945 ;
        RECT 62.820 177.900 63.325 178.275 ;
        RECT 64.170 177.900 64.745 179.400 ;
        RECT 65.520 178.275 66.560 178.750 ;
        RECT 65.520 177.900 66.025 178.275 ;
        RECT 66.870 177.900 67.445 179.400 ;
        RECT 68.410 177.900 68.780 183.925 ;
        RECT 69.200 177.900 69.570 183.925 ;
        RECT 71.110 177.900 71.480 183.925 ;
        RECT 61.100 177.875 63.325 177.900 ;
        RECT 61.100 176.930 63.345 177.875 ;
        RECT 61.100 176.900 63.325 176.930 ;
        RECT 63.705 176.900 66.025 177.900 ;
        RECT 66.450 176.900 68.780 177.900 ;
        RECT 69.155 176.900 70.245 177.900 ;
        RECT 61.100 176.855 62.100 176.900 ;
        RECT 61.100 172.700 61.470 176.855 ;
        RECT 62.820 176.525 63.325 176.900 ;
        RECT 62.820 176.030 63.860 176.525 ;
        RECT 64.170 175.625 64.745 176.900 ;
        RECT 65.520 176.525 66.025 176.900 ;
        RECT 65.520 176.030 66.560 176.525 ;
        RECT 66.870 175.625 67.445 176.900 ;
        RECT 62.325 175.250 63.380 175.625 ;
        RECT 63.800 175.250 64.745 175.625 ;
        RECT 65.025 175.250 66.080 175.625 ;
        RECT 66.500 175.250 67.445 175.625 ;
        RECT 62.325 174.375 63.325 175.250 ;
        RECT 65.025 174.375 66.025 175.250 ;
        RECT 62.325 173.375 66.025 174.375 ;
        RECT 66.600 173.700 67.600 173.745 ;
        RECT 67.780 173.700 68.780 176.900 ;
        RECT 62.325 171.860 63.325 173.375 ;
        RECT 66.600 172.700 68.780 173.700 ;
        RECT 69.200 172.700 69.570 176.900 ;
        RECT 70.475 175.900 71.480 177.900 ;
        RECT 71.900 177.925 72.270 183.925 ;
        RECT 82.325 180.400 83.325 186.545 ;
        RECT 88.925 185.250 89.925 186.625 ;
        RECT 92.450 186.550 113.725 187.650 ;
        RECT 115.275 187.625 116.275 188.600 ;
        RECT 122.075 188.580 123.025 188.600 ;
        RECT 136.700 188.580 137.650 188.600 ;
        RECT 131.050 187.655 132.105 187.675 ;
        RECT 130.700 187.650 133.125 187.655 ;
        RECT 114.350 186.625 116.275 187.625 ;
        RECT 93.165 186.545 95.675 186.550 ;
        RECT 95.865 186.545 112.990 186.550 ;
        RECT 105.625 186.530 106.680 186.545 ;
        RECT 88.905 184.300 89.945 185.250 ;
        RECT 88.925 184.275 89.925 184.300 ;
        RECT 90.680 184.275 91.770 185.275 ;
        RECT 82.325 179.400 83.350 180.400 ;
        RECT 83.825 179.400 84.770 179.925 ;
        RECT 82.845 178.275 83.885 178.750 ;
        RECT 78.175 177.925 79.175 177.930 ;
        RECT 71.900 177.900 73.225 177.925 ;
        RECT 78.145 177.900 79.205 177.925 ;
        RECT 82.845 177.900 83.350 178.275 ;
        RECT 84.195 177.945 84.770 179.400 ;
        RECT 71.900 176.900 77.100 177.900 ;
        RECT 78.125 177.875 83.350 177.900 ;
        RECT 78.125 176.925 83.370 177.875 ;
        RECT 78.125 176.900 83.350 176.925 ;
        RECT 71.900 176.885 73.225 176.900 ;
        RECT 70.455 174.950 71.495 175.900 ;
        RECT 70.475 174.925 71.480 174.950 ;
        RECT 71.110 172.700 71.480 174.925 ;
        RECT 71.900 172.700 72.270 176.885 ;
        RECT 74.005 173.775 75.005 176.900 ;
        RECT 78.175 176.870 79.175 176.900 ;
        RECT 82.845 176.525 83.350 176.900 ;
        RECT 83.775 176.855 84.775 177.945 ;
        RECT 85.735 177.900 86.105 183.925 ;
        RECT 85.100 176.900 86.105 177.900 ;
        RECT 82.845 176.030 83.885 176.525 ;
        RECT 84.195 175.625 84.770 176.855 ;
        RECT 82.350 175.250 83.405 175.625 ;
        RECT 83.825 175.250 84.770 175.625 ;
        RECT 73.985 172.825 75.025 173.775 ;
        RECT 74.005 172.800 75.005 172.825 ;
        RECT 66.600 172.655 67.600 172.700 ;
        RECT 73.965 171.860 75.080 171.890 ;
        RECT 80.180 171.860 81.295 171.885 ;
        RECT 82.350 171.860 83.350 175.250 ;
        RECT 85.105 173.700 86.105 176.900 ;
        RECT 83.905 172.700 86.105 173.700 ;
        RECT 86.525 177.945 86.895 183.925 ;
        RECT 90.725 183.500 91.725 183.530 ;
        RECT 90.725 182.500 93.495 183.500 ;
        RECT 90.725 182.470 91.725 182.500 ;
        RECT 87.750 179.400 88.750 181.850 ;
        RECT 89.225 179.400 90.170 179.925 ;
        RECT 90.450 179.400 91.450 181.850 ;
        RECT 91.925 179.400 92.870 179.925 ;
        RECT 88.245 178.275 89.285 178.750 ;
        RECT 86.525 177.900 87.525 177.945 ;
        RECT 88.245 177.900 88.750 178.275 ;
        RECT 89.595 177.900 90.170 179.400 ;
        RECT 90.945 178.275 91.985 178.750 ;
        RECT 90.945 177.900 91.450 178.275 ;
        RECT 92.295 177.900 92.870 179.400 ;
        RECT 93.835 177.900 94.205 183.925 ;
        RECT 94.625 177.900 94.995 183.925 ;
        RECT 96.535 177.900 96.905 183.925 ;
        RECT 86.525 177.875 88.750 177.900 ;
        RECT 86.525 176.930 88.770 177.875 ;
        RECT 86.525 176.900 88.750 176.930 ;
        RECT 89.130 176.900 91.450 177.900 ;
        RECT 91.875 176.900 94.205 177.900 ;
        RECT 94.580 176.900 95.670 177.900 ;
        RECT 86.525 176.855 87.525 176.900 ;
        RECT 86.525 172.700 86.895 176.855 ;
        RECT 88.245 176.525 88.750 176.900 ;
        RECT 88.245 176.030 89.285 176.525 ;
        RECT 89.595 175.625 90.170 176.900 ;
        RECT 90.945 176.525 91.450 176.900 ;
        RECT 90.945 176.030 91.985 176.525 ;
        RECT 92.295 175.625 92.870 176.900 ;
        RECT 87.750 175.250 88.805 175.625 ;
        RECT 89.225 175.250 90.170 175.625 ;
        RECT 90.450 175.250 91.505 175.625 ;
        RECT 91.925 175.250 92.870 175.625 ;
        RECT 87.750 174.375 88.750 175.250 ;
        RECT 90.450 174.375 91.450 175.250 ;
        RECT 87.750 173.375 91.450 174.375 ;
        RECT 92.025 173.700 93.025 173.745 ;
        RECT 93.205 173.700 94.205 176.900 ;
        RECT 87.750 171.860 88.750 173.375 ;
        RECT 92.025 172.700 94.205 173.700 ;
        RECT 94.625 172.700 94.995 176.900 ;
        RECT 95.900 175.900 96.905 177.900 ;
        RECT 97.325 177.900 97.695 183.925 ;
        RECT 107.750 180.400 108.750 186.545 ;
        RECT 114.350 185.250 115.350 186.625 ;
        RECT 117.875 186.550 139.150 187.650 ;
        RECT 140.700 187.625 141.700 188.600 ;
        RECT 147.500 188.580 148.450 188.600 ;
        RECT 139.775 186.625 141.700 187.625 ;
        RECT 118.590 186.545 121.100 186.550 ;
        RECT 121.290 186.545 138.415 186.550 ;
        RECT 131.050 186.530 132.105 186.545 ;
        RECT 114.330 184.300 115.370 185.250 ;
        RECT 114.350 184.275 115.350 184.300 ;
        RECT 116.105 184.275 117.195 185.275 ;
        RECT 107.750 179.400 108.775 180.400 ;
        RECT 109.250 179.400 110.195 179.925 ;
        RECT 108.270 178.275 109.310 178.750 ;
        RECT 103.600 177.925 104.600 177.930 ;
        RECT 103.570 177.900 104.630 177.925 ;
        RECT 108.270 177.900 108.775 178.275 ;
        RECT 109.620 177.945 110.195 179.400 ;
        RECT 97.325 176.900 102.570 177.900 ;
        RECT 103.550 177.875 108.775 177.900 ;
        RECT 103.550 176.925 108.795 177.875 ;
        RECT 103.550 176.900 108.775 176.925 ;
        RECT 95.880 174.950 96.920 175.900 ;
        RECT 95.900 174.925 96.905 174.950 ;
        RECT 96.535 172.700 96.905 174.925 ;
        RECT 97.325 172.700 97.695 176.900 ;
        RECT 99.430 173.775 100.430 176.900 ;
        RECT 103.600 176.870 104.600 176.900 ;
        RECT 108.270 176.525 108.775 176.900 ;
        RECT 109.200 176.855 110.200 177.945 ;
        RECT 111.160 177.900 111.530 183.925 ;
        RECT 110.525 176.900 111.530 177.900 ;
        RECT 108.270 176.030 109.310 176.525 ;
        RECT 109.620 175.625 110.195 176.855 ;
        RECT 107.775 175.250 108.830 175.625 ;
        RECT 109.250 175.250 110.195 175.625 ;
        RECT 99.410 172.825 100.450 173.775 ;
        RECT 99.430 172.800 100.430 172.825 ;
        RECT 92.025 172.655 93.025 172.700 ;
        RECT 99.390 171.860 100.505 171.890 ;
        RECT 105.605 171.860 106.720 171.885 ;
        RECT 107.775 171.860 108.775 175.250 ;
        RECT 110.530 173.700 111.530 176.900 ;
        RECT 109.330 172.700 111.530 173.700 ;
        RECT 111.950 177.945 112.320 183.925 ;
        RECT 116.150 183.500 117.150 183.530 ;
        RECT 116.150 182.500 118.920 183.500 ;
        RECT 116.150 182.470 117.150 182.500 ;
        RECT 113.175 179.400 114.175 181.850 ;
        RECT 114.650 179.400 115.595 179.925 ;
        RECT 115.875 179.400 116.875 181.850 ;
        RECT 117.350 179.400 118.295 179.925 ;
        RECT 113.670 178.275 114.710 178.750 ;
        RECT 111.950 177.900 112.950 177.945 ;
        RECT 113.670 177.900 114.175 178.275 ;
        RECT 115.020 177.900 115.595 179.400 ;
        RECT 116.370 178.275 117.410 178.750 ;
        RECT 116.370 177.900 116.875 178.275 ;
        RECT 117.720 177.900 118.295 179.400 ;
        RECT 119.260 177.900 119.630 183.925 ;
        RECT 120.050 177.900 120.420 183.925 ;
        RECT 121.960 177.900 122.330 183.925 ;
        RECT 111.950 177.875 114.175 177.900 ;
        RECT 111.950 176.930 114.195 177.875 ;
        RECT 111.950 176.900 114.175 176.930 ;
        RECT 114.555 176.900 116.875 177.900 ;
        RECT 117.300 176.900 119.630 177.900 ;
        RECT 120.005 176.900 121.095 177.900 ;
        RECT 111.950 176.855 112.950 176.900 ;
        RECT 111.950 172.700 112.320 176.855 ;
        RECT 113.670 176.525 114.175 176.900 ;
        RECT 113.670 176.030 114.710 176.525 ;
        RECT 115.020 175.625 115.595 176.900 ;
        RECT 116.370 176.525 116.875 176.900 ;
        RECT 116.370 176.030 117.410 176.525 ;
        RECT 117.720 175.625 118.295 176.900 ;
        RECT 113.175 175.250 114.230 175.625 ;
        RECT 114.650 175.250 115.595 175.625 ;
        RECT 115.875 175.250 116.930 175.625 ;
        RECT 117.350 175.250 118.295 175.625 ;
        RECT 113.175 174.375 114.175 175.250 ;
        RECT 115.875 174.375 116.875 175.250 ;
        RECT 113.175 173.375 116.875 174.375 ;
        RECT 117.450 173.700 118.450 173.745 ;
        RECT 118.630 173.700 119.630 176.900 ;
        RECT 113.175 171.860 114.175 173.375 ;
        RECT 117.450 172.700 119.630 173.700 ;
        RECT 120.050 172.700 120.420 176.900 ;
        RECT 121.325 175.900 122.330 177.900 ;
        RECT 122.750 177.925 123.120 183.925 ;
        RECT 133.175 180.400 134.175 186.545 ;
        RECT 139.775 185.250 140.775 186.625 ;
        RECT 143.300 186.550 149.225 187.650 ;
        RECT 144.015 186.545 146.525 186.550 ;
        RECT 146.715 186.545 149.215 186.550 ;
        RECT 139.755 184.300 140.795 185.250 ;
        RECT 139.775 184.275 140.775 184.300 ;
        RECT 141.530 184.275 142.620 185.275 ;
        RECT 133.175 179.400 134.200 180.400 ;
        RECT 134.675 179.400 135.620 179.925 ;
        RECT 133.695 178.275 134.735 178.750 ;
        RECT 129.025 177.925 130.025 177.930 ;
        RECT 122.750 177.900 124.075 177.925 ;
        RECT 128.995 177.900 130.055 177.925 ;
        RECT 133.695 177.900 134.200 178.275 ;
        RECT 135.045 177.945 135.620 179.400 ;
        RECT 122.750 176.900 127.950 177.900 ;
        RECT 128.975 177.875 134.200 177.900 ;
        RECT 128.975 176.925 134.220 177.875 ;
        RECT 128.975 176.900 134.200 176.925 ;
        RECT 122.750 176.885 124.075 176.900 ;
        RECT 121.305 174.950 122.345 175.900 ;
        RECT 121.325 174.925 122.330 174.950 ;
        RECT 121.960 172.700 122.330 174.925 ;
        RECT 122.750 172.700 123.120 176.885 ;
        RECT 124.855 173.775 125.855 176.900 ;
        RECT 129.025 176.870 130.025 176.900 ;
        RECT 133.695 176.525 134.200 176.900 ;
        RECT 134.625 176.855 135.625 177.945 ;
        RECT 136.585 177.900 136.955 183.925 ;
        RECT 135.950 176.900 136.955 177.900 ;
        RECT 133.695 176.030 134.735 176.525 ;
        RECT 135.045 175.625 135.620 176.855 ;
        RECT 133.200 175.250 134.255 175.625 ;
        RECT 134.675 175.250 135.620 175.625 ;
        RECT 124.835 172.825 125.875 173.775 ;
        RECT 124.855 172.800 125.855 172.825 ;
        RECT 117.450 172.655 118.450 172.700 ;
        RECT 124.815 171.860 125.930 171.890 ;
        RECT 131.030 171.860 132.145 171.885 ;
        RECT 133.200 171.860 134.200 175.250 ;
        RECT 135.955 173.700 136.955 176.900 ;
        RECT 134.755 172.700 136.955 173.700 ;
        RECT 137.375 177.945 137.745 183.925 ;
        RECT 141.575 183.500 142.575 183.530 ;
        RECT 141.575 182.500 144.345 183.500 ;
        RECT 141.575 182.470 142.575 182.500 ;
        RECT 138.600 179.400 139.600 181.850 ;
        RECT 140.075 179.400 141.020 179.925 ;
        RECT 141.300 179.400 142.300 181.850 ;
        RECT 142.775 179.400 143.720 179.925 ;
        RECT 139.095 178.275 140.135 178.750 ;
        RECT 137.375 177.900 138.375 177.945 ;
        RECT 139.095 177.900 139.600 178.275 ;
        RECT 140.445 177.900 141.020 179.400 ;
        RECT 141.795 178.275 142.835 178.750 ;
        RECT 141.795 177.900 142.300 178.275 ;
        RECT 143.145 177.900 143.720 179.400 ;
        RECT 144.685 177.900 145.055 183.925 ;
        RECT 145.475 177.900 145.845 183.925 ;
        RECT 147.385 177.900 147.755 183.925 ;
        RECT 137.375 177.875 139.600 177.900 ;
        RECT 137.375 176.930 139.620 177.875 ;
        RECT 137.375 176.900 139.600 176.930 ;
        RECT 139.980 176.900 142.300 177.900 ;
        RECT 142.725 176.900 145.055 177.900 ;
        RECT 145.430 176.900 146.520 177.900 ;
        RECT 137.375 176.855 138.375 176.900 ;
        RECT 137.375 172.700 137.745 176.855 ;
        RECT 139.095 176.525 139.600 176.900 ;
        RECT 139.095 176.030 140.135 176.525 ;
        RECT 140.445 175.625 141.020 176.900 ;
        RECT 141.795 176.525 142.300 176.900 ;
        RECT 141.795 176.030 142.835 176.525 ;
        RECT 143.145 175.625 143.720 176.900 ;
        RECT 138.600 175.250 139.655 175.625 ;
        RECT 140.075 175.250 141.020 175.625 ;
        RECT 141.300 175.250 142.355 175.625 ;
        RECT 142.775 175.250 143.720 175.625 ;
        RECT 138.600 174.375 139.600 175.250 ;
        RECT 141.300 174.375 142.300 175.250 ;
        RECT 138.600 173.375 142.300 174.375 ;
        RECT 142.875 173.700 143.875 173.745 ;
        RECT 144.055 173.700 145.055 176.900 ;
        RECT 138.600 171.860 139.600 173.375 ;
        RECT 142.875 172.700 145.055 173.700 ;
        RECT 145.475 172.700 145.845 176.900 ;
        RECT 146.750 175.900 147.755 177.900 ;
        RECT 148.175 177.900 148.545 183.925 ;
        RECT 156.525 177.900 157.525 177.945 ;
        RECT 148.175 176.900 157.525 177.900 ;
        RECT 146.730 174.950 147.770 175.900 ;
        RECT 146.750 174.925 147.755 174.950 ;
        RECT 147.385 172.700 147.755 174.925 ;
        RECT 148.175 172.700 148.545 176.900 ;
        RECT 150.280 173.775 151.280 176.900 ;
        RECT 156.525 176.855 157.525 176.900 ;
        RECT 150.260 172.825 151.300 173.775 ;
        RECT 150.280 172.800 151.280 172.825 ;
        RECT 142.875 172.655 143.875 172.700 ;
        RECT 150.240 171.860 151.355 171.890 ;
        RECT 1.850 171.850 14.575 171.860 ;
        RECT 15.350 171.850 19.390 171.860 ;
        RECT 19.590 171.850 40.000 171.860 ;
        RECT 40.775 171.850 44.815 171.860 ;
        RECT 45.015 171.850 65.425 171.860 ;
        RECT 66.200 171.850 70.240 171.860 ;
        RECT 70.440 171.850 90.850 171.860 ;
        RECT 91.625 171.850 95.665 171.860 ;
        RECT 95.865 171.850 116.275 171.860 ;
        RECT 117.050 171.850 121.090 171.860 ;
        RECT 121.290 171.850 141.700 171.860 ;
        RECT 142.475 171.850 146.515 171.860 ;
        RECT 146.715 171.850 151.355 171.860 ;
        RECT 1.850 170.750 151.355 171.850 ;
        RECT 1.850 170.745 19.390 170.750 ;
        RECT 19.590 170.745 44.815 170.750 ;
        RECT 45.015 170.745 70.240 170.750 ;
        RECT 70.440 170.745 95.665 170.750 ;
        RECT 95.865 170.745 121.090 170.750 ;
        RECT 121.290 170.745 146.515 170.750 ;
        RECT 146.715 170.745 151.355 170.750 ;
        RECT 3.875 170.740 7.105 170.745 ;
        RECT 3.905 170.710 5.020 170.740 ;
        RECT 23.115 170.715 24.230 170.745 ;
        RECT 29.300 170.740 32.530 170.745 ;
        RECT 29.330 170.710 30.445 170.740 ;
        RECT 48.540 170.715 49.655 170.745 ;
        RECT 54.725 170.740 57.955 170.745 ;
        RECT 54.755 170.710 55.870 170.740 ;
        RECT 73.965 170.715 75.080 170.745 ;
        RECT 80.150 170.740 83.380 170.745 ;
        RECT 80.180 170.710 81.295 170.740 ;
        RECT 99.390 170.715 100.505 170.745 ;
        RECT 105.575 170.740 108.805 170.745 ;
        RECT 105.605 170.710 106.720 170.740 ;
        RECT 124.815 170.715 125.930 170.745 ;
        RECT 131.000 170.740 134.230 170.745 ;
        RECT 131.030 170.710 132.145 170.740 ;
        RECT 150.240 170.715 151.355 170.745 ;
        RECT 19.370 169.800 21.325 169.820 ;
        RECT 44.795 169.800 46.750 169.820 ;
        RECT 70.220 169.800 72.175 169.820 ;
        RECT 95.645 169.800 97.600 169.820 ;
        RECT 121.070 169.800 123.025 169.820 ;
        RECT 146.495 169.800 148.450 169.820 ;
        RECT 9.550 169.775 10.550 169.800 ;
        RECT 15.750 169.775 16.750 169.800 ;
        RECT 17.650 169.775 18.650 169.800 ;
        RECT 9.530 168.825 10.570 169.775 ;
        RECT 15.730 168.825 16.770 169.775 ;
        RECT 17.630 168.825 18.670 169.775 ;
        RECT 9.550 168.800 10.550 168.825 ;
        RECT 15.750 168.800 16.750 168.825 ;
        RECT 17.650 168.800 18.650 168.825 ;
        RECT 19.365 168.800 21.350 169.800 ;
        RECT 34.975 169.775 35.975 169.800 ;
        RECT 41.175 169.775 42.175 169.800 ;
        RECT 43.075 169.775 44.075 169.800 ;
        RECT 34.955 168.825 35.995 169.775 ;
        RECT 41.155 168.825 42.195 169.775 ;
        RECT 43.055 168.825 44.095 169.775 ;
        RECT 34.975 168.800 35.975 168.825 ;
        RECT 41.175 168.800 42.175 168.825 ;
        RECT 43.075 168.800 44.075 168.825 ;
        RECT 44.790 168.800 46.775 169.800 ;
        RECT 60.400 169.775 61.400 169.800 ;
        RECT 66.600 169.775 67.600 169.800 ;
        RECT 68.500 169.775 69.500 169.800 ;
        RECT 60.380 168.825 61.420 169.775 ;
        RECT 66.580 168.825 67.620 169.775 ;
        RECT 68.480 168.825 69.520 169.775 ;
        RECT 60.400 168.800 61.400 168.825 ;
        RECT 66.600 168.800 67.600 168.825 ;
        RECT 68.500 168.800 69.500 168.825 ;
        RECT 70.215 168.800 72.200 169.800 ;
        RECT 85.825 169.775 86.825 169.800 ;
        RECT 92.025 169.775 93.025 169.800 ;
        RECT 93.925 169.775 94.925 169.800 ;
        RECT 85.805 168.825 86.845 169.775 ;
        RECT 92.005 168.825 93.045 169.775 ;
        RECT 93.905 168.825 94.945 169.775 ;
        RECT 85.825 168.800 86.825 168.825 ;
        RECT 92.025 168.800 93.025 168.825 ;
        RECT 93.925 168.800 94.925 168.825 ;
        RECT 95.640 168.800 97.625 169.800 ;
        RECT 111.250 169.775 112.250 169.800 ;
        RECT 117.450 169.775 118.450 169.800 ;
        RECT 119.350 169.775 120.350 169.800 ;
        RECT 111.230 168.825 112.270 169.775 ;
        RECT 117.430 168.825 118.470 169.775 ;
        RECT 119.330 168.825 120.370 169.775 ;
        RECT 111.250 168.800 112.250 168.825 ;
        RECT 117.450 168.800 118.450 168.825 ;
        RECT 119.350 168.800 120.350 168.825 ;
        RECT 121.065 168.800 123.050 169.800 ;
        RECT 136.675 169.775 137.675 169.800 ;
        RECT 142.875 169.775 143.875 169.800 ;
        RECT 144.775 169.775 145.775 169.800 ;
        RECT 136.655 168.825 137.695 169.775 ;
        RECT 142.855 168.825 143.895 169.775 ;
        RECT 144.755 168.825 145.795 169.775 ;
        RECT 136.675 168.800 137.675 168.825 ;
        RECT 142.875 168.800 143.875 168.825 ;
        RECT 144.775 168.800 145.775 168.825 ;
        RECT 146.490 168.800 148.475 169.800 ;
        RECT 19.370 168.780 21.325 168.800 ;
        RECT 44.795 168.780 46.750 168.800 ;
        RECT 70.220 168.780 72.175 168.800 ;
        RECT 95.645 168.780 97.600 168.800 ;
        RECT 121.070 168.780 123.025 168.800 ;
        RECT 146.495 168.780 148.450 168.800 ;
        RECT 9.575 167.025 10.525 167.045 ;
        RECT 20.375 167.025 21.325 167.045 ;
        RECT 35.000 167.025 35.950 167.045 ;
        RECT 45.800 167.025 46.750 167.045 ;
        RECT 60.425 167.025 61.375 167.045 ;
        RECT 71.225 167.025 72.175 167.045 ;
        RECT 85.850 167.025 86.800 167.045 ;
        RECT 96.650 167.025 97.600 167.045 ;
        RECT 111.275 167.025 112.225 167.045 ;
        RECT 122.075 167.025 123.025 167.045 ;
        RECT 136.700 167.025 137.650 167.045 ;
        RECT 147.500 167.025 148.450 167.045 ;
        RECT 9.550 166.025 12.755 167.025 ;
        RECT 13.530 166.025 14.620 167.025 ;
        RECT 15.370 166.025 18.650 167.025 ;
        RECT 20.350 166.025 21.350 167.025 ;
        RECT 9.575 166.005 10.525 166.025 ;
        RECT 2.900 165.075 7.100 165.080 ;
        RECT 1.850 163.975 12.025 165.075 ;
        RECT 13.575 165.050 14.575 166.025 ;
        RECT 20.375 166.005 21.325 166.025 ;
        RECT 23.155 165.730 24.155 166.825 ;
        RECT 34.975 166.025 38.180 167.025 ;
        RECT 38.955 166.025 40.045 167.025 ;
        RECT 40.795 166.025 44.075 167.025 ;
        RECT 45.775 166.025 46.775 167.025 ;
        RECT 35.000 166.005 35.950 166.025 ;
        RECT 23.430 165.115 23.880 165.730 ;
        RECT 28.325 165.075 32.525 165.080 ;
        RECT 12.650 164.050 14.575 165.050 ;
        RECT 16.175 164.155 22.100 165.075 ;
        RECT 27.275 164.155 37.450 165.075 ;
        RECT 39.000 165.050 40.000 166.025 ;
        RECT 45.800 166.005 46.750 166.025 ;
        RECT 48.580 165.730 49.580 166.825 ;
        RECT 60.400 166.025 63.605 167.025 ;
        RECT 64.380 166.025 65.470 167.025 ;
        RECT 66.220 166.025 69.500 167.025 ;
        RECT 71.200 166.025 72.200 167.025 ;
        RECT 60.425 166.005 61.375 166.025 ;
        RECT 48.855 165.115 49.305 165.730 ;
        RECT 53.750 165.075 57.950 165.080 ;
        RECT 1.850 163.970 11.290 163.975 ;
        RECT 6.050 157.825 7.050 163.970 ;
        RECT 12.650 162.675 13.650 164.050 ;
        RECT 16.175 163.975 37.450 164.155 ;
        RECT 38.075 164.050 40.000 165.050 ;
        RECT 41.600 164.155 47.525 165.075 ;
        RECT 52.700 164.155 62.875 165.075 ;
        RECT 64.425 165.050 65.425 166.025 ;
        RECT 71.225 166.005 72.175 166.025 ;
        RECT 74.005 165.730 75.005 166.825 ;
        RECT 85.825 166.025 89.030 167.025 ;
        RECT 89.805 166.025 90.895 167.025 ;
        RECT 91.645 166.025 94.925 167.025 ;
        RECT 96.625 166.025 97.625 167.025 ;
        RECT 85.850 166.005 86.800 166.025 ;
        RECT 74.280 165.115 74.730 165.730 ;
        RECT 79.175 165.075 83.375 165.080 ;
        RECT 16.890 163.970 19.400 163.975 ;
        RECT 19.590 163.970 36.715 163.975 ;
        RECT 20.320 163.050 28.380 163.970 ;
        RECT 12.630 161.725 13.670 162.675 ;
        RECT 12.650 161.700 13.650 161.725 ;
        RECT 14.405 161.700 15.495 162.700 ;
        RECT 6.050 156.825 7.075 157.825 ;
        RECT 7.550 156.825 8.495 157.350 ;
        RECT 6.570 155.700 7.610 156.175 ;
        RECT 1.900 155.325 2.900 155.355 ;
        RECT 6.570 155.325 7.075 155.700 ;
        RECT 7.920 155.370 8.495 156.825 ;
        RECT 1.850 155.300 7.075 155.325 ;
        RECT 1.850 154.350 7.095 155.300 ;
        RECT 1.850 154.325 7.075 154.350 ;
        RECT 1.900 154.295 2.900 154.325 ;
        RECT 6.570 153.950 7.075 154.325 ;
        RECT 7.500 154.280 8.500 155.370 ;
        RECT 9.460 155.325 9.830 161.350 ;
        RECT 8.825 154.325 9.830 155.325 ;
        RECT 6.570 153.455 7.610 153.950 ;
        RECT 7.920 153.050 8.495 154.280 ;
        RECT 6.075 152.675 7.130 153.050 ;
        RECT 7.550 152.675 8.495 153.050 ;
        RECT 3.890 149.285 5.030 149.315 ;
        RECT 6.075 149.285 7.075 152.675 ;
        RECT 8.830 151.125 9.830 154.325 ;
        RECT 7.630 150.125 9.830 151.125 ;
        RECT 10.250 155.370 10.620 161.350 ;
        RECT 14.450 160.925 15.450 160.955 ;
        RECT 14.450 159.925 17.220 160.925 ;
        RECT 14.450 159.895 15.450 159.925 ;
        RECT 11.475 156.825 12.475 159.275 ;
        RECT 12.950 156.825 13.895 157.350 ;
        RECT 14.175 156.825 15.175 159.275 ;
        RECT 15.650 156.825 16.595 157.350 ;
        RECT 11.970 155.700 13.010 156.175 ;
        RECT 10.250 155.325 11.250 155.370 ;
        RECT 11.970 155.325 12.475 155.700 ;
        RECT 13.320 155.325 13.895 156.825 ;
        RECT 14.670 155.700 15.710 156.175 ;
        RECT 14.670 155.325 15.175 155.700 ;
        RECT 16.020 155.325 16.595 156.825 ;
        RECT 17.560 155.325 17.930 161.350 ;
        RECT 18.350 155.325 18.720 161.350 ;
        RECT 20.260 155.325 20.630 161.350 ;
        RECT 10.250 155.300 12.475 155.325 ;
        RECT 10.250 154.355 12.495 155.300 ;
        RECT 10.250 154.325 12.475 154.355 ;
        RECT 12.855 154.325 15.175 155.325 ;
        RECT 15.600 154.325 17.930 155.325 ;
        RECT 18.305 154.325 19.395 155.325 ;
        RECT 19.625 154.325 20.630 155.325 ;
        RECT 10.250 154.280 11.250 154.325 ;
        RECT 10.250 150.125 10.620 154.280 ;
        RECT 11.970 153.950 12.475 154.325 ;
        RECT 11.970 153.455 13.010 153.950 ;
        RECT 13.320 153.050 13.895 154.325 ;
        RECT 14.670 153.950 15.175 154.325 ;
        RECT 14.670 153.455 15.710 153.950 ;
        RECT 16.020 153.050 16.595 154.325 ;
        RECT 11.475 152.675 12.530 153.050 ;
        RECT 12.950 152.675 13.895 153.050 ;
        RECT 14.175 152.675 15.230 153.050 ;
        RECT 15.650 152.675 16.595 153.050 ;
        RECT 11.475 151.800 12.475 152.675 ;
        RECT 14.175 151.800 15.175 152.675 ;
        RECT 11.475 150.800 15.175 151.800 ;
        RECT 15.750 151.125 16.750 151.170 ;
        RECT 16.930 151.125 17.930 154.325 ;
        RECT 11.475 149.285 12.475 150.800 ;
        RECT 15.750 150.125 17.930 151.125 ;
        RECT 18.350 150.125 18.720 154.325 ;
        RECT 19.630 153.325 20.630 154.325 ;
        RECT 21.050 155.325 21.420 161.350 ;
        RECT 31.475 157.825 32.475 163.970 ;
        RECT 38.075 162.675 39.075 164.050 ;
        RECT 41.600 163.975 62.875 164.155 ;
        RECT 63.500 164.050 65.425 165.050 ;
        RECT 67.025 164.155 72.950 165.075 ;
        RECT 78.125 164.155 88.300 165.075 ;
        RECT 89.850 165.050 90.850 166.025 ;
        RECT 96.650 166.005 97.600 166.025 ;
        RECT 99.430 165.730 100.430 166.825 ;
        RECT 111.250 166.025 114.455 167.025 ;
        RECT 115.230 166.025 116.320 167.025 ;
        RECT 117.070 166.025 120.350 167.025 ;
        RECT 122.050 166.025 123.050 167.025 ;
        RECT 111.275 166.005 112.225 166.025 ;
        RECT 99.705 165.115 100.155 165.730 ;
        RECT 104.600 165.075 108.800 165.080 ;
        RECT 42.315 163.970 44.825 163.975 ;
        RECT 45.015 163.970 62.140 163.975 ;
        RECT 45.745 163.050 53.805 163.970 ;
        RECT 38.055 161.725 39.095 162.675 ;
        RECT 38.075 161.700 39.075 161.725 ;
        RECT 39.830 161.700 40.920 162.700 ;
        RECT 31.475 156.825 32.500 157.825 ;
        RECT 32.975 156.825 33.920 157.350 ;
        RECT 23.430 155.875 23.880 156.515 ;
        RECT 23.150 155.325 24.150 155.875 ;
        RECT 31.995 155.700 33.035 156.175 ;
        RECT 27.325 155.325 28.325 155.355 ;
        RECT 31.995 155.325 32.500 155.700 ;
        RECT 33.345 155.370 33.920 156.825 ;
        RECT 21.050 154.325 24.150 155.325 ;
        RECT 27.275 155.300 32.500 155.325 ;
        RECT 27.275 154.350 32.520 155.300 ;
        RECT 27.275 154.325 32.500 154.350 ;
        RECT 19.585 152.325 20.675 153.325 ;
        RECT 20.260 150.125 20.630 152.325 ;
        RECT 21.050 150.125 21.420 154.325 ;
        RECT 23.430 154.205 23.880 154.325 ;
        RECT 27.325 154.295 28.325 154.325 ;
        RECT 31.995 153.950 32.500 154.325 ;
        RECT 32.925 154.280 33.925 155.370 ;
        RECT 34.885 155.325 35.255 161.350 ;
        RECT 34.250 154.325 35.255 155.325 ;
        RECT 31.995 153.455 33.035 153.950 ;
        RECT 33.345 153.050 33.920 154.280 ;
        RECT 31.500 152.675 32.555 153.050 ;
        RECT 32.975 152.675 33.920 153.050 ;
        RECT 15.750 150.080 16.750 150.125 ;
        RECT 29.315 149.285 30.455 149.315 ;
        RECT 31.500 149.285 32.500 152.675 ;
        RECT 34.255 151.125 35.255 154.325 ;
        RECT 33.055 150.125 35.255 151.125 ;
        RECT 35.675 155.370 36.045 161.350 ;
        RECT 39.875 160.925 40.875 160.955 ;
        RECT 39.875 159.925 42.645 160.925 ;
        RECT 39.875 159.895 40.875 159.925 ;
        RECT 36.900 156.825 37.900 159.275 ;
        RECT 38.375 156.825 39.320 157.350 ;
        RECT 39.600 156.825 40.600 159.275 ;
        RECT 41.075 156.825 42.020 157.350 ;
        RECT 37.395 155.700 38.435 156.175 ;
        RECT 35.675 155.325 36.675 155.370 ;
        RECT 37.395 155.325 37.900 155.700 ;
        RECT 38.745 155.325 39.320 156.825 ;
        RECT 40.095 155.700 41.135 156.175 ;
        RECT 40.095 155.325 40.600 155.700 ;
        RECT 41.445 155.325 42.020 156.825 ;
        RECT 42.985 155.325 43.355 161.350 ;
        RECT 43.775 155.325 44.145 161.350 ;
        RECT 45.685 155.325 46.055 161.350 ;
        RECT 35.675 155.300 37.900 155.325 ;
        RECT 35.675 154.355 37.920 155.300 ;
        RECT 35.675 154.325 37.900 154.355 ;
        RECT 38.280 154.325 40.600 155.325 ;
        RECT 41.025 154.325 43.355 155.325 ;
        RECT 43.730 154.325 44.820 155.325 ;
        RECT 45.050 154.325 46.055 155.325 ;
        RECT 35.675 154.280 36.675 154.325 ;
        RECT 35.675 150.125 36.045 154.280 ;
        RECT 37.395 153.950 37.900 154.325 ;
        RECT 37.395 153.455 38.435 153.950 ;
        RECT 38.745 153.050 39.320 154.325 ;
        RECT 40.095 153.950 40.600 154.325 ;
        RECT 40.095 153.455 41.135 153.950 ;
        RECT 41.445 153.050 42.020 154.325 ;
        RECT 36.900 152.675 37.955 153.050 ;
        RECT 38.375 152.675 39.320 153.050 ;
        RECT 39.600 152.675 40.655 153.050 ;
        RECT 41.075 152.675 42.020 153.050 ;
        RECT 36.900 151.800 37.900 152.675 ;
        RECT 39.600 151.800 40.600 152.675 ;
        RECT 36.900 150.800 40.600 151.800 ;
        RECT 41.175 151.125 42.175 151.170 ;
        RECT 42.355 151.125 43.355 154.325 ;
        RECT 36.900 149.285 37.900 150.800 ;
        RECT 41.175 150.125 43.355 151.125 ;
        RECT 43.775 150.125 44.145 154.325 ;
        RECT 45.055 153.325 46.055 154.325 ;
        RECT 46.475 155.325 46.845 161.350 ;
        RECT 56.900 157.825 57.900 163.970 ;
        RECT 63.500 162.675 64.500 164.050 ;
        RECT 67.025 163.975 88.300 164.155 ;
        RECT 88.925 164.050 90.850 165.050 ;
        RECT 92.450 164.155 98.375 165.075 ;
        RECT 103.550 164.155 113.725 165.075 ;
        RECT 115.275 165.050 116.275 166.025 ;
        RECT 122.075 166.005 123.025 166.025 ;
        RECT 124.855 165.730 125.855 166.825 ;
        RECT 136.675 166.025 139.880 167.025 ;
        RECT 140.655 166.025 141.745 167.025 ;
        RECT 142.495 166.025 145.775 167.025 ;
        RECT 147.475 166.025 148.475 167.025 ;
        RECT 136.700 166.005 137.650 166.025 ;
        RECT 125.130 165.115 125.580 165.730 ;
        RECT 130.025 165.075 134.225 165.080 ;
        RECT 67.740 163.970 70.250 163.975 ;
        RECT 70.440 163.970 87.565 163.975 ;
        RECT 71.170 163.050 79.230 163.970 ;
        RECT 63.480 161.725 64.520 162.675 ;
        RECT 63.500 161.700 64.500 161.725 ;
        RECT 65.255 161.700 66.345 162.700 ;
        RECT 56.900 156.825 57.925 157.825 ;
        RECT 58.400 156.825 59.345 157.350 ;
        RECT 48.855 155.875 49.305 156.515 ;
        RECT 48.575 155.325 49.575 155.875 ;
        RECT 57.420 155.700 58.460 156.175 ;
        RECT 52.750 155.325 53.750 155.355 ;
        RECT 57.420 155.325 57.925 155.700 ;
        RECT 58.770 155.370 59.345 156.825 ;
        RECT 46.475 154.325 49.575 155.325 ;
        RECT 52.700 155.300 57.925 155.325 ;
        RECT 52.700 154.350 57.945 155.300 ;
        RECT 52.700 154.325 57.925 154.350 ;
        RECT 45.010 152.325 46.100 153.325 ;
        RECT 45.685 150.125 46.055 152.325 ;
        RECT 46.475 150.125 46.845 154.325 ;
        RECT 48.855 154.205 49.305 154.325 ;
        RECT 52.750 154.295 53.750 154.325 ;
        RECT 57.420 153.950 57.925 154.325 ;
        RECT 58.350 154.280 59.350 155.370 ;
        RECT 60.310 155.325 60.680 161.350 ;
        RECT 59.675 154.325 60.680 155.325 ;
        RECT 57.420 153.455 58.460 153.950 ;
        RECT 58.770 153.050 59.345 154.280 ;
        RECT 56.925 152.675 57.980 153.050 ;
        RECT 58.400 152.675 59.345 153.050 ;
        RECT 41.175 150.080 42.175 150.125 ;
        RECT 54.740 149.285 55.880 149.315 ;
        RECT 56.925 149.285 57.925 152.675 ;
        RECT 59.680 151.125 60.680 154.325 ;
        RECT 58.480 150.125 60.680 151.125 ;
        RECT 61.100 155.370 61.470 161.350 ;
        RECT 65.300 160.925 66.300 160.955 ;
        RECT 65.300 159.925 68.070 160.925 ;
        RECT 65.300 159.895 66.300 159.925 ;
        RECT 62.325 156.825 63.325 159.275 ;
        RECT 63.800 156.825 64.745 157.350 ;
        RECT 65.025 156.825 66.025 159.275 ;
        RECT 66.500 156.825 67.445 157.350 ;
        RECT 62.820 155.700 63.860 156.175 ;
        RECT 61.100 155.325 62.100 155.370 ;
        RECT 62.820 155.325 63.325 155.700 ;
        RECT 64.170 155.325 64.745 156.825 ;
        RECT 65.520 155.700 66.560 156.175 ;
        RECT 65.520 155.325 66.025 155.700 ;
        RECT 66.870 155.325 67.445 156.825 ;
        RECT 68.410 155.325 68.780 161.350 ;
        RECT 69.200 155.325 69.570 161.350 ;
        RECT 71.110 155.325 71.480 161.350 ;
        RECT 61.100 155.300 63.325 155.325 ;
        RECT 61.100 154.355 63.345 155.300 ;
        RECT 61.100 154.325 63.325 154.355 ;
        RECT 63.705 154.325 66.025 155.325 ;
        RECT 66.450 154.325 68.780 155.325 ;
        RECT 69.155 154.325 70.245 155.325 ;
        RECT 70.475 154.325 71.480 155.325 ;
        RECT 61.100 154.280 62.100 154.325 ;
        RECT 61.100 150.125 61.470 154.280 ;
        RECT 62.820 153.950 63.325 154.325 ;
        RECT 62.820 153.455 63.860 153.950 ;
        RECT 64.170 153.050 64.745 154.325 ;
        RECT 65.520 153.950 66.025 154.325 ;
        RECT 65.520 153.455 66.560 153.950 ;
        RECT 66.870 153.050 67.445 154.325 ;
        RECT 62.325 152.675 63.380 153.050 ;
        RECT 63.800 152.675 64.745 153.050 ;
        RECT 65.025 152.675 66.080 153.050 ;
        RECT 66.500 152.675 67.445 153.050 ;
        RECT 62.325 151.800 63.325 152.675 ;
        RECT 65.025 151.800 66.025 152.675 ;
        RECT 62.325 150.800 66.025 151.800 ;
        RECT 66.600 151.125 67.600 151.170 ;
        RECT 67.780 151.125 68.780 154.325 ;
        RECT 62.325 149.285 63.325 150.800 ;
        RECT 66.600 150.125 68.780 151.125 ;
        RECT 69.200 150.125 69.570 154.325 ;
        RECT 70.480 153.325 71.480 154.325 ;
        RECT 71.900 155.325 72.270 161.350 ;
        RECT 82.325 157.825 83.325 163.970 ;
        RECT 88.925 162.675 89.925 164.050 ;
        RECT 92.450 163.975 113.725 164.155 ;
        RECT 114.350 164.050 116.275 165.050 ;
        RECT 117.875 164.155 123.800 165.075 ;
        RECT 128.975 164.155 139.150 165.075 ;
        RECT 140.700 165.050 141.700 166.025 ;
        RECT 147.500 166.005 148.450 166.025 ;
        RECT 150.280 165.730 151.280 166.825 ;
        RECT 150.555 165.115 151.005 165.730 ;
        RECT 93.165 163.970 95.675 163.975 ;
        RECT 95.865 163.970 112.990 163.975 ;
        RECT 96.595 163.050 104.655 163.970 ;
        RECT 88.905 161.725 89.945 162.675 ;
        RECT 88.925 161.700 89.925 161.725 ;
        RECT 90.680 161.700 91.770 162.700 ;
        RECT 82.325 156.825 83.350 157.825 ;
        RECT 83.825 156.825 84.770 157.350 ;
        RECT 74.280 155.875 74.730 156.515 ;
        RECT 74.000 155.325 75.000 155.875 ;
        RECT 82.845 155.700 83.885 156.175 ;
        RECT 78.175 155.325 79.175 155.355 ;
        RECT 82.845 155.325 83.350 155.700 ;
        RECT 84.195 155.370 84.770 156.825 ;
        RECT 71.900 154.325 75.000 155.325 ;
        RECT 78.125 155.300 83.350 155.325 ;
        RECT 78.125 154.350 83.370 155.300 ;
        RECT 78.125 154.325 83.350 154.350 ;
        RECT 70.435 152.325 71.525 153.325 ;
        RECT 71.110 150.125 71.480 152.325 ;
        RECT 71.900 150.125 72.270 154.325 ;
        RECT 74.280 154.205 74.730 154.325 ;
        RECT 78.175 154.295 79.175 154.325 ;
        RECT 82.845 153.950 83.350 154.325 ;
        RECT 83.775 154.280 84.775 155.370 ;
        RECT 85.735 155.325 86.105 161.350 ;
        RECT 85.100 154.325 86.105 155.325 ;
        RECT 82.845 153.455 83.885 153.950 ;
        RECT 84.195 153.050 84.770 154.280 ;
        RECT 82.350 152.675 83.405 153.050 ;
        RECT 83.825 152.675 84.770 153.050 ;
        RECT 66.600 150.080 67.600 150.125 ;
        RECT 80.165 149.285 81.305 149.315 ;
        RECT 82.350 149.285 83.350 152.675 ;
        RECT 85.105 151.125 86.105 154.325 ;
        RECT 83.905 150.125 86.105 151.125 ;
        RECT 86.525 155.370 86.895 161.350 ;
        RECT 90.725 160.925 91.725 160.955 ;
        RECT 90.725 159.925 93.495 160.925 ;
        RECT 90.725 159.895 91.725 159.925 ;
        RECT 87.750 156.825 88.750 159.275 ;
        RECT 89.225 156.825 90.170 157.350 ;
        RECT 90.450 156.825 91.450 159.275 ;
        RECT 91.925 156.825 92.870 157.350 ;
        RECT 88.245 155.700 89.285 156.175 ;
        RECT 86.525 155.325 87.525 155.370 ;
        RECT 88.245 155.325 88.750 155.700 ;
        RECT 89.595 155.325 90.170 156.825 ;
        RECT 90.945 155.700 91.985 156.175 ;
        RECT 90.945 155.325 91.450 155.700 ;
        RECT 92.295 155.325 92.870 156.825 ;
        RECT 93.835 155.325 94.205 161.350 ;
        RECT 94.625 155.325 94.995 161.350 ;
        RECT 96.535 155.325 96.905 161.350 ;
        RECT 86.525 155.300 88.750 155.325 ;
        RECT 86.525 154.355 88.770 155.300 ;
        RECT 86.525 154.325 88.750 154.355 ;
        RECT 89.130 154.325 91.450 155.325 ;
        RECT 91.875 154.325 94.205 155.325 ;
        RECT 94.580 154.325 95.670 155.325 ;
        RECT 95.900 154.325 96.905 155.325 ;
        RECT 86.525 154.280 87.525 154.325 ;
        RECT 86.525 150.125 86.895 154.280 ;
        RECT 88.245 153.950 88.750 154.325 ;
        RECT 88.245 153.455 89.285 153.950 ;
        RECT 89.595 153.050 90.170 154.325 ;
        RECT 90.945 153.950 91.450 154.325 ;
        RECT 90.945 153.455 91.985 153.950 ;
        RECT 92.295 153.050 92.870 154.325 ;
        RECT 87.750 152.675 88.805 153.050 ;
        RECT 89.225 152.675 90.170 153.050 ;
        RECT 90.450 152.675 91.505 153.050 ;
        RECT 91.925 152.675 92.870 153.050 ;
        RECT 87.750 151.800 88.750 152.675 ;
        RECT 90.450 151.800 91.450 152.675 ;
        RECT 87.750 150.800 91.450 151.800 ;
        RECT 92.025 151.125 93.025 151.170 ;
        RECT 93.205 151.125 94.205 154.325 ;
        RECT 87.750 149.285 88.750 150.800 ;
        RECT 92.025 150.125 94.205 151.125 ;
        RECT 94.625 150.125 94.995 154.325 ;
        RECT 95.905 153.325 96.905 154.325 ;
        RECT 97.325 155.325 97.695 161.350 ;
        RECT 107.750 157.825 108.750 163.970 ;
        RECT 114.350 162.675 115.350 164.050 ;
        RECT 117.875 163.975 139.150 164.155 ;
        RECT 139.775 164.050 141.700 165.050 ;
        RECT 118.590 163.970 121.100 163.975 ;
        RECT 121.290 163.970 138.415 163.975 ;
        RECT 122.020 163.050 130.080 163.970 ;
        RECT 114.330 161.725 115.370 162.675 ;
        RECT 114.350 161.700 115.350 161.725 ;
        RECT 116.105 161.700 117.195 162.700 ;
        RECT 107.750 156.825 108.775 157.825 ;
        RECT 109.250 156.825 110.195 157.350 ;
        RECT 99.705 155.875 100.155 156.515 ;
        RECT 99.425 155.325 100.425 155.875 ;
        RECT 108.270 155.700 109.310 156.175 ;
        RECT 103.600 155.325 104.600 155.355 ;
        RECT 108.270 155.325 108.775 155.700 ;
        RECT 109.620 155.370 110.195 156.825 ;
        RECT 97.325 154.325 100.425 155.325 ;
        RECT 103.550 155.300 108.775 155.325 ;
        RECT 103.550 154.350 108.795 155.300 ;
        RECT 103.550 154.325 108.775 154.350 ;
        RECT 95.860 152.325 96.950 153.325 ;
        RECT 96.535 150.125 96.905 152.325 ;
        RECT 97.325 150.125 97.695 154.325 ;
        RECT 99.705 154.205 100.155 154.325 ;
        RECT 103.600 154.295 104.600 154.325 ;
        RECT 108.270 153.950 108.775 154.325 ;
        RECT 109.200 154.280 110.200 155.370 ;
        RECT 111.160 155.325 111.530 161.350 ;
        RECT 110.525 154.325 111.530 155.325 ;
        RECT 108.270 153.455 109.310 153.950 ;
        RECT 109.620 153.050 110.195 154.280 ;
        RECT 107.775 152.675 108.830 153.050 ;
        RECT 109.250 152.675 110.195 153.050 ;
        RECT 92.025 150.080 93.025 150.125 ;
        RECT 105.590 149.285 106.730 149.315 ;
        RECT 107.775 149.285 108.775 152.675 ;
        RECT 110.530 151.125 111.530 154.325 ;
        RECT 109.330 150.125 111.530 151.125 ;
        RECT 111.950 155.370 112.320 161.350 ;
        RECT 116.150 160.925 117.150 160.955 ;
        RECT 116.150 159.925 118.920 160.925 ;
        RECT 116.150 159.895 117.150 159.925 ;
        RECT 113.175 156.825 114.175 159.275 ;
        RECT 114.650 156.825 115.595 157.350 ;
        RECT 115.875 156.825 116.875 159.275 ;
        RECT 117.350 156.825 118.295 157.350 ;
        RECT 113.670 155.700 114.710 156.175 ;
        RECT 111.950 155.325 112.950 155.370 ;
        RECT 113.670 155.325 114.175 155.700 ;
        RECT 115.020 155.325 115.595 156.825 ;
        RECT 116.370 155.700 117.410 156.175 ;
        RECT 116.370 155.325 116.875 155.700 ;
        RECT 117.720 155.325 118.295 156.825 ;
        RECT 119.260 155.325 119.630 161.350 ;
        RECT 120.050 155.325 120.420 161.350 ;
        RECT 121.960 155.325 122.330 161.350 ;
        RECT 111.950 155.300 114.175 155.325 ;
        RECT 111.950 154.355 114.195 155.300 ;
        RECT 111.950 154.325 114.175 154.355 ;
        RECT 114.555 154.325 116.875 155.325 ;
        RECT 117.300 154.325 119.630 155.325 ;
        RECT 120.005 154.325 121.095 155.325 ;
        RECT 121.325 154.325 122.330 155.325 ;
        RECT 111.950 154.280 112.950 154.325 ;
        RECT 111.950 150.125 112.320 154.280 ;
        RECT 113.670 153.950 114.175 154.325 ;
        RECT 113.670 153.455 114.710 153.950 ;
        RECT 115.020 153.050 115.595 154.325 ;
        RECT 116.370 153.950 116.875 154.325 ;
        RECT 116.370 153.455 117.410 153.950 ;
        RECT 117.720 153.050 118.295 154.325 ;
        RECT 113.175 152.675 114.230 153.050 ;
        RECT 114.650 152.675 115.595 153.050 ;
        RECT 115.875 152.675 116.930 153.050 ;
        RECT 117.350 152.675 118.295 153.050 ;
        RECT 113.175 151.800 114.175 152.675 ;
        RECT 115.875 151.800 116.875 152.675 ;
        RECT 113.175 150.800 116.875 151.800 ;
        RECT 117.450 151.125 118.450 151.170 ;
        RECT 118.630 151.125 119.630 154.325 ;
        RECT 113.175 149.285 114.175 150.800 ;
        RECT 117.450 150.125 119.630 151.125 ;
        RECT 120.050 150.125 120.420 154.325 ;
        RECT 121.330 153.325 122.330 154.325 ;
        RECT 122.750 155.325 123.120 161.350 ;
        RECT 133.175 157.825 134.175 163.970 ;
        RECT 139.775 162.675 140.775 164.050 ;
        RECT 143.300 163.975 149.225 165.075 ;
        RECT 144.015 163.970 146.525 163.975 ;
        RECT 146.715 163.970 149.215 163.975 ;
        RECT 139.755 161.725 140.795 162.675 ;
        RECT 139.775 161.700 140.775 161.725 ;
        RECT 141.530 161.700 142.620 162.700 ;
        RECT 133.175 156.825 134.200 157.825 ;
        RECT 134.675 156.825 135.620 157.350 ;
        RECT 125.130 155.875 125.580 156.515 ;
        RECT 124.850 155.325 125.850 155.875 ;
        RECT 133.695 155.700 134.735 156.175 ;
        RECT 129.025 155.325 130.025 155.355 ;
        RECT 133.695 155.325 134.200 155.700 ;
        RECT 135.045 155.370 135.620 156.825 ;
        RECT 122.750 154.325 125.850 155.325 ;
        RECT 128.975 155.300 134.200 155.325 ;
        RECT 128.975 154.350 134.220 155.300 ;
        RECT 128.975 154.325 134.200 154.350 ;
        RECT 121.285 152.325 122.375 153.325 ;
        RECT 121.960 150.125 122.330 152.325 ;
        RECT 122.750 150.125 123.120 154.325 ;
        RECT 125.130 154.205 125.580 154.325 ;
        RECT 129.025 154.295 130.025 154.325 ;
        RECT 133.695 153.950 134.200 154.325 ;
        RECT 134.625 154.280 135.625 155.370 ;
        RECT 136.585 155.325 136.955 161.350 ;
        RECT 135.950 154.325 136.955 155.325 ;
        RECT 133.695 153.455 134.735 153.950 ;
        RECT 135.045 153.050 135.620 154.280 ;
        RECT 133.200 152.675 134.255 153.050 ;
        RECT 134.675 152.675 135.620 153.050 ;
        RECT 117.450 150.080 118.450 150.125 ;
        RECT 131.015 149.285 132.155 149.315 ;
        RECT 133.200 149.285 134.200 152.675 ;
        RECT 135.955 151.125 136.955 154.325 ;
        RECT 134.755 150.125 136.955 151.125 ;
        RECT 137.375 155.370 137.745 161.350 ;
        RECT 141.575 160.925 142.575 160.955 ;
        RECT 141.575 159.925 144.345 160.925 ;
        RECT 141.575 159.895 142.575 159.925 ;
        RECT 138.600 156.825 139.600 159.275 ;
        RECT 140.075 156.825 141.020 157.350 ;
        RECT 141.300 156.825 142.300 159.275 ;
        RECT 142.775 156.825 143.720 157.350 ;
        RECT 139.095 155.700 140.135 156.175 ;
        RECT 137.375 155.325 138.375 155.370 ;
        RECT 139.095 155.325 139.600 155.700 ;
        RECT 140.445 155.325 141.020 156.825 ;
        RECT 141.795 155.700 142.835 156.175 ;
        RECT 141.795 155.325 142.300 155.700 ;
        RECT 143.145 155.325 143.720 156.825 ;
        RECT 144.685 155.325 145.055 161.350 ;
        RECT 145.475 155.325 145.845 161.350 ;
        RECT 147.385 155.325 147.755 161.350 ;
        RECT 137.375 155.300 139.600 155.325 ;
        RECT 137.375 154.355 139.620 155.300 ;
        RECT 137.375 154.325 139.600 154.355 ;
        RECT 139.980 154.325 142.300 155.325 ;
        RECT 142.725 154.325 145.055 155.325 ;
        RECT 145.430 154.325 146.520 155.325 ;
        RECT 146.750 154.325 147.755 155.325 ;
        RECT 137.375 154.280 138.375 154.325 ;
        RECT 137.375 150.125 137.745 154.280 ;
        RECT 139.095 153.950 139.600 154.325 ;
        RECT 139.095 153.455 140.135 153.950 ;
        RECT 140.445 153.050 141.020 154.325 ;
        RECT 141.795 153.950 142.300 154.325 ;
        RECT 141.795 153.455 142.835 153.950 ;
        RECT 143.145 153.050 143.720 154.325 ;
        RECT 138.600 152.675 139.655 153.050 ;
        RECT 140.075 152.675 141.020 153.050 ;
        RECT 141.300 152.675 142.355 153.050 ;
        RECT 142.775 152.675 143.720 153.050 ;
        RECT 138.600 151.800 139.600 152.675 ;
        RECT 141.300 151.800 142.300 152.675 ;
        RECT 138.600 150.800 142.300 151.800 ;
        RECT 142.875 151.125 143.875 151.170 ;
        RECT 144.055 151.125 145.055 154.325 ;
        RECT 138.600 149.285 139.600 150.800 ;
        RECT 142.875 150.125 145.055 151.125 ;
        RECT 145.475 150.125 145.845 154.325 ;
        RECT 146.755 153.325 147.755 154.325 ;
        RECT 148.175 155.325 148.545 161.350 ;
        RECT 150.555 155.875 151.005 156.515 ;
        RECT 150.275 155.325 151.275 155.875 ;
        RECT 148.175 154.325 151.275 155.325 ;
        RECT 146.710 152.325 147.800 153.325 ;
        RECT 147.385 150.125 147.755 152.325 ;
        RECT 148.175 150.125 148.545 154.325 ;
        RECT 150.555 154.205 151.005 154.325 ;
        RECT 142.875 150.080 143.875 150.125 ;
        RECT 1.850 149.275 14.575 149.285 ;
        RECT 15.350 149.275 19.390 149.285 ;
        RECT 19.590 149.275 40.000 149.285 ;
        RECT 40.775 149.275 44.815 149.285 ;
        RECT 45.015 149.275 65.425 149.285 ;
        RECT 66.200 149.275 70.240 149.285 ;
        RECT 70.440 149.275 90.850 149.285 ;
        RECT 91.625 149.275 95.665 149.285 ;
        RECT 95.865 149.275 116.275 149.285 ;
        RECT 117.050 149.275 121.090 149.285 ;
        RECT 121.290 149.275 141.700 149.285 ;
        RECT 142.475 149.275 146.515 149.285 ;
        RECT 146.715 149.275 151.360 149.285 ;
        RECT 1.850 148.175 151.360 149.275 ;
        RECT 1.850 148.170 19.390 148.175 ;
        RECT 19.590 148.170 44.815 148.175 ;
        RECT 45.015 148.170 70.240 148.175 ;
        RECT 70.440 148.170 95.665 148.175 ;
        RECT 95.865 148.170 121.090 148.175 ;
        RECT 121.290 148.170 146.515 148.175 ;
        RECT 146.715 148.170 151.360 148.175 ;
        RECT 3.890 148.140 5.030 148.170 ;
        RECT 29.315 148.140 30.455 148.170 ;
        RECT 54.740 148.140 55.880 148.170 ;
        RECT 80.165 148.140 81.305 148.170 ;
        RECT 105.590 148.140 106.730 148.170 ;
        RECT 131.015 148.140 132.155 148.170 ;
        RECT 19.370 147.225 21.325 147.245 ;
        RECT 44.795 147.225 46.750 147.245 ;
        RECT 70.220 147.225 72.175 147.245 ;
        RECT 95.645 147.225 97.600 147.245 ;
        RECT 121.070 147.225 123.025 147.245 ;
        RECT 146.495 147.225 148.450 147.245 ;
        RECT 9.550 147.200 10.550 147.225 ;
        RECT 15.750 147.200 16.750 147.225 ;
        RECT 17.650 147.200 18.650 147.225 ;
        RECT 9.530 146.250 10.570 147.200 ;
        RECT 15.730 146.250 16.770 147.200 ;
        RECT 17.630 146.250 18.670 147.200 ;
        RECT 9.550 146.225 10.550 146.250 ;
        RECT 15.750 146.225 16.750 146.250 ;
        RECT 17.650 146.225 18.650 146.250 ;
        RECT 19.365 146.225 21.350 147.225 ;
        RECT 34.975 147.200 35.975 147.225 ;
        RECT 41.175 147.200 42.175 147.225 ;
        RECT 43.075 147.200 44.075 147.225 ;
        RECT 34.955 146.250 35.995 147.200 ;
        RECT 41.155 146.250 42.195 147.200 ;
        RECT 43.055 146.250 44.095 147.200 ;
        RECT 34.975 146.225 35.975 146.250 ;
        RECT 41.175 146.225 42.175 146.250 ;
        RECT 43.075 146.225 44.075 146.250 ;
        RECT 44.790 146.225 46.775 147.225 ;
        RECT 60.400 147.200 61.400 147.225 ;
        RECT 66.600 147.200 67.600 147.225 ;
        RECT 68.500 147.200 69.500 147.225 ;
        RECT 60.380 146.250 61.420 147.200 ;
        RECT 66.580 146.250 67.620 147.200 ;
        RECT 68.480 146.250 69.520 147.200 ;
        RECT 60.400 146.225 61.400 146.250 ;
        RECT 66.600 146.225 67.600 146.250 ;
        RECT 68.500 146.225 69.500 146.250 ;
        RECT 70.215 146.225 72.200 147.225 ;
        RECT 85.825 147.200 86.825 147.225 ;
        RECT 92.025 147.200 93.025 147.225 ;
        RECT 93.925 147.200 94.925 147.225 ;
        RECT 85.805 146.250 86.845 147.200 ;
        RECT 92.005 146.250 93.045 147.200 ;
        RECT 93.905 146.250 94.945 147.200 ;
        RECT 85.825 146.225 86.825 146.250 ;
        RECT 92.025 146.225 93.025 146.250 ;
        RECT 93.925 146.225 94.925 146.250 ;
        RECT 95.640 146.225 97.625 147.225 ;
        RECT 111.250 147.200 112.250 147.225 ;
        RECT 117.450 147.200 118.450 147.225 ;
        RECT 119.350 147.200 120.350 147.225 ;
        RECT 111.230 146.250 112.270 147.200 ;
        RECT 117.430 146.250 118.470 147.200 ;
        RECT 119.330 146.250 120.370 147.200 ;
        RECT 111.250 146.225 112.250 146.250 ;
        RECT 117.450 146.225 118.450 146.250 ;
        RECT 119.350 146.225 120.350 146.250 ;
        RECT 121.065 146.225 123.050 147.225 ;
        RECT 136.675 147.200 137.675 147.225 ;
        RECT 142.875 147.200 143.875 147.225 ;
        RECT 144.775 147.200 145.775 147.225 ;
        RECT 136.655 146.250 137.695 147.200 ;
        RECT 142.855 146.250 143.895 147.200 ;
        RECT 144.755 146.250 145.795 147.200 ;
        RECT 136.675 146.225 137.675 146.250 ;
        RECT 142.875 146.225 143.875 146.250 ;
        RECT 144.775 146.225 145.775 146.250 ;
        RECT 146.490 146.225 148.475 147.225 ;
        RECT 19.370 146.205 21.325 146.225 ;
        RECT 44.795 146.205 46.750 146.225 ;
        RECT 70.220 146.205 72.175 146.225 ;
        RECT 95.645 146.205 97.600 146.225 ;
        RECT 121.070 146.205 123.025 146.225 ;
        RECT 146.495 146.205 148.450 146.225 ;
        RECT 23.545 142.550 24.495 142.570 ;
        RECT 74.395 142.550 75.345 142.570 ;
        RECT 99.700 142.550 100.650 142.570 ;
        RECT 125.245 142.550 126.195 142.570 ;
        RECT 23.525 141.550 126.215 142.550 ;
        RECT 23.545 141.530 24.495 141.550 ;
        RECT 74.395 141.530 75.345 141.550 ;
        RECT 99.700 141.530 100.650 141.550 ;
        RECT 125.245 141.530 126.195 141.550 ;
        RECT 9.575 140.175 10.525 140.195 ;
        RECT 20.375 140.175 21.325 140.195 ;
        RECT 9.550 139.175 12.755 140.175 ;
        RECT 13.530 139.175 14.620 140.175 ;
        RECT 15.370 139.175 18.650 140.175 ;
        RECT 20.350 139.175 21.350 140.175 ;
        RECT 21.795 140.000 32.470 141.000 ;
        RECT 35.000 140.175 35.950 140.195 ;
        RECT 45.800 140.175 46.750 140.195 ;
        RECT 60.425 140.175 61.375 140.195 ;
        RECT 71.225 140.175 72.175 140.195 ;
        RECT 9.575 139.155 10.525 139.175 ;
        RECT 5.995 138.225 7.100 138.270 ;
        RECT 5.965 137.125 12.025 138.225 ;
        RECT 13.575 138.200 14.575 139.175 ;
        RECT 20.375 139.155 21.325 139.175 ;
        RECT 21.795 138.225 22.795 140.000 ;
        RECT 23.520 138.325 24.520 139.220 ;
        RECT 12.650 137.200 14.575 138.200 ;
        RECT 5.965 137.120 11.290 137.125 ;
        RECT 5.995 137.075 7.100 137.120 ;
        RECT 6.050 130.975 7.050 137.075 ;
        RECT 12.650 135.825 13.650 137.200 ;
        RECT 16.175 137.150 22.795 138.225 ;
        RECT 23.490 137.325 24.550 138.325 ;
        RECT 16.175 137.125 22.100 137.150 ;
        RECT 16.890 137.120 19.400 137.125 ;
        RECT 19.590 137.120 22.090 137.125 ;
        RECT 24.870 136.575 25.870 139.525 ;
        RECT 27.145 138.975 29.170 140.000 ;
        RECT 29.645 138.975 30.590 139.500 ;
        RECT 27.145 138.945 28.145 138.975 ;
        RECT 26.245 138.295 27.245 138.340 ;
        RECT 26.215 137.295 27.275 138.295 ;
        RECT 28.665 137.850 29.705 138.325 ;
        RECT 28.665 137.475 29.170 137.850 ;
        RECT 30.015 137.475 30.590 138.975 ;
        RECT 31.470 138.270 32.470 140.000 ;
        RECT 34.975 139.175 38.180 140.175 ;
        RECT 38.955 139.175 40.045 140.175 ;
        RECT 40.795 139.175 44.075 140.175 ;
        RECT 45.775 139.175 46.775 140.175 ;
        RECT 60.400 139.175 63.605 140.175 ;
        RECT 64.380 139.175 65.470 140.175 ;
        RECT 66.220 139.175 69.500 140.175 ;
        RECT 71.200 139.175 72.200 140.175 ;
        RECT 72.645 140.000 83.320 141.000 ;
        RECT 85.850 140.175 86.800 140.195 ;
        RECT 96.650 140.175 97.600 140.195 ;
        RECT 111.275 140.175 112.225 140.195 ;
        RECT 122.075 140.175 123.025 140.195 ;
        RECT 35.000 139.155 35.950 139.175 ;
        RECT 31.420 138.225 32.525 138.270 ;
        RECT 26.245 137.250 27.245 137.295 ;
        RECT 28.170 136.575 29.170 137.475 ;
        RECT 16.175 136.340 17.175 136.385 ;
        RECT 20.370 136.340 21.320 136.360 ;
        RECT 12.630 134.875 13.670 135.825 ;
        RECT 12.650 134.850 13.650 134.875 ;
        RECT 14.405 134.850 15.495 135.850 ;
        RECT 16.175 135.340 21.345 136.340 ;
        RECT 24.870 136.100 29.170 136.575 ;
        RECT 29.550 136.475 30.640 137.475 ;
        RECT 31.390 137.125 37.450 138.225 ;
        RECT 39.000 138.200 40.000 139.175 ;
        RECT 45.800 139.155 46.750 139.175 ;
        RECT 60.425 139.155 61.375 139.175 ;
        RECT 56.845 138.225 57.950 138.270 ;
        RECT 38.075 137.200 40.000 138.200 ;
        RECT 31.390 137.120 36.715 137.125 ;
        RECT 31.420 137.075 32.525 137.120 ;
        RECT 24.870 135.650 29.705 136.100 ;
        RECT 23.020 135.605 29.705 135.650 ;
        RECT 23.020 135.575 29.170 135.605 ;
        RECT 16.175 135.295 17.175 135.340 ;
        RECT 20.370 135.320 21.320 135.340 ;
        RECT 23.020 134.650 25.870 135.575 ;
        RECT 27.145 135.200 28.145 135.230 ;
        RECT 30.015 135.200 30.590 136.475 ;
        RECT 27.145 134.825 29.225 135.200 ;
        RECT 29.645 134.825 30.590 135.200 ;
        RECT 6.050 129.975 7.075 130.975 ;
        RECT 7.550 129.975 8.495 130.500 ;
        RECT 6.570 128.850 7.610 129.325 ;
        RECT 3.950 128.500 4.950 128.505 ;
        RECT 3.920 128.475 4.980 128.500 ;
        RECT 6.570 128.475 7.075 128.850 ;
        RECT 7.920 128.520 8.495 129.975 ;
        RECT 3.875 128.450 7.075 128.475 ;
        RECT 3.875 127.500 7.095 128.450 ;
        RECT 3.875 127.475 7.075 127.500 ;
        RECT 3.950 127.445 4.950 127.475 ;
        RECT 6.570 127.100 7.075 127.475 ;
        RECT 7.500 127.430 8.500 128.520 ;
        RECT 9.460 128.475 9.830 134.500 ;
        RECT 8.825 127.475 9.830 128.475 ;
        RECT 6.570 126.605 7.610 127.100 ;
        RECT 7.920 126.200 8.495 127.430 ;
        RECT 6.075 125.825 7.130 126.200 ;
        RECT 7.550 125.825 8.495 126.200 ;
        RECT 3.905 122.455 5.020 122.460 ;
        RECT 3.875 122.435 5.050 122.455 ;
        RECT 6.075 122.435 7.075 125.825 ;
        RECT 8.830 124.275 9.830 127.475 ;
        RECT 7.630 123.275 9.830 124.275 ;
        RECT 10.250 128.520 10.620 134.500 ;
        RECT 14.450 134.075 15.450 134.105 ;
        RECT 14.450 133.075 17.220 134.075 ;
        RECT 14.450 133.045 15.450 133.075 ;
        RECT 11.475 129.975 12.475 132.425 ;
        RECT 12.950 129.975 13.895 130.500 ;
        RECT 14.175 129.975 15.175 132.425 ;
        RECT 15.650 129.975 16.595 130.500 ;
        RECT 11.970 128.850 13.010 129.325 ;
        RECT 10.250 128.475 11.250 128.520 ;
        RECT 11.970 128.475 12.475 128.850 ;
        RECT 13.320 128.475 13.895 129.975 ;
        RECT 14.670 128.850 15.710 129.325 ;
        RECT 14.670 128.475 15.175 128.850 ;
        RECT 16.020 128.475 16.595 129.975 ;
        RECT 17.560 128.475 17.930 134.500 ;
        RECT 18.350 128.475 18.720 134.500 ;
        RECT 20.260 128.475 20.630 134.500 ;
        RECT 10.250 128.450 12.475 128.475 ;
        RECT 10.250 127.505 12.495 128.450 ;
        RECT 10.250 127.475 12.475 127.505 ;
        RECT 12.855 127.475 15.175 128.475 ;
        RECT 15.600 127.475 17.930 128.475 ;
        RECT 18.305 127.475 19.395 128.475 ;
        RECT 10.250 127.430 11.250 127.475 ;
        RECT 10.250 123.275 10.620 127.430 ;
        RECT 11.970 127.100 12.475 127.475 ;
        RECT 11.970 126.605 13.010 127.100 ;
        RECT 13.320 126.200 13.895 127.475 ;
        RECT 14.670 127.100 15.175 127.475 ;
        RECT 14.670 126.605 15.710 127.100 ;
        RECT 16.020 126.200 16.595 127.475 ;
        RECT 11.475 125.825 12.530 126.200 ;
        RECT 12.950 125.825 13.895 126.200 ;
        RECT 14.175 125.825 15.230 126.200 ;
        RECT 15.650 125.825 16.595 126.200 ;
        RECT 11.475 124.950 12.475 125.825 ;
        RECT 14.175 124.950 15.175 125.825 ;
        RECT 11.475 123.950 15.175 124.950 ;
        RECT 15.750 124.275 16.750 124.320 ;
        RECT 16.930 124.275 17.930 127.475 ;
        RECT 11.475 122.435 12.475 123.950 ;
        RECT 15.750 123.275 17.930 124.275 ;
        RECT 18.350 123.275 18.720 127.475 ;
        RECT 19.625 125.975 20.630 128.475 ;
        RECT 21.050 128.475 21.420 134.500 ;
        RECT 27.145 134.200 29.170 134.825 ;
        RECT 27.145 134.170 28.370 134.200 ;
        RECT 24.820 133.155 25.925 133.200 ;
        RECT 24.775 132.050 25.970 133.155 ;
        RECT 24.790 132.045 25.955 132.050 ;
        RECT 23.425 128.475 24.375 128.500 ;
        RECT 21.050 127.475 26.300 128.475 ;
        RECT 19.605 125.025 20.645 125.975 ;
        RECT 19.625 125.000 20.630 125.025 ;
        RECT 20.260 123.275 20.630 125.000 ;
        RECT 21.050 123.275 21.420 127.475 ;
        RECT 23.425 127.460 24.375 127.475 ;
        RECT 15.750 123.230 16.750 123.275 ;
        RECT 27.370 122.435 28.370 134.170 ;
        RECT 31.475 130.975 32.475 137.075 ;
        RECT 38.075 135.825 39.075 137.200 ;
        RECT 41.600 137.125 62.875 138.225 ;
        RECT 64.425 138.200 65.425 139.175 ;
        RECT 71.225 139.155 72.175 139.175 ;
        RECT 72.645 138.225 73.645 140.000 ;
        RECT 74.370 138.325 75.370 139.220 ;
        RECT 63.500 137.200 65.425 138.200 ;
        RECT 42.315 137.120 44.825 137.125 ;
        RECT 45.015 137.120 62.140 137.125 ;
        RECT 56.845 137.075 57.950 137.120 ;
        RECT 38.055 134.875 39.095 135.825 ;
        RECT 38.075 134.850 39.075 134.875 ;
        RECT 39.830 134.850 40.920 135.850 ;
        RECT 31.475 129.975 32.500 130.975 ;
        RECT 32.975 129.975 33.920 130.500 ;
        RECT 31.995 128.850 33.035 129.325 ;
        RECT 29.375 128.500 30.375 128.505 ;
        RECT 29.345 128.475 30.405 128.500 ;
        RECT 31.995 128.475 32.500 128.850 ;
        RECT 33.345 128.520 33.920 129.975 ;
        RECT 29.300 128.450 32.500 128.475 ;
        RECT 29.300 127.500 32.520 128.450 ;
        RECT 29.300 127.475 32.500 127.500 ;
        RECT 29.375 127.445 30.375 127.475 ;
        RECT 31.995 127.100 32.500 127.475 ;
        RECT 32.925 127.430 33.925 128.520 ;
        RECT 34.885 128.475 35.255 134.500 ;
        RECT 34.250 127.475 35.255 128.475 ;
        RECT 31.995 126.605 33.035 127.100 ;
        RECT 33.345 126.200 33.920 127.430 ;
        RECT 31.500 125.825 32.555 126.200 ;
        RECT 32.975 125.825 33.920 126.200 ;
        RECT 29.330 122.455 30.445 122.460 ;
        RECT 29.300 122.435 30.475 122.455 ;
        RECT 31.500 122.435 32.500 125.825 ;
        RECT 34.255 124.275 35.255 127.475 ;
        RECT 33.055 123.275 35.255 124.275 ;
        RECT 35.675 128.520 36.045 134.500 ;
        RECT 39.875 134.075 40.875 134.105 ;
        RECT 39.875 133.075 42.645 134.075 ;
        RECT 39.875 133.045 40.875 133.075 ;
        RECT 36.900 129.975 37.900 132.425 ;
        RECT 38.375 129.975 39.320 130.500 ;
        RECT 39.600 129.975 40.600 132.425 ;
        RECT 41.075 129.975 42.020 130.500 ;
        RECT 37.395 128.850 38.435 129.325 ;
        RECT 35.675 128.475 36.675 128.520 ;
        RECT 37.395 128.475 37.900 128.850 ;
        RECT 38.745 128.475 39.320 129.975 ;
        RECT 40.095 128.850 41.135 129.325 ;
        RECT 40.095 128.475 40.600 128.850 ;
        RECT 41.445 128.475 42.020 129.975 ;
        RECT 42.985 128.475 43.355 134.500 ;
        RECT 43.775 128.475 44.145 134.500 ;
        RECT 45.685 128.475 46.055 134.500 ;
        RECT 35.675 128.450 37.900 128.475 ;
        RECT 35.675 127.505 37.920 128.450 ;
        RECT 35.675 127.475 37.900 127.505 ;
        RECT 38.280 127.475 40.600 128.475 ;
        RECT 41.025 127.475 43.355 128.475 ;
        RECT 43.730 127.475 44.820 128.475 ;
        RECT 35.675 127.430 36.675 127.475 ;
        RECT 35.675 123.275 36.045 127.430 ;
        RECT 37.395 127.100 37.900 127.475 ;
        RECT 37.395 126.605 38.435 127.100 ;
        RECT 38.745 126.200 39.320 127.475 ;
        RECT 40.095 127.100 40.600 127.475 ;
        RECT 40.095 126.605 41.135 127.100 ;
        RECT 41.445 126.200 42.020 127.475 ;
        RECT 36.900 125.825 37.955 126.200 ;
        RECT 38.375 125.825 39.320 126.200 ;
        RECT 39.600 125.825 40.655 126.200 ;
        RECT 41.075 125.825 42.020 126.200 ;
        RECT 36.900 124.950 37.900 125.825 ;
        RECT 39.600 124.950 40.600 125.825 ;
        RECT 36.900 123.950 40.600 124.950 ;
        RECT 41.175 124.275 42.175 124.320 ;
        RECT 42.355 124.275 43.355 127.475 ;
        RECT 36.900 122.435 37.900 123.950 ;
        RECT 41.175 123.275 43.355 124.275 ;
        RECT 43.775 123.275 44.145 127.475 ;
        RECT 45.050 125.975 46.055 128.475 ;
        RECT 46.475 128.475 46.845 134.500 ;
        RECT 56.900 130.975 57.900 137.075 ;
        RECT 63.500 135.825 64.500 137.200 ;
        RECT 67.025 137.150 73.645 138.225 ;
        RECT 74.340 137.325 75.400 138.325 ;
        RECT 67.025 137.125 72.950 137.150 ;
        RECT 67.740 137.120 70.250 137.125 ;
        RECT 70.440 137.120 72.940 137.125 ;
        RECT 75.720 136.575 76.720 139.525 ;
        RECT 77.995 138.975 80.020 140.000 ;
        RECT 80.495 138.975 81.440 139.500 ;
        RECT 77.995 138.945 78.995 138.975 ;
        RECT 77.095 138.295 78.095 138.340 ;
        RECT 77.065 137.295 78.125 138.295 ;
        RECT 79.515 137.850 80.555 138.325 ;
        RECT 79.515 137.475 80.020 137.850 ;
        RECT 80.865 137.475 81.440 138.975 ;
        RECT 82.320 138.270 83.320 140.000 ;
        RECT 85.825 139.175 89.030 140.175 ;
        RECT 89.805 139.175 90.895 140.175 ;
        RECT 91.645 139.175 94.925 140.175 ;
        RECT 96.625 139.175 97.625 140.175 ;
        RECT 111.250 139.175 114.455 140.175 ;
        RECT 115.230 139.175 116.320 140.175 ;
        RECT 117.070 139.175 120.350 140.175 ;
        RECT 122.050 139.175 123.050 140.175 ;
        RECT 123.495 140.000 134.170 141.000 ;
        RECT 136.700 140.175 137.650 140.195 ;
        RECT 147.500 140.175 148.450 140.195 ;
        RECT 85.850 139.155 86.800 139.175 ;
        RECT 82.270 138.225 83.375 138.270 ;
        RECT 77.095 137.250 78.095 137.295 ;
        RECT 79.020 136.575 80.020 137.475 ;
        RECT 67.025 136.340 68.025 136.385 ;
        RECT 71.220 136.340 72.170 136.360 ;
        RECT 63.480 134.875 64.520 135.825 ;
        RECT 63.500 134.850 64.500 134.875 ;
        RECT 65.255 134.850 66.345 135.850 ;
        RECT 67.025 135.340 72.195 136.340 ;
        RECT 75.720 136.100 80.020 136.575 ;
        RECT 80.400 136.475 81.490 137.475 ;
        RECT 82.240 137.125 88.300 138.225 ;
        RECT 89.850 138.200 90.850 139.175 ;
        RECT 96.650 139.155 97.600 139.175 ;
        RECT 111.275 139.155 112.225 139.175 ;
        RECT 107.695 138.225 108.800 138.270 ;
        RECT 88.925 137.200 90.850 138.200 ;
        RECT 82.240 137.120 87.565 137.125 ;
        RECT 82.270 137.075 83.375 137.120 ;
        RECT 75.720 135.650 80.555 136.100 ;
        RECT 73.870 135.605 80.555 135.650 ;
        RECT 73.870 135.575 80.020 135.605 ;
        RECT 67.025 135.295 68.025 135.340 ;
        RECT 71.220 135.320 72.170 135.340 ;
        RECT 73.870 134.650 76.720 135.575 ;
        RECT 77.995 135.200 78.995 135.230 ;
        RECT 80.865 135.200 81.440 136.475 ;
        RECT 77.995 134.825 80.075 135.200 ;
        RECT 80.495 134.825 81.440 135.200 ;
        RECT 56.900 129.975 57.925 130.975 ;
        RECT 58.400 129.975 59.345 130.500 ;
        RECT 57.420 128.850 58.460 129.325 ;
        RECT 50.725 128.475 51.725 128.505 ;
        RECT 54.800 128.500 55.800 128.505 ;
        RECT 54.770 128.475 55.830 128.500 ;
        RECT 57.420 128.475 57.925 128.850 ;
        RECT 58.770 128.520 59.345 129.975 ;
        RECT 46.475 127.475 51.725 128.475 ;
        RECT 54.725 128.450 57.925 128.475 ;
        RECT 54.725 127.500 57.945 128.450 ;
        RECT 54.725 127.475 57.925 127.500 ;
        RECT 45.030 125.025 46.070 125.975 ;
        RECT 45.050 125.000 46.055 125.025 ;
        RECT 45.685 123.275 46.055 125.000 ;
        RECT 46.475 123.275 46.845 127.475 ;
        RECT 50.725 127.445 51.725 127.475 ;
        RECT 54.800 127.445 55.800 127.475 ;
        RECT 57.420 127.100 57.925 127.475 ;
        RECT 58.350 127.430 59.350 128.520 ;
        RECT 60.310 128.475 60.680 134.500 ;
        RECT 59.675 127.475 60.680 128.475 ;
        RECT 57.420 126.605 58.460 127.100 ;
        RECT 58.770 126.200 59.345 127.430 ;
        RECT 56.925 125.825 57.980 126.200 ;
        RECT 58.400 125.825 59.345 126.200 ;
        RECT 41.175 123.230 42.175 123.275 ;
        RECT 54.755 122.455 55.870 122.460 ;
        RECT 54.725 122.435 55.900 122.455 ;
        RECT 56.925 122.435 57.925 125.825 ;
        RECT 59.680 124.275 60.680 127.475 ;
        RECT 58.480 123.275 60.680 124.275 ;
        RECT 61.100 128.520 61.470 134.500 ;
        RECT 65.300 134.075 66.300 134.105 ;
        RECT 65.300 133.075 68.070 134.075 ;
        RECT 65.300 133.045 66.300 133.075 ;
        RECT 62.325 129.975 63.325 132.425 ;
        RECT 63.800 129.975 64.745 130.500 ;
        RECT 65.025 129.975 66.025 132.425 ;
        RECT 66.500 129.975 67.445 130.500 ;
        RECT 62.820 128.850 63.860 129.325 ;
        RECT 61.100 128.475 62.100 128.520 ;
        RECT 62.820 128.475 63.325 128.850 ;
        RECT 64.170 128.475 64.745 129.975 ;
        RECT 65.520 128.850 66.560 129.325 ;
        RECT 65.520 128.475 66.025 128.850 ;
        RECT 66.870 128.475 67.445 129.975 ;
        RECT 68.410 128.475 68.780 134.500 ;
        RECT 69.200 128.475 69.570 134.500 ;
        RECT 71.110 128.475 71.480 134.500 ;
        RECT 61.100 128.450 63.325 128.475 ;
        RECT 61.100 127.505 63.345 128.450 ;
        RECT 61.100 127.475 63.325 127.505 ;
        RECT 63.705 127.475 66.025 128.475 ;
        RECT 66.450 127.475 68.780 128.475 ;
        RECT 69.155 127.475 70.245 128.475 ;
        RECT 61.100 127.430 62.100 127.475 ;
        RECT 61.100 123.275 61.470 127.430 ;
        RECT 62.820 127.100 63.325 127.475 ;
        RECT 62.820 126.605 63.860 127.100 ;
        RECT 64.170 126.200 64.745 127.475 ;
        RECT 65.520 127.100 66.025 127.475 ;
        RECT 65.520 126.605 66.560 127.100 ;
        RECT 66.870 126.200 67.445 127.475 ;
        RECT 62.325 125.825 63.380 126.200 ;
        RECT 63.800 125.825 64.745 126.200 ;
        RECT 65.025 125.825 66.080 126.200 ;
        RECT 66.500 125.825 67.445 126.200 ;
        RECT 62.325 124.950 63.325 125.825 ;
        RECT 65.025 124.950 66.025 125.825 ;
        RECT 62.325 123.950 66.025 124.950 ;
        RECT 66.600 124.275 67.600 124.320 ;
        RECT 67.780 124.275 68.780 127.475 ;
        RECT 62.325 122.435 63.325 123.950 ;
        RECT 66.600 123.275 68.780 124.275 ;
        RECT 69.200 123.275 69.570 127.475 ;
        RECT 70.475 125.975 71.480 128.475 ;
        RECT 71.900 128.475 72.270 134.500 ;
        RECT 77.995 134.200 80.020 134.825 ;
        RECT 77.995 134.170 79.220 134.200 ;
        RECT 75.670 133.155 76.775 133.200 ;
        RECT 75.625 132.050 76.820 133.155 ;
        RECT 75.640 132.045 76.805 132.050 ;
        RECT 74.275 128.475 75.225 128.500 ;
        RECT 71.900 127.475 77.150 128.475 ;
        RECT 70.455 125.025 71.495 125.975 ;
        RECT 70.475 125.000 71.480 125.025 ;
        RECT 71.110 123.275 71.480 125.000 ;
        RECT 71.900 123.275 72.270 127.475 ;
        RECT 74.275 127.460 75.225 127.475 ;
        RECT 66.600 123.230 67.600 123.275 ;
        RECT 78.220 122.435 79.220 134.170 ;
        RECT 82.325 130.975 83.325 137.075 ;
        RECT 88.925 135.825 89.925 137.200 ;
        RECT 92.450 137.125 113.725 138.225 ;
        RECT 115.275 138.200 116.275 139.175 ;
        RECT 122.075 139.155 123.025 139.175 ;
        RECT 123.495 138.225 124.495 140.000 ;
        RECT 125.220 138.325 126.220 139.220 ;
        RECT 114.350 137.200 116.275 138.200 ;
        RECT 93.165 137.120 95.675 137.125 ;
        RECT 95.865 137.120 112.990 137.125 ;
        RECT 107.695 137.075 108.800 137.120 ;
        RECT 88.905 134.875 89.945 135.825 ;
        RECT 88.925 134.850 89.925 134.875 ;
        RECT 90.680 134.850 91.770 135.850 ;
        RECT 82.325 129.975 83.350 130.975 ;
        RECT 83.825 129.975 84.770 130.500 ;
        RECT 82.845 128.850 83.885 129.325 ;
        RECT 80.225 128.500 81.225 128.505 ;
        RECT 80.195 128.475 81.255 128.500 ;
        RECT 82.845 128.475 83.350 128.850 ;
        RECT 84.195 128.520 84.770 129.975 ;
        RECT 80.150 128.450 83.350 128.475 ;
        RECT 80.150 127.500 83.370 128.450 ;
        RECT 80.150 127.475 83.350 127.500 ;
        RECT 80.225 127.445 81.225 127.475 ;
        RECT 82.845 127.100 83.350 127.475 ;
        RECT 83.775 127.430 84.775 128.520 ;
        RECT 85.735 128.475 86.105 134.500 ;
        RECT 85.100 127.475 86.105 128.475 ;
        RECT 82.845 126.605 83.885 127.100 ;
        RECT 84.195 126.200 84.770 127.430 ;
        RECT 82.350 125.825 83.405 126.200 ;
        RECT 83.825 125.825 84.770 126.200 ;
        RECT 80.180 122.455 81.295 122.460 ;
        RECT 80.150 122.435 81.325 122.455 ;
        RECT 82.350 122.435 83.350 125.825 ;
        RECT 85.105 124.275 86.105 127.475 ;
        RECT 83.905 123.275 86.105 124.275 ;
        RECT 86.525 128.520 86.895 134.500 ;
        RECT 90.725 134.075 91.725 134.105 ;
        RECT 90.725 133.075 93.495 134.075 ;
        RECT 90.725 133.045 91.725 133.075 ;
        RECT 87.750 129.975 88.750 132.425 ;
        RECT 89.225 129.975 90.170 130.500 ;
        RECT 90.450 129.975 91.450 132.425 ;
        RECT 91.925 129.975 92.870 130.500 ;
        RECT 88.245 128.850 89.285 129.325 ;
        RECT 86.525 128.475 87.525 128.520 ;
        RECT 88.245 128.475 88.750 128.850 ;
        RECT 89.595 128.475 90.170 129.975 ;
        RECT 90.945 128.850 91.985 129.325 ;
        RECT 90.945 128.475 91.450 128.850 ;
        RECT 92.295 128.475 92.870 129.975 ;
        RECT 93.835 128.475 94.205 134.500 ;
        RECT 94.625 128.475 94.995 134.500 ;
        RECT 96.535 128.475 96.905 134.500 ;
        RECT 86.525 128.450 88.750 128.475 ;
        RECT 86.525 127.505 88.770 128.450 ;
        RECT 86.525 127.475 88.750 127.505 ;
        RECT 89.130 127.475 91.450 128.475 ;
        RECT 91.875 127.475 94.205 128.475 ;
        RECT 94.580 127.475 95.670 128.475 ;
        RECT 86.525 127.430 87.525 127.475 ;
        RECT 86.525 123.275 86.895 127.430 ;
        RECT 88.245 127.100 88.750 127.475 ;
        RECT 88.245 126.605 89.285 127.100 ;
        RECT 89.595 126.200 90.170 127.475 ;
        RECT 90.945 127.100 91.450 127.475 ;
        RECT 90.945 126.605 91.985 127.100 ;
        RECT 92.295 126.200 92.870 127.475 ;
        RECT 87.750 125.825 88.805 126.200 ;
        RECT 89.225 125.825 90.170 126.200 ;
        RECT 90.450 125.825 91.505 126.200 ;
        RECT 91.925 125.825 92.870 126.200 ;
        RECT 87.750 124.950 88.750 125.825 ;
        RECT 90.450 124.950 91.450 125.825 ;
        RECT 87.750 123.950 91.450 124.950 ;
        RECT 92.025 124.275 93.025 124.320 ;
        RECT 93.205 124.275 94.205 127.475 ;
        RECT 87.750 122.435 88.750 123.950 ;
        RECT 92.025 123.275 94.205 124.275 ;
        RECT 94.625 123.275 94.995 127.475 ;
        RECT 95.900 125.975 96.905 128.475 ;
        RECT 97.325 128.475 97.695 134.500 ;
        RECT 107.750 130.975 108.750 137.075 ;
        RECT 114.350 135.825 115.350 137.200 ;
        RECT 117.875 137.150 124.495 138.225 ;
        RECT 125.190 137.325 126.250 138.325 ;
        RECT 117.875 137.125 123.800 137.150 ;
        RECT 118.590 137.120 121.100 137.125 ;
        RECT 121.290 137.120 123.790 137.125 ;
        RECT 126.570 136.575 127.570 139.525 ;
        RECT 128.845 138.975 130.870 140.000 ;
        RECT 131.345 138.975 132.290 139.500 ;
        RECT 128.845 138.945 129.845 138.975 ;
        RECT 127.945 138.295 128.945 138.340 ;
        RECT 127.915 137.295 128.975 138.295 ;
        RECT 130.365 137.850 131.405 138.325 ;
        RECT 130.365 137.475 130.870 137.850 ;
        RECT 131.715 137.475 132.290 138.975 ;
        RECT 133.170 138.270 134.170 140.000 ;
        RECT 136.675 139.175 139.880 140.175 ;
        RECT 140.655 139.175 141.745 140.175 ;
        RECT 142.495 139.175 145.775 140.175 ;
        RECT 147.475 139.175 148.475 140.175 ;
        RECT 136.700 139.155 137.650 139.175 ;
        RECT 133.120 138.225 134.225 138.270 ;
        RECT 127.945 137.250 128.945 137.295 ;
        RECT 129.870 136.575 130.870 137.475 ;
        RECT 117.875 136.340 118.875 136.385 ;
        RECT 122.070 136.340 123.020 136.360 ;
        RECT 114.330 134.875 115.370 135.825 ;
        RECT 114.350 134.850 115.350 134.875 ;
        RECT 116.105 134.850 117.195 135.850 ;
        RECT 117.875 135.340 123.045 136.340 ;
        RECT 126.570 136.100 130.870 136.575 ;
        RECT 131.250 136.475 132.340 137.475 ;
        RECT 133.090 137.125 139.150 138.225 ;
        RECT 140.700 138.200 141.700 139.175 ;
        RECT 147.500 139.155 148.450 139.175 ;
        RECT 139.775 137.200 141.700 138.200 ;
        RECT 133.090 137.120 138.415 137.125 ;
        RECT 133.120 137.075 134.225 137.120 ;
        RECT 126.570 135.650 131.405 136.100 ;
        RECT 124.720 135.605 131.405 135.650 ;
        RECT 124.720 135.575 130.870 135.605 ;
        RECT 117.875 135.295 118.875 135.340 ;
        RECT 122.070 135.320 123.020 135.340 ;
        RECT 124.720 134.650 127.570 135.575 ;
        RECT 128.845 135.200 129.845 135.230 ;
        RECT 131.715 135.200 132.290 136.475 ;
        RECT 128.845 134.825 130.925 135.200 ;
        RECT 131.345 134.825 132.290 135.200 ;
        RECT 107.750 129.975 108.775 130.975 ;
        RECT 109.250 129.975 110.195 130.500 ;
        RECT 108.270 128.850 109.310 129.325 ;
        RECT 101.575 128.475 102.575 128.505 ;
        RECT 105.650 128.500 106.650 128.505 ;
        RECT 105.620 128.475 106.680 128.500 ;
        RECT 108.270 128.475 108.775 128.850 ;
        RECT 109.620 128.520 110.195 129.975 ;
        RECT 97.325 127.475 102.575 128.475 ;
        RECT 105.575 128.450 108.775 128.475 ;
        RECT 105.575 127.500 108.795 128.450 ;
        RECT 105.575 127.475 108.775 127.500 ;
        RECT 95.880 125.025 96.920 125.975 ;
        RECT 95.900 125.000 96.905 125.025 ;
        RECT 96.535 123.275 96.905 125.000 ;
        RECT 97.325 123.275 97.695 127.475 ;
        RECT 101.575 127.445 102.575 127.475 ;
        RECT 105.650 127.445 106.650 127.475 ;
        RECT 108.270 127.100 108.775 127.475 ;
        RECT 109.200 127.430 110.200 128.520 ;
        RECT 111.160 128.475 111.530 134.500 ;
        RECT 110.525 127.475 111.530 128.475 ;
        RECT 108.270 126.605 109.310 127.100 ;
        RECT 109.620 126.200 110.195 127.430 ;
        RECT 107.775 125.825 108.830 126.200 ;
        RECT 109.250 125.825 110.195 126.200 ;
        RECT 92.025 123.230 93.025 123.275 ;
        RECT 105.605 122.455 106.720 122.460 ;
        RECT 105.575 122.435 106.750 122.455 ;
        RECT 107.775 122.435 108.775 125.825 ;
        RECT 110.530 124.275 111.530 127.475 ;
        RECT 109.330 123.275 111.530 124.275 ;
        RECT 111.950 128.520 112.320 134.500 ;
        RECT 116.150 134.075 117.150 134.105 ;
        RECT 116.150 133.075 118.920 134.075 ;
        RECT 116.150 133.045 117.150 133.075 ;
        RECT 113.175 129.975 114.175 132.425 ;
        RECT 114.650 129.975 115.595 130.500 ;
        RECT 115.875 129.975 116.875 132.425 ;
        RECT 117.350 129.975 118.295 130.500 ;
        RECT 113.670 128.850 114.710 129.325 ;
        RECT 111.950 128.475 112.950 128.520 ;
        RECT 113.670 128.475 114.175 128.850 ;
        RECT 115.020 128.475 115.595 129.975 ;
        RECT 116.370 128.850 117.410 129.325 ;
        RECT 116.370 128.475 116.875 128.850 ;
        RECT 117.720 128.475 118.295 129.975 ;
        RECT 119.260 128.475 119.630 134.500 ;
        RECT 120.050 128.475 120.420 134.500 ;
        RECT 121.960 128.475 122.330 134.500 ;
        RECT 111.950 128.450 114.175 128.475 ;
        RECT 111.950 127.505 114.195 128.450 ;
        RECT 111.950 127.475 114.175 127.505 ;
        RECT 114.555 127.475 116.875 128.475 ;
        RECT 117.300 127.475 119.630 128.475 ;
        RECT 120.005 127.475 121.095 128.475 ;
        RECT 111.950 127.430 112.950 127.475 ;
        RECT 111.950 123.275 112.320 127.430 ;
        RECT 113.670 127.100 114.175 127.475 ;
        RECT 113.670 126.605 114.710 127.100 ;
        RECT 115.020 126.200 115.595 127.475 ;
        RECT 116.370 127.100 116.875 127.475 ;
        RECT 116.370 126.605 117.410 127.100 ;
        RECT 117.720 126.200 118.295 127.475 ;
        RECT 113.175 125.825 114.230 126.200 ;
        RECT 114.650 125.825 115.595 126.200 ;
        RECT 115.875 125.825 116.930 126.200 ;
        RECT 117.350 125.825 118.295 126.200 ;
        RECT 113.175 124.950 114.175 125.825 ;
        RECT 115.875 124.950 116.875 125.825 ;
        RECT 113.175 123.950 116.875 124.950 ;
        RECT 117.450 124.275 118.450 124.320 ;
        RECT 118.630 124.275 119.630 127.475 ;
        RECT 113.175 122.435 114.175 123.950 ;
        RECT 117.450 123.275 119.630 124.275 ;
        RECT 120.050 123.275 120.420 127.475 ;
        RECT 121.325 125.975 122.330 128.475 ;
        RECT 122.750 128.475 123.120 134.500 ;
        RECT 128.845 134.200 130.870 134.825 ;
        RECT 128.845 134.170 130.070 134.200 ;
        RECT 126.520 133.155 127.625 133.200 ;
        RECT 126.475 132.050 127.670 133.155 ;
        RECT 126.490 132.045 127.655 132.050 ;
        RECT 125.125 128.475 126.075 128.500 ;
        RECT 122.750 127.475 128.000 128.475 ;
        RECT 121.305 125.025 122.345 125.975 ;
        RECT 121.325 125.000 122.330 125.025 ;
        RECT 121.960 123.275 122.330 125.000 ;
        RECT 122.750 123.275 123.120 127.475 ;
        RECT 125.125 127.460 126.075 127.475 ;
        RECT 117.450 123.230 118.450 123.275 ;
        RECT 129.070 122.435 130.070 134.170 ;
        RECT 133.175 130.975 134.175 137.075 ;
        RECT 139.775 135.825 140.775 137.200 ;
        RECT 143.300 137.125 149.225 138.225 ;
        RECT 144.015 137.120 146.525 137.125 ;
        RECT 146.715 137.120 149.215 137.125 ;
        RECT 139.755 134.875 140.795 135.825 ;
        RECT 139.775 134.850 140.775 134.875 ;
        RECT 141.530 134.850 142.620 135.850 ;
        RECT 133.175 129.975 134.200 130.975 ;
        RECT 134.675 129.975 135.620 130.500 ;
        RECT 133.695 128.850 134.735 129.325 ;
        RECT 131.075 128.500 132.075 128.505 ;
        RECT 131.045 128.475 132.105 128.500 ;
        RECT 133.695 128.475 134.200 128.850 ;
        RECT 135.045 128.520 135.620 129.975 ;
        RECT 131.000 128.450 134.200 128.475 ;
        RECT 131.000 127.500 134.220 128.450 ;
        RECT 131.000 127.475 134.200 127.500 ;
        RECT 131.075 127.445 132.075 127.475 ;
        RECT 133.695 127.100 134.200 127.475 ;
        RECT 134.625 127.430 135.625 128.520 ;
        RECT 136.585 128.475 136.955 134.500 ;
        RECT 135.950 127.475 136.955 128.475 ;
        RECT 133.695 126.605 134.735 127.100 ;
        RECT 135.045 126.200 135.620 127.430 ;
        RECT 133.200 125.825 134.255 126.200 ;
        RECT 134.675 125.825 135.620 126.200 ;
        RECT 131.030 122.455 132.145 122.460 ;
        RECT 131.000 122.435 132.175 122.455 ;
        RECT 133.200 122.435 134.200 125.825 ;
        RECT 135.955 124.275 136.955 127.475 ;
        RECT 134.755 123.275 136.955 124.275 ;
        RECT 137.375 128.520 137.745 134.500 ;
        RECT 141.575 134.075 142.575 134.105 ;
        RECT 141.575 133.075 144.345 134.075 ;
        RECT 141.575 133.045 142.575 133.075 ;
        RECT 138.600 129.975 139.600 132.425 ;
        RECT 140.075 129.975 141.020 130.500 ;
        RECT 141.300 129.975 142.300 132.425 ;
        RECT 142.775 129.975 143.720 130.500 ;
        RECT 139.095 128.850 140.135 129.325 ;
        RECT 137.375 128.475 138.375 128.520 ;
        RECT 139.095 128.475 139.600 128.850 ;
        RECT 140.445 128.475 141.020 129.975 ;
        RECT 141.795 128.850 142.835 129.325 ;
        RECT 141.795 128.475 142.300 128.850 ;
        RECT 143.145 128.475 143.720 129.975 ;
        RECT 144.685 128.475 145.055 134.500 ;
        RECT 145.475 128.475 145.845 134.500 ;
        RECT 147.385 128.475 147.755 134.500 ;
        RECT 137.375 128.450 139.600 128.475 ;
        RECT 137.375 127.505 139.620 128.450 ;
        RECT 137.375 127.475 139.600 127.505 ;
        RECT 139.980 127.475 142.300 128.475 ;
        RECT 142.725 127.475 145.055 128.475 ;
        RECT 145.430 127.475 146.520 128.475 ;
        RECT 137.375 127.430 138.375 127.475 ;
        RECT 137.375 123.275 137.745 127.430 ;
        RECT 139.095 127.100 139.600 127.475 ;
        RECT 139.095 126.605 140.135 127.100 ;
        RECT 140.445 126.200 141.020 127.475 ;
        RECT 141.795 127.100 142.300 127.475 ;
        RECT 141.795 126.605 142.835 127.100 ;
        RECT 143.145 126.200 143.720 127.475 ;
        RECT 138.600 125.825 139.655 126.200 ;
        RECT 140.075 125.825 141.020 126.200 ;
        RECT 141.300 125.825 142.355 126.200 ;
        RECT 142.775 125.825 143.720 126.200 ;
        RECT 138.600 124.950 139.600 125.825 ;
        RECT 141.300 124.950 142.300 125.825 ;
        RECT 138.600 123.950 142.300 124.950 ;
        RECT 142.875 124.275 143.875 124.320 ;
        RECT 144.055 124.275 145.055 127.475 ;
        RECT 138.600 122.435 139.600 123.950 ;
        RECT 142.875 123.275 145.055 124.275 ;
        RECT 145.475 123.275 145.845 127.475 ;
        RECT 146.750 125.975 147.755 128.475 ;
        RECT 148.175 128.475 148.545 134.500 ;
        RECT 152.425 128.475 153.425 128.505 ;
        RECT 148.175 127.475 153.425 128.475 ;
        RECT 146.730 125.025 147.770 125.975 ;
        RECT 146.750 125.000 147.755 125.025 ;
        RECT 147.385 123.275 147.755 125.000 ;
        RECT 148.175 123.275 148.545 127.475 ;
        RECT 152.425 127.445 153.425 127.475 ;
        RECT 142.875 123.230 143.875 123.275 ;
        RECT 1.850 122.425 14.575 122.435 ;
        RECT 15.350 122.425 19.390 122.435 ;
        RECT 19.590 122.425 40.000 122.435 ;
        RECT 40.775 122.425 44.815 122.435 ;
        RECT 45.015 122.425 65.425 122.435 ;
        RECT 66.200 122.425 70.240 122.435 ;
        RECT 70.440 122.425 90.850 122.435 ;
        RECT 91.625 122.425 95.665 122.435 ;
        RECT 95.865 122.425 116.275 122.435 ;
        RECT 117.050 122.425 121.090 122.435 ;
        RECT 121.290 122.425 141.700 122.435 ;
        RECT 142.475 122.425 146.515 122.435 ;
        RECT 146.715 122.425 149.215 122.435 ;
        RECT 1.850 121.325 149.215 122.425 ;
        RECT 1.850 121.320 19.390 121.325 ;
        RECT 19.590 121.320 44.815 121.325 ;
        RECT 45.015 121.320 70.240 121.325 ;
        RECT 70.440 121.320 95.665 121.325 ;
        RECT 95.865 121.320 121.090 121.325 ;
        RECT 121.290 121.320 146.515 121.325 ;
        RECT 146.715 121.320 149.215 121.325 ;
        RECT 3.905 121.315 6.480 121.320 ;
        RECT 29.330 121.315 31.905 121.320 ;
        RECT 54.755 121.315 57.330 121.320 ;
        RECT 80.180 121.315 82.755 121.320 ;
        RECT 105.605 121.315 108.180 121.320 ;
        RECT 131.030 121.315 133.605 121.320 ;
        RECT 3.905 121.285 5.020 121.315 ;
        RECT 29.330 121.285 30.445 121.315 ;
        RECT 54.755 121.285 55.870 121.315 ;
        RECT 80.180 121.285 81.295 121.315 ;
        RECT 105.605 121.285 106.720 121.315 ;
        RECT 131.030 121.285 132.145 121.315 ;
        RECT 19.370 120.375 21.325 120.395 ;
        RECT 44.795 120.375 46.750 120.395 ;
        RECT 70.220 120.375 72.175 120.395 ;
        RECT 95.645 120.375 97.600 120.395 ;
        RECT 121.070 120.375 123.025 120.395 ;
        RECT 146.495 120.375 148.450 120.395 ;
        RECT 9.550 120.350 10.550 120.375 ;
        RECT 15.750 120.350 16.750 120.375 ;
        RECT 17.650 120.350 18.650 120.375 ;
        RECT 9.530 119.400 10.570 120.350 ;
        RECT 15.730 119.400 16.770 120.350 ;
        RECT 17.630 119.400 18.670 120.350 ;
        RECT 9.550 119.375 10.550 119.400 ;
        RECT 15.750 119.375 16.750 119.400 ;
        RECT 17.650 119.375 18.650 119.400 ;
        RECT 19.365 119.375 21.350 120.375 ;
        RECT 34.975 120.350 35.975 120.375 ;
        RECT 41.175 120.350 42.175 120.375 ;
        RECT 43.075 120.350 44.075 120.375 ;
        RECT 34.955 119.400 35.995 120.350 ;
        RECT 41.155 119.400 42.195 120.350 ;
        RECT 43.055 119.400 44.095 120.350 ;
        RECT 34.975 119.375 35.975 119.400 ;
        RECT 41.175 119.375 42.175 119.400 ;
        RECT 43.075 119.375 44.075 119.400 ;
        RECT 44.790 119.375 46.775 120.375 ;
        RECT 60.400 120.350 61.400 120.375 ;
        RECT 66.600 120.350 67.600 120.375 ;
        RECT 68.500 120.350 69.500 120.375 ;
        RECT 60.380 119.400 61.420 120.350 ;
        RECT 66.580 119.400 67.620 120.350 ;
        RECT 68.480 119.400 69.520 120.350 ;
        RECT 60.400 119.375 61.400 119.400 ;
        RECT 66.600 119.375 67.600 119.400 ;
        RECT 68.500 119.375 69.500 119.400 ;
        RECT 70.215 119.375 72.200 120.375 ;
        RECT 85.825 120.350 86.825 120.375 ;
        RECT 92.025 120.350 93.025 120.375 ;
        RECT 93.925 120.350 94.925 120.375 ;
        RECT 85.805 119.400 86.845 120.350 ;
        RECT 92.005 119.400 93.045 120.350 ;
        RECT 93.905 119.400 94.945 120.350 ;
        RECT 85.825 119.375 86.825 119.400 ;
        RECT 92.025 119.375 93.025 119.400 ;
        RECT 93.925 119.375 94.925 119.400 ;
        RECT 95.640 119.375 97.625 120.375 ;
        RECT 111.250 120.350 112.250 120.375 ;
        RECT 117.450 120.350 118.450 120.375 ;
        RECT 119.350 120.350 120.350 120.375 ;
        RECT 111.230 119.400 112.270 120.350 ;
        RECT 117.430 119.400 118.470 120.350 ;
        RECT 119.330 119.400 120.370 120.350 ;
        RECT 111.250 119.375 112.250 119.400 ;
        RECT 117.450 119.375 118.450 119.400 ;
        RECT 119.350 119.375 120.350 119.400 ;
        RECT 121.065 119.375 123.050 120.375 ;
        RECT 136.675 120.350 137.675 120.375 ;
        RECT 142.875 120.350 143.875 120.375 ;
        RECT 144.775 120.350 145.775 120.375 ;
        RECT 136.655 119.400 137.695 120.350 ;
        RECT 142.855 119.400 143.895 120.350 ;
        RECT 144.755 119.400 145.795 120.350 ;
        RECT 136.675 119.375 137.675 119.400 ;
        RECT 142.875 119.375 143.875 119.400 ;
        RECT 144.775 119.375 145.775 119.400 ;
        RECT 146.490 119.375 148.475 120.375 ;
        RECT 19.370 119.355 21.325 119.375 ;
        RECT 44.795 119.355 46.750 119.375 ;
        RECT 70.220 119.355 72.175 119.375 ;
        RECT 95.645 119.355 97.600 119.375 ;
        RECT 121.070 119.355 123.025 119.375 ;
        RECT 146.495 119.355 148.450 119.375 ;
        RECT 9.575 117.600 10.525 117.620 ;
        RECT 20.375 117.600 21.325 117.620 ;
        RECT 35.000 117.600 35.950 117.620 ;
        RECT 45.800 117.600 46.750 117.620 ;
        RECT 60.425 117.600 61.375 117.620 ;
        RECT 71.225 117.600 72.175 117.620 ;
        RECT 85.850 117.600 86.800 117.620 ;
        RECT 96.650 117.600 97.600 117.620 ;
        RECT 111.275 117.600 112.225 117.620 ;
        RECT 122.075 117.600 123.025 117.620 ;
        RECT 136.700 117.600 137.650 117.620 ;
        RECT 147.500 117.600 148.450 117.620 ;
        RECT 9.550 116.600 12.755 117.600 ;
        RECT 13.530 116.600 14.620 117.600 ;
        RECT 15.370 116.600 18.650 117.600 ;
        RECT 20.350 116.600 21.350 117.600 ;
        RECT 34.975 116.600 38.180 117.600 ;
        RECT 38.955 116.600 40.045 117.600 ;
        RECT 40.795 116.600 44.075 117.600 ;
        RECT 45.775 116.600 46.775 117.600 ;
        RECT 60.400 116.600 63.605 117.600 ;
        RECT 64.380 116.600 65.470 117.600 ;
        RECT 66.220 116.600 69.500 117.600 ;
        RECT 71.200 116.600 72.200 117.600 ;
        RECT 85.825 116.600 89.030 117.600 ;
        RECT 89.805 116.600 90.895 117.600 ;
        RECT 91.645 116.600 94.925 117.600 ;
        RECT 96.625 116.600 97.625 117.600 ;
        RECT 111.250 116.600 114.455 117.600 ;
        RECT 115.230 116.600 116.320 117.600 ;
        RECT 117.070 116.600 120.350 117.600 ;
        RECT 122.050 116.600 123.050 117.600 ;
        RECT 136.675 116.600 139.880 117.600 ;
        RECT 140.655 116.600 141.745 117.600 ;
        RECT 142.495 116.600 145.775 117.600 ;
        RECT 147.475 116.600 148.475 117.600 ;
        RECT 9.575 116.580 10.525 116.600 ;
        RECT 3.925 115.655 4.980 115.675 ;
        RECT 3.575 115.650 6.000 115.655 ;
        RECT 1.850 114.550 12.025 115.650 ;
        RECT 13.575 115.625 14.575 116.600 ;
        RECT 20.375 116.580 21.325 116.600 ;
        RECT 35.000 116.580 35.950 116.600 ;
        RECT 29.350 115.655 30.405 115.675 ;
        RECT 29.000 115.650 31.425 115.655 ;
        RECT 12.650 114.625 14.575 115.625 ;
        RECT 1.850 114.545 11.290 114.550 ;
        RECT 3.925 114.530 4.980 114.545 ;
        RECT 6.050 108.400 7.050 114.545 ;
        RECT 12.650 113.250 13.650 114.625 ;
        RECT 16.175 114.550 37.450 115.650 ;
        RECT 39.000 115.625 40.000 116.600 ;
        RECT 45.800 116.580 46.750 116.600 ;
        RECT 60.425 116.580 61.375 116.600 ;
        RECT 54.775 115.655 55.830 115.675 ;
        RECT 54.425 115.650 56.850 115.655 ;
        RECT 38.075 114.625 40.000 115.625 ;
        RECT 16.890 114.545 19.400 114.550 ;
        RECT 19.590 114.545 36.715 114.550 ;
        RECT 29.350 114.530 30.405 114.545 ;
        RECT 12.630 112.300 13.670 113.250 ;
        RECT 12.650 112.275 13.650 112.300 ;
        RECT 14.405 112.275 15.495 113.275 ;
        RECT 6.050 107.400 7.075 108.400 ;
        RECT 7.550 107.400 8.495 107.925 ;
        RECT 6.570 106.275 7.610 106.750 ;
        RECT 1.900 105.925 2.900 105.930 ;
        RECT 1.870 105.900 2.930 105.925 ;
        RECT 6.570 105.900 7.075 106.275 ;
        RECT 7.920 105.945 8.495 107.400 ;
        RECT 1.850 105.875 7.075 105.900 ;
        RECT 1.850 104.925 7.095 105.875 ;
        RECT 1.850 104.900 7.075 104.925 ;
        RECT 1.900 104.870 2.900 104.900 ;
        RECT 6.570 104.525 7.075 104.900 ;
        RECT 7.500 104.855 8.500 105.945 ;
        RECT 9.460 105.900 9.830 111.925 ;
        RECT 8.825 104.900 9.830 105.900 ;
        RECT 6.570 104.030 7.610 104.525 ;
        RECT 7.920 103.625 8.495 104.855 ;
        RECT 6.075 103.250 7.130 103.625 ;
        RECT 7.550 103.250 8.495 103.625 ;
        RECT 3.905 99.860 5.020 99.885 ;
        RECT 6.075 99.860 7.075 103.250 ;
        RECT 8.830 101.700 9.830 104.900 ;
        RECT 7.630 100.700 9.830 101.700 ;
        RECT 10.250 105.945 10.620 111.925 ;
        RECT 14.450 111.500 15.450 111.530 ;
        RECT 14.450 110.500 17.220 111.500 ;
        RECT 14.450 110.470 15.450 110.500 ;
        RECT 11.475 107.400 12.475 109.850 ;
        RECT 12.950 107.400 13.895 107.925 ;
        RECT 14.175 107.400 15.175 109.850 ;
        RECT 15.650 107.400 16.595 107.925 ;
        RECT 11.970 106.275 13.010 106.750 ;
        RECT 10.250 105.900 11.250 105.945 ;
        RECT 11.970 105.900 12.475 106.275 ;
        RECT 13.320 105.900 13.895 107.400 ;
        RECT 14.670 106.275 15.710 106.750 ;
        RECT 14.670 105.900 15.175 106.275 ;
        RECT 16.020 105.900 16.595 107.400 ;
        RECT 17.560 105.900 17.930 111.925 ;
        RECT 18.350 105.900 18.720 111.925 ;
        RECT 20.260 105.900 20.630 111.925 ;
        RECT 10.250 105.875 12.475 105.900 ;
        RECT 10.250 104.930 12.495 105.875 ;
        RECT 10.250 104.900 12.475 104.930 ;
        RECT 12.855 104.900 15.175 105.900 ;
        RECT 15.600 104.900 17.930 105.900 ;
        RECT 18.305 104.900 19.395 105.900 ;
        RECT 10.250 104.855 11.250 104.900 ;
        RECT 10.250 100.700 10.620 104.855 ;
        RECT 11.970 104.525 12.475 104.900 ;
        RECT 11.970 104.030 13.010 104.525 ;
        RECT 13.320 103.625 13.895 104.900 ;
        RECT 14.670 104.525 15.175 104.900 ;
        RECT 14.670 104.030 15.710 104.525 ;
        RECT 16.020 103.625 16.595 104.900 ;
        RECT 11.475 103.250 12.530 103.625 ;
        RECT 12.950 103.250 13.895 103.625 ;
        RECT 14.175 103.250 15.230 103.625 ;
        RECT 15.650 103.250 16.595 103.625 ;
        RECT 11.475 102.375 12.475 103.250 ;
        RECT 14.175 102.375 15.175 103.250 ;
        RECT 11.475 101.375 15.175 102.375 ;
        RECT 15.750 101.700 16.750 101.745 ;
        RECT 16.930 101.700 17.930 104.900 ;
        RECT 11.475 99.860 12.475 101.375 ;
        RECT 15.750 100.700 17.930 101.700 ;
        RECT 18.350 100.700 18.720 104.900 ;
        RECT 19.625 103.900 20.630 105.900 ;
        RECT 21.050 105.925 21.420 111.925 ;
        RECT 31.475 108.400 32.475 114.545 ;
        RECT 38.075 113.250 39.075 114.625 ;
        RECT 41.600 114.550 62.875 115.650 ;
        RECT 64.425 115.625 65.425 116.600 ;
        RECT 71.225 116.580 72.175 116.600 ;
        RECT 85.850 116.580 86.800 116.600 ;
        RECT 80.200 115.655 81.255 115.675 ;
        RECT 79.850 115.650 82.275 115.655 ;
        RECT 63.500 114.625 65.425 115.625 ;
        RECT 42.315 114.545 44.825 114.550 ;
        RECT 45.015 114.545 62.140 114.550 ;
        RECT 54.775 114.530 55.830 114.545 ;
        RECT 38.055 112.300 39.095 113.250 ;
        RECT 38.075 112.275 39.075 112.300 ;
        RECT 39.830 112.275 40.920 113.275 ;
        RECT 31.475 107.400 32.500 108.400 ;
        RECT 32.975 107.400 33.920 107.925 ;
        RECT 31.995 106.275 33.035 106.750 ;
        RECT 27.325 105.925 28.325 105.930 ;
        RECT 21.050 105.900 22.375 105.925 ;
        RECT 27.295 105.900 28.355 105.925 ;
        RECT 31.995 105.900 32.500 106.275 ;
        RECT 33.345 105.945 33.920 107.400 ;
        RECT 21.050 104.900 26.250 105.900 ;
        RECT 27.275 105.875 32.500 105.900 ;
        RECT 27.275 104.925 32.520 105.875 ;
        RECT 27.275 104.900 32.500 104.925 ;
        RECT 21.050 104.885 22.375 104.900 ;
        RECT 19.605 102.950 20.645 103.900 ;
        RECT 19.625 102.925 20.630 102.950 ;
        RECT 20.260 100.700 20.630 102.925 ;
        RECT 21.050 100.700 21.420 104.885 ;
        RECT 23.155 101.775 24.155 104.900 ;
        RECT 27.325 104.870 28.325 104.900 ;
        RECT 31.995 104.525 32.500 104.900 ;
        RECT 32.925 104.855 33.925 105.945 ;
        RECT 34.885 105.900 35.255 111.925 ;
        RECT 34.250 104.900 35.255 105.900 ;
        RECT 31.995 104.030 33.035 104.525 ;
        RECT 33.345 103.625 33.920 104.855 ;
        RECT 31.500 103.250 32.555 103.625 ;
        RECT 32.975 103.250 33.920 103.625 ;
        RECT 23.135 100.825 24.175 101.775 ;
        RECT 23.155 100.800 24.155 100.825 ;
        RECT 15.750 100.655 16.750 100.700 ;
        RECT 23.115 99.860 24.230 99.890 ;
        RECT 29.330 99.860 30.445 99.885 ;
        RECT 31.500 99.860 32.500 103.250 ;
        RECT 34.255 101.700 35.255 104.900 ;
        RECT 33.055 100.700 35.255 101.700 ;
        RECT 35.675 105.945 36.045 111.925 ;
        RECT 39.875 111.500 40.875 111.530 ;
        RECT 39.875 110.500 42.645 111.500 ;
        RECT 39.875 110.470 40.875 110.500 ;
        RECT 36.900 107.400 37.900 109.850 ;
        RECT 38.375 107.400 39.320 107.925 ;
        RECT 39.600 107.400 40.600 109.850 ;
        RECT 41.075 107.400 42.020 107.925 ;
        RECT 37.395 106.275 38.435 106.750 ;
        RECT 35.675 105.900 36.675 105.945 ;
        RECT 37.395 105.900 37.900 106.275 ;
        RECT 38.745 105.900 39.320 107.400 ;
        RECT 40.095 106.275 41.135 106.750 ;
        RECT 40.095 105.900 40.600 106.275 ;
        RECT 41.445 105.900 42.020 107.400 ;
        RECT 42.985 105.900 43.355 111.925 ;
        RECT 43.775 105.900 44.145 111.925 ;
        RECT 45.685 105.900 46.055 111.925 ;
        RECT 35.675 105.875 37.900 105.900 ;
        RECT 35.675 104.930 37.920 105.875 ;
        RECT 35.675 104.900 37.900 104.930 ;
        RECT 38.280 104.900 40.600 105.900 ;
        RECT 41.025 104.900 43.355 105.900 ;
        RECT 43.730 104.900 44.820 105.900 ;
        RECT 35.675 104.855 36.675 104.900 ;
        RECT 35.675 100.700 36.045 104.855 ;
        RECT 37.395 104.525 37.900 104.900 ;
        RECT 37.395 104.030 38.435 104.525 ;
        RECT 38.745 103.625 39.320 104.900 ;
        RECT 40.095 104.525 40.600 104.900 ;
        RECT 40.095 104.030 41.135 104.525 ;
        RECT 41.445 103.625 42.020 104.900 ;
        RECT 36.900 103.250 37.955 103.625 ;
        RECT 38.375 103.250 39.320 103.625 ;
        RECT 39.600 103.250 40.655 103.625 ;
        RECT 41.075 103.250 42.020 103.625 ;
        RECT 36.900 102.375 37.900 103.250 ;
        RECT 39.600 102.375 40.600 103.250 ;
        RECT 36.900 101.375 40.600 102.375 ;
        RECT 41.175 101.700 42.175 101.745 ;
        RECT 42.355 101.700 43.355 104.900 ;
        RECT 36.900 99.860 37.900 101.375 ;
        RECT 41.175 100.700 43.355 101.700 ;
        RECT 43.775 100.700 44.145 104.900 ;
        RECT 45.050 103.900 46.055 105.900 ;
        RECT 46.475 105.900 46.845 111.925 ;
        RECT 56.900 108.400 57.900 114.545 ;
        RECT 63.500 113.250 64.500 114.625 ;
        RECT 67.025 114.550 88.300 115.650 ;
        RECT 89.850 115.625 90.850 116.600 ;
        RECT 96.650 116.580 97.600 116.600 ;
        RECT 111.275 116.580 112.225 116.600 ;
        RECT 105.625 115.655 106.680 115.675 ;
        RECT 105.275 115.650 107.700 115.655 ;
        RECT 88.925 114.625 90.850 115.625 ;
        RECT 67.740 114.545 70.250 114.550 ;
        RECT 70.440 114.545 87.565 114.550 ;
        RECT 80.200 114.530 81.255 114.545 ;
        RECT 63.480 112.300 64.520 113.250 ;
        RECT 63.500 112.275 64.500 112.300 ;
        RECT 65.255 112.275 66.345 113.275 ;
        RECT 56.900 107.400 57.925 108.400 ;
        RECT 58.400 107.400 59.345 107.925 ;
        RECT 57.420 106.275 58.460 106.750 ;
        RECT 52.750 105.925 53.750 105.930 ;
        RECT 52.720 105.900 53.780 105.925 ;
        RECT 57.420 105.900 57.925 106.275 ;
        RECT 58.770 105.945 59.345 107.400 ;
        RECT 46.475 104.900 51.720 105.900 ;
        RECT 52.700 105.875 57.925 105.900 ;
        RECT 52.700 104.925 57.945 105.875 ;
        RECT 52.700 104.900 57.925 104.925 ;
        RECT 45.030 102.950 46.070 103.900 ;
        RECT 45.050 102.925 46.055 102.950 ;
        RECT 45.685 100.700 46.055 102.925 ;
        RECT 46.475 100.700 46.845 104.900 ;
        RECT 48.580 101.775 49.580 104.900 ;
        RECT 52.750 104.870 53.750 104.900 ;
        RECT 57.420 104.525 57.925 104.900 ;
        RECT 58.350 104.855 59.350 105.945 ;
        RECT 60.310 105.900 60.680 111.925 ;
        RECT 59.675 104.900 60.680 105.900 ;
        RECT 57.420 104.030 58.460 104.525 ;
        RECT 58.770 103.625 59.345 104.855 ;
        RECT 56.925 103.250 57.980 103.625 ;
        RECT 58.400 103.250 59.345 103.625 ;
        RECT 48.560 100.825 49.600 101.775 ;
        RECT 48.580 100.800 49.580 100.825 ;
        RECT 41.175 100.655 42.175 100.700 ;
        RECT 48.540 99.860 49.655 99.890 ;
        RECT 54.755 99.860 55.870 99.885 ;
        RECT 56.925 99.860 57.925 103.250 ;
        RECT 59.680 101.700 60.680 104.900 ;
        RECT 58.480 100.700 60.680 101.700 ;
        RECT 61.100 105.945 61.470 111.925 ;
        RECT 65.300 111.500 66.300 111.530 ;
        RECT 65.300 110.500 68.070 111.500 ;
        RECT 65.300 110.470 66.300 110.500 ;
        RECT 62.325 107.400 63.325 109.850 ;
        RECT 63.800 107.400 64.745 107.925 ;
        RECT 65.025 107.400 66.025 109.850 ;
        RECT 66.500 107.400 67.445 107.925 ;
        RECT 62.820 106.275 63.860 106.750 ;
        RECT 61.100 105.900 62.100 105.945 ;
        RECT 62.820 105.900 63.325 106.275 ;
        RECT 64.170 105.900 64.745 107.400 ;
        RECT 65.520 106.275 66.560 106.750 ;
        RECT 65.520 105.900 66.025 106.275 ;
        RECT 66.870 105.900 67.445 107.400 ;
        RECT 68.410 105.900 68.780 111.925 ;
        RECT 69.200 105.900 69.570 111.925 ;
        RECT 71.110 105.900 71.480 111.925 ;
        RECT 61.100 105.875 63.325 105.900 ;
        RECT 61.100 104.930 63.345 105.875 ;
        RECT 61.100 104.900 63.325 104.930 ;
        RECT 63.705 104.900 66.025 105.900 ;
        RECT 66.450 104.900 68.780 105.900 ;
        RECT 69.155 104.900 70.245 105.900 ;
        RECT 61.100 104.855 62.100 104.900 ;
        RECT 61.100 100.700 61.470 104.855 ;
        RECT 62.820 104.525 63.325 104.900 ;
        RECT 62.820 104.030 63.860 104.525 ;
        RECT 64.170 103.625 64.745 104.900 ;
        RECT 65.520 104.525 66.025 104.900 ;
        RECT 65.520 104.030 66.560 104.525 ;
        RECT 66.870 103.625 67.445 104.900 ;
        RECT 62.325 103.250 63.380 103.625 ;
        RECT 63.800 103.250 64.745 103.625 ;
        RECT 65.025 103.250 66.080 103.625 ;
        RECT 66.500 103.250 67.445 103.625 ;
        RECT 62.325 102.375 63.325 103.250 ;
        RECT 65.025 102.375 66.025 103.250 ;
        RECT 62.325 101.375 66.025 102.375 ;
        RECT 66.600 101.700 67.600 101.745 ;
        RECT 67.780 101.700 68.780 104.900 ;
        RECT 62.325 99.860 63.325 101.375 ;
        RECT 66.600 100.700 68.780 101.700 ;
        RECT 69.200 100.700 69.570 104.900 ;
        RECT 70.475 103.900 71.480 105.900 ;
        RECT 71.900 105.925 72.270 111.925 ;
        RECT 82.325 108.400 83.325 114.545 ;
        RECT 88.925 113.250 89.925 114.625 ;
        RECT 92.450 114.550 113.725 115.650 ;
        RECT 115.275 115.625 116.275 116.600 ;
        RECT 122.075 116.580 123.025 116.600 ;
        RECT 136.700 116.580 137.650 116.600 ;
        RECT 131.050 115.655 132.105 115.675 ;
        RECT 130.700 115.650 133.125 115.655 ;
        RECT 114.350 114.625 116.275 115.625 ;
        RECT 93.165 114.545 95.675 114.550 ;
        RECT 95.865 114.545 112.990 114.550 ;
        RECT 105.625 114.530 106.680 114.545 ;
        RECT 88.905 112.300 89.945 113.250 ;
        RECT 88.925 112.275 89.925 112.300 ;
        RECT 90.680 112.275 91.770 113.275 ;
        RECT 82.325 107.400 83.350 108.400 ;
        RECT 83.825 107.400 84.770 107.925 ;
        RECT 82.845 106.275 83.885 106.750 ;
        RECT 78.175 105.925 79.175 105.930 ;
        RECT 71.900 105.900 73.225 105.925 ;
        RECT 78.145 105.900 79.205 105.925 ;
        RECT 82.845 105.900 83.350 106.275 ;
        RECT 84.195 105.945 84.770 107.400 ;
        RECT 71.900 104.900 77.100 105.900 ;
        RECT 78.125 105.875 83.350 105.900 ;
        RECT 78.125 104.925 83.370 105.875 ;
        RECT 78.125 104.900 83.350 104.925 ;
        RECT 71.900 104.885 73.225 104.900 ;
        RECT 70.455 102.950 71.495 103.900 ;
        RECT 70.475 102.925 71.480 102.950 ;
        RECT 71.110 100.700 71.480 102.925 ;
        RECT 71.900 100.700 72.270 104.885 ;
        RECT 74.005 101.775 75.005 104.900 ;
        RECT 78.175 104.870 79.175 104.900 ;
        RECT 82.845 104.525 83.350 104.900 ;
        RECT 83.775 104.855 84.775 105.945 ;
        RECT 85.735 105.900 86.105 111.925 ;
        RECT 85.100 104.900 86.105 105.900 ;
        RECT 82.845 104.030 83.885 104.525 ;
        RECT 84.195 103.625 84.770 104.855 ;
        RECT 82.350 103.250 83.405 103.625 ;
        RECT 83.825 103.250 84.770 103.625 ;
        RECT 73.985 100.825 75.025 101.775 ;
        RECT 74.005 100.800 75.005 100.825 ;
        RECT 66.600 100.655 67.600 100.700 ;
        RECT 73.965 99.860 75.080 99.890 ;
        RECT 80.180 99.860 81.295 99.885 ;
        RECT 82.350 99.860 83.350 103.250 ;
        RECT 85.105 101.700 86.105 104.900 ;
        RECT 83.905 100.700 86.105 101.700 ;
        RECT 86.525 105.945 86.895 111.925 ;
        RECT 90.725 111.500 91.725 111.530 ;
        RECT 90.725 110.500 93.495 111.500 ;
        RECT 90.725 110.470 91.725 110.500 ;
        RECT 87.750 107.400 88.750 109.850 ;
        RECT 89.225 107.400 90.170 107.925 ;
        RECT 90.450 107.400 91.450 109.850 ;
        RECT 91.925 107.400 92.870 107.925 ;
        RECT 88.245 106.275 89.285 106.750 ;
        RECT 86.525 105.900 87.525 105.945 ;
        RECT 88.245 105.900 88.750 106.275 ;
        RECT 89.595 105.900 90.170 107.400 ;
        RECT 90.945 106.275 91.985 106.750 ;
        RECT 90.945 105.900 91.450 106.275 ;
        RECT 92.295 105.900 92.870 107.400 ;
        RECT 93.835 105.900 94.205 111.925 ;
        RECT 94.625 105.900 94.995 111.925 ;
        RECT 96.535 105.900 96.905 111.925 ;
        RECT 86.525 105.875 88.750 105.900 ;
        RECT 86.525 104.930 88.770 105.875 ;
        RECT 86.525 104.900 88.750 104.930 ;
        RECT 89.130 104.900 91.450 105.900 ;
        RECT 91.875 104.900 94.205 105.900 ;
        RECT 94.580 104.900 95.670 105.900 ;
        RECT 86.525 104.855 87.525 104.900 ;
        RECT 86.525 100.700 86.895 104.855 ;
        RECT 88.245 104.525 88.750 104.900 ;
        RECT 88.245 104.030 89.285 104.525 ;
        RECT 89.595 103.625 90.170 104.900 ;
        RECT 90.945 104.525 91.450 104.900 ;
        RECT 90.945 104.030 91.985 104.525 ;
        RECT 92.295 103.625 92.870 104.900 ;
        RECT 87.750 103.250 88.805 103.625 ;
        RECT 89.225 103.250 90.170 103.625 ;
        RECT 90.450 103.250 91.505 103.625 ;
        RECT 91.925 103.250 92.870 103.625 ;
        RECT 87.750 102.375 88.750 103.250 ;
        RECT 90.450 102.375 91.450 103.250 ;
        RECT 87.750 101.375 91.450 102.375 ;
        RECT 92.025 101.700 93.025 101.745 ;
        RECT 93.205 101.700 94.205 104.900 ;
        RECT 87.750 99.860 88.750 101.375 ;
        RECT 92.025 100.700 94.205 101.700 ;
        RECT 94.625 100.700 94.995 104.900 ;
        RECT 95.900 103.900 96.905 105.900 ;
        RECT 97.325 105.900 97.695 111.925 ;
        RECT 107.750 108.400 108.750 114.545 ;
        RECT 114.350 113.250 115.350 114.625 ;
        RECT 117.875 114.550 139.150 115.650 ;
        RECT 140.700 115.625 141.700 116.600 ;
        RECT 147.500 116.580 148.450 116.600 ;
        RECT 139.775 114.625 141.700 115.625 ;
        RECT 118.590 114.545 121.100 114.550 ;
        RECT 121.290 114.545 138.415 114.550 ;
        RECT 131.050 114.530 132.105 114.545 ;
        RECT 114.330 112.300 115.370 113.250 ;
        RECT 114.350 112.275 115.350 112.300 ;
        RECT 116.105 112.275 117.195 113.275 ;
        RECT 107.750 107.400 108.775 108.400 ;
        RECT 109.250 107.400 110.195 107.925 ;
        RECT 108.270 106.275 109.310 106.750 ;
        RECT 103.600 105.925 104.600 105.930 ;
        RECT 103.570 105.900 104.630 105.925 ;
        RECT 108.270 105.900 108.775 106.275 ;
        RECT 109.620 105.945 110.195 107.400 ;
        RECT 97.325 104.900 102.570 105.900 ;
        RECT 103.550 105.875 108.775 105.900 ;
        RECT 103.550 104.925 108.795 105.875 ;
        RECT 103.550 104.900 108.775 104.925 ;
        RECT 95.880 102.950 96.920 103.900 ;
        RECT 95.900 102.925 96.905 102.950 ;
        RECT 96.535 100.700 96.905 102.925 ;
        RECT 97.325 100.700 97.695 104.900 ;
        RECT 99.430 101.775 100.430 104.900 ;
        RECT 103.600 104.870 104.600 104.900 ;
        RECT 108.270 104.525 108.775 104.900 ;
        RECT 109.200 104.855 110.200 105.945 ;
        RECT 111.160 105.900 111.530 111.925 ;
        RECT 110.525 104.900 111.530 105.900 ;
        RECT 108.270 104.030 109.310 104.525 ;
        RECT 109.620 103.625 110.195 104.855 ;
        RECT 107.775 103.250 108.830 103.625 ;
        RECT 109.250 103.250 110.195 103.625 ;
        RECT 99.410 100.825 100.450 101.775 ;
        RECT 99.430 100.800 100.430 100.825 ;
        RECT 92.025 100.655 93.025 100.700 ;
        RECT 99.390 99.860 100.505 99.890 ;
        RECT 105.605 99.860 106.720 99.885 ;
        RECT 107.775 99.860 108.775 103.250 ;
        RECT 110.530 101.700 111.530 104.900 ;
        RECT 109.330 100.700 111.530 101.700 ;
        RECT 111.950 105.945 112.320 111.925 ;
        RECT 116.150 111.500 117.150 111.530 ;
        RECT 116.150 110.500 118.920 111.500 ;
        RECT 116.150 110.470 117.150 110.500 ;
        RECT 113.175 107.400 114.175 109.850 ;
        RECT 114.650 107.400 115.595 107.925 ;
        RECT 115.875 107.400 116.875 109.850 ;
        RECT 117.350 107.400 118.295 107.925 ;
        RECT 113.670 106.275 114.710 106.750 ;
        RECT 111.950 105.900 112.950 105.945 ;
        RECT 113.670 105.900 114.175 106.275 ;
        RECT 115.020 105.900 115.595 107.400 ;
        RECT 116.370 106.275 117.410 106.750 ;
        RECT 116.370 105.900 116.875 106.275 ;
        RECT 117.720 105.900 118.295 107.400 ;
        RECT 119.260 105.900 119.630 111.925 ;
        RECT 120.050 105.900 120.420 111.925 ;
        RECT 121.960 105.900 122.330 111.925 ;
        RECT 111.950 105.875 114.175 105.900 ;
        RECT 111.950 104.930 114.195 105.875 ;
        RECT 111.950 104.900 114.175 104.930 ;
        RECT 114.555 104.900 116.875 105.900 ;
        RECT 117.300 104.900 119.630 105.900 ;
        RECT 120.005 104.900 121.095 105.900 ;
        RECT 111.950 104.855 112.950 104.900 ;
        RECT 111.950 100.700 112.320 104.855 ;
        RECT 113.670 104.525 114.175 104.900 ;
        RECT 113.670 104.030 114.710 104.525 ;
        RECT 115.020 103.625 115.595 104.900 ;
        RECT 116.370 104.525 116.875 104.900 ;
        RECT 116.370 104.030 117.410 104.525 ;
        RECT 117.720 103.625 118.295 104.900 ;
        RECT 113.175 103.250 114.230 103.625 ;
        RECT 114.650 103.250 115.595 103.625 ;
        RECT 115.875 103.250 116.930 103.625 ;
        RECT 117.350 103.250 118.295 103.625 ;
        RECT 113.175 102.375 114.175 103.250 ;
        RECT 115.875 102.375 116.875 103.250 ;
        RECT 113.175 101.375 116.875 102.375 ;
        RECT 117.450 101.700 118.450 101.745 ;
        RECT 118.630 101.700 119.630 104.900 ;
        RECT 113.175 99.860 114.175 101.375 ;
        RECT 117.450 100.700 119.630 101.700 ;
        RECT 120.050 100.700 120.420 104.900 ;
        RECT 121.325 103.900 122.330 105.900 ;
        RECT 122.750 105.925 123.120 111.925 ;
        RECT 133.175 108.400 134.175 114.545 ;
        RECT 139.775 113.250 140.775 114.625 ;
        RECT 143.300 114.550 149.225 115.650 ;
        RECT 144.015 114.545 146.525 114.550 ;
        RECT 146.715 114.545 149.215 114.550 ;
        RECT 139.755 112.300 140.795 113.250 ;
        RECT 139.775 112.275 140.775 112.300 ;
        RECT 141.530 112.275 142.620 113.275 ;
        RECT 133.175 107.400 134.200 108.400 ;
        RECT 134.675 107.400 135.620 107.925 ;
        RECT 133.695 106.275 134.735 106.750 ;
        RECT 129.025 105.925 130.025 105.930 ;
        RECT 122.750 105.900 124.075 105.925 ;
        RECT 128.995 105.900 130.055 105.925 ;
        RECT 133.695 105.900 134.200 106.275 ;
        RECT 135.045 105.945 135.620 107.400 ;
        RECT 122.750 104.900 127.950 105.900 ;
        RECT 128.975 105.875 134.200 105.900 ;
        RECT 128.975 104.925 134.220 105.875 ;
        RECT 128.975 104.900 134.200 104.925 ;
        RECT 122.750 104.885 124.075 104.900 ;
        RECT 121.305 102.950 122.345 103.900 ;
        RECT 121.325 102.925 122.330 102.950 ;
        RECT 121.960 100.700 122.330 102.925 ;
        RECT 122.750 100.700 123.120 104.885 ;
        RECT 124.855 101.775 125.855 104.900 ;
        RECT 129.025 104.870 130.025 104.900 ;
        RECT 133.695 104.525 134.200 104.900 ;
        RECT 134.625 104.855 135.625 105.945 ;
        RECT 136.585 105.900 136.955 111.925 ;
        RECT 135.950 104.900 136.955 105.900 ;
        RECT 133.695 104.030 134.735 104.525 ;
        RECT 135.045 103.625 135.620 104.855 ;
        RECT 133.200 103.250 134.255 103.625 ;
        RECT 134.675 103.250 135.620 103.625 ;
        RECT 124.835 100.825 125.875 101.775 ;
        RECT 124.855 100.800 125.855 100.825 ;
        RECT 117.450 100.655 118.450 100.700 ;
        RECT 124.815 99.860 125.930 99.890 ;
        RECT 131.030 99.860 132.145 99.885 ;
        RECT 133.200 99.860 134.200 103.250 ;
        RECT 135.955 101.700 136.955 104.900 ;
        RECT 134.755 100.700 136.955 101.700 ;
        RECT 137.375 105.945 137.745 111.925 ;
        RECT 141.575 111.500 142.575 111.530 ;
        RECT 141.575 110.500 144.345 111.500 ;
        RECT 141.575 110.470 142.575 110.500 ;
        RECT 138.600 107.400 139.600 109.850 ;
        RECT 140.075 107.400 141.020 107.925 ;
        RECT 141.300 107.400 142.300 109.850 ;
        RECT 142.775 107.400 143.720 107.925 ;
        RECT 139.095 106.275 140.135 106.750 ;
        RECT 137.375 105.900 138.375 105.945 ;
        RECT 139.095 105.900 139.600 106.275 ;
        RECT 140.445 105.900 141.020 107.400 ;
        RECT 141.795 106.275 142.835 106.750 ;
        RECT 141.795 105.900 142.300 106.275 ;
        RECT 143.145 105.900 143.720 107.400 ;
        RECT 144.685 105.900 145.055 111.925 ;
        RECT 145.475 105.900 145.845 111.925 ;
        RECT 147.385 105.900 147.755 111.925 ;
        RECT 137.375 105.875 139.600 105.900 ;
        RECT 137.375 104.930 139.620 105.875 ;
        RECT 137.375 104.900 139.600 104.930 ;
        RECT 139.980 104.900 142.300 105.900 ;
        RECT 142.725 104.900 145.055 105.900 ;
        RECT 145.430 104.900 146.520 105.900 ;
        RECT 137.375 104.855 138.375 104.900 ;
        RECT 137.375 100.700 137.745 104.855 ;
        RECT 139.095 104.525 139.600 104.900 ;
        RECT 139.095 104.030 140.135 104.525 ;
        RECT 140.445 103.625 141.020 104.900 ;
        RECT 141.795 104.525 142.300 104.900 ;
        RECT 141.795 104.030 142.835 104.525 ;
        RECT 143.145 103.625 143.720 104.900 ;
        RECT 138.600 103.250 139.655 103.625 ;
        RECT 140.075 103.250 141.020 103.625 ;
        RECT 141.300 103.250 142.355 103.625 ;
        RECT 142.775 103.250 143.720 103.625 ;
        RECT 138.600 102.375 139.600 103.250 ;
        RECT 141.300 102.375 142.300 103.250 ;
        RECT 138.600 101.375 142.300 102.375 ;
        RECT 142.875 101.700 143.875 101.745 ;
        RECT 144.055 101.700 145.055 104.900 ;
        RECT 138.600 99.860 139.600 101.375 ;
        RECT 142.875 100.700 145.055 101.700 ;
        RECT 145.475 100.700 145.845 104.900 ;
        RECT 146.750 103.900 147.755 105.900 ;
        RECT 148.175 105.900 148.545 111.925 ;
        RECT 154.525 105.900 155.525 105.945 ;
        RECT 148.175 104.900 155.525 105.900 ;
        RECT 146.730 102.950 147.770 103.900 ;
        RECT 146.750 102.925 147.755 102.950 ;
        RECT 147.385 100.700 147.755 102.925 ;
        RECT 148.175 100.700 148.545 104.900 ;
        RECT 150.280 101.775 151.280 104.900 ;
        RECT 154.525 104.855 155.525 104.900 ;
        RECT 150.260 100.825 151.300 101.775 ;
        RECT 150.280 100.800 151.280 100.825 ;
        RECT 142.875 100.655 143.875 100.700 ;
        RECT 150.240 99.860 151.355 99.890 ;
        RECT 1.850 99.850 14.575 99.860 ;
        RECT 15.350 99.850 19.390 99.860 ;
        RECT 19.590 99.850 40.000 99.860 ;
        RECT 40.775 99.850 44.815 99.860 ;
        RECT 45.015 99.850 65.425 99.860 ;
        RECT 66.200 99.850 70.240 99.860 ;
        RECT 70.440 99.850 90.850 99.860 ;
        RECT 91.625 99.850 95.665 99.860 ;
        RECT 95.865 99.850 116.275 99.860 ;
        RECT 117.050 99.850 121.090 99.860 ;
        RECT 121.290 99.850 141.700 99.860 ;
        RECT 142.475 99.850 146.515 99.860 ;
        RECT 146.715 99.850 151.355 99.860 ;
        RECT 1.850 98.750 151.355 99.850 ;
        RECT 1.850 98.745 19.390 98.750 ;
        RECT 19.590 98.745 44.815 98.750 ;
        RECT 45.015 98.745 70.240 98.750 ;
        RECT 70.440 98.745 95.665 98.750 ;
        RECT 95.865 98.745 121.090 98.750 ;
        RECT 121.290 98.745 146.515 98.750 ;
        RECT 146.715 98.745 151.355 98.750 ;
        RECT 3.875 98.740 7.105 98.745 ;
        RECT 3.905 98.710 5.020 98.740 ;
        RECT 23.115 98.715 24.230 98.745 ;
        RECT 29.300 98.740 32.530 98.745 ;
        RECT 29.330 98.710 30.445 98.740 ;
        RECT 48.540 98.715 49.655 98.745 ;
        RECT 54.725 98.740 57.955 98.745 ;
        RECT 54.755 98.710 55.870 98.740 ;
        RECT 73.965 98.715 75.080 98.745 ;
        RECT 80.150 98.740 83.380 98.745 ;
        RECT 80.180 98.710 81.295 98.740 ;
        RECT 99.390 98.715 100.505 98.745 ;
        RECT 105.575 98.740 108.805 98.745 ;
        RECT 105.605 98.710 106.720 98.740 ;
        RECT 124.815 98.715 125.930 98.745 ;
        RECT 131.000 98.740 134.230 98.745 ;
        RECT 131.030 98.710 132.145 98.740 ;
        RECT 150.240 98.715 151.355 98.745 ;
        RECT 19.370 97.800 21.325 97.820 ;
        RECT 44.795 97.800 46.750 97.820 ;
        RECT 70.220 97.800 72.175 97.820 ;
        RECT 95.645 97.800 97.600 97.820 ;
        RECT 121.070 97.800 123.025 97.820 ;
        RECT 146.495 97.800 148.450 97.820 ;
        RECT 9.550 97.775 10.550 97.800 ;
        RECT 15.750 97.775 16.750 97.800 ;
        RECT 17.650 97.775 18.650 97.800 ;
        RECT 9.530 96.825 10.570 97.775 ;
        RECT 15.730 96.825 16.770 97.775 ;
        RECT 17.630 96.825 18.670 97.775 ;
        RECT 9.550 96.800 10.550 96.825 ;
        RECT 15.750 96.800 16.750 96.825 ;
        RECT 17.650 96.800 18.650 96.825 ;
        RECT 19.365 96.800 21.350 97.800 ;
        RECT 34.975 97.775 35.975 97.800 ;
        RECT 41.175 97.775 42.175 97.800 ;
        RECT 43.075 97.775 44.075 97.800 ;
        RECT 34.955 96.825 35.995 97.775 ;
        RECT 41.155 96.825 42.195 97.775 ;
        RECT 43.055 96.825 44.095 97.775 ;
        RECT 34.975 96.800 35.975 96.825 ;
        RECT 41.175 96.800 42.175 96.825 ;
        RECT 43.075 96.800 44.075 96.825 ;
        RECT 44.790 96.800 46.775 97.800 ;
        RECT 60.400 97.775 61.400 97.800 ;
        RECT 66.600 97.775 67.600 97.800 ;
        RECT 68.500 97.775 69.500 97.800 ;
        RECT 60.380 96.825 61.420 97.775 ;
        RECT 66.580 96.825 67.620 97.775 ;
        RECT 68.480 96.825 69.520 97.775 ;
        RECT 60.400 96.800 61.400 96.825 ;
        RECT 66.600 96.800 67.600 96.825 ;
        RECT 68.500 96.800 69.500 96.825 ;
        RECT 70.215 96.800 72.200 97.800 ;
        RECT 85.825 97.775 86.825 97.800 ;
        RECT 92.025 97.775 93.025 97.800 ;
        RECT 93.925 97.775 94.925 97.800 ;
        RECT 85.805 96.825 86.845 97.775 ;
        RECT 92.005 96.825 93.045 97.775 ;
        RECT 93.905 96.825 94.945 97.775 ;
        RECT 85.825 96.800 86.825 96.825 ;
        RECT 92.025 96.800 93.025 96.825 ;
        RECT 93.925 96.800 94.925 96.825 ;
        RECT 95.640 96.800 97.625 97.800 ;
        RECT 111.250 97.775 112.250 97.800 ;
        RECT 117.450 97.775 118.450 97.800 ;
        RECT 119.350 97.775 120.350 97.800 ;
        RECT 111.230 96.825 112.270 97.775 ;
        RECT 117.430 96.825 118.470 97.775 ;
        RECT 119.330 96.825 120.370 97.775 ;
        RECT 111.250 96.800 112.250 96.825 ;
        RECT 117.450 96.800 118.450 96.825 ;
        RECT 119.350 96.800 120.350 96.825 ;
        RECT 121.065 96.800 123.050 97.800 ;
        RECT 136.675 97.775 137.675 97.800 ;
        RECT 142.875 97.775 143.875 97.800 ;
        RECT 144.775 97.775 145.775 97.800 ;
        RECT 136.655 96.825 137.695 97.775 ;
        RECT 142.855 96.825 143.895 97.775 ;
        RECT 144.755 96.825 145.795 97.775 ;
        RECT 136.675 96.800 137.675 96.825 ;
        RECT 142.875 96.800 143.875 96.825 ;
        RECT 144.775 96.800 145.775 96.825 ;
        RECT 146.490 96.800 148.475 97.800 ;
        RECT 19.370 96.780 21.325 96.800 ;
        RECT 44.795 96.780 46.750 96.800 ;
        RECT 70.220 96.780 72.175 96.800 ;
        RECT 95.645 96.780 97.600 96.800 ;
        RECT 121.070 96.780 123.025 96.800 ;
        RECT 146.495 96.780 148.450 96.800 ;
        RECT 9.575 95.025 10.525 95.045 ;
        RECT 20.375 95.025 21.325 95.045 ;
        RECT 35.000 95.025 35.950 95.045 ;
        RECT 45.800 95.025 46.750 95.045 ;
        RECT 60.425 95.025 61.375 95.045 ;
        RECT 71.225 95.025 72.175 95.045 ;
        RECT 85.850 95.025 86.800 95.045 ;
        RECT 96.650 95.025 97.600 95.045 ;
        RECT 111.275 95.025 112.225 95.045 ;
        RECT 122.075 95.025 123.025 95.045 ;
        RECT 136.700 95.025 137.650 95.045 ;
        RECT 147.500 95.025 148.450 95.045 ;
        RECT 9.550 94.025 12.755 95.025 ;
        RECT 13.530 94.025 14.620 95.025 ;
        RECT 15.370 94.025 18.650 95.025 ;
        RECT 20.350 94.025 21.350 95.025 ;
        RECT 9.575 94.005 10.525 94.025 ;
        RECT 2.900 93.075 7.100 93.080 ;
        RECT 1.850 91.975 12.025 93.075 ;
        RECT 13.575 93.050 14.575 94.025 ;
        RECT 20.375 94.005 21.325 94.025 ;
        RECT 23.155 93.730 24.155 94.825 ;
        RECT 34.975 94.025 38.180 95.025 ;
        RECT 38.955 94.025 40.045 95.025 ;
        RECT 40.795 94.025 44.075 95.025 ;
        RECT 45.775 94.025 46.775 95.025 ;
        RECT 35.000 94.005 35.950 94.025 ;
        RECT 23.430 93.115 23.880 93.730 ;
        RECT 28.325 93.075 32.525 93.080 ;
        RECT 12.650 92.050 14.575 93.050 ;
        RECT 16.175 92.155 22.100 93.075 ;
        RECT 27.275 92.155 37.450 93.075 ;
        RECT 39.000 93.050 40.000 94.025 ;
        RECT 45.800 94.005 46.750 94.025 ;
        RECT 48.580 93.730 49.580 94.825 ;
        RECT 60.400 94.025 63.605 95.025 ;
        RECT 64.380 94.025 65.470 95.025 ;
        RECT 66.220 94.025 69.500 95.025 ;
        RECT 71.200 94.025 72.200 95.025 ;
        RECT 60.425 94.005 61.375 94.025 ;
        RECT 48.855 93.115 49.305 93.730 ;
        RECT 53.750 93.075 57.950 93.080 ;
        RECT 1.850 91.970 11.290 91.975 ;
        RECT 6.050 85.825 7.050 91.970 ;
        RECT 12.650 90.675 13.650 92.050 ;
        RECT 16.175 91.975 37.450 92.155 ;
        RECT 38.075 92.050 40.000 93.050 ;
        RECT 41.600 92.155 47.525 93.075 ;
        RECT 52.700 92.155 62.875 93.075 ;
        RECT 64.425 93.050 65.425 94.025 ;
        RECT 71.225 94.005 72.175 94.025 ;
        RECT 74.005 93.730 75.005 94.825 ;
        RECT 85.825 94.025 89.030 95.025 ;
        RECT 89.805 94.025 90.895 95.025 ;
        RECT 91.645 94.025 94.925 95.025 ;
        RECT 96.625 94.025 97.625 95.025 ;
        RECT 85.850 94.005 86.800 94.025 ;
        RECT 74.280 93.115 74.730 93.730 ;
        RECT 79.175 93.075 83.375 93.080 ;
        RECT 16.890 91.970 19.400 91.975 ;
        RECT 19.590 91.970 36.715 91.975 ;
        RECT 20.320 91.050 28.380 91.970 ;
        RECT 12.630 89.725 13.670 90.675 ;
        RECT 12.650 89.700 13.650 89.725 ;
        RECT 14.405 89.700 15.495 90.700 ;
        RECT 6.050 84.825 7.075 85.825 ;
        RECT 7.550 84.825 8.495 85.350 ;
        RECT 6.570 83.700 7.610 84.175 ;
        RECT 1.900 83.325 2.900 83.355 ;
        RECT 6.570 83.325 7.075 83.700 ;
        RECT 7.920 83.370 8.495 84.825 ;
        RECT 1.850 83.300 7.075 83.325 ;
        RECT 1.850 82.350 7.095 83.300 ;
        RECT 1.850 82.325 7.075 82.350 ;
        RECT 1.900 82.295 2.900 82.325 ;
        RECT 6.570 81.950 7.075 82.325 ;
        RECT 7.500 82.280 8.500 83.370 ;
        RECT 9.460 83.325 9.830 89.350 ;
        RECT 8.825 82.325 9.830 83.325 ;
        RECT 6.570 81.455 7.610 81.950 ;
        RECT 7.920 81.050 8.495 82.280 ;
        RECT 6.075 80.675 7.130 81.050 ;
        RECT 7.550 80.675 8.495 81.050 ;
        RECT 3.890 77.285 5.030 77.315 ;
        RECT 6.075 77.285 7.075 80.675 ;
        RECT 8.830 79.125 9.830 82.325 ;
        RECT 7.630 78.125 9.830 79.125 ;
        RECT 10.250 83.370 10.620 89.350 ;
        RECT 14.450 88.925 15.450 88.955 ;
        RECT 14.450 87.925 17.220 88.925 ;
        RECT 14.450 87.895 15.450 87.925 ;
        RECT 11.475 84.825 12.475 87.275 ;
        RECT 12.950 84.825 13.895 85.350 ;
        RECT 14.175 84.825 15.175 87.275 ;
        RECT 15.650 84.825 16.595 85.350 ;
        RECT 11.970 83.700 13.010 84.175 ;
        RECT 10.250 83.325 11.250 83.370 ;
        RECT 11.970 83.325 12.475 83.700 ;
        RECT 13.320 83.325 13.895 84.825 ;
        RECT 14.670 83.700 15.710 84.175 ;
        RECT 14.670 83.325 15.175 83.700 ;
        RECT 16.020 83.325 16.595 84.825 ;
        RECT 17.560 83.325 17.930 89.350 ;
        RECT 18.350 83.325 18.720 89.350 ;
        RECT 20.260 83.325 20.630 89.350 ;
        RECT 10.250 83.300 12.475 83.325 ;
        RECT 10.250 82.355 12.495 83.300 ;
        RECT 10.250 82.325 12.475 82.355 ;
        RECT 12.855 82.325 15.175 83.325 ;
        RECT 15.600 82.325 17.930 83.325 ;
        RECT 18.305 82.325 19.395 83.325 ;
        RECT 19.625 82.325 20.630 83.325 ;
        RECT 10.250 82.280 11.250 82.325 ;
        RECT 10.250 78.125 10.620 82.280 ;
        RECT 11.970 81.950 12.475 82.325 ;
        RECT 11.970 81.455 13.010 81.950 ;
        RECT 13.320 81.050 13.895 82.325 ;
        RECT 14.670 81.950 15.175 82.325 ;
        RECT 14.670 81.455 15.710 81.950 ;
        RECT 16.020 81.050 16.595 82.325 ;
        RECT 11.475 80.675 12.530 81.050 ;
        RECT 12.950 80.675 13.895 81.050 ;
        RECT 14.175 80.675 15.230 81.050 ;
        RECT 15.650 80.675 16.595 81.050 ;
        RECT 11.475 79.800 12.475 80.675 ;
        RECT 14.175 79.800 15.175 80.675 ;
        RECT 11.475 78.800 15.175 79.800 ;
        RECT 15.750 79.125 16.750 79.170 ;
        RECT 16.930 79.125 17.930 82.325 ;
        RECT 11.475 77.285 12.475 78.800 ;
        RECT 15.750 78.125 17.930 79.125 ;
        RECT 18.350 78.125 18.720 82.325 ;
        RECT 19.630 81.325 20.630 82.325 ;
        RECT 21.050 83.325 21.420 89.350 ;
        RECT 31.475 85.825 32.475 91.970 ;
        RECT 38.075 90.675 39.075 92.050 ;
        RECT 41.600 91.975 62.875 92.155 ;
        RECT 63.500 92.050 65.425 93.050 ;
        RECT 67.025 92.155 72.950 93.075 ;
        RECT 78.125 92.155 88.300 93.075 ;
        RECT 89.850 93.050 90.850 94.025 ;
        RECT 96.650 94.005 97.600 94.025 ;
        RECT 99.430 93.730 100.430 94.825 ;
        RECT 111.250 94.025 114.455 95.025 ;
        RECT 115.230 94.025 116.320 95.025 ;
        RECT 117.070 94.025 120.350 95.025 ;
        RECT 122.050 94.025 123.050 95.025 ;
        RECT 111.275 94.005 112.225 94.025 ;
        RECT 99.705 93.115 100.155 93.730 ;
        RECT 104.600 93.075 108.800 93.080 ;
        RECT 42.315 91.970 44.825 91.975 ;
        RECT 45.015 91.970 62.140 91.975 ;
        RECT 45.745 91.050 53.805 91.970 ;
        RECT 38.055 89.725 39.095 90.675 ;
        RECT 38.075 89.700 39.075 89.725 ;
        RECT 39.830 89.700 40.920 90.700 ;
        RECT 31.475 84.825 32.500 85.825 ;
        RECT 32.975 84.825 33.920 85.350 ;
        RECT 23.430 83.875 23.880 84.515 ;
        RECT 23.150 83.325 24.150 83.875 ;
        RECT 31.995 83.700 33.035 84.175 ;
        RECT 27.325 83.325 28.325 83.355 ;
        RECT 31.995 83.325 32.500 83.700 ;
        RECT 33.345 83.370 33.920 84.825 ;
        RECT 21.050 82.325 24.150 83.325 ;
        RECT 27.275 83.300 32.500 83.325 ;
        RECT 27.275 82.350 32.520 83.300 ;
        RECT 27.275 82.325 32.500 82.350 ;
        RECT 19.585 80.325 20.675 81.325 ;
        RECT 20.260 78.125 20.630 80.325 ;
        RECT 21.050 78.125 21.420 82.325 ;
        RECT 23.430 82.205 23.880 82.325 ;
        RECT 27.325 82.295 28.325 82.325 ;
        RECT 31.995 81.950 32.500 82.325 ;
        RECT 32.925 82.280 33.925 83.370 ;
        RECT 34.885 83.325 35.255 89.350 ;
        RECT 34.250 82.325 35.255 83.325 ;
        RECT 31.995 81.455 33.035 81.950 ;
        RECT 33.345 81.050 33.920 82.280 ;
        RECT 31.500 80.675 32.555 81.050 ;
        RECT 32.975 80.675 33.920 81.050 ;
        RECT 15.750 78.080 16.750 78.125 ;
        RECT 29.315 77.285 30.455 77.315 ;
        RECT 31.500 77.285 32.500 80.675 ;
        RECT 34.255 79.125 35.255 82.325 ;
        RECT 33.055 78.125 35.255 79.125 ;
        RECT 35.675 83.370 36.045 89.350 ;
        RECT 39.875 88.925 40.875 88.955 ;
        RECT 39.875 87.925 42.645 88.925 ;
        RECT 39.875 87.895 40.875 87.925 ;
        RECT 36.900 84.825 37.900 87.275 ;
        RECT 38.375 84.825 39.320 85.350 ;
        RECT 39.600 84.825 40.600 87.275 ;
        RECT 41.075 84.825 42.020 85.350 ;
        RECT 37.395 83.700 38.435 84.175 ;
        RECT 35.675 83.325 36.675 83.370 ;
        RECT 37.395 83.325 37.900 83.700 ;
        RECT 38.745 83.325 39.320 84.825 ;
        RECT 40.095 83.700 41.135 84.175 ;
        RECT 40.095 83.325 40.600 83.700 ;
        RECT 41.445 83.325 42.020 84.825 ;
        RECT 42.985 83.325 43.355 89.350 ;
        RECT 43.775 83.325 44.145 89.350 ;
        RECT 45.685 83.325 46.055 89.350 ;
        RECT 35.675 83.300 37.900 83.325 ;
        RECT 35.675 82.355 37.920 83.300 ;
        RECT 35.675 82.325 37.900 82.355 ;
        RECT 38.280 82.325 40.600 83.325 ;
        RECT 41.025 82.325 43.355 83.325 ;
        RECT 43.730 82.325 44.820 83.325 ;
        RECT 45.050 82.325 46.055 83.325 ;
        RECT 35.675 82.280 36.675 82.325 ;
        RECT 35.675 78.125 36.045 82.280 ;
        RECT 37.395 81.950 37.900 82.325 ;
        RECT 37.395 81.455 38.435 81.950 ;
        RECT 38.745 81.050 39.320 82.325 ;
        RECT 40.095 81.950 40.600 82.325 ;
        RECT 40.095 81.455 41.135 81.950 ;
        RECT 41.445 81.050 42.020 82.325 ;
        RECT 36.900 80.675 37.955 81.050 ;
        RECT 38.375 80.675 39.320 81.050 ;
        RECT 39.600 80.675 40.655 81.050 ;
        RECT 41.075 80.675 42.020 81.050 ;
        RECT 36.900 79.800 37.900 80.675 ;
        RECT 39.600 79.800 40.600 80.675 ;
        RECT 36.900 78.800 40.600 79.800 ;
        RECT 41.175 79.125 42.175 79.170 ;
        RECT 42.355 79.125 43.355 82.325 ;
        RECT 36.900 77.285 37.900 78.800 ;
        RECT 41.175 78.125 43.355 79.125 ;
        RECT 43.775 78.125 44.145 82.325 ;
        RECT 45.055 81.325 46.055 82.325 ;
        RECT 46.475 83.325 46.845 89.350 ;
        RECT 56.900 85.825 57.900 91.970 ;
        RECT 63.500 90.675 64.500 92.050 ;
        RECT 67.025 91.975 88.300 92.155 ;
        RECT 88.925 92.050 90.850 93.050 ;
        RECT 92.450 92.155 98.375 93.075 ;
        RECT 103.550 92.155 113.725 93.075 ;
        RECT 115.275 93.050 116.275 94.025 ;
        RECT 122.075 94.005 123.025 94.025 ;
        RECT 124.855 93.730 125.855 94.825 ;
        RECT 136.675 94.025 139.880 95.025 ;
        RECT 140.655 94.025 141.745 95.025 ;
        RECT 142.495 94.025 145.775 95.025 ;
        RECT 147.475 94.025 148.475 95.025 ;
        RECT 136.700 94.005 137.650 94.025 ;
        RECT 125.130 93.115 125.580 93.730 ;
        RECT 130.025 93.075 134.225 93.080 ;
        RECT 67.740 91.970 70.250 91.975 ;
        RECT 70.440 91.970 87.565 91.975 ;
        RECT 71.170 91.050 79.230 91.970 ;
        RECT 63.480 89.725 64.520 90.675 ;
        RECT 63.500 89.700 64.500 89.725 ;
        RECT 65.255 89.700 66.345 90.700 ;
        RECT 56.900 84.825 57.925 85.825 ;
        RECT 58.400 84.825 59.345 85.350 ;
        RECT 48.855 83.875 49.305 84.515 ;
        RECT 48.575 83.325 49.575 83.875 ;
        RECT 57.420 83.700 58.460 84.175 ;
        RECT 52.750 83.325 53.750 83.355 ;
        RECT 57.420 83.325 57.925 83.700 ;
        RECT 58.770 83.370 59.345 84.825 ;
        RECT 46.475 82.325 49.575 83.325 ;
        RECT 52.700 83.300 57.925 83.325 ;
        RECT 52.700 82.350 57.945 83.300 ;
        RECT 52.700 82.325 57.925 82.350 ;
        RECT 45.010 80.325 46.100 81.325 ;
        RECT 45.685 78.125 46.055 80.325 ;
        RECT 46.475 78.125 46.845 82.325 ;
        RECT 48.855 82.205 49.305 82.325 ;
        RECT 52.750 82.295 53.750 82.325 ;
        RECT 57.420 81.950 57.925 82.325 ;
        RECT 58.350 82.280 59.350 83.370 ;
        RECT 60.310 83.325 60.680 89.350 ;
        RECT 59.675 82.325 60.680 83.325 ;
        RECT 57.420 81.455 58.460 81.950 ;
        RECT 58.770 81.050 59.345 82.280 ;
        RECT 56.925 80.675 57.980 81.050 ;
        RECT 58.400 80.675 59.345 81.050 ;
        RECT 41.175 78.080 42.175 78.125 ;
        RECT 54.740 77.285 55.880 77.315 ;
        RECT 56.925 77.285 57.925 80.675 ;
        RECT 59.680 79.125 60.680 82.325 ;
        RECT 58.480 78.125 60.680 79.125 ;
        RECT 61.100 83.370 61.470 89.350 ;
        RECT 65.300 88.925 66.300 88.955 ;
        RECT 65.300 87.925 68.070 88.925 ;
        RECT 65.300 87.895 66.300 87.925 ;
        RECT 62.325 84.825 63.325 87.275 ;
        RECT 63.800 84.825 64.745 85.350 ;
        RECT 65.025 84.825 66.025 87.275 ;
        RECT 66.500 84.825 67.445 85.350 ;
        RECT 62.820 83.700 63.860 84.175 ;
        RECT 61.100 83.325 62.100 83.370 ;
        RECT 62.820 83.325 63.325 83.700 ;
        RECT 64.170 83.325 64.745 84.825 ;
        RECT 65.520 83.700 66.560 84.175 ;
        RECT 65.520 83.325 66.025 83.700 ;
        RECT 66.870 83.325 67.445 84.825 ;
        RECT 68.410 83.325 68.780 89.350 ;
        RECT 69.200 83.325 69.570 89.350 ;
        RECT 71.110 83.325 71.480 89.350 ;
        RECT 61.100 83.300 63.325 83.325 ;
        RECT 61.100 82.355 63.345 83.300 ;
        RECT 61.100 82.325 63.325 82.355 ;
        RECT 63.705 82.325 66.025 83.325 ;
        RECT 66.450 82.325 68.780 83.325 ;
        RECT 69.155 82.325 70.245 83.325 ;
        RECT 70.475 82.325 71.480 83.325 ;
        RECT 61.100 82.280 62.100 82.325 ;
        RECT 61.100 78.125 61.470 82.280 ;
        RECT 62.820 81.950 63.325 82.325 ;
        RECT 62.820 81.455 63.860 81.950 ;
        RECT 64.170 81.050 64.745 82.325 ;
        RECT 65.520 81.950 66.025 82.325 ;
        RECT 65.520 81.455 66.560 81.950 ;
        RECT 66.870 81.050 67.445 82.325 ;
        RECT 62.325 80.675 63.380 81.050 ;
        RECT 63.800 80.675 64.745 81.050 ;
        RECT 65.025 80.675 66.080 81.050 ;
        RECT 66.500 80.675 67.445 81.050 ;
        RECT 62.325 79.800 63.325 80.675 ;
        RECT 65.025 79.800 66.025 80.675 ;
        RECT 62.325 78.800 66.025 79.800 ;
        RECT 66.600 79.125 67.600 79.170 ;
        RECT 67.780 79.125 68.780 82.325 ;
        RECT 62.325 77.285 63.325 78.800 ;
        RECT 66.600 78.125 68.780 79.125 ;
        RECT 69.200 78.125 69.570 82.325 ;
        RECT 70.480 81.325 71.480 82.325 ;
        RECT 71.900 83.325 72.270 89.350 ;
        RECT 82.325 85.825 83.325 91.970 ;
        RECT 88.925 90.675 89.925 92.050 ;
        RECT 92.450 91.975 113.725 92.155 ;
        RECT 114.350 92.050 116.275 93.050 ;
        RECT 117.875 92.155 123.800 93.075 ;
        RECT 128.975 92.155 139.150 93.075 ;
        RECT 140.700 93.050 141.700 94.025 ;
        RECT 147.500 94.005 148.450 94.025 ;
        RECT 150.280 93.730 151.280 94.825 ;
        RECT 150.555 93.115 151.005 93.730 ;
        RECT 93.165 91.970 95.675 91.975 ;
        RECT 95.865 91.970 112.990 91.975 ;
        RECT 96.595 91.050 104.655 91.970 ;
        RECT 88.905 89.725 89.945 90.675 ;
        RECT 88.925 89.700 89.925 89.725 ;
        RECT 90.680 89.700 91.770 90.700 ;
        RECT 82.325 84.825 83.350 85.825 ;
        RECT 83.825 84.825 84.770 85.350 ;
        RECT 74.280 83.875 74.730 84.515 ;
        RECT 74.000 83.325 75.000 83.875 ;
        RECT 82.845 83.700 83.885 84.175 ;
        RECT 78.175 83.325 79.175 83.355 ;
        RECT 82.845 83.325 83.350 83.700 ;
        RECT 84.195 83.370 84.770 84.825 ;
        RECT 71.900 82.325 75.000 83.325 ;
        RECT 78.125 83.300 83.350 83.325 ;
        RECT 78.125 82.350 83.370 83.300 ;
        RECT 78.125 82.325 83.350 82.350 ;
        RECT 70.435 80.325 71.525 81.325 ;
        RECT 71.110 78.125 71.480 80.325 ;
        RECT 71.900 78.125 72.270 82.325 ;
        RECT 74.280 82.205 74.730 82.325 ;
        RECT 78.175 82.295 79.175 82.325 ;
        RECT 82.845 81.950 83.350 82.325 ;
        RECT 83.775 82.280 84.775 83.370 ;
        RECT 85.735 83.325 86.105 89.350 ;
        RECT 85.100 82.325 86.105 83.325 ;
        RECT 82.845 81.455 83.885 81.950 ;
        RECT 84.195 81.050 84.770 82.280 ;
        RECT 82.350 80.675 83.405 81.050 ;
        RECT 83.825 80.675 84.770 81.050 ;
        RECT 66.600 78.080 67.600 78.125 ;
        RECT 80.165 77.285 81.305 77.315 ;
        RECT 82.350 77.285 83.350 80.675 ;
        RECT 85.105 79.125 86.105 82.325 ;
        RECT 83.905 78.125 86.105 79.125 ;
        RECT 86.525 83.370 86.895 89.350 ;
        RECT 90.725 88.925 91.725 88.955 ;
        RECT 90.725 87.925 93.495 88.925 ;
        RECT 90.725 87.895 91.725 87.925 ;
        RECT 87.750 84.825 88.750 87.275 ;
        RECT 89.225 84.825 90.170 85.350 ;
        RECT 90.450 84.825 91.450 87.275 ;
        RECT 91.925 84.825 92.870 85.350 ;
        RECT 88.245 83.700 89.285 84.175 ;
        RECT 86.525 83.325 87.525 83.370 ;
        RECT 88.245 83.325 88.750 83.700 ;
        RECT 89.595 83.325 90.170 84.825 ;
        RECT 90.945 83.700 91.985 84.175 ;
        RECT 90.945 83.325 91.450 83.700 ;
        RECT 92.295 83.325 92.870 84.825 ;
        RECT 93.835 83.325 94.205 89.350 ;
        RECT 94.625 83.325 94.995 89.350 ;
        RECT 96.535 83.325 96.905 89.350 ;
        RECT 86.525 83.300 88.750 83.325 ;
        RECT 86.525 82.355 88.770 83.300 ;
        RECT 86.525 82.325 88.750 82.355 ;
        RECT 89.130 82.325 91.450 83.325 ;
        RECT 91.875 82.325 94.205 83.325 ;
        RECT 94.580 82.325 95.670 83.325 ;
        RECT 95.900 82.325 96.905 83.325 ;
        RECT 86.525 82.280 87.525 82.325 ;
        RECT 86.525 78.125 86.895 82.280 ;
        RECT 88.245 81.950 88.750 82.325 ;
        RECT 88.245 81.455 89.285 81.950 ;
        RECT 89.595 81.050 90.170 82.325 ;
        RECT 90.945 81.950 91.450 82.325 ;
        RECT 90.945 81.455 91.985 81.950 ;
        RECT 92.295 81.050 92.870 82.325 ;
        RECT 87.750 80.675 88.805 81.050 ;
        RECT 89.225 80.675 90.170 81.050 ;
        RECT 90.450 80.675 91.505 81.050 ;
        RECT 91.925 80.675 92.870 81.050 ;
        RECT 87.750 79.800 88.750 80.675 ;
        RECT 90.450 79.800 91.450 80.675 ;
        RECT 87.750 78.800 91.450 79.800 ;
        RECT 92.025 79.125 93.025 79.170 ;
        RECT 93.205 79.125 94.205 82.325 ;
        RECT 87.750 77.285 88.750 78.800 ;
        RECT 92.025 78.125 94.205 79.125 ;
        RECT 94.625 78.125 94.995 82.325 ;
        RECT 95.905 81.325 96.905 82.325 ;
        RECT 97.325 83.325 97.695 89.350 ;
        RECT 107.750 85.825 108.750 91.970 ;
        RECT 114.350 90.675 115.350 92.050 ;
        RECT 117.875 91.975 139.150 92.155 ;
        RECT 139.775 92.050 141.700 93.050 ;
        RECT 118.590 91.970 121.100 91.975 ;
        RECT 121.290 91.970 138.415 91.975 ;
        RECT 122.020 91.050 130.080 91.970 ;
        RECT 114.330 89.725 115.370 90.675 ;
        RECT 114.350 89.700 115.350 89.725 ;
        RECT 116.105 89.700 117.195 90.700 ;
        RECT 107.750 84.825 108.775 85.825 ;
        RECT 109.250 84.825 110.195 85.350 ;
        RECT 99.705 83.875 100.155 84.515 ;
        RECT 99.425 83.325 100.425 83.875 ;
        RECT 108.270 83.700 109.310 84.175 ;
        RECT 103.600 83.325 104.600 83.355 ;
        RECT 108.270 83.325 108.775 83.700 ;
        RECT 109.620 83.370 110.195 84.825 ;
        RECT 97.325 82.325 100.425 83.325 ;
        RECT 103.550 83.300 108.775 83.325 ;
        RECT 103.550 82.350 108.795 83.300 ;
        RECT 103.550 82.325 108.775 82.350 ;
        RECT 95.860 80.325 96.950 81.325 ;
        RECT 96.535 78.125 96.905 80.325 ;
        RECT 97.325 78.125 97.695 82.325 ;
        RECT 99.705 82.205 100.155 82.325 ;
        RECT 103.600 82.295 104.600 82.325 ;
        RECT 108.270 81.950 108.775 82.325 ;
        RECT 109.200 82.280 110.200 83.370 ;
        RECT 111.160 83.325 111.530 89.350 ;
        RECT 110.525 82.325 111.530 83.325 ;
        RECT 108.270 81.455 109.310 81.950 ;
        RECT 109.620 81.050 110.195 82.280 ;
        RECT 107.775 80.675 108.830 81.050 ;
        RECT 109.250 80.675 110.195 81.050 ;
        RECT 92.025 78.080 93.025 78.125 ;
        RECT 105.590 77.285 106.730 77.315 ;
        RECT 107.775 77.285 108.775 80.675 ;
        RECT 110.530 79.125 111.530 82.325 ;
        RECT 109.330 78.125 111.530 79.125 ;
        RECT 111.950 83.370 112.320 89.350 ;
        RECT 116.150 88.925 117.150 88.955 ;
        RECT 116.150 87.925 118.920 88.925 ;
        RECT 116.150 87.895 117.150 87.925 ;
        RECT 113.175 84.825 114.175 87.275 ;
        RECT 114.650 84.825 115.595 85.350 ;
        RECT 115.875 84.825 116.875 87.275 ;
        RECT 117.350 84.825 118.295 85.350 ;
        RECT 113.670 83.700 114.710 84.175 ;
        RECT 111.950 83.325 112.950 83.370 ;
        RECT 113.670 83.325 114.175 83.700 ;
        RECT 115.020 83.325 115.595 84.825 ;
        RECT 116.370 83.700 117.410 84.175 ;
        RECT 116.370 83.325 116.875 83.700 ;
        RECT 117.720 83.325 118.295 84.825 ;
        RECT 119.260 83.325 119.630 89.350 ;
        RECT 120.050 83.325 120.420 89.350 ;
        RECT 121.960 83.325 122.330 89.350 ;
        RECT 111.950 83.300 114.175 83.325 ;
        RECT 111.950 82.355 114.195 83.300 ;
        RECT 111.950 82.325 114.175 82.355 ;
        RECT 114.555 82.325 116.875 83.325 ;
        RECT 117.300 82.325 119.630 83.325 ;
        RECT 120.005 82.325 121.095 83.325 ;
        RECT 121.325 82.325 122.330 83.325 ;
        RECT 111.950 82.280 112.950 82.325 ;
        RECT 111.950 78.125 112.320 82.280 ;
        RECT 113.670 81.950 114.175 82.325 ;
        RECT 113.670 81.455 114.710 81.950 ;
        RECT 115.020 81.050 115.595 82.325 ;
        RECT 116.370 81.950 116.875 82.325 ;
        RECT 116.370 81.455 117.410 81.950 ;
        RECT 117.720 81.050 118.295 82.325 ;
        RECT 113.175 80.675 114.230 81.050 ;
        RECT 114.650 80.675 115.595 81.050 ;
        RECT 115.875 80.675 116.930 81.050 ;
        RECT 117.350 80.675 118.295 81.050 ;
        RECT 113.175 79.800 114.175 80.675 ;
        RECT 115.875 79.800 116.875 80.675 ;
        RECT 113.175 78.800 116.875 79.800 ;
        RECT 117.450 79.125 118.450 79.170 ;
        RECT 118.630 79.125 119.630 82.325 ;
        RECT 113.175 77.285 114.175 78.800 ;
        RECT 117.450 78.125 119.630 79.125 ;
        RECT 120.050 78.125 120.420 82.325 ;
        RECT 121.330 81.325 122.330 82.325 ;
        RECT 122.750 83.325 123.120 89.350 ;
        RECT 133.175 85.825 134.175 91.970 ;
        RECT 139.775 90.675 140.775 92.050 ;
        RECT 143.300 91.975 149.225 93.075 ;
        RECT 144.015 91.970 146.525 91.975 ;
        RECT 146.715 91.970 149.215 91.975 ;
        RECT 139.755 89.725 140.795 90.675 ;
        RECT 139.775 89.700 140.775 89.725 ;
        RECT 141.530 89.700 142.620 90.700 ;
        RECT 133.175 84.825 134.200 85.825 ;
        RECT 134.675 84.825 135.620 85.350 ;
        RECT 125.130 83.875 125.580 84.515 ;
        RECT 124.850 83.325 125.850 83.875 ;
        RECT 133.695 83.700 134.735 84.175 ;
        RECT 129.025 83.325 130.025 83.355 ;
        RECT 133.695 83.325 134.200 83.700 ;
        RECT 135.045 83.370 135.620 84.825 ;
        RECT 122.750 82.325 125.850 83.325 ;
        RECT 128.975 83.300 134.200 83.325 ;
        RECT 128.975 82.350 134.220 83.300 ;
        RECT 128.975 82.325 134.200 82.350 ;
        RECT 121.285 80.325 122.375 81.325 ;
        RECT 121.960 78.125 122.330 80.325 ;
        RECT 122.750 78.125 123.120 82.325 ;
        RECT 125.130 82.205 125.580 82.325 ;
        RECT 129.025 82.295 130.025 82.325 ;
        RECT 133.695 81.950 134.200 82.325 ;
        RECT 134.625 82.280 135.625 83.370 ;
        RECT 136.585 83.325 136.955 89.350 ;
        RECT 135.950 82.325 136.955 83.325 ;
        RECT 133.695 81.455 134.735 81.950 ;
        RECT 135.045 81.050 135.620 82.280 ;
        RECT 133.200 80.675 134.255 81.050 ;
        RECT 134.675 80.675 135.620 81.050 ;
        RECT 117.450 78.080 118.450 78.125 ;
        RECT 131.015 77.285 132.155 77.315 ;
        RECT 133.200 77.285 134.200 80.675 ;
        RECT 135.955 79.125 136.955 82.325 ;
        RECT 134.755 78.125 136.955 79.125 ;
        RECT 137.375 83.370 137.745 89.350 ;
        RECT 141.575 88.925 142.575 88.955 ;
        RECT 141.575 87.925 144.345 88.925 ;
        RECT 141.575 87.895 142.575 87.925 ;
        RECT 138.600 84.825 139.600 87.275 ;
        RECT 140.075 84.825 141.020 85.350 ;
        RECT 141.300 84.825 142.300 87.275 ;
        RECT 142.775 84.825 143.720 85.350 ;
        RECT 139.095 83.700 140.135 84.175 ;
        RECT 137.375 83.325 138.375 83.370 ;
        RECT 139.095 83.325 139.600 83.700 ;
        RECT 140.445 83.325 141.020 84.825 ;
        RECT 141.795 83.700 142.835 84.175 ;
        RECT 141.795 83.325 142.300 83.700 ;
        RECT 143.145 83.325 143.720 84.825 ;
        RECT 144.685 83.325 145.055 89.350 ;
        RECT 145.475 83.325 145.845 89.350 ;
        RECT 147.385 83.325 147.755 89.350 ;
        RECT 137.375 83.300 139.600 83.325 ;
        RECT 137.375 82.355 139.620 83.300 ;
        RECT 137.375 82.325 139.600 82.355 ;
        RECT 139.980 82.325 142.300 83.325 ;
        RECT 142.725 82.325 145.055 83.325 ;
        RECT 145.430 82.325 146.520 83.325 ;
        RECT 146.750 82.325 147.755 83.325 ;
        RECT 137.375 82.280 138.375 82.325 ;
        RECT 137.375 78.125 137.745 82.280 ;
        RECT 139.095 81.950 139.600 82.325 ;
        RECT 139.095 81.455 140.135 81.950 ;
        RECT 140.445 81.050 141.020 82.325 ;
        RECT 141.795 81.950 142.300 82.325 ;
        RECT 141.795 81.455 142.835 81.950 ;
        RECT 143.145 81.050 143.720 82.325 ;
        RECT 138.600 80.675 139.655 81.050 ;
        RECT 140.075 80.675 141.020 81.050 ;
        RECT 141.300 80.675 142.355 81.050 ;
        RECT 142.775 80.675 143.720 81.050 ;
        RECT 138.600 79.800 139.600 80.675 ;
        RECT 141.300 79.800 142.300 80.675 ;
        RECT 138.600 78.800 142.300 79.800 ;
        RECT 142.875 79.125 143.875 79.170 ;
        RECT 144.055 79.125 145.055 82.325 ;
        RECT 138.600 77.285 139.600 78.800 ;
        RECT 142.875 78.125 145.055 79.125 ;
        RECT 145.475 78.125 145.845 82.325 ;
        RECT 146.755 81.325 147.755 82.325 ;
        RECT 148.175 83.325 148.545 89.350 ;
        RECT 150.555 83.875 151.005 84.515 ;
        RECT 150.275 83.325 151.275 83.875 ;
        RECT 148.175 82.325 151.275 83.325 ;
        RECT 146.710 80.325 147.800 81.325 ;
        RECT 147.385 78.125 147.755 80.325 ;
        RECT 148.175 78.125 148.545 82.325 ;
        RECT 150.555 82.205 151.005 82.325 ;
        RECT 142.875 78.080 143.875 78.125 ;
        RECT 1.850 77.275 14.575 77.285 ;
        RECT 15.350 77.275 19.390 77.285 ;
        RECT 19.590 77.275 40.000 77.285 ;
        RECT 40.775 77.275 44.815 77.285 ;
        RECT 45.015 77.275 65.425 77.285 ;
        RECT 66.200 77.275 70.240 77.285 ;
        RECT 70.440 77.275 90.850 77.285 ;
        RECT 91.625 77.275 95.665 77.285 ;
        RECT 95.865 77.275 116.275 77.285 ;
        RECT 117.050 77.275 121.090 77.285 ;
        RECT 121.290 77.275 141.700 77.285 ;
        RECT 142.475 77.275 146.515 77.285 ;
        RECT 146.715 77.275 151.360 77.285 ;
        RECT 1.850 76.175 151.360 77.275 ;
        RECT 1.850 76.170 19.390 76.175 ;
        RECT 19.590 76.170 44.815 76.175 ;
        RECT 45.015 76.170 70.240 76.175 ;
        RECT 70.440 76.170 95.665 76.175 ;
        RECT 95.865 76.170 121.090 76.175 ;
        RECT 121.290 76.170 146.515 76.175 ;
        RECT 146.715 76.170 151.360 76.175 ;
        RECT 3.890 76.140 5.030 76.170 ;
        RECT 29.315 76.140 30.455 76.170 ;
        RECT 54.740 76.140 55.880 76.170 ;
        RECT 80.165 76.140 81.305 76.170 ;
        RECT 105.590 76.140 106.730 76.170 ;
        RECT 131.015 76.140 132.155 76.170 ;
        RECT 19.370 75.225 21.325 75.245 ;
        RECT 44.795 75.225 46.750 75.245 ;
        RECT 70.220 75.225 72.175 75.245 ;
        RECT 95.645 75.225 97.600 75.245 ;
        RECT 121.070 75.225 123.025 75.245 ;
        RECT 146.495 75.225 148.450 75.245 ;
        RECT 9.550 75.200 10.550 75.225 ;
        RECT 15.750 75.200 16.750 75.225 ;
        RECT 17.650 75.200 18.650 75.225 ;
        RECT 9.530 74.250 10.570 75.200 ;
        RECT 15.730 74.250 16.770 75.200 ;
        RECT 17.630 74.250 18.670 75.200 ;
        RECT 9.550 74.225 10.550 74.250 ;
        RECT 15.750 74.225 16.750 74.250 ;
        RECT 17.650 74.225 18.650 74.250 ;
        RECT 19.365 74.225 21.350 75.225 ;
        RECT 34.975 75.200 35.975 75.225 ;
        RECT 41.175 75.200 42.175 75.225 ;
        RECT 43.075 75.200 44.075 75.225 ;
        RECT 34.955 74.250 35.995 75.200 ;
        RECT 41.155 74.250 42.195 75.200 ;
        RECT 43.055 74.250 44.095 75.200 ;
        RECT 34.975 74.225 35.975 74.250 ;
        RECT 41.175 74.225 42.175 74.250 ;
        RECT 43.075 74.225 44.075 74.250 ;
        RECT 44.790 74.225 46.775 75.225 ;
        RECT 60.400 75.200 61.400 75.225 ;
        RECT 66.600 75.200 67.600 75.225 ;
        RECT 68.500 75.200 69.500 75.225 ;
        RECT 60.380 74.250 61.420 75.200 ;
        RECT 66.580 74.250 67.620 75.200 ;
        RECT 68.480 74.250 69.520 75.200 ;
        RECT 60.400 74.225 61.400 74.250 ;
        RECT 66.600 74.225 67.600 74.250 ;
        RECT 68.500 74.225 69.500 74.250 ;
        RECT 70.215 74.225 72.200 75.225 ;
        RECT 85.825 75.200 86.825 75.225 ;
        RECT 92.025 75.200 93.025 75.225 ;
        RECT 93.925 75.200 94.925 75.225 ;
        RECT 85.805 74.250 86.845 75.200 ;
        RECT 92.005 74.250 93.045 75.200 ;
        RECT 93.905 74.250 94.945 75.200 ;
        RECT 85.825 74.225 86.825 74.250 ;
        RECT 92.025 74.225 93.025 74.250 ;
        RECT 93.925 74.225 94.925 74.250 ;
        RECT 95.640 74.225 97.625 75.225 ;
        RECT 111.250 75.200 112.250 75.225 ;
        RECT 117.450 75.200 118.450 75.225 ;
        RECT 119.350 75.200 120.350 75.225 ;
        RECT 111.230 74.250 112.270 75.200 ;
        RECT 117.430 74.250 118.470 75.200 ;
        RECT 119.330 74.250 120.370 75.200 ;
        RECT 111.250 74.225 112.250 74.250 ;
        RECT 117.450 74.225 118.450 74.250 ;
        RECT 119.350 74.225 120.350 74.250 ;
        RECT 121.065 74.225 123.050 75.225 ;
        RECT 136.675 75.200 137.675 75.225 ;
        RECT 142.875 75.200 143.875 75.225 ;
        RECT 144.775 75.200 145.775 75.225 ;
        RECT 136.655 74.250 137.695 75.200 ;
        RECT 142.855 74.250 143.895 75.200 ;
        RECT 144.755 74.250 145.795 75.200 ;
        RECT 136.675 74.225 137.675 74.250 ;
        RECT 142.875 74.225 143.875 74.250 ;
        RECT 144.775 74.225 145.775 74.250 ;
        RECT 146.490 74.225 148.475 75.225 ;
        RECT 19.370 74.205 21.325 74.225 ;
        RECT 44.795 74.205 46.750 74.225 ;
        RECT 70.220 74.205 72.175 74.225 ;
        RECT 95.645 74.205 97.600 74.225 ;
        RECT 121.070 74.205 123.025 74.225 ;
        RECT 146.495 74.205 148.450 74.225 ;
        RECT 23.545 70.550 24.495 70.570 ;
        RECT 48.850 70.550 49.800 70.570 ;
        RECT 74.395 70.550 75.345 70.570 ;
        RECT 125.245 70.550 126.195 70.570 ;
        RECT 23.525 69.550 126.215 70.550 ;
        RECT 23.545 69.530 24.495 69.550 ;
        RECT 48.850 69.530 49.800 69.550 ;
        RECT 74.395 69.530 75.345 69.550 ;
        RECT 125.245 69.530 126.195 69.550 ;
        RECT 9.575 68.175 10.525 68.195 ;
        RECT 20.375 68.175 21.325 68.195 ;
        RECT 9.550 67.175 12.755 68.175 ;
        RECT 13.530 67.175 14.620 68.175 ;
        RECT 15.370 67.175 18.650 68.175 ;
        RECT 20.350 67.175 21.350 68.175 ;
        RECT 21.795 68.000 32.470 69.000 ;
        RECT 35.000 68.175 35.950 68.195 ;
        RECT 45.800 68.175 46.750 68.195 ;
        RECT 60.425 68.175 61.375 68.195 ;
        RECT 71.225 68.175 72.175 68.195 ;
        RECT 9.575 67.155 10.525 67.175 ;
        RECT 5.995 66.225 7.100 66.270 ;
        RECT 5.965 65.125 12.025 66.225 ;
        RECT 13.575 66.200 14.575 67.175 ;
        RECT 20.375 67.155 21.325 67.175 ;
        RECT 21.795 66.225 22.795 68.000 ;
        RECT 23.520 66.325 24.520 67.220 ;
        RECT 12.650 65.200 14.575 66.200 ;
        RECT 5.965 65.120 11.290 65.125 ;
        RECT 5.995 65.075 7.100 65.120 ;
        RECT 6.050 58.975 7.050 65.075 ;
        RECT 12.650 63.825 13.650 65.200 ;
        RECT 16.175 65.150 22.795 66.225 ;
        RECT 23.490 65.325 24.550 66.325 ;
        RECT 16.175 65.125 22.100 65.150 ;
        RECT 16.890 65.120 19.400 65.125 ;
        RECT 19.590 65.120 22.090 65.125 ;
        RECT 24.870 64.575 25.870 67.525 ;
        RECT 27.145 66.975 29.170 68.000 ;
        RECT 29.645 66.975 30.590 67.500 ;
        RECT 27.145 66.945 28.145 66.975 ;
        RECT 26.245 66.295 27.245 66.340 ;
        RECT 26.215 65.295 27.275 66.295 ;
        RECT 28.665 65.850 29.705 66.325 ;
        RECT 28.665 65.475 29.170 65.850 ;
        RECT 30.015 65.475 30.590 66.975 ;
        RECT 31.470 66.270 32.470 68.000 ;
        RECT 34.975 67.175 38.180 68.175 ;
        RECT 38.955 67.175 40.045 68.175 ;
        RECT 40.795 67.175 44.075 68.175 ;
        RECT 45.775 67.175 46.775 68.175 ;
        RECT 60.400 67.175 63.605 68.175 ;
        RECT 64.380 67.175 65.470 68.175 ;
        RECT 66.220 67.175 69.500 68.175 ;
        RECT 71.200 67.175 72.200 68.175 ;
        RECT 72.645 68.000 83.320 69.000 ;
        RECT 85.850 68.175 86.800 68.195 ;
        RECT 96.650 68.175 97.600 68.195 ;
        RECT 111.275 68.175 112.225 68.195 ;
        RECT 122.075 68.175 123.025 68.195 ;
        RECT 35.000 67.155 35.950 67.175 ;
        RECT 31.420 66.225 32.525 66.270 ;
        RECT 26.245 65.250 27.245 65.295 ;
        RECT 28.170 64.575 29.170 65.475 ;
        RECT 16.175 64.340 17.175 64.385 ;
        RECT 20.370 64.340 21.320 64.360 ;
        RECT 12.630 62.875 13.670 63.825 ;
        RECT 12.650 62.850 13.650 62.875 ;
        RECT 14.405 62.850 15.495 63.850 ;
        RECT 16.175 63.340 21.345 64.340 ;
        RECT 24.870 64.100 29.170 64.575 ;
        RECT 29.550 64.475 30.640 65.475 ;
        RECT 31.390 65.125 37.450 66.225 ;
        RECT 39.000 66.200 40.000 67.175 ;
        RECT 45.800 67.155 46.750 67.175 ;
        RECT 60.425 67.155 61.375 67.175 ;
        RECT 56.845 66.225 57.950 66.270 ;
        RECT 38.075 65.200 40.000 66.200 ;
        RECT 31.390 65.120 36.715 65.125 ;
        RECT 31.420 65.075 32.525 65.120 ;
        RECT 24.870 63.650 29.705 64.100 ;
        RECT 23.020 63.605 29.705 63.650 ;
        RECT 23.020 63.575 29.170 63.605 ;
        RECT 16.175 63.295 17.175 63.340 ;
        RECT 20.370 63.320 21.320 63.340 ;
        RECT 23.020 62.650 25.870 63.575 ;
        RECT 27.145 63.200 28.145 63.230 ;
        RECT 30.015 63.200 30.590 64.475 ;
        RECT 27.145 62.825 29.225 63.200 ;
        RECT 29.645 62.825 30.590 63.200 ;
        RECT 6.050 57.975 7.075 58.975 ;
        RECT 7.550 57.975 8.495 58.500 ;
        RECT 6.570 56.850 7.610 57.325 ;
        RECT 3.950 56.500 4.950 56.505 ;
        RECT 3.920 56.475 4.980 56.500 ;
        RECT 6.570 56.475 7.075 56.850 ;
        RECT 7.920 56.520 8.495 57.975 ;
        RECT 3.875 56.450 7.075 56.475 ;
        RECT 3.875 55.500 7.095 56.450 ;
        RECT 3.875 55.475 7.075 55.500 ;
        RECT 3.950 55.445 4.950 55.475 ;
        RECT 6.570 55.100 7.075 55.475 ;
        RECT 7.500 55.430 8.500 56.520 ;
        RECT 9.460 56.475 9.830 62.500 ;
        RECT 8.825 55.475 9.830 56.475 ;
        RECT 6.570 54.605 7.610 55.100 ;
        RECT 7.920 54.200 8.495 55.430 ;
        RECT 6.075 53.825 7.130 54.200 ;
        RECT 7.550 53.825 8.495 54.200 ;
        RECT 3.905 50.455 5.020 50.460 ;
        RECT 3.875 50.435 5.050 50.455 ;
        RECT 6.075 50.435 7.075 53.825 ;
        RECT 8.830 52.275 9.830 55.475 ;
        RECT 7.630 51.275 9.830 52.275 ;
        RECT 10.250 56.520 10.620 62.500 ;
        RECT 14.450 62.075 15.450 62.105 ;
        RECT 14.450 61.075 17.220 62.075 ;
        RECT 14.450 61.045 15.450 61.075 ;
        RECT 11.475 57.975 12.475 60.425 ;
        RECT 12.950 57.975 13.895 58.500 ;
        RECT 14.175 57.975 15.175 60.425 ;
        RECT 15.650 57.975 16.595 58.500 ;
        RECT 11.970 56.850 13.010 57.325 ;
        RECT 10.250 56.475 11.250 56.520 ;
        RECT 11.970 56.475 12.475 56.850 ;
        RECT 13.320 56.475 13.895 57.975 ;
        RECT 14.670 56.850 15.710 57.325 ;
        RECT 14.670 56.475 15.175 56.850 ;
        RECT 16.020 56.475 16.595 57.975 ;
        RECT 17.560 56.475 17.930 62.500 ;
        RECT 18.350 56.475 18.720 62.500 ;
        RECT 20.260 56.475 20.630 62.500 ;
        RECT 10.250 56.450 12.475 56.475 ;
        RECT 10.250 55.505 12.495 56.450 ;
        RECT 10.250 55.475 12.475 55.505 ;
        RECT 12.855 55.475 15.175 56.475 ;
        RECT 15.600 55.475 17.930 56.475 ;
        RECT 18.305 55.475 19.395 56.475 ;
        RECT 10.250 55.430 11.250 55.475 ;
        RECT 10.250 51.275 10.620 55.430 ;
        RECT 11.970 55.100 12.475 55.475 ;
        RECT 11.970 54.605 13.010 55.100 ;
        RECT 13.320 54.200 13.895 55.475 ;
        RECT 14.670 55.100 15.175 55.475 ;
        RECT 14.670 54.605 15.710 55.100 ;
        RECT 16.020 54.200 16.595 55.475 ;
        RECT 11.475 53.825 12.530 54.200 ;
        RECT 12.950 53.825 13.895 54.200 ;
        RECT 14.175 53.825 15.230 54.200 ;
        RECT 15.650 53.825 16.595 54.200 ;
        RECT 11.475 52.950 12.475 53.825 ;
        RECT 14.175 52.950 15.175 53.825 ;
        RECT 11.475 51.950 15.175 52.950 ;
        RECT 15.750 52.275 16.750 52.320 ;
        RECT 16.930 52.275 17.930 55.475 ;
        RECT 11.475 50.435 12.475 51.950 ;
        RECT 15.750 51.275 17.930 52.275 ;
        RECT 18.350 51.275 18.720 55.475 ;
        RECT 19.625 53.975 20.630 56.475 ;
        RECT 21.050 56.475 21.420 62.500 ;
        RECT 27.145 62.200 29.170 62.825 ;
        RECT 27.145 62.170 28.370 62.200 ;
        RECT 24.820 61.155 25.925 61.200 ;
        RECT 24.775 60.050 25.970 61.155 ;
        RECT 24.790 60.045 25.955 60.050 ;
        RECT 23.425 56.475 24.375 56.500 ;
        RECT 21.050 55.475 26.300 56.475 ;
        RECT 19.605 53.025 20.645 53.975 ;
        RECT 19.625 53.000 20.630 53.025 ;
        RECT 20.260 51.275 20.630 53.000 ;
        RECT 21.050 51.275 21.420 55.475 ;
        RECT 23.425 55.460 24.375 55.475 ;
        RECT 15.750 51.230 16.750 51.275 ;
        RECT 27.370 50.435 28.370 62.170 ;
        RECT 31.475 58.975 32.475 65.075 ;
        RECT 38.075 63.825 39.075 65.200 ;
        RECT 41.600 65.125 62.875 66.225 ;
        RECT 64.425 66.200 65.425 67.175 ;
        RECT 71.225 67.155 72.175 67.175 ;
        RECT 72.645 66.225 73.645 68.000 ;
        RECT 74.370 66.325 75.370 67.220 ;
        RECT 63.500 65.200 65.425 66.200 ;
        RECT 42.315 65.120 44.825 65.125 ;
        RECT 45.015 65.120 62.140 65.125 ;
        RECT 56.845 65.075 57.950 65.120 ;
        RECT 38.055 62.875 39.095 63.825 ;
        RECT 38.075 62.850 39.075 62.875 ;
        RECT 39.830 62.850 40.920 63.850 ;
        RECT 31.475 57.975 32.500 58.975 ;
        RECT 32.975 57.975 33.920 58.500 ;
        RECT 31.995 56.850 33.035 57.325 ;
        RECT 29.375 56.500 30.375 56.505 ;
        RECT 29.345 56.475 30.405 56.500 ;
        RECT 31.995 56.475 32.500 56.850 ;
        RECT 33.345 56.520 33.920 57.975 ;
        RECT 29.300 56.450 32.500 56.475 ;
        RECT 29.300 55.500 32.520 56.450 ;
        RECT 29.300 55.475 32.500 55.500 ;
        RECT 29.375 55.445 30.375 55.475 ;
        RECT 31.995 55.100 32.500 55.475 ;
        RECT 32.925 55.430 33.925 56.520 ;
        RECT 34.885 56.475 35.255 62.500 ;
        RECT 34.250 55.475 35.255 56.475 ;
        RECT 31.995 54.605 33.035 55.100 ;
        RECT 33.345 54.200 33.920 55.430 ;
        RECT 31.500 53.825 32.555 54.200 ;
        RECT 32.975 53.825 33.920 54.200 ;
        RECT 29.330 50.455 30.445 50.460 ;
        RECT 29.300 50.435 30.475 50.455 ;
        RECT 31.500 50.435 32.500 53.825 ;
        RECT 34.255 52.275 35.255 55.475 ;
        RECT 33.055 51.275 35.255 52.275 ;
        RECT 35.675 56.520 36.045 62.500 ;
        RECT 39.875 62.075 40.875 62.105 ;
        RECT 39.875 61.075 42.645 62.075 ;
        RECT 39.875 61.045 40.875 61.075 ;
        RECT 36.900 57.975 37.900 60.425 ;
        RECT 38.375 57.975 39.320 58.500 ;
        RECT 39.600 57.975 40.600 60.425 ;
        RECT 41.075 57.975 42.020 58.500 ;
        RECT 37.395 56.850 38.435 57.325 ;
        RECT 35.675 56.475 36.675 56.520 ;
        RECT 37.395 56.475 37.900 56.850 ;
        RECT 38.745 56.475 39.320 57.975 ;
        RECT 40.095 56.850 41.135 57.325 ;
        RECT 40.095 56.475 40.600 56.850 ;
        RECT 41.445 56.475 42.020 57.975 ;
        RECT 42.985 56.475 43.355 62.500 ;
        RECT 43.775 56.475 44.145 62.500 ;
        RECT 45.685 56.475 46.055 62.500 ;
        RECT 35.675 56.450 37.900 56.475 ;
        RECT 35.675 55.505 37.920 56.450 ;
        RECT 35.675 55.475 37.900 55.505 ;
        RECT 38.280 55.475 40.600 56.475 ;
        RECT 41.025 55.475 43.355 56.475 ;
        RECT 43.730 55.475 44.820 56.475 ;
        RECT 35.675 55.430 36.675 55.475 ;
        RECT 35.675 51.275 36.045 55.430 ;
        RECT 37.395 55.100 37.900 55.475 ;
        RECT 37.395 54.605 38.435 55.100 ;
        RECT 38.745 54.200 39.320 55.475 ;
        RECT 40.095 55.100 40.600 55.475 ;
        RECT 40.095 54.605 41.135 55.100 ;
        RECT 41.445 54.200 42.020 55.475 ;
        RECT 36.900 53.825 37.955 54.200 ;
        RECT 38.375 53.825 39.320 54.200 ;
        RECT 39.600 53.825 40.655 54.200 ;
        RECT 41.075 53.825 42.020 54.200 ;
        RECT 36.900 52.950 37.900 53.825 ;
        RECT 39.600 52.950 40.600 53.825 ;
        RECT 36.900 51.950 40.600 52.950 ;
        RECT 41.175 52.275 42.175 52.320 ;
        RECT 42.355 52.275 43.355 55.475 ;
        RECT 36.900 50.435 37.900 51.950 ;
        RECT 41.175 51.275 43.355 52.275 ;
        RECT 43.775 51.275 44.145 55.475 ;
        RECT 45.050 53.975 46.055 56.475 ;
        RECT 46.475 56.475 46.845 62.500 ;
        RECT 56.900 58.975 57.900 65.075 ;
        RECT 63.500 63.825 64.500 65.200 ;
        RECT 67.025 65.150 73.645 66.225 ;
        RECT 74.340 65.325 75.400 66.325 ;
        RECT 67.025 65.125 72.950 65.150 ;
        RECT 67.740 65.120 70.250 65.125 ;
        RECT 70.440 65.120 72.940 65.125 ;
        RECT 75.720 64.575 76.720 67.525 ;
        RECT 77.995 66.975 80.020 68.000 ;
        RECT 80.495 66.975 81.440 67.500 ;
        RECT 77.995 66.945 78.995 66.975 ;
        RECT 77.095 66.295 78.095 66.340 ;
        RECT 77.065 65.295 78.125 66.295 ;
        RECT 79.515 65.850 80.555 66.325 ;
        RECT 79.515 65.475 80.020 65.850 ;
        RECT 80.865 65.475 81.440 66.975 ;
        RECT 82.320 66.270 83.320 68.000 ;
        RECT 85.825 67.175 89.030 68.175 ;
        RECT 89.805 67.175 90.895 68.175 ;
        RECT 91.645 67.175 94.925 68.175 ;
        RECT 96.625 67.175 97.625 68.175 ;
        RECT 111.250 67.175 114.455 68.175 ;
        RECT 115.230 67.175 116.320 68.175 ;
        RECT 117.070 67.175 120.350 68.175 ;
        RECT 122.050 67.175 123.050 68.175 ;
        RECT 123.495 68.000 134.170 69.000 ;
        RECT 136.700 68.175 137.650 68.195 ;
        RECT 147.500 68.175 148.450 68.195 ;
        RECT 85.850 67.155 86.800 67.175 ;
        RECT 82.270 66.225 83.375 66.270 ;
        RECT 77.095 65.250 78.095 65.295 ;
        RECT 79.020 64.575 80.020 65.475 ;
        RECT 67.025 64.340 68.025 64.385 ;
        RECT 71.220 64.340 72.170 64.360 ;
        RECT 63.480 62.875 64.520 63.825 ;
        RECT 63.500 62.850 64.500 62.875 ;
        RECT 65.255 62.850 66.345 63.850 ;
        RECT 67.025 63.340 72.195 64.340 ;
        RECT 75.720 64.100 80.020 64.575 ;
        RECT 80.400 64.475 81.490 65.475 ;
        RECT 82.240 65.125 88.300 66.225 ;
        RECT 89.850 66.200 90.850 67.175 ;
        RECT 96.650 67.155 97.600 67.175 ;
        RECT 111.275 67.155 112.225 67.175 ;
        RECT 107.695 66.225 108.800 66.270 ;
        RECT 88.925 65.200 90.850 66.200 ;
        RECT 82.240 65.120 87.565 65.125 ;
        RECT 82.270 65.075 83.375 65.120 ;
        RECT 75.720 63.650 80.555 64.100 ;
        RECT 73.870 63.605 80.555 63.650 ;
        RECT 73.870 63.575 80.020 63.605 ;
        RECT 67.025 63.295 68.025 63.340 ;
        RECT 71.220 63.320 72.170 63.340 ;
        RECT 73.870 62.650 76.720 63.575 ;
        RECT 77.995 63.200 78.995 63.230 ;
        RECT 80.865 63.200 81.440 64.475 ;
        RECT 77.995 62.825 80.075 63.200 ;
        RECT 80.495 62.825 81.440 63.200 ;
        RECT 56.900 57.975 57.925 58.975 ;
        RECT 58.400 57.975 59.345 58.500 ;
        RECT 57.420 56.850 58.460 57.325 ;
        RECT 50.725 56.475 51.725 56.505 ;
        RECT 54.800 56.500 55.800 56.505 ;
        RECT 54.770 56.475 55.830 56.500 ;
        RECT 57.420 56.475 57.925 56.850 ;
        RECT 58.770 56.520 59.345 57.975 ;
        RECT 46.475 55.475 51.725 56.475 ;
        RECT 54.725 56.450 57.925 56.475 ;
        RECT 54.725 55.500 57.945 56.450 ;
        RECT 54.725 55.475 57.925 55.500 ;
        RECT 45.030 53.025 46.070 53.975 ;
        RECT 45.050 53.000 46.055 53.025 ;
        RECT 45.685 51.275 46.055 53.000 ;
        RECT 46.475 51.275 46.845 55.475 ;
        RECT 50.725 55.445 51.725 55.475 ;
        RECT 54.800 55.445 55.800 55.475 ;
        RECT 57.420 55.100 57.925 55.475 ;
        RECT 58.350 55.430 59.350 56.520 ;
        RECT 60.310 56.475 60.680 62.500 ;
        RECT 59.675 55.475 60.680 56.475 ;
        RECT 57.420 54.605 58.460 55.100 ;
        RECT 58.770 54.200 59.345 55.430 ;
        RECT 56.925 53.825 57.980 54.200 ;
        RECT 58.400 53.825 59.345 54.200 ;
        RECT 41.175 51.230 42.175 51.275 ;
        RECT 54.755 50.455 55.870 50.460 ;
        RECT 54.725 50.435 55.900 50.455 ;
        RECT 56.925 50.435 57.925 53.825 ;
        RECT 59.680 52.275 60.680 55.475 ;
        RECT 58.480 51.275 60.680 52.275 ;
        RECT 61.100 56.520 61.470 62.500 ;
        RECT 65.300 62.075 66.300 62.105 ;
        RECT 65.300 61.075 68.070 62.075 ;
        RECT 65.300 61.045 66.300 61.075 ;
        RECT 62.325 57.975 63.325 60.425 ;
        RECT 63.800 57.975 64.745 58.500 ;
        RECT 65.025 57.975 66.025 60.425 ;
        RECT 66.500 57.975 67.445 58.500 ;
        RECT 62.820 56.850 63.860 57.325 ;
        RECT 61.100 56.475 62.100 56.520 ;
        RECT 62.820 56.475 63.325 56.850 ;
        RECT 64.170 56.475 64.745 57.975 ;
        RECT 65.520 56.850 66.560 57.325 ;
        RECT 65.520 56.475 66.025 56.850 ;
        RECT 66.870 56.475 67.445 57.975 ;
        RECT 68.410 56.475 68.780 62.500 ;
        RECT 69.200 56.475 69.570 62.500 ;
        RECT 71.110 56.475 71.480 62.500 ;
        RECT 61.100 56.450 63.325 56.475 ;
        RECT 61.100 55.505 63.345 56.450 ;
        RECT 61.100 55.475 63.325 55.505 ;
        RECT 63.705 55.475 66.025 56.475 ;
        RECT 66.450 55.475 68.780 56.475 ;
        RECT 69.155 55.475 70.245 56.475 ;
        RECT 61.100 55.430 62.100 55.475 ;
        RECT 61.100 51.275 61.470 55.430 ;
        RECT 62.820 55.100 63.325 55.475 ;
        RECT 62.820 54.605 63.860 55.100 ;
        RECT 64.170 54.200 64.745 55.475 ;
        RECT 65.520 55.100 66.025 55.475 ;
        RECT 65.520 54.605 66.560 55.100 ;
        RECT 66.870 54.200 67.445 55.475 ;
        RECT 62.325 53.825 63.380 54.200 ;
        RECT 63.800 53.825 64.745 54.200 ;
        RECT 65.025 53.825 66.080 54.200 ;
        RECT 66.500 53.825 67.445 54.200 ;
        RECT 62.325 52.950 63.325 53.825 ;
        RECT 65.025 52.950 66.025 53.825 ;
        RECT 62.325 51.950 66.025 52.950 ;
        RECT 66.600 52.275 67.600 52.320 ;
        RECT 67.780 52.275 68.780 55.475 ;
        RECT 62.325 50.435 63.325 51.950 ;
        RECT 66.600 51.275 68.780 52.275 ;
        RECT 69.200 51.275 69.570 55.475 ;
        RECT 70.475 53.975 71.480 56.475 ;
        RECT 71.900 56.475 72.270 62.500 ;
        RECT 77.995 62.200 80.020 62.825 ;
        RECT 77.995 62.170 79.220 62.200 ;
        RECT 75.670 61.155 76.775 61.200 ;
        RECT 75.625 60.050 76.820 61.155 ;
        RECT 75.640 60.045 76.805 60.050 ;
        RECT 74.275 56.475 75.225 56.500 ;
        RECT 71.900 55.475 77.150 56.475 ;
        RECT 70.455 53.025 71.495 53.975 ;
        RECT 70.475 53.000 71.480 53.025 ;
        RECT 71.110 51.275 71.480 53.000 ;
        RECT 71.900 51.275 72.270 55.475 ;
        RECT 74.275 55.460 75.225 55.475 ;
        RECT 66.600 51.230 67.600 51.275 ;
        RECT 78.220 50.435 79.220 62.170 ;
        RECT 82.325 58.975 83.325 65.075 ;
        RECT 88.925 63.825 89.925 65.200 ;
        RECT 92.450 65.125 113.725 66.225 ;
        RECT 115.275 66.200 116.275 67.175 ;
        RECT 122.075 67.155 123.025 67.175 ;
        RECT 123.495 66.225 124.495 68.000 ;
        RECT 125.220 66.325 126.220 67.220 ;
        RECT 114.350 65.200 116.275 66.200 ;
        RECT 93.165 65.120 95.675 65.125 ;
        RECT 95.865 65.120 112.990 65.125 ;
        RECT 107.695 65.075 108.800 65.120 ;
        RECT 88.905 62.875 89.945 63.825 ;
        RECT 88.925 62.850 89.925 62.875 ;
        RECT 90.680 62.850 91.770 63.850 ;
        RECT 82.325 57.975 83.350 58.975 ;
        RECT 83.825 57.975 84.770 58.500 ;
        RECT 82.845 56.850 83.885 57.325 ;
        RECT 80.225 56.500 81.225 56.505 ;
        RECT 80.195 56.475 81.255 56.500 ;
        RECT 82.845 56.475 83.350 56.850 ;
        RECT 84.195 56.520 84.770 57.975 ;
        RECT 80.150 56.450 83.350 56.475 ;
        RECT 80.150 55.500 83.370 56.450 ;
        RECT 80.150 55.475 83.350 55.500 ;
        RECT 80.225 55.445 81.225 55.475 ;
        RECT 82.845 55.100 83.350 55.475 ;
        RECT 83.775 55.430 84.775 56.520 ;
        RECT 85.735 56.475 86.105 62.500 ;
        RECT 85.100 55.475 86.105 56.475 ;
        RECT 82.845 54.605 83.885 55.100 ;
        RECT 84.195 54.200 84.770 55.430 ;
        RECT 82.350 53.825 83.405 54.200 ;
        RECT 83.825 53.825 84.770 54.200 ;
        RECT 80.180 50.455 81.295 50.460 ;
        RECT 80.150 50.435 81.325 50.455 ;
        RECT 82.350 50.435 83.350 53.825 ;
        RECT 85.105 52.275 86.105 55.475 ;
        RECT 83.905 51.275 86.105 52.275 ;
        RECT 86.525 56.520 86.895 62.500 ;
        RECT 90.725 62.075 91.725 62.105 ;
        RECT 90.725 61.075 93.495 62.075 ;
        RECT 90.725 61.045 91.725 61.075 ;
        RECT 87.750 57.975 88.750 60.425 ;
        RECT 89.225 57.975 90.170 58.500 ;
        RECT 90.450 57.975 91.450 60.425 ;
        RECT 91.925 57.975 92.870 58.500 ;
        RECT 88.245 56.850 89.285 57.325 ;
        RECT 86.525 56.475 87.525 56.520 ;
        RECT 88.245 56.475 88.750 56.850 ;
        RECT 89.595 56.475 90.170 57.975 ;
        RECT 90.945 56.850 91.985 57.325 ;
        RECT 90.945 56.475 91.450 56.850 ;
        RECT 92.295 56.475 92.870 57.975 ;
        RECT 93.835 56.475 94.205 62.500 ;
        RECT 94.625 56.475 94.995 62.500 ;
        RECT 96.535 56.475 96.905 62.500 ;
        RECT 86.525 56.450 88.750 56.475 ;
        RECT 86.525 55.505 88.770 56.450 ;
        RECT 86.525 55.475 88.750 55.505 ;
        RECT 89.130 55.475 91.450 56.475 ;
        RECT 91.875 55.475 94.205 56.475 ;
        RECT 94.580 55.475 95.670 56.475 ;
        RECT 86.525 55.430 87.525 55.475 ;
        RECT 86.525 51.275 86.895 55.430 ;
        RECT 88.245 55.100 88.750 55.475 ;
        RECT 88.245 54.605 89.285 55.100 ;
        RECT 89.595 54.200 90.170 55.475 ;
        RECT 90.945 55.100 91.450 55.475 ;
        RECT 90.945 54.605 91.985 55.100 ;
        RECT 92.295 54.200 92.870 55.475 ;
        RECT 87.750 53.825 88.805 54.200 ;
        RECT 89.225 53.825 90.170 54.200 ;
        RECT 90.450 53.825 91.505 54.200 ;
        RECT 91.925 53.825 92.870 54.200 ;
        RECT 87.750 52.950 88.750 53.825 ;
        RECT 90.450 52.950 91.450 53.825 ;
        RECT 87.750 51.950 91.450 52.950 ;
        RECT 92.025 52.275 93.025 52.320 ;
        RECT 93.205 52.275 94.205 55.475 ;
        RECT 87.750 50.435 88.750 51.950 ;
        RECT 92.025 51.275 94.205 52.275 ;
        RECT 94.625 51.275 94.995 55.475 ;
        RECT 95.900 53.975 96.905 56.475 ;
        RECT 97.325 56.475 97.695 62.500 ;
        RECT 107.750 58.975 108.750 65.075 ;
        RECT 114.350 63.825 115.350 65.200 ;
        RECT 117.875 65.150 124.495 66.225 ;
        RECT 125.190 65.325 126.250 66.325 ;
        RECT 117.875 65.125 123.800 65.150 ;
        RECT 118.590 65.120 121.100 65.125 ;
        RECT 121.290 65.120 123.790 65.125 ;
        RECT 126.570 64.575 127.570 67.525 ;
        RECT 128.845 66.975 130.870 68.000 ;
        RECT 131.345 66.975 132.290 67.500 ;
        RECT 128.845 66.945 129.845 66.975 ;
        RECT 127.945 66.295 128.945 66.340 ;
        RECT 127.915 65.295 128.975 66.295 ;
        RECT 130.365 65.850 131.405 66.325 ;
        RECT 130.365 65.475 130.870 65.850 ;
        RECT 131.715 65.475 132.290 66.975 ;
        RECT 133.170 66.270 134.170 68.000 ;
        RECT 136.675 67.175 139.880 68.175 ;
        RECT 140.655 67.175 141.745 68.175 ;
        RECT 142.495 67.175 145.775 68.175 ;
        RECT 147.475 67.175 148.475 68.175 ;
        RECT 136.700 67.155 137.650 67.175 ;
        RECT 133.120 66.225 134.225 66.270 ;
        RECT 127.945 65.250 128.945 65.295 ;
        RECT 129.870 64.575 130.870 65.475 ;
        RECT 117.875 64.340 118.875 64.385 ;
        RECT 122.070 64.340 123.020 64.360 ;
        RECT 114.330 62.875 115.370 63.825 ;
        RECT 114.350 62.850 115.350 62.875 ;
        RECT 116.105 62.850 117.195 63.850 ;
        RECT 117.875 63.340 123.045 64.340 ;
        RECT 126.570 64.100 130.870 64.575 ;
        RECT 131.250 64.475 132.340 65.475 ;
        RECT 133.090 65.125 139.150 66.225 ;
        RECT 140.700 66.200 141.700 67.175 ;
        RECT 147.500 67.155 148.450 67.175 ;
        RECT 139.775 65.200 141.700 66.200 ;
        RECT 133.090 65.120 138.415 65.125 ;
        RECT 133.120 65.075 134.225 65.120 ;
        RECT 126.570 63.650 131.405 64.100 ;
        RECT 124.720 63.605 131.405 63.650 ;
        RECT 124.720 63.575 130.870 63.605 ;
        RECT 117.875 63.295 118.875 63.340 ;
        RECT 122.070 63.320 123.020 63.340 ;
        RECT 124.720 62.650 127.570 63.575 ;
        RECT 128.845 63.200 129.845 63.230 ;
        RECT 131.715 63.200 132.290 64.475 ;
        RECT 128.845 62.825 130.925 63.200 ;
        RECT 131.345 62.825 132.290 63.200 ;
        RECT 107.750 57.975 108.775 58.975 ;
        RECT 109.250 57.975 110.195 58.500 ;
        RECT 108.270 56.850 109.310 57.325 ;
        RECT 101.575 56.475 102.575 56.505 ;
        RECT 105.650 56.500 106.650 56.505 ;
        RECT 105.620 56.475 106.680 56.500 ;
        RECT 108.270 56.475 108.775 56.850 ;
        RECT 109.620 56.520 110.195 57.975 ;
        RECT 97.325 55.475 102.575 56.475 ;
        RECT 105.575 56.450 108.775 56.475 ;
        RECT 105.575 55.500 108.795 56.450 ;
        RECT 105.575 55.475 108.775 55.500 ;
        RECT 95.880 53.025 96.920 53.975 ;
        RECT 95.900 53.000 96.905 53.025 ;
        RECT 96.535 51.275 96.905 53.000 ;
        RECT 97.325 51.275 97.695 55.475 ;
        RECT 101.575 55.445 102.575 55.475 ;
        RECT 105.650 55.445 106.650 55.475 ;
        RECT 108.270 55.100 108.775 55.475 ;
        RECT 109.200 55.430 110.200 56.520 ;
        RECT 111.160 56.475 111.530 62.500 ;
        RECT 110.525 55.475 111.530 56.475 ;
        RECT 108.270 54.605 109.310 55.100 ;
        RECT 109.620 54.200 110.195 55.430 ;
        RECT 107.775 53.825 108.830 54.200 ;
        RECT 109.250 53.825 110.195 54.200 ;
        RECT 92.025 51.230 93.025 51.275 ;
        RECT 105.605 50.455 106.720 50.460 ;
        RECT 105.575 50.435 106.750 50.455 ;
        RECT 107.775 50.435 108.775 53.825 ;
        RECT 110.530 52.275 111.530 55.475 ;
        RECT 109.330 51.275 111.530 52.275 ;
        RECT 111.950 56.520 112.320 62.500 ;
        RECT 116.150 62.075 117.150 62.105 ;
        RECT 116.150 61.075 118.920 62.075 ;
        RECT 116.150 61.045 117.150 61.075 ;
        RECT 113.175 57.975 114.175 60.425 ;
        RECT 114.650 57.975 115.595 58.500 ;
        RECT 115.875 57.975 116.875 60.425 ;
        RECT 117.350 57.975 118.295 58.500 ;
        RECT 113.670 56.850 114.710 57.325 ;
        RECT 111.950 56.475 112.950 56.520 ;
        RECT 113.670 56.475 114.175 56.850 ;
        RECT 115.020 56.475 115.595 57.975 ;
        RECT 116.370 56.850 117.410 57.325 ;
        RECT 116.370 56.475 116.875 56.850 ;
        RECT 117.720 56.475 118.295 57.975 ;
        RECT 119.260 56.475 119.630 62.500 ;
        RECT 120.050 56.475 120.420 62.500 ;
        RECT 121.960 56.475 122.330 62.500 ;
        RECT 111.950 56.450 114.175 56.475 ;
        RECT 111.950 55.505 114.195 56.450 ;
        RECT 111.950 55.475 114.175 55.505 ;
        RECT 114.555 55.475 116.875 56.475 ;
        RECT 117.300 55.475 119.630 56.475 ;
        RECT 120.005 55.475 121.095 56.475 ;
        RECT 111.950 55.430 112.950 55.475 ;
        RECT 111.950 51.275 112.320 55.430 ;
        RECT 113.670 55.100 114.175 55.475 ;
        RECT 113.670 54.605 114.710 55.100 ;
        RECT 115.020 54.200 115.595 55.475 ;
        RECT 116.370 55.100 116.875 55.475 ;
        RECT 116.370 54.605 117.410 55.100 ;
        RECT 117.720 54.200 118.295 55.475 ;
        RECT 113.175 53.825 114.230 54.200 ;
        RECT 114.650 53.825 115.595 54.200 ;
        RECT 115.875 53.825 116.930 54.200 ;
        RECT 117.350 53.825 118.295 54.200 ;
        RECT 113.175 52.950 114.175 53.825 ;
        RECT 115.875 52.950 116.875 53.825 ;
        RECT 113.175 51.950 116.875 52.950 ;
        RECT 117.450 52.275 118.450 52.320 ;
        RECT 118.630 52.275 119.630 55.475 ;
        RECT 113.175 50.435 114.175 51.950 ;
        RECT 117.450 51.275 119.630 52.275 ;
        RECT 120.050 51.275 120.420 55.475 ;
        RECT 121.325 53.975 122.330 56.475 ;
        RECT 122.750 56.475 123.120 62.500 ;
        RECT 128.845 62.200 130.870 62.825 ;
        RECT 128.845 62.170 130.070 62.200 ;
        RECT 126.520 61.155 127.625 61.200 ;
        RECT 126.475 60.050 127.670 61.155 ;
        RECT 126.490 60.045 127.655 60.050 ;
        RECT 125.125 56.475 126.075 56.500 ;
        RECT 122.750 55.475 128.000 56.475 ;
        RECT 121.305 53.025 122.345 53.975 ;
        RECT 121.325 53.000 122.330 53.025 ;
        RECT 121.960 51.275 122.330 53.000 ;
        RECT 122.750 51.275 123.120 55.475 ;
        RECT 125.125 55.460 126.075 55.475 ;
        RECT 117.450 51.230 118.450 51.275 ;
        RECT 129.070 50.435 130.070 62.170 ;
        RECT 133.175 58.975 134.175 65.075 ;
        RECT 139.775 63.825 140.775 65.200 ;
        RECT 143.300 65.125 149.225 66.225 ;
        RECT 144.015 65.120 146.525 65.125 ;
        RECT 146.715 65.120 149.215 65.125 ;
        RECT 139.755 62.875 140.795 63.825 ;
        RECT 139.775 62.850 140.775 62.875 ;
        RECT 141.530 62.850 142.620 63.850 ;
        RECT 133.175 57.975 134.200 58.975 ;
        RECT 134.675 57.975 135.620 58.500 ;
        RECT 133.695 56.850 134.735 57.325 ;
        RECT 131.075 56.500 132.075 56.505 ;
        RECT 131.045 56.475 132.105 56.500 ;
        RECT 133.695 56.475 134.200 56.850 ;
        RECT 135.045 56.520 135.620 57.975 ;
        RECT 131.000 56.450 134.200 56.475 ;
        RECT 131.000 55.500 134.220 56.450 ;
        RECT 131.000 55.475 134.200 55.500 ;
        RECT 131.075 55.445 132.075 55.475 ;
        RECT 133.695 55.100 134.200 55.475 ;
        RECT 134.625 55.430 135.625 56.520 ;
        RECT 136.585 56.475 136.955 62.500 ;
        RECT 135.950 55.475 136.955 56.475 ;
        RECT 133.695 54.605 134.735 55.100 ;
        RECT 135.045 54.200 135.620 55.430 ;
        RECT 133.200 53.825 134.255 54.200 ;
        RECT 134.675 53.825 135.620 54.200 ;
        RECT 131.030 50.455 132.145 50.460 ;
        RECT 131.000 50.435 132.175 50.455 ;
        RECT 133.200 50.435 134.200 53.825 ;
        RECT 135.955 52.275 136.955 55.475 ;
        RECT 134.755 51.275 136.955 52.275 ;
        RECT 137.375 56.520 137.745 62.500 ;
        RECT 141.575 62.075 142.575 62.105 ;
        RECT 141.575 61.075 144.345 62.075 ;
        RECT 141.575 61.045 142.575 61.075 ;
        RECT 138.600 57.975 139.600 60.425 ;
        RECT 140.075 57.975 141.020 58.500 ;
        RECT 141.300 57.975 142.300 60.425 ;
        RECT 142.775 57.975 143.720 58.500 ;
        RECT 139.095 56.850 140.135 57.325 ;
        RECT 137.375 56.475 138.375 56.520 ;
        RECT 139.095 56.475 139.600 56.850 ;
        RECT 140.445 56.475 141.020 57.975 ;
        RECT 141.795 56.850 142.835 57.325 ;
        RECT 141.795 56.475 142.300 56.850 ;
        RECT 143.145 56.475 143.720 57.975 ;
        RECT 144.685 56.475 145.055 62.500 ;
        RECT 145.475 56.475 145.845 62.500 ;
        RECT 147.385 56.475 147.755 62.500 ;
        RECT 137.375 56.450 139.600 56.475 ;
        RECT 137.375 55.505 139.620 56.450 ;
        RECT 137.375 55.475 139.600 55.505 ;
        RECT 139.980 55.475 142.300 56.475 ;
        RECT 142.725 55.475 145.055 56.475 ;
        RECT 145.430 55.475 146.520 56.475 ;
        RECT 137.375 55.430 138.375 55.475 ;
        RECT 137.375 51.275 137.745 55.430 ;
        RECT 139.095 55.100 139.600 55.475 ;
        RECT 139.095 54.605 140.135 55.100 ;
        RECT 140.445 54.200 141.020 55.475 ;
        RECT 141.795 55.100 142.300 55.475 ;
        RECT 141.795 54.605 142.835 55.100 ;
        RECT 143.145 54.200 143.720 55.475 ;
        RECT 138.600 53.825 139.655 54.200 ;
        RECT 140.075 53.825 141.020 54.200 ;
        RECT 141.300 53.825 142.355 54.200 ;
        RECT 142.775 53.825 143.720 54.200 ;
        RECT 138.600 52.950 139.600 53.825 ;
        RECT 141.300 52.950 142.300 53.825 ;
        RECT 138.600 51.950 142.300 52.950 ;
        RECT 142.875 52.275 143.875 52.320 ;
        RECT 144.055 52.275 145.055 55.475 ;
        RECT 138.600 50.435 139.600 51.950 ;
        RECT 142.875 51.275 145.055 52.275 ;
        RECT 145.475 51.275 145.845 55.475 ;
        RECT 146.750 53.975 147.755 56.475 ;
        RECT 148.175 56.475 148.545 62.500 ;
        RECT 152.425 56.475 153.425 56.505 ;
        RECT 148.175 55.475 153.425 56.475 ;
        RECT 146.730 53.025 147.770 53.975 ;
        RECT 146.750 53.000 147.755 53.025 ;
        RECT 147.385 51.275 147.755 53.000 ;
        RECT 148.175 51.275 148.545 55.475 ;
        RECT 152.425 55.445 153.425 55.475 ;
        RECT 142.875 51.230 143.875 51.275 ;
        RECT 1.850 50.425 14.575 50.435 ;
        RECT 15.350 50.425 19.390 50.435 ;
        RECT 19.590 50.425 40.000 50.435 ;
        RECT 40.775 50.425 44.815 50.435 ;
        RECT 45.015 50.425 65.425 50.435 ;
        RECT 66.200 50.425 70.240 50.435 ;
        RECT 70.440 50.425 90.850 50.435 ;
        RECT 91.625 50.425 95.665 50.435 ;
        RECT 95.865 50.425 116.275 50.435 ;
        RECT 117.050 50.425 121.090 50.435 ;
        RECT 121.290 50.425 141.700 50.435 ;
        RECT 142.475 50.425 146.515 50.435 ;
        RECT 146.715 50.425 149.215 50.435 ;
        RECT 1.850 49.325 149.215 50.425 ;
        RECT 1.850 49.320 19.390 49.325 ;
        RECT 19.590 49.320 44.815 49.325 ;
        RECT 45.015 49.320 70.240 49.325 ;
        RECT 70.440 49.320 95.665 49.325 ;
        RECT 95.865 49.320 121.090 49.325 ;
        RECT 121.290 49.320 146.515 49.325 ;
        RECT 146.715 49.320 149.215 49.325 ;
        RECT 3.905 49.315 6.480 49.320 ;
        RECT 29.330 49.315 31.905 49.320 ;
        RECT 54.755 49.315 57.330 49.320 ;
        RECT 80.180 49.315 82.755 49.320 ;
        RECT 105.605 49.315 108.180 49.320 ;
        RECT 131.030 49.315 133.605 49.320 ;
        RECT 3.905 49.285 5.020 49.315 ;
        RECT 29.330 49.285 30.445 49.315 ;
        RECT 54.755 49.285 55.870 49.315 ;
        RECT 80.180 49.285 81.295 49.315 ;
        RECT 105.605 49.285 106.720 49.315 ;
        RECT 131.030 49.285 132.145 49.315 ;
        RECT 19.370 48.375 21.325 48.395 ;
        RECT 44.795 48.375 46.750 48.395 ;
        RECT 70.220 48.375 72.175 48.395 ;
        RECT 95.645 48.375 97.600 48.395 ;
        RECT 121.070 48.375 123.025 48.395 ;
        RECT 146.495 48.375 148.450 48.395 ;
        RECT 9.550 48.350 10.550 48.375 ;
        RECT 15.750 48.350 16.750 48.375 ;
        RECT 17.650 48.350 18.650 48.375 ;
        RECT 9.530 47.400 10.570 48.350 ;
        RECT 15.730 47.400 16.770 48.350 ;
        RECT 17.630 47.400 18.670 48.350 ;
        RECT 9.550 47.375 10.550 47.400 ;
        RECT 15.750 47.375 16.750 47.400 ;
        RECT 17.650 47.375 18.650 47.400 ;
        RECT 19.365 47.375 21.350 48.375 ;
        RECT 34.975 48.350 35.975 48.375 ;
        RECT 41.175 48.350 42.175 48.375 ;
        RECT 43.075 48.350 44.075 48.375 ;
        RECT 34.955 47.400 35.995 48.350 ;
        RECT 41.155 47.400 42.195 48.350 ;
        RECT 43.055 47.400 44.095 48.350 ;
        RECT 34.975 47.375 35.975 47.400 ;
        RECT 41.175 47.375 42.175 47.400 ;
        RECT 43.075 47.375 44.075 47.400 ;
        RECT 44.790 47.375 46.775 48.375 ;
        RECT 60.400 48.350 61.400 48.375 ;
        RECT 66.600 48.350 67.600 48.375 ;
        RECT 68.500 48.350 69.500 48.375 ;
        RECT 60.380 47.400 61.420 48.350 ;
        RECT 66.580 47.400 67.620 48.350 ;
        RECT 68.480 47.400 69.520 48.350 ;
        RECT 60.400 47.375 61.400 47.400 ;
        RECT 66.600 47.375 67.600 47.400 ;
        RECT 68.500 47.375 69.500 47.400 ;
        RECT 70.215 47.375 72.200 48.375 ;
        RECT 85.825 48.350 86.825 48.375 ;
        RECT 92.025 48.350 93.025 48.375 ;
        RECT 93.925 48.350 94.925 48.375 ;
        RECT 85.805 47.400 86.845 48.350 ;
        RECT 92.005 47.400 93.045 48.350 ;
        RECT 93.905 47.400 94.945 48.350 ;
        RECT 85.825 47.375 86.825 47.400 ;
        RECT 92.025 47.375 93.025 47.400 ;
        RECT 93.925 47.375 94.925 47.400 ;
        RECT 95.640 47.375 97.625 48.375 ;
        RECT 111.250 48.350 112.250 48.375 ;
        RECT 117.450 48.350 118.450 48.375 ;
        RECT 119.350 48.350 120.350 48.375 ;
        RECT 111.230 47.400 112.270 48.350 ;
        RECT 117.430 47.400 118.470 48.350 ;
        RECT 119.330 47.400 120.370 48.350 ;
        RECT 111.250 47.375 112.250 47.400 ;
        RECT 117.450 47.375 118.450 47.400 ;
        RECT 119.350 47.375 120.350 47.400 ;
        RECT 121.065 47.375 123.050 48.375 ;
        RECT 136.675 48.350 137.675 48.375 ;
        RECT 142.875 48.350 143.875 48.375 ;
        RECT 144.775 48.350 145.775 48.375 ;
        RECT 136.655 47.400 137.695 48.350 ;
        RECT 142.855 47.400 143.895 48.350 ;
        RECT 144.755 47.400 145.795 48.350 ;
        RECT 136.675 47.375 137.675 47.400 ;
        RECT 142.875 47.375 143.875 47.400 ;
        RECT 144.775 47.375 145.775 47.400 ;
        RECT 146.490 47.375 148.475 48.375 ;
        RECT 19.370 47.355 21.325 47.375 ;
        RECT 44.795 47.355 46.750 47.375 ;
        RECT 70.220 47.355 72.175 47.375 ;
        RECT 95.645 47.355 97.600 47.375 ;
        RECT 121.070 47.355 123.025 47.375 ;
        RECT 146.495 47.355 148.450 47.375 ;
        RECT 9.575 45.600 10.525 45.620 ;
        RECT 20.375 45.600 21.325 45.620 ;
        RECT 35.000 45.600 35.950 45.620 ;
        RECT 45.800 45.600 46.750 45.620 ;
        RECT 60.425 45.600 61.375 45.620 ;
        RECT 71.225 45.600 72.175 45.620 ;
        RECT 85.850 45.600 86.800 45.620 ;
        RECT 96.650 45.600 97.600 45.620 ;
        RECT 111.275 45.600 112.225 45.620 ;
        RECT 122.075 45.600 123.025 45.620 ;
        RECT 136.700 45.600 137.650 45.620 ;
        RECT 147.500 45.600 148.450 45.620 ;
        RECT 9.550 44.600 12.755 45.600 ;
        RECT 13.530 44.600 14.620 45.600 ;
        RECT 15.370 44.600 18.650 45.600 ;
        RECT 20.350 44.600 21.350 45.600 ;
        RECT 34.975 44.600 38.180 45.600 ;
        RECT 38.955 44.600 40.045 45.600 ;
        RECT 40.795 44.600 44.075 45.600 ;
        RECT 45.775 44.600 46.775 45.600 ;
        RECT 60.400 44.600 63.605 45.600 ;
        RECT 64.380 44.600 65.470 45.600 ;
        RECT 66.220 44.600 69.500 45.600 ;
        RECT 71.200 44.600 72.200 45.600 ;
        RECT 85.825 44.600 89.030 45.600 ;
        RECT 89.805 44.600 90.895 45.600 ;
        RECT 91.645 44.600 94.925 45.600 ;
        RECT 96.625 44.600 97.625 45.600 ;
        RECT 111.250 44.600 114.455 45.600 ;
        RECT 115.230 44.600 116.320 45.600 ;
        RECT 117.070 44.600 120.350 45.600 ;
        RECT 122.050 44.600 123.050 45.600 ;
        RECT 136.675 44.600 139.880 45.600 ;
        RECT 140.655 44.600 141.745 45.600 ;
        RECT 142.495 44.600 145.775 45.600 ;
        RECT 147.475 44.600 148.475 45.600 ;
        RECT 9.575 44.580 10.525 44.600 ;
        RECT 3.925 43.655 4.980 43.675 ;
        RECT 3.575 43.650 6.000 43.655 ;
        RECT 1.850 42.550 12.025 43.650 ;
        RECT 13.575 43.625 14.575 44.600 ;
        RECT 20.375 44.580 21.325 44.600 ;
        RECT 35.000 44.580 35.950 44.600 ;
        RECT 29.350 43.655 30.405 43.675 ;
        RECT 29.000 43.650 31.425 43.655 ;
        RECT 12.650 42.625 14.575 43.625 ;
        RECT 1.850 42.545 11.290 42.550 ;
        RECT 3.925 42.530 4.980 42.545 ;
        RECT 6.050 36.400 7.050 42.545 ;
        RECT 12.650 41.250 13.650 42.625 ;
        RECT 16.175 42.550 37.450 43.650 ;
        RECT 39.000 43.625 40.000 44.600 ;
        RECT 45.800 44.580 46.750 44.600 ;
        RECT 60.425 44.580 61.375 44.600 ;
        RECT 54.775 43.655 55.830 43.675 ;
        RECT 54.425 43.650 56.850 43.655 ;
        RECT 38.075 42.625 40.000 43.625 ;
        RECT 16.890 42.545 19.400 42.550 ;
        RECT 19.590 42.545 36.715 42.550 ;
        RECT 29.350 42.530 30.405 42.545 ;
        RECT 12.630 40.300 13.670 41.250 ;
        RECT 12.650 40.275 13.650 40.300 ;
        RECT 14.405 40.275 15.495 41.275 ;
        RECT 6.050 35.400 7.075 36.400 ;
        RECT 7.550 35.400 8.495 35.925 ;
        RECT 6.570 34.275 7.610 34.750 ;
        RECT 1.900 33.925 2.900 33.930 ;
        RECT 1.870 33.900 2.930 33.925 ;
        RECT 6.570 33.900 7.075 34.275 ;
        RECT 7.920 33.945 8.495 35.400 ;
        RECT 1.850 33.875 7.075 33.900 ;
        RECT 1.850 32.925 7.095 33.875 ;
        RECT 1.850 32.900 7.075 32.925 ;
        RECT 1.900 32.870 2.900 32.900 ;
        RECT 6.570 32.525 7.075 32.900 ;
        RECT 7.500 32.855 8.500 33.945 ;
        RECT 9.460 33.900 9.830 39.925 ;
        RECT 8.825 32.900 9.830 33.900 ;
        RECT 6.570 32.030 7.610 32.525 ;
        RECT 7.920 31.625 8.495 32.855 ;
        RECT 6.075 31.250 7.130 31.625 ;
        RECT 7.550 31.250 8.495 31.625 ;
        RECT 3.905 27.860 5.020 27.885 ;
        RECT 6.075 27.860 7.075 31.250 ;
        RECT 8.830 29.700 9.830 32.900 ;
        RECT 7.630 28.700 9.830 29.700 ;
        RECT 10.250 33.945 10.620 39.925 ;
        RECT 14.450 39.500 15.450 39.530 ;
        RECT 14.450 38.500 17.220 39.500 ;
        RECT 14.450 38.470 15.450 38.500 ;
        RECT 11.475 35.400 12.475 37.850 ;
        RECT 12.950 35.400 13.895 35.925 ;
        RECT 14.175 35.400 15.175 37.850 ;
        RECT 15.650 35.400 16.595 35.925 ;
        RECT 11.970 34.275 13.010 34.750 ;
        RECT 10.250 33.900 11.250 33.945 ;
        RECT 11.970 33.900 12.475 34.275 ;
        RECT 13.320 33.900 13.895 35.400 ;
        RECT 14.670 34.275 15.710 34.750 ;
        RECT 14.670 33.900 15.175 34.275 ;
        RECT 16.020 33.900 16.595 35.400 ;
        RECT 17.560 33.900 17.930 39.925 ;
        RECT 18.350 33.900 18.720 39.925 ;
        RECT 20.260 33.900 20.630 39.925 ;
        RECT 10.250 33.875 12.475 33.900 ;
        RECT 10.250 32.930 12.495 33.875 ;
        RECT 10.250 32.900 12.475 32.930 ;
        RECT 12.855 32.900 15.175 33.900 ;
        RECT 15.600 32.900 17.930 33.900 ;
        RECT 18.305 32.900 19.395 33.900 ;
        RECT 10.250 32.855 11.250 32.900 ;
        RECT 10.250 28.700 10.620 32.855 ;
        RECT 11.970 32.525 12.475 32.900 ;
        RECT 11.970 32.030 13.010 32.525 ;
        RECT 13.320 31.625 13.895 32.900 ;
        RECT 14.670 32.525 15.175 32.900 ;
        RECT 14.670 32.030 15.710 32.525 ;
        RECT 16.020 31.625 16.595 32.900 ;
        RECT 11.475 31.250 12.530 31.625 ;
        RECT 12.950 31.250 13.895 31.625 ;
        RECT 14.175 31.250 15.230 31.625 ;
        RECT 15.650 31.250 16.595 31.625 ;
        RECT 11.475 30.375 12.475 31.250 ;
        RECT 14.175 30.375 15.175 31.250 ;
        RECT 11.475 29.375 15.175 30.375 ;
        RECT 15.750 29.700 16.750 29.745 ;
        RECT 16.930 29.700 17.930 32.900 ;
        RECT 11.475 27.860 12.475 29.375 ;
        RECT 15.750 28.700 17.930 29.700 ;
        RECT 18.350 28.700 18.720 32.900 ;
        RECT 19.625 31.900 20.630 33.900 ;
        RECT 21.050 33.925 21.420 39.925 ;
        RECT 31.475 36.400 32.475 42.545 ;
        RECT 38.075 41.250 39.075 42.625 ;
        RECT 41.600 42.550 62.875 43.650 ;
        RECT 64.425 43.625 65.425 44.600 ;
        RECT 71.225 44.580 72.175 44.600 ;
        RECT 85.850 44.580 86.800 44.600 ;
        RECT 80.200 43.655 81.255 43.675 ;
        RECT 79.850 43.650 82.275 43.655 ;
        RECT 63.500 42.625 65.425 43.625 ;
        RECT 42.315 42.545 44.825 42.550 ;
        RECT 45.015 42.545 62.140 42.550 ;
        RECT 54.775 42.530 55.830 42.545 ;
        RECT 38.055 40.300 39.095 41.250 ;
        RECT 38.075 40.275 39.075 40.300 ;
        RECT 39.830 40.275 40.920 41.275 ;
        RECT 31.475 35.400 32.500 36.400 ;
        RECT 32.975 35.400 33.920 35.925 ;
        RECT 31.995 34.275 33.035 34.750 ;
        RECT 27.325 33.925 28.325 33.930 ;
        RECT 21.050 33.900 22.375 33.925 ;
        RECT 27.295 33.900 28.355 33.925 ;
        RECT 31.995 33.900 32.500 34.275 ;
        RECT 33.345 33.945 33.920 35.400 ;
        RECT 21.050 32.900 26.250 33.900 ;
        RECT 27.275 33.875 32.500 33.900 ;
        RECT 27.275 32.925 32.520 33.875 ;
        RECT 27.275 32.900 32.500 32.925 ;
        RECT 21.050 32.885 22.375 32.900 ;
        RECT 19.605 30.950 20.645 31.900 ;
        RECT 19.625 30.925 20.630 30.950 ;
        RECT 20.260 28.700 20.630 30.925 ;
        RECT 21.050 28.700 21.420 32.885 ;
        RECT 23.155 29.775 24.155 32.900 ;
        RECT 27.325 32.870 28.325 32.900 ;
        RECT 31.995 32.525 32.500 32.900 ;
        RECT 32.925 32.855 33.925 33.945 ;
        RECT 34.885 33.900 35.255 39.925 ;
        RECT 34.250 32.900 35.255 33.900 ;
        RECT 31.995 32.030 33.035 32.525 ;
        RECT 33.345 31.625 33.920 32.855 ;
        RECT 31.500 31.250 32.555 31.625 ;
        RECT 32.975 31.250 33.920 31.625 ;
        RECT 23.135 28.825 24.175 29.775 ;
        RECT 23.155 28.800 24.155 28.825 ;
        RECT 15.750 28.655 16.750 28.700 ;
        RECT 23.115 27.860 24.230 27.890 ;
        RECT 29.330 27.860 30.445 27.885 ;
        RECT 31.500 27.860 32.500 31.250 ;
        RECT 34.255 29.700 35.255 32.900 ;
        RECT 33.055 28.700 35.255 29.700 ;
        RECT 35.675 33.945 36.045 39.925 ;
        RECT 39.875 39.500 40.875 39.530 ;
        RECT 39.875 38.500 42.645 39.500 ;
        RECT 39.875 38.470 40.875 38.500 ;
        RECT 36.900 35.400 37.900 37.850 ;
        RECT 38.375 35.400 39.320 35.925 ;
        RECT 39.600 35.400 40.600 37.850 ;
        RECT 41.075 35.400 42.020 35.925 ;
        RECT 37.395 34.275 38.435 34.750 ;
        RECT 35.675 33.900 36.675 33.945 ;
        RECT 37.395 33.900 37.900 34.275 ;
        RECT 38.745 33.900 39.320 35.400 ;
        RECT 40.095 34.275 41.135 34.750 ;
        RECT 40.095 33.900 40.600 34.275 ;
        RECT 41.445 33.900 42.020 35.400 ;
        RECT 42.985 33.900 43.355 39.925 ;
        RECT 43.775 33.900 44.145 39.925 ;
        RECT 45.685 33.900 46.055 39.925 ;
        RECT 35.675 33.875 37.900 33.900 ;
        RECT 35.675 32.930 37.920 33.875 ;
        RECT 35.675 32.900 37.900 32.930 ;
        RECT 38.280 32.900 40.600 33.900 ;
        RECT 41.025 32.900 43.355 33.900 ;
        RECT 43.730 32.900 44.820 33.900 ;
        RECT 35.675 32.855 36.675 32.900 ;
        RECT 35.675 28.700 36.045 32.855 ;
        RECT 37.395 32.525 37.900 32.900 ;
        RECT 37.395 32.030 38.435 32.525 ;
        RECT 38.745 31.625 39.320 32.900 ;
        RECT 40.095 32.525 40.600 32.900 ;
        RECT 40.095 32.030 41.135 32.525 ;
        RECT 41.445 31.625 42.020 32.900 ;
        RECT 36.900 31.250 37.955 31.625 ;
        RECT 38.375 31.250 39.320 31.625 ;
        RECT 39.600 31.250 40.655 31.625 ;
        RECT 41.075 31.250 42.020 31.625 ;
        RECT 36.900 30.375 37.900 31.250 ;
        RECT 39.600 30.375 40.600 31.250 ;
        RECT 36.900 29.375 40.600 30.375 ;
        RECT 41.175 29.700 42.175 29.745 ;
        RECT 42.355 29.700 43.355 32.900 ;
        RECT 36.900 27.860 37.900 29.375 ;
        RECT 41.175 28.700 43.355 29.700 ;
        RECT 43.775 28.700 44.145 32.900 ;
        RECT 45.050 31.900 46.055 33.900 ;
        RECT 46.475 33.900 46.845 39.925 ;
        RECT 56.900 36.400 57.900 42.545 ;
        RECT 63.500 41.250 64.500 42.625 ;
        RECT 67.025 42.550 88.300 43.650 ;
        RECT 89.850 43.625 90.850 44.600 ;
        RECT 96.650 44.580 97.600 44.600 ;
        RECT 111.275 44.580 112.225 44.600 ;
        RECT 105.625 43.655 106.680 43.675 ;
        RECT 105.275 43.650 107.700 43.655 ;
        RECT 88.925 42.625 90.850 43.625 ;
        RECT 67.740 42.545 70.250 42.550 ;
        RECT 70.440 42.545 87.565 42.550 ;
        RECT 80.200 42.530 81.255 42.545 ;
        RECT 63.480 40.300 64.520 41.250 ;
        RECT 63.500 40.275 64.500 40.300 ;
        RECT 65.255 40.275 66.345 41.275 ;
        RECT 56.900 35.400 57.925 36.400 ;
        RECT 58.400 35.400 59.345 35.925 ;
        RECT 57.420 34.275 58.460 34.750 ;
        RECT 52.750 33.925 53.750 33.930 ;
        RECT 52.720 33.900 53.780 33.925 ;
        RECT 57.420 33.900 57.925 34.275 ;
        RECT 58.770 33.945 59.345 35.400 ;
        RECT 46.475 32.900 51.720 33.900 ;
        RECT 52.700 33.875 57.925 33.900 ;
        RECT 52.700 32.925 57.945 33.875 ;
        RECT 52.700 32.900 57.925 32.925 ;
        RECT 45.030 30.950 46.070 31.900 ;
        RECT 45.050 30.925 46.055 30.950 ;
        RECT 45.685 28.700 46.055 30.925 ;
        RECT 46.475 28.700 46.845 32.900 ;
        RECT 48.580 29.775 49.580 32.900 ;
        RECT 52.750 32.870 53.750 32.900 ;
        RECT 57.420 32.525 57.925 32.900 ;
        RECT 58.350 32.855 59.350 33.945 ;
        RECT 60.310 33.900 60.680 39.925 ;
        RECT 59.675 32.900 60.680 33.900 ;
        RECT 57.420 32.030 58.460 32.525 ;
        RECT 58.770 31.625 59.345 32.855 ;
        RECT 56.925 31.250 57.980 31.625 ;
        RECT 58.400 31.250 59.345 31.625 ;
        RECT 48.560 28.825 49.600 29.775 ;
        RECT 48.580 28.800 49.580 28.825 ;
        RECT 41.175 28.655 42.175 28.700 ;
        RECT 48.540 27.860 49.655 27.890 ;
        RECT 54.755 27.860 55.870 27.885 ;
        RECT 56.925 27.860 57.925 31.250 ;
        RECT 59.680 29.700 60.680 32.900 ;
        RECT 58.480 28.700 60.680 29.700 ;
        RECT 61.100 33.945 61.470 39.925 ;
        RECT 65.300 39.500 66.300 39.530 ;
        RECT 65.300 38.500 68.070 39.500 ;
        RECT 65.300 38.470 66.300 38.500 ;
        RECT 62.325 35.400 63.325 37.850 ;
        RECT 63.800 35.400 64.745 35.925 ;
        RECT 65.025 35.400 66.025 37.850 ;
        RECT 66.500 35.400 67.445 35.925 ;
        RECT 62.820 34.275 63.860 34.750 ;
        RECT 61.100 33.900 62.100 33.945 ;
        RECT 62.820 33.900 63.325 34.275 ;
        RECT 64.170 33.900 64.745 35.400 ;
        RECT 65.520 34.275 66.560 34.750 ;
        RECT 65.520 33.900 66.025 34.275 ;
        RECT 66.870 33.900 67.445 35.400 ;
        RECT 68.410 33.900 68.780 39.925 ;
        RECT 69.200 33.900 69.570 39.925 ;
        RECT 71.110 33.900 71.480 39.925 ;
        RECT 61.100 33.875 63.325 33.900 ;
        RECT 61.100 32.930 63.345 33.875 ;
        RECT 61.100 32.900 63.325 32.930 ;
        RECT 63.705 32.900 66.025 33.900 ;
        RECT 66.450 32.900 68.780 33.900 ;
        RECT 69.155 32.900 70.245 33.900 ;
        RECT 61.100 32.855 62.100 32.900 ;
        RECT 61.100 28.700 61.470 32.855 ;
        RECT 62.820 32.525 63.325 32.900 ;
        RECT 62.820 32.030 63.860 32.525 ;
        RECT 64.170 31.625 64.745 32.900 ;
        RECT 65.520 32.525 66.025 32.900 ;
        RECT 65.520 32.030 66.560 32.525 ;
        RECT 66.870 31.625 67.445 32.900 ;
        RECT 62.325 31.250 63.380 31.625 ;
        RECT 63.800 31.250 64.745 31.625 ;
        RECT 65.025 31.250 66.080 31.625 ;
        RECT 66.500 31.250 67.445 31.625 ;
        RECT 62.325 30.375 63.325 31.250 ;
        RECT 65.025 30.375 66.025 31.250 ;
        RECT 62.325 29.375 66.025 30.375 ;
        RECT 66.600 29.700 67.600 29.745 ;
        RECT 67.780 29.700 68.780 32.900 ;
        RECT 62.325 27.860 63.325 29.375 ;
        RECT 66.600 28.700 68.780 29.700 ;
        RECT 69.200 28.700 69.570 32.900 ;
        RECT 70.475 31.900 71.480 33.900 ;
        RECT 71.900 33.925 72.270 39.925 ;
        RECT 82.325 36.400 83.325 42.545 ;
        RECT 88.925 41.250 89.925 42.625 ;
        RECT 92.450 42.550 113.725 43.650 ;
        RECT 115.275 43.625 116.275 44.600 ;
        RECT 122.075 44.580 123.025 44.600 ;
        RECT 136.700 44.580 137.650 44.600 ;
        RECT 131.050 43.655 132.105 43.675 ;
        RECT 130.700 43.650 133.125 43.655 ;
        RECT 114.350 42.625 116.275 43.625 ;
        RECT 93.165 42.545 95.675 42.550 ;
        RECT 95.865 42.545 112.990 42.550 ;
        RECT 105.625 42.530 106.680 42.545 ;
        RECT 88.905 40.300 89.945 41.250 ;
        RECT 88.925 40.275 89.925 40.300 ;
        RECT 90.680 40.275 91.770 41.275 ;
        RECT 82.325 35.400 83.350 36.400 ;
        RECT 83.825 35.400 84.770 35.925 ;
        RECT 82.845 34.275 83.885 34.750 ;
        RECT 78.175 33.925 79.175 33.930 ;
        RECT 71.900 33.900 73.225 33.925 ;
        RECT 78.145 33.900 79.205 33.925 ;
        RECT 82.845 33.900 83.350 34.275 ;
        RECT 84.195 33.945 84.770 35.400 ;
        RECT 71.900 32.900 77.100 33.900 ;
        RECT 78.125 33.875 83.350 33.900 ;
        RECT 78.125 32.925 83.370 33.875 ;
        RECT 78.125 32.900 83.350 32.925 ;
        RECT 71.900 32.885 73.225 32.900 ;
        RECT 70.455 30.950 71.495 31.900 ;
        RECT 70.475 30.925 71.480 30.950 ;
        RECT 71.110 28.700 71.480 30.925 ;
        RECT 71.900 28.700 72.270 32.885 ;
        RECT 74.005 29.775 75.005 32.900 ;
        RECT 78.175 32.870 79.175 32.900 ;
        RECT 82.845 32.525 83.350 32.900 ;
        RECT 83.775 32.855 84.775 33.945 ;
        RECT 85.735 33.900 86.105 39.925 ;
        RECT 85.100 32.900 86.105 33.900 ;
        RECT 82.845 32.030 83.885 32.525 ;
        RECT 84.195 31.625 84.770 32.855 ;
        RECT 82.350 31.250 83.405 31.625 ;
        RECT 83.825 31.250 84.770 31.625 ;
        RECT 73.985 28.825 75.025 29.775 ;
        RECT 74.005 28.800 75.005 28.825 ;
        RECT 66.600 28.655 67.600 28.700 ;
        RECT 73.965 27.860 75.080 27.890 ;
        RECT 80.180 27.860 81.295 27.885 ;
        RECT 82.350 27.860 83.350 31.250 ;
        RECT 85.105 29.700 86.105 32.900 ;
        RECT 83.905 28.700 86.105 29.700 ;
        RECT 86.525 33.945 86.895 39.925 ;
        RECT 90.725 39.500 91.725 39.530 ;
        RECT 90.725 38.500 93.495 39.500 ;
        RECT 90.725 38.470 91.725 38.500 ;
        RECT 87.750 35.400 88.750 37.850 ;
        RECT 89.225 35.400 90.170 35.925 ;
        RECT 90.450 35.400 91.450 37.850 ;
        RECT 91.925 35.400 92.870 35.925 ;
        RECT 88.245 34.275 89.285 34.750 ;
        RECT 86.525 33.900 87.525 33.945 ;
        RECT 88.245 33.900 88.750 34.275 ;
        RECT 89.595 33.900 90.170 35.400 ;
        RECT 90.945 34.275 91.985 34.750 ;
        RECT 90.945 33.900 91.450 34.275 ;
        RECT 92.295 33.900 92.870 35.400 ;
        RECT 93.835 33.900 94.205 39.925 ;
        RECT 94.625 33.900 94.995 39.925 ;
        RECT 96.535 33.900 96.905 39.925 ;
        RECT 86.525 33.875 88.750 33.900 ;
        RECT 86.525 32.930 88.770 33.875 ;
        RECT 86.525 32.900 88.750 32.930 ;
        RECT 89.130 32.900 91.450 33.900 ;
        RECT 91.875 32.900 94.205 33.900 ;
        RECT 94.580 32.900 95.670 33.900 ;
        RECT 86.525 32.855 87.525 32.900 ;
        RECT 86.525 28.700 86.895 32.855 ;
        RECT 88.245 32.525 88.750 32.900 ;
        RECT 88.245 32.030 89.285 32.525 ;
        RECT 89.595 31.625 90.170 32.900 ;
        RECT 90.945 32.525 91.450 32.900 ;
        RECT 90.945 32.030 91.985 32.525 ;
        RECT 92.295 31.625 92.870 32.900 ;
        RECT 87.750 31.250 88.805 31.625 ;
        RECT 89.225 31.250 90.170 31.625 ;
        RECT 90.450 31.250 91.505 31.625 ;
        RECT 91.925 31.250 92.870 31.625 ;
        RECT 87.750 30.375 88.750 31.250 ;
        RECT 90.450 30.375 91.450 31.250 ;
        RECT 87.750 29.375 91.450 30.375 ;
        RECT 92.025 29.700 93.025 29.745 ;
        RECT 93.205 29.700 94.205 32.900 ;
        RECT 87.750 27.860 88.750 29.375 ;
        RECT 92.025 28.700 94.205 29.700 ;
        RECT 94.625 28.700 94.995 32.900 ;
        RECT 95.900 31.900 96.905 33.900 ;
        RECT 97.325 33.900 97.695 39.925 ;
        RECT 107.750 36.400 108.750 42.545 ;
        RECT 114.350 41.250 115.350 42.625 ;
        RECT 117.875 42.550 139.150 43.650 ;
        RECT 140.700 43.625 141.700 44.600 ;
        RECT 147.500 44.580 148.450 44.600 ;
        RECT 139.775 42.625 141.700 43.625 ;
        RECT 118.590 42.545 121.100 42.550 ;
        RECT 121.290 42.545 138.415 42.550 ;
        RECT 131.050 42.530 132.105 42.545 ;
        RECT 114.330 40.300 115.370 41.250 ;
        RECT 114.350 40.275 115.350 40.300 ;
        RECT 116.105 40.275 117.195 41.275 ;
        RECT 107.750 35.400 108.775 36.400 ;
        RECT 109.250 35.400 110.195 35.925 ;
        RECT 108.270 34.275 109.310 34.750 ;
        RECT 103.600 33.925 104.600 33.930 ;
        RECT 103.570 33.900 104.630 33.925 ;
        RECT 108.270 33.900 108.775 34.275 ;
        RECT 109.620 33.945 110.195 35.400 ;
        RECT 97.325 32.900 102.570 33.900 ;
        RECT 103.550 33.875 108.775 33.900 ;
        RECT 103.550 32.925 108.795 33.875 ;
        RECT 103.550 32.900 108.775 32.925 ;
        RECT 95.880 30.950 96.920 31.900 ;
        RECT 95.900 30.925 96.905 30.950 ;
        RECT 96.535 28.700 96.905 30.925 ;
        RECT 97.325 28.700 97.695 32.900 ;
        RECT 99.430 29.775 100.430 32.900 ;
        RECT 103.600 32.870 104.600 32.900 ;
        RECT 108.270 32.525 108.775 32.900 ;
        RECT 109.200 32.855 110.200 33.945 ;
        RECT 111.160 33.900 111.530 39.925 ;
        RECT 110.525 32.900 111.530 33.900 ;
        RECT 108.270 32.030 109.310 32.525 ;
        RECT 109.620 31.625 110.195 32.855 ;
        RECT 107.775 31.250 108.830 31.625 ;
        RECT 109.250 31.250 110.195 31.625 ;
        RECT 99.410 28.825 100.450 29.775 ;
        RECT 99.430 28.800 100.430 28.825 ;
        RECT 92.025 28.655 93.025 28.700 ;
        RECT 99.390 27.860 100.505 27.890 ;
        RECT 105.605 27.860 106.720 27.885 ;
        RECT 107.775 27.860 108.775 31.250 ;
        RECT 110.530 29.700 111.530 32.900 ;
        RECT 109.330 28.700 111.530 29.700 ;
        RECT 111.950 33.945 112.320 39.925 ;
        RECT 116.150 39.500 117.150 39.530 ;
        RECT 116.150 38.500 118.920 39.500 ;
        RECT 116.150 38.470 117.150 38.500 ;
        RECT 113.175 35.400 114.175 37.850 ;
        RECT 114.650 35.400 115.595 35.925 ;
        RECT 115.875 35.400 116.875 37.850 ;
        RECT 117.350 35.400 118.295 35.925 ;
        RECT 113.670 34.275 114.710 34.750 ;
        RECT 111.950 33.900 112.950 33.945 ;
        RECT 113.670 33.900 114.175 34.275 ;
        RECT 115.020 33.900 115.595 35.400 ;
        RECT 116.370 34.275 117.410 34.750 ;
        RECT 116.370 33.900 116.875 34.275 ;
        RECT 117.720 33.900 118.295 35.400 ;
        RECT 119.260 33.900 119.630 39.925 ;
        RECT 120.050 33.900 120.420 39.925 ;
        RECT 121.960 33.900 122.330 39.925 ;
        RECT 111.950 33.875 114.175 33.900 ;
        RECT 111.950 32.930 114.195 33.875 ;
        RECT 111.950 32.900 114.175 32.930 ;
        RECT 114.555 32.900 116.875 33.900 ;
        RECT 117.300 32.900 119.630 33.900 ;
        RECT 120.005 32.900 121.095 33.900 ;
        RECT 111.950 32.855 112.950 32.900 ;
        RECT 111.950 28.700 112.320 32.855 ;
        RECT 113.670 32.525 114.175 32.900 ;
        RECT 113.670 32.030 114.710 32.525 ;
        RECT 115.020 31.625 115.595 32.900 ;
        RECT 116.370 32.525 116.875 32.900 ;
        RECT 116.370 32.030 117.410 32.525 ;
        RECT 117.720 31.625 118.295 32.900 ;
        RECT 113.175 31.250 114.230 31.625 ;
        RECT 114.650 31.250 115.595 31.625 ;
        RECT 115.875 31.250 116.930 31.625 ;
        RECT 117.350 31.250 118.295 31.625 ;
        RECT 113.175 30.375 114.175 31.250 ;
        RECT 115.875 30.375 116.875 31.250 ;
        RECT 113.175 29.375 116.875 30.375 ;
        RECT 117.450 29.700 118.450 29.745 ;
        RECT 118.630 29.700 119.630 32.900 ;
        RECT 113.175 27.860 114.175 29.375 ;
        RECT 117.450 28.700 119.630 29.700 ;
        RECT 120.050 28.700 120.420 32.900 ;
        RECT 121.325 31.900 122.330 33.900 ;
        RECT 122.750 33.925 123.120 39.925 ;
        RECT 133.175 36.400 134.175 42.545 ;
        RECT 139.775 41.250 140.775 42.625 ;
        RECT 143.300 42.550 149.225 43.650 ;
        RECT 144.015 42.545 146.525 42.550 ;
        RECT 146.715 42.545 149.215 42.550 ;
        RECT 139.755 40.300 140.795 41.250 ;
        RECT 139.775 40.275 140.775 40.300 ;
        RECT 141.530 40.275 142.620 41.275 ;
        RECT 133.175 35.400 134.200 36.400 ;
        RECT 134.675 35.400 135.620 35.925 ;
        RECT 133.695 34.275 134.735 34.750 ;
        RECT 129.025 33.925 130.025 33.930 ;
        RECT 122.750 33.900 124.075 33.925 ;
        RECT 128.995 33.900 130.055 33.925 ;
        RECT 133.695 33.900 134.200 34.275 ;
        RECT 135.045 33.945 135.620 35.400 ;
        RECT 122.750 32.900 127.950 33.900 ;
        RECT 128.975 33.875 134.200 33.900 ;
        RECT 128.975 32.925 134.220 33.875 ;
        RECT 128.975 32.900 134.200 32.925 ;
        RECT 122.750 32.885 124.075 32.900 ;
        RECT 121.305 30.950 122.345 31.900 ;
        RECT 121.325 30.925 122.330 30.950 ;
        RECT 121.960 28.700 122.330 30.925 ;
        RECT 122.750 28.700 123.120 32.885 ;
        RECT 124.855 29.775 125.855 32.900 ;
        RECT 129.025 32.870 130.025 32.900 ;
        RECT 133.695 32.525 134.200 32.900 ;
        RECT 134.625 32.855 135.625 33.945 ;
        RECT 136.585 33.900 136.955 39.925 ;
        RECT 135.950 32.900 136.955 33.900 ;
        RECT 133.695 32.030 134.735 32.525 ;
        RECT 135.045 31.625 135.620 32.855 ;
        RECT 133.200 31.250 134.255 31.625 ;
        RECT 134.675 31.250 135.620 31.625 ;
        RECT 124.835 28.825 125.875 29.775 ;
        RECT 124.855 28.800 125.855 28.825 ;
        RECT 117.450 28.655 118.450 28.700 ;
        RECT 124.815 27.860 125.930 27.890 ;
        RECT 131.030 27.860 132.145 27.885 ;
        RECT 133.200 27.860 134.200 31.250 ;
        RECT 135.955 29.700 136.955 32.900 ;
        RECT 134.755 28.700 136.955 29.700 ;
        RECT 137.375 33.945 137.745 39.925 ;
        RECT 141.575 39.500 142.575 39.530 ;
        RECT 141.575 38.500 144.345 39.500 ;
        RECT 141.575 38.470 142.575 38.500 ;
        RECT 138.600 35.400 139.600 37.850 ;
        RECT 140.075 35.400 141.020 35.925 ;
        RECT 141.300 35.400 142.300 37.850 ;
        RECT 142.775 35.400 143.720 35.925 ;
        RECT 139.095 34.275 140.135 34.750 ;
        RECT 137.375 33.900 138.375 33.945 ;
        RECT 139.095 33.900 139.600 34.275 ;
        RECT 140.445 33.900 141.020 35.400 ;
        RECT 141.795 34.275 142.835 34.750 ;
        RECT 141.795 33.900 142.300 34.275 ;
        RECT 143.145 33.900 143.720 35.400 ;
        RECT 144.685 33.900 145.055 39.925 ;
        RECT 145.475 33.900 145.845 39.925 ;
        RECT 147.385 33.900 147.755 39.925 ;
        RECT 137.375 33.875 139.600 33.900 ;
        RECT 137.375 32.930 139.620 33.875 ;
        RECT 137.375 32.900 139.600 32.930 ;
        RECT 139.980 32.900 142.300 33.900 ;
        RECT 142.725 32.900 145.055 33.900 ;
        RECT 145.430 32.900 146.520 33.900 ;
        RECT 137.375 32.855 138.375 32.900 ;
        RECT 137.375 28.700 137.745 32.855 ;
        RECT 139.095 32.525 139.600 32.900 ;
        RECT 139.095 32.030 140.135 32.525 ;
        RECT 140.445 31.625 141.020 32.900 ;
        RECT 141.795 32.525 142.300 32.900 ;
        RECT 141.795 32.030 142.835 32.525 ;
        RECT 143.145 31.625 143.720 32.900 ;
        RECT 138.600 31.250 139.655 31.625 ;
        RECT 140.075 31.250 141.020 31.625 ;
        RECT 141.300 31.250 142.355 31.625 ;
        RECT 142.775 31.250 143.720 31.625 ;
        RECT 138.600 30.375 139.600 31.250 ;
        RECT 141.300 30.375 142.300 31.250 ;
        RECT 138.600 29.375 142.300 30.375 ;
        RECT 142.875 29.700 143.875 29.745 ;
        RECT 144.055 29.700 145.055 32.900 ;
        RECT 138.600 27.860 139.600 29.375 ;
        RECT 142.875 28.700 145.055 29.700 ;
        RECT 145.475 28.700 145.845 32.900 ;
        RECT 146.750 31.900 147.755 33.900 ;
        RECT 148.175 33.900 148.545 39.925 ;
        RECT 152.525 33.900 153.525 33.945 ;
        RECT 148.175 32.900 153.525 33.900 ;
        RECT 146.730 30.950 147.770 31.900 ;
        RECT 146.750 30.925 147.755 30.950 ;
        RECT 147.385 28.700 147.755 30.925 ;
        RECT 148.175 28.700 148.545 32.900 ;
        RECT 150.280 29.775 151.280 32.900 ;
        RECT 152.525 32.855 153.525 32.900 ;
        RECT 150.260 28.825 151.300 29.775 ;
        RECT 150.280 28.800 151.280 28.825 ;
        RECT 142.875 28.655 143.875 28.700 ;
        RECT 150.240 27.860 151.355 27.890 ;
        RECT 1.850 27.850 14.575 27.860 ;
        RECT 15.350 27.850 19.390 27.860 ;
        RECT 19.590 27.850 40.000 27.860 ;
        RECT 40.775 27.850 44.815 27.860 ;
        RECT 45.015 27.850 65.425 27.860 ;
        RECT 66.200 27.850 70.240 27.860 ;
        RECT 70.440 27.850 90.850 27.860 ;
        RECT 91.625 27.850 95.665 27.860 ;
        RECT 95.865 27.850 116.275 27.860 ;
        RECT 117.050 27.850 121.090 27.860 ;
        RECT 121.290 27.850 141.700 27.860 ;
        RECT 142.475 27.850 146.515 27.860 ;
        RECT 146.715 27.850 151.355 27.860 ;
        RECT 1.850 26.750 151.355 27.850 ;
        RECT 1.850 26.745 19.390 26.750 ;
        RECT 19.590 26.745 44.815 26.750 ;
        RECT 45.015 26.745 70.240 26.750 ;
        RECT 70.440 26.745 95.665 26.750 ;
        RECT 95.865 26.745 121.090 26.750 ;
        RECT 121.290 26.745 146.515 26.750 ;
        RECT 146.715 26.745 151.355 26.750 ;
        RECT 3.875 26.740 7.105 26.745 ;
        RECT 3.905 26.710 5.020 26.740 ;
        RECT 23.115 26.715 24.230 26.745 ;
        RECT 29.300 26.740 32.530 26.745 ;
        RECT 29.330 26.710 30.445 26.740 ;
        RECT 48.540 26.715 49.655 26.745 ;
        RECT 54.725 26.740 57.955 26.745 ;
        RECT 54.755 26.710 55.870 26.740 ;
        RECT 73.965 26.715 75.080 26.745 ;
        RECT 80.150 26.740 83.380 26.745 ;
        RECT 80.180 26.710 81.295 26.740 ;
        RECT 99.390 26.715 100.505 26.745 ;
        RECT 105.575 26.740 108.805 26.745 ;
        RECT 105.605 26.710 106.720 26.740 ;
        RECT 124.815 26.715 125.930 26.745 ;
        RECT 131.000 26.740 134.230 26.745 ;
        RECT 131.030 26.710 132.145 26.740 ;
        RECT 150.240 26.715 151.355 26.745 ;
        RECT 19.370 25.800 21.325 25.820 ;
        RECT 44.795 25.800 46.750 25.820 ;
        RECT 70.220 25.800 72.175 25.820 ;
        RECT 95.645 25.800 97.600 25.820 ;
        RECT 121.070 25.800 123.025 25.820 ;
        RECT 146.495 25.800 148.450 25.820 ;
        RECT 9.550 25.775 10.550 25.800 ;
        RECT 15.750 25.775 16.750 25.800 ;
        RECT 17.650 25.775 18.650 25.800 ;
        RECT 9.530 24.825 10.570 25.775 ;
        RECT 15.730 24.825 16.770 25.775 ;
        RECT 17.630 24.825 18.670 25.775 ;
        RECT 9.550 24.800 10.550 24.825 ;
        RECT 15.750 24.800 16.750 24.825 ;
        RECT 17.650 24.800 18.650 24.825 ;
        RECT 19.365 24.800 21.350 25.800 ;
        RECT 34.975 25.775 35.975 25.800 ;
        RECT 41.175 25.775 42.175 25.800 ;
        RECT 43.075 25.775 44.075 25.800 ;
        RECT 34.955 24.825 35.995 25.775 ;
        RECT 41.155 24.825 42.195 25.775 ;
        RECT 43.055 24.825 44.095 25.775 ;
        RECT 34.975 24.800 35.975 24.825 ;
        RECT 41.175 24.800 42.175 24.825 ;
        RECT 43.075 24.800 44.075 24.825 ;
        RECT 44.790 24.800 46.775 25.800 ;
        RECT 60.400 25.775 61.400 25.800 ;
        RECT 66.600 25.775 67.600 25.800 ;
        RECT 68.500 25.775 69.500 25.800 ;
        RECT 60.380 24.825 61.420 25.775 ;
        RECT 66.580 24.825 67.620 25.775 ;
        RECT 68.480 24.825 69.520 25.775 ;
        RECT 60.400 24.800 61.400 24.825 ;
        RECT 66.600 24.800 67.600 24.825 ;
        RECT 68.500 24.800 69.500 24.825 ;
        RECT 70.215 24.800 72.200 25.800 ;
        RECT 85.825 25.775 86.825 25.800 ;
        RECT 92.025 25.775 93.025 25.800 ;
        RECT 93.925 25.775 94.925 25.800 ;
        RECT 85.805 24.825 86.845 25.775 ;
        RECT 92.005 24.825 93.045 25.775 ;
        RECT 93.905 24.825 94.945 25.775 ;
        RECT 85.825 24.800 86.825 24.825 ;
        RECT 92.025 24.800 93.025 24.825 ;
        RECT 93.925 24.800 94.925 24.825 ;
        RECT 95.640 24.800 97.625 25.800 ;
        RECT 111.250 25.775 112.250 25.800 ;
        RECT 117.450 25.775 118.450 25.800 ;
        RECT 119.350 25.775 120.350 25.800 ;
        RECT 111.230 24.825 112.270 25.775 ;
        RECT 117.430 24.825 118.470 25.775 ;
        RECT 119.330 24.825 120.370 25.775 ;
        RECT 111.250 24.800 112.250 24.825 ;
        RECT 117.450 24.800 118.450 24.825 ;
        RECT 119.350 24.800 120.350 24.825 ;
        RECT 121.065 24.800 123.050 25.800 ;
        RECT 136.675 25.775 137.675 25.800 ;
        RECT 142.875 25.775 143.875 25.800 ;
        RECT 144.775 25.775 145.775 25.800 ;
        RECT 136.655 24.825 137.695 25.775 ;
        RECT 142.855 24.825 143.895 25.775 ;
        RECT 144.755 24.825 145.795 25.775 ;
        RECT 136.675 24.800 137.675 24.825 ;
        RECT 142.875 24.800 143.875 24.825 ;
        RECT 144.775 24.800 145.775 24.825 ;
        RECT 146.490 24.800 148.475 25.800 ;
        RECT 19.370 24.780 21.325 24.800 ;
        RECT 44.795 24.780 46.750 24.800 ;
        RECT 70.220 24.780 72.175 24.800 ;
        RECT 95.645 24.780 97.600 24.800 ;
        RECT 121.070 24.780 123.025 24.800 ;
        RECT 146.495 24.780 148.450 24.800 ;
        RECT 9.575 23.025 10.525 23.045 ;
        RECT 20.375 23.025 21.325 23.045 ;
        RECT 35.000 23.025 35.950 23.045 ;
        RECT 45.800 23.025 46.750 23.045 ;
        RECT 60.425 23.025 61.375 23.045 ;
        RECT 71.225 23.025 72.175 23.045 ;
        RECT 85.850 23.025 86.800 23.045 ;
        RECT 96.650 23.025 97.600 23.045 ;
        RECT 111.275 23.025 112.225 23.045 ;
        RECT 122.075 23.025 123.025 23.045 ;
        RECT 136.700 23.025 137.650 23.045 ;
        RECT 147.500 23.025 148.450 23.045 ;
        RECT 9.550 22.025 12.755 23.025 ;
        RECT 13.530 22.025 14.620 23.025 ;
        RECT 15.370 22.025 18.650 23.025 ;
        RECT 20.350 22.025 21.350 23.025 ;
        RECT 9.575 22.005 10.525 22.025 ;
        RECT 2.900 21.075 7.100 21.080 ;
        RECT 1.850 19.975 12.025 21.075 ;
        RECT 13.575 21.050 14.575 22.025 ;
        RECT 20.375 22.005 21.325 22.025 ;
        RECT 23.155 21.730 24.155 22.825 ;
        RECT 34.975 22.025 38.180 23.025 ;
        RECT 38.955 22.025 40.045 23.025 ;
        RECT 40.795 22.025 44.075 23.025 ;
        RECT 45.775 22.025 46.775 23.025 ;
        RECT 35.000 22.005 35.950 22.025 ;
        RECT 23.430 21.115 23.880 21.730 ;
        RECT 28.325 21.075 32.525 21.080 ;
        RECT 12.650 20.050 14.575 21.050 ;
        RECT 16.175 20.155 22.100 21.075 ;
        RECT 27.275 20.155 37.450 21.075 ;
        RECT 39.000 21.050 40.000 22.025 ;
        RECT 45.800 22.005 46.750 22.025 ;
        RECT 48.580 21.730 49.580 22.825 ;
        RECT 60.400 22.025 63.605 23.025 ;
        RECT 64.380 22.025 65.470 23.025 ;
        RECT 66.220 22.025 69.500 23.025 ;
        RECT 71.200 22.025 72.200 23.025 ;
        RECT 60.425 22.005 61.375 22.025 ;
        RECT 48.855 21.115 49.305 21.730 ;
        RECT 53.750 21.075 57.950 21.080 ;
        RECT 1.850 19.970 11.290 19.975 ;
        RECT 6.050 13.825 7.050 19.970 ;
        RECT 12.650 18.675 13.650 20.050 ;
        RECT 16.175 19.975 37.450 20.155 ;
        RECT 38.075 20.050 40.000 21.050 ;
        RECT 41.600 20.155 47.525 21.075 ;
        RECT 52.700 20.155 62.875 21.075 ;
        RECT 64.425 21.050 65.425 22.025 ;
        RECT 71.225 22.005 72.175 22.025 ;
        RECT 74.005 21.730 75.005 22.825 ;
        RECT 85.825 22.025 89.030 23.025 ;
        RECT 89.805 22.025 90.895 23.025 ;
        RECT 91.645 22.025 94.925 23.025 ;
        RECT 96.625 22.025 97.625 23.025 ;
        RECT 85.850 22.005 86.800 22.025 ;
        RECT 74.280 21.115 74.730 21.730 ;
        RECT 79.175 21.075 83.375 21.080 ;
        RECT 16.890 19.970 19.400 19.975 ;
        RECT 19.590 19.970 36.715 19.975 ;
        RECT 20.320 19.050 28.380 19.970 ;
        RECT 12.630 17.725 13.670 18.675 ;
        RECT 12.650 17.700 13.650 17.725 ;
        RECT 14.405 17.700 15.495 18.700 ;
        RECT 6.050 12.825 7.075 13.825 ;
        RECT 7.550 12.825 8.495 13.350 ;
        RECT 6.570 11.700 7.610 12.175 ;
        RECT 1.900 11.325 2.900 11.355 ;
        RECT 6.570 11.325 7.075 11.700 ;
        RECT 7.920 11.370 8.495 12.825 ;
        RECT 1.850 11.300 7.075 11.325 ;
        RECT 1.850 10.350 7.095 11.300 ;
        RECT 1.850 10.325 7.075 10.350 ;
        RECT 1.900 10.295 2.900 10.325 ;
        RECT 6.570 9.950 7.075 10.325 ;
        RECT 7.500 10.280 8.500 11.370 ;
        RECT 9.460 11.325 9.830 17.350 ;
        RECT 8.825 10.325 9.830 11.325 ;
        RECT 6.570 9.455 7.610 9.950 ;
        RECT 7.920 9.050 8.495 10.280 ;
        RECT 6.075 8.675 7.130 9.050 ;
        RECT 7.550 8.675 8.495 9.050 ;
        RECT 3.890 5.285 5.030 5.315 ;
        RECT 6.075 5.285 7.075 8.675 ;
        RECT 8.830 7.125 9.830 10.325 ;
        RECT 7.630 6.125 9.830 7.125 ;
        RECT 10.250 11.370 10.620 17.350 ;
        RECT 14.450 16.925 15.450 16.955 ;
        RECT 14.450 15.925 17.220 16.925 ;
        RECT 14.450 15.895 15.450 15.925 ;
        RECT 11.475 12.825 12.475 15.275 ;
        RECT 12.950 12.825 13.895 13.350 ;
        RECT 14.175 12.825 15.175 15.275 ;
        RECT 15.650 12.825 16.595 13.350 ;
        RECT 11.970 11.700 13.010 12.175 ;
        RECT 10.250 11.325 11.250 11.370 ;
        RECT 11.970 11.325 12.475 11.700 ;
        RECT 13.320 11.325 13.895 12.825 ;
        RECT 14.670 11.700 15.710 12.175 ;
        RECT 14.670 11.325 15.175 11.700 ;
        RECT 16.020 11.325 16.595 12.825 ;
        RECT 17.560 11.325 17.930 17.350 ;
        RECT 18.350 11.325 18.720 17.350 ;
        RECT 20.260 11.325 20.630 17.350 ;
        RECT 10.250 11.300 12.475 11.325 ;
        RECT 10.250 10.355 12.495 11.300 ;
        RECT 10.250 10.325 12.475 10.355 ;
        RECT 12.855 10.325 15.175 11.325 ;
        RECT 15.600 10.325 17.930 11.325 ;
        RECT 18.305 10.325 19.395 11.325 ;
        RECT 19.625 10.325 20.630 11.325 ;
        RECT 10.250 10.280 11.250 10.325 ;
        RECT 10.250 6.125 10.620 10.280 ;
        RECT 11.970 9.950 12.475 10.325 ;
        RECT 11.970 9.455 13.010 9.950 ;
        RECT 13.320 9.050 13.895 10.325 ;
        RECT 14.670 9.950 15.175 10.325 ;
        RECT 14.670 9.455 15.710 9.950 ;
        RECT 16.020 9.050 16.595 10.325 ;
        RECT 11.475 8.675 12.530 9.050 ;
        RECT 12.950 8.675 13.895 9.050 ;
        RECT 14.175 8.675 15.230 9.050 ;
        RECT 15.650 8.675 16.595 9.050 ;
        RECT 11.475 7.800 12.475 8.675 ;
        RECT 14.175 7.800 15.175 8.675 ;
        RECT 11.475 6.800 15.175 7.800 ;
        RECT 15.750 7.125 16.750 7.170 ;
        RECT 16.930 7.125 17.930 10.325 ;
        RECT 11.475 5.285 12.475 6.800 ;
        RECT 15.750 6.125 17.930 7.125 ;
        RECT 18.350 6.125 18.720 10.325 ;
        RECT 19.630 9.325 20.630 10.325 ;
        RECT 21.050 11.325 21.420 17.350 ;
        RECT 31.475 13.825 32.475 19.970 ;
        RECT 38.075 18.675 39.075 20.050 ;
        RECT 41.600 19.975 62.875 20.155 ;
        RECT 63.500 20.050 65.425 21.050 ;
        RECT 67.025 20.155 72.950 21.075 ;
        RECT 78.125 20.155 88.300 21.075 ;
        RECT 89.850 21.050 90.850 22.025 ;
        RECT 96.650 22.005 97.600 22.025 ;
        RECT 99.430 21.730 100.430 22.825 ;
        RECT 111.250 22.025 114.455 23.025 ;
        RECT 115.230 22.025 116.320 23.025 ;
        RECT 117.070 22.025 120.350 23.025 ;
        RECT 122.050 22.025 123.050 23.025 ;
        RECT 111.275 22.005 112.225 22.025 ;
        RECT 99.705 21.115 100.155 21.730 ;
        RECT 104.600 21.075 108.800 21.080 ;
        RECT 42.315 19.970 44.825 19.975 ;
        RECT 45.015 19.970 62.140 19.975 ;
        RECT 45.745 19.050 53.805 19.970 ;
        RECT 38.055 17.725 39.095 18.675 ;
        RECT 38.075 17.700 39.075 17.725 ;
        RECT 39.830 17.700 40.920 18.700 ;
        RECT 31.475 12.825 32.500 13.825 ;
        RECT 32.975 12.825 33.920 13.350 ;
        RECT 23.430 11.875 23.880 12.515 ;
        RECT 23.150 11.325 24.150 11.875 ;
        RECT 31.995 11.700 33.035 12.175 ;
        RECT 27.325 11.325 28.325 11.355 ;
        RECT 31.995 11.325 32.500 11.700 ;
        RECT 33.345 11.370 33.920 12.825 ;
        RECT 21.050 10.325 24.150 11.325 ;
        RECT 27.275 11.300 32.500 11.325 ;
        RECT 27.275 10.350 32.520 11.300 ;
        RECT 27.275 10.325 32.500 10.350 ;
        RECT 19.585 8.325 20.675 9.325 ;
        RECT 20.260 6.125 20.630 8.325 ;
        RECT 21.050 6.125 21.420 10.325 ;
        RECT 23.430 10.205 23.880 10.325 ;
        RECT 27.325 10.295 28.325 10.325 ;
        RECT 31.995 9.950 32.500 10.325 ;
        RECT 32.925 10.280 33.925 11.370 ;
        RECT 34.885 11.325 35.255 17.350 ;
        RECT 34.250 10.325 35.255 11.325 ;
        RECT 31.995 9.455 33.035 9.950 ;
        RECT 33.345 9.050 33.920 10.280 ;
        RECT 31.500 8.675 32.555 9.050 ;
        RECT 32.975 8.675 33.920 9.050 ;
        RECT 15.750 6.080 16.750 6.125 ;
        RECT 29.315 5.285 30.455 5.315 ;
        RECT 31.500 5.285 32.500 8.675 ;
        RECT 34.255 7.125 35.255 10.325 ;
        RECT 33.055 6.125 35.255 7.125 ;
        RECT 35.675 11.370 36.045 17.350 ;
        RECT 39.875 16.925 40.875 16.955 ;
        RECT 39.875 15.925 42.645 16.925 ;
        RECT 39.875 15.895 40.875 15.925 ;
        RECT 36.900 12.825 37.900 15.275 ;
        RECT 38.375 12.825 39.320 13.350 ;
        RECT 39.600 12.825 40.600 15.275 ;
        RECT 41.075 12.825 42.020 13.350 ;
        RECT 37.395 11.700 38.435 12.175 ;
        RECT 35.675 11.325 36.675 11.370 ;
        RECT 37.395 11.325 37.900 11.700 ;
        RECT 38.745 11.325 39.320 12.825 ;
        RECT 40.095 11.700 41.135 12.175 ;
        RECT 40.095 11.325 40.600 11.700 ;
        RECT 41.445 11.325 42.020 12.825 ;
        RECT 42.985 11.325 43.355 17.350 ;
        RECT 43.775 11.325 44.145 17.350 ;
        RECT 45.685 11.325 46.055 17.350 ;
        RECT 35.675 11.300 37.900 11.325 ;
        RECT 35.675 10.355 37.920 11.300 ;
        RECT 35.675 10.325 37.900 10.355 ;
        RECT 38.280 10.325 40.600 11.325 ;
        RECT 41.025 10.325 43.355 11.325 ;
        RECT 43.730 10.325 44.820 11.325 ;
        RECT 45.050 10.325 46.055 11.325 ;
        RECT 35.675 10.280 36.675 10.325 ;
        RECT 35.675 6.125 36.045 10.280 ;
        RECT 37.395 9.950 37.900 10.325 ;
        RECT 37.395 9.455 38.435 9.950 ;
        RECT 38.745 9.050 39.320 10.325 ;
        RECT 40.095 9.950 40.600 10.325 ;
        RECT 40.095 9.455 41.135 9.950 ;
        RECT 41.445 9.050 42.020 10.325 ;
        RECT 36.900 8.675 37.955 9.050 ;
        RECT 38.375 8.675 39.320 9.050 ;
        RECT 39.600 8.675 40.655 9.050 ;
        RECT 41.075 8.675 42.020 9.050 ;
        RECT 36.900 7.800 37.900 8.675 ;
        RECT 39.600 7.800 40.600 8.675 ;
        RECT 36.900 6.800 40.600 7.800 ;
        RECT 41.175 7.125 42.175 7.170 ;
        RECT 42.355 7.125 43.355 10.325 ;
        RECT 36.900 5.285 37.900 6.800 ;
        RECT 41.175 6.125 43.355 7.125 ;
        RECT 43.775 6.125 44.145 10.325 ;
        RECT 45.055 9.325 46.055 10.325 ;
        RECT 46.475 11.325 46.845 17.350 ;
        RECT 56.900 13.825 57.900 19.970 ;
        RECT 63.500 18.675 64.500 20.050 ;
        RECT 67.025 19.975 88.300 20.155 ;
        RECT 88.925 20.050 90.850 21.050 ;
        RECT 92.450 20.155 98.375 21.075 ;
        RECT 103.550 20.155 113.725 21.075 ;
        RECT 115.275 21.050 116.275 22.025 ;
        RECT 122.075 22.005 123.025 22.025 ;
        RECT 124.855 21.730 125.855 22.825 ;
        RECT 136.675 22.025 139.880 23.025 ;
        RECT 140.655 22.025 141.745 23.025 ;
        RECT 142.495 22.025 145.775 23.025 ;
        RECT 147.475 22.025 148.475 23.025 ;
        RECT 136.700 22.005 137.650 22.025 ;
        RECT 125.130 21.115 125.580 21.730 ;
        RECT 130.025 21.075 134.225 21.080 ;
        RECT 67.740 19.970 70.250 19.975 ;
        RECT 70.440 19.970 87.565 19.975 ;
        RECT 71.170 19.050 79.230 19.970 ;
        RECT 63.480 17.725 64.520 18.675 ;
        RECT 63.500 17.700 64.500 17.725 ;
        RECT 65.255 17.700 66.345 18.700 ;
        RECT 56.900 12.825 57.925 13.825 ;
        RECT 58.400 12.825 59.345 13.350 ;
        RECT 48.855 11.875 49.305 12.515 ;
        RECT 48.575 11.325 49.575 11.875 ;
        RECT 57.420 11.700 58.460 12.175 ;
        RECT 52.750 11.325 53.750 11.355 ;
        RECT 57.420 11.325 57.925 11.700 ;
        RECT 58.770 11.370 59.345 12.825 ;
        RECT 46.475 10.325 49.575 11.325 ;
        RECT 52.700 11.300 57.925 11.325 ;
        RECT 52.700 10.350 57.945 11.300 ;
        RECT 52.700 10.325 57.925 10.350 ;
        RECT 45.010 8.325 46.100 9.325 ;
        RECT 45.685 6.125 46.055 8.325 ;
        RECT 46.475 6.125 46.845 10.325 ;
        RECT 48.855 10.205 49.305 10.325 ;
        RECT 52.750 10.295 53.750 10.325 ;
        RECT 57.420 9.950 57.925 10.325 ;
        RECT 58.350 10.280 59.350 11.370 ;
        RECT 60.310 11.325 60.680 17.350 ;
        RECT 59.675 10.325 60.680 11.325 ;
        RECT 57.420 9.455 58.460 9.950 ;
        RECT 58.770 9.050 59.345 10.280 ;
        RECT 56.925 8.675 57.980 9.050 ;
        RECT 58.400 8.675 59.345 9.050 ;
        RECT 41.175 6.080 42.175 6.125 ;
        RECT 54.740 5.285 55.880 5.315 ;
        RECT 56.925 5.285 57.925 8.675 ;
        RECT 59.680 7.125 60.680 10.325 ;
        RECT 58.480 6.125 60.680 7.125 ;
        RECT 61.100 11.370 61.470 17.350 ;
        RECT 65.300 16.925 66.300 16.955 ;
        RECT 65.300 15.925 68.070 16.925 ;
        RECT 65.300 15.895 66.300 15.925 ;
        RECT 62.325 12.825 63.325 15.275 ;
        RECT 63.800 12.825 64.745 13.350 ;
        RECT 65.025 12.825 66.025 15.275 ;
        RECT 66.500 12.825 67.445 13.350 ;
        RECT 62.820 11.700 63.860 12.175 ;
        RECT 61.100 11.325 62.100 11.370 ;
        RECT 62.820 11.325 63.325 11.700 ;
        RECT 64.170 11.325 64.745 12.825 ;
        RECT 65.520 11.700 66.560 12.175 ;
        RECT 65.520 11.325 66.025 11.700 ;
        RECT 66.870 11.325 67.445 12.825 ;
        RECT 68.410 11.325 68.780 17.350 ;
        RECT 69.200 11.325 69.570 17.350 ;
        RECT 71.110 11.325 71.480 17.350 ;
        RECT 61.100 11.300 63.325 11.325 ;
        RECT 61.100 10.355 63.345 11.300 ;
        RECT 61.100 10.325 63.325 10.355 ;
        RECT 63.705 10.325 66.025 11.325 ;
        RECT 66.450 10.325 68.780 11.325 ;
        RECT 69.155 10.325 70.245 11.325 ;
        RECT 70.475 10.325 71.480 11.325 ;
        RECT 61.100 10.280 62.100 10.325 ;
        RECT 61.100 6.125 61.470 10.280 ;
        RECT 62.820 9.950 63.325 10.325 ;
        RECT 62.820 9.455 63.860 9.950 ;
        RECT 64.170 9.050 64.745 10.325 ;
        RECT 65.520 9.950 66.025 10.325 ;
        RECT 65.520 9.455 66.560 9.950 ;
        RECT 66.870 9.050 67.445 10.325 ;
        RECT 62.325 8.675 63.380 9.050 ;
        RECT 63.800 8.675 64.745 9.050 ;
        RECT 65.025 8.675 66.080 9.050 ;
        RECT 66.500 8.675 67.445 9.050 ;
        RECT 62.325 7.800 63.325 8.675 ;
        RECT 65.025 7.800 66.025 8.675 ;
        RECT 62.325 6.800 66.025 7.800 ;
        RECT 66.600 7.125 67.600 7.170 ;
        RECT 67.780 7.125 68.780 10.325 ;
        RECT 62.325 5.285 63.325 6.800 ;
        RECT 66.600 6.125 68.780 7.125 ;
        RECT 69.200 6.125 69.570 10.325 ;
        RECT 70.480 9.325 71.480 10.325 ;
        RECT 71.900 11.325 72.270 17.350 ;
        RECT 82.325 13.825 83.325 19.970 ;
        RECT 88.925 18.675 89.925 20.050 ;
        RECT 92.450 19.975 113.725 20.155 ;
        RECT 114.350 20.050 116.275 21.050 ;
        RECT 117.875 20.155 123.800 21.075 ;
        RECT 128.975 20.155 139.150 21.075 ;
        RECT 140.700 21.050 141.700 22.025 ;
        RECT 147.500 22.005 148.450 22.025 ;
        RECT 150.280 21.730 151.280 22.825 ;
        RECT 150.555 21.115 151.005 21.730 ;
        RECT 93.165 19.970 95.675 19.975 ;
        RECT 95.865 19.970 112.990 19.975 ;
        RECT 96.595 19.050 104.655 19.970 ;
        RECT 88.905 17.725 89.945 18.675 ;
        RECT 88.925 17.700 89.925 17.725 ;
        RECT 90.680 17.700 91.770 18.700 ;
        RECT 82.325 12.825 83.350 13.825 ;
        RECT 83.825 12.825 84.770 13.350 ;
        RECT 74.280 11.875 74.730 12.515 ;
        RECT 74.000 11.325 75.000 11.875 ;
        RECT 82.845 11.700 83.885 12.175 ;
        RECT 78.175 11.325 79.175 11.355 ;
        RECT 82.845 11.325 83.350 11.700 ;
        RECT 84.195 11.370 84.770 12.825 ;
        RECT 71.900 10.325 75.000 11.325 ;
        RECT 78.125 11.300 83.350 11.325 ;
        RECT 78.125 10.350 83.370 11.300 ;
        RECT 78.125 10.325 83.350 10.350 ;
        RECT 70.435 8.325 71.525 9.325 ;
        RECT 71.110 6.125 71.480 8.325 ;
        RECT 71.900 6.125 72.270 10.325 ;
        RECT 74.280 10.205 74.730 10.325 ;
        RECT 78.175 10.295 79.175 10.325 ;
        RECT 82.845 9.950 83.350 10.325 ;
        RECT 83.775 10.280 84.775 11.370 ;
        RECT 85.735 11.325 86.105 17.350 ;
        RECT 85.100 10.325 86.105 11.325 ;
        RECT 82.845 9.455 83.885 9.950 ;
        RECT 84.195 9.050 84.770 10.280 ;
        RECT 82.350 8.675 83.405 9.050 ;
        RECT 83.825 8.675 84.770 9.050 ;
        RECT 66.600 6.080 67.600 6.125 ;
        RECT 80.165 5.285 81.305 5.315 ;
        RECT 82.350 5.285 83.350 8.675 ;
        RECT 85.105 7.125 86.105 10.325 ;
        RECT 83.905 6.125 86.105 7.125 ;
        RECT 86.525 11.370 86.895 17.350 ;
        RECT 90.725 16.925 91.725 16.955 ;
        RECT 90.725 15.925 93.495 16.925 ;
        RECT 90.725 15.895 91.725 15.925 ;
        RECT 87.750 12.825 88.750 15.275 ;
        RECT 89.225 12.825 90.170 13.350 ;
        RECT 90.450 12.825 91.450 15.275 ;
        RECT 91.925 12.825 92.870 13.350 ;
        RECT 88.245 11.700 89.285 12.175 ;
        RECT 86.525 11.325 87.525 11.370 ;
        RECT 88.245 11.325 88.750 11.700 ;
        RECT 89.595 11.325 90.170 12.825 ;
        RECT 90.945 11.700 91.985 12.175 ;
        RECT 90.945 11.325 91.450 11.700 ;
        RECT 92.295 11.325 92.870 12.825 ;
        RECT 93.835 11.325 94.205 17.350 ;
        RECT 94.625 11.325 94.995 17.350 ;
        RECT 96.535 11.325 96.905 17.350 ;
        RECT 86.525 11.300 88.750 11.325 ;
        RECT 86.525 10.355 88.770 11.300 ;
        RECT 86.525 10.325 88.750 10.355 ;
        RECT 89.130 10.325 91.450 11.325 ;
        RECT 91.875 10.325 94.205 11.325 ;
        RECT 94.580 10.325 95.670 11.325 ;
        RECT 95.900 10.325 96.905 11.325 ;
        RECT 86.525 10.280 87.525 10.325 ;
        RECT 86.525 6.125 86.895 10.280 ;
        RECT 88.245 9.950 88.750 10.325 ;
        RECT 88.245 9.455 89.285 9.950 ;
        RECT 89.595 9.050 90.170 10.325 ;
        RECT 90.945 9.950 91.450 10.325 ;
        RECT 90.945 9.455 91.985 9.950 ;
        RECT 92.295 9.050 92.870 10.325 ;
        RECT 87.750 8.675 88.805 9.050 ;
        RECT 89.225 8.675 90.170 9.050 ;
        RECT 90.450 8.675 91.505 9.050 ;
        RECT 91.925 8.675 92.870 9.050 ;
        RECT 87.750 7.800 88.750 8.675 ;
        RECT 90.450 7.800 91.450 8.675 ;
        RECT 87.750 6.800 91.450 7.800 ;
        RECT 92.025 7.125 93.025 7.170 ;
        RECT 93.205 7.125 94.205 10.325 ;
        RECT 87.750 5.285 88.750 6.800 ;
        RECT 92.025 6.125 94.205 7.125 ;
        RECT 94.625 6.125 94.995 10.325 ;
        RECT 95.905 9.325 96.905 10.325 ;
        RECT 97.325 11.325 97.695 17.350 ;
        RECT 107.750 13.825 108.750 19.970 ;
        RECT 114.350 18.675 115.350 20.050 ;
        RECT 117.875 19.975 139.150 20.155 ;
        RECT 139.775 20.050 141.700 21.050 ;
        RECT 118.590 19.970 121.100 19.975 ;
        RECT 121.290 19.970 138.415 19.975 ;
        RECT 122.020 19.050 130.080 19.970 ;
        RECT 114.330 17.725 115.370 18.675 ;
        RECT 114.350 17.700 115.350 17.725 ;
        RECT 116.105 17.700 117.195 18.700 ;
        RECT 107.750 12.825 108.775 13.825 ;
        RECT 109.250 12.825 110.195 13.350 ;
        RECT 99.705 11.875 100.155 12.515 ;
        RECT 99.425 11.325 100.425 11.875 ;
        RECT 108.270 11.700 109.310 12.175 ;
        RECT 103.600 11.325 104.600 11.355 ;
        RECT 108.270 11.325 108.775 11.700 ;
        RECT 109.620 11.370 110.195 12.825 ;
        RECT 97.325 10.325 100.425 11.325 ;
        RECT 103.550 11.300 108.775 11.325 ;
        RECT 103.550 10.350 108.795 11.300 ;
        RECT 103.550 10.325 108.775 10.350 ;
        RECT 95.860 8.325 96.950 9.325 ;
        RECT 96.535 6.125 96.905 8.325 ;
        RECT 97.325 6.125 97.695 10.325 ;
        RECT 99.705 10.205 100.155 10.325 ;
        RECT 103.600 10.295 104.600 10.325 ;
        RECT 108.270 9.950 108.775 10.325 ;
        RECT 109.200 10.280 110.200 11.370 ;
        RECT 111.160 11.325 111.530 17.350 ;
        RECT 110.525 10.325 111.530 11.325 ;
        RECT 108.270 9.455 109.310 9.950 ;
        RECT 109.620 9.050 110.195 10.280 ;
        RECT 107.775 8.675 108.830 9.050 ;
        RECT 109.250 8.675 110.195 9.050 ;
        RECT 92.025 6.080 93.025 6.125 ;
        RECT 105.590 5.285 106.730 5.315 ;
        RECT 107.775 5.285 108.775 8.675 ;
        RECT 110.530 7.125 111.530 10.325 ;
        RECT 109.330 6.125 111.530 7.125 ;
        RECT 111.950 11.370 112.320 17.350 ;
        RECT 116.150 16.925 117.150 16.955 ;
        RECT 116.150 15.925 118.920 16.925 ;
        RECT 116.150 15.895 117.150 15.925 ;
        RECT 113.175 12.825 114.175 15.275 ;
        RECT 114.650 12.825 115.595 13.350 ;
        RECT 115.875 12.825 116.875 15.275 ;
        RECT 117.350 12.825 118.295 13.350 ;
        RECT 113.670 11.700 114.710 12.175 ;
        RECT 111.950 11.325 112.950 11.370 ;
        RECT 113.670 11.325 114.175 11.700 ;
        RECT 115.020 11.325 115.595 12.825 ;
        RECT 116.370 11.700 117.410 12.175 ;
        RECT 116.370 11.325 116.875 11.700 ;
        RECT 117.720 11.325 118.295 12.825 ;
        RECT 119.260 11.325 119.630 17.350 ;
        RECT 120.050 11.325 120.420 17.350 ;
        RECT 121.960 11.325 122.330 17.350 ;
        RECT 111.950 11.300 114.175 11.325 ;
        RECT 111.950 10.355 114.195 11.300 ;
        RECT 111.950 10.325 114.175 10.355 ;
        RECT 114.555 10.325 116.875 11.325 ;
        RECT 117.300 10.325 119.630 11.325 ;
        RECT 120.005 10.325 121.095 11.325 ;
        RECT 121.325 10.325 122.330 11.325 ;
        RECT 111.950 10.280 112.950 10.325 ;
        RECT 111.950 6.125 112.320 10.280 ;
        RECT 113.670 9.950 114.175 10.325 ;
        RECT 113.670 9.455 114.710 9.950 ;
        RECT 115.020 9.050 115.595 10.325 ;
        RECT 116.370 9.950 116.875 10.325 ;
        RECT 116.370 9.455 117.410 9.950 ;
        RECT 117.720 9.050 118.295 10.325 ;
        RECT 113.175 8.675 114.230 9.050 ;
        RECT 114.650 8.675 115.595 9.050 ;
        RECT 115.875 8.675 116.930 9.050 ;
        RECT 117.350 8.675 118.295 9.050 ;
        RECT 113.175 7.800 114.175 8.675 ;
        RECT 115.875 7.800 116.875 8.675 ;
        RECT 113.175 6.800 116.875 7.800 ;
        RECT 117.450 7.125 118.450 7.170 ;
        RECT 118.630 7.125 119.630 10.325 ;
        RECT 113.175 5.285 114.175 6.800 ;
        RECT 117.450 6.125 119.630 7.125 ;
        RECT 120.050 6.125 120.420 10.325 ;
        RECT 121.330 9.325 122.330 10.325 ;
        RECT 122.750 11.325 123.120 17.350 ;
        RECT 133.175 13.825 134.175 19.970 ;
        RECT 139.775 18.675 140.775 20.050 ;
        RECT 143.300 19.975 149.225 21.075 ;
        RECT 144.015 19.970 146.525 19.975 ;
        RECT 146.715 19.970 149.215 19.975 ;
        RECT 139.755 17.725 140.795 18.675 ;
        RECT 139.775 17.700 140.775 17.725 ;
        RECT 141.530 17.700 142.620 18.700 ;
        RECT 133.175 12.825 134.200 13.825 ;
        RECT 134.675 12.825 135.620 13.350 ;
        RECT 125.130 11.875 125.580 12.515 ;
        RECT 124.850 11.325 125.850 11.875 ;
        RECT 133.695 11.700 134.735 12.175 ;
        RECT 129.025 11.325 130.025 11.355 ;
        RECT 133.695 11.325 134.200 11.700 ;
        RECT 135.045 11.370 135.620 12.825 ;
        RECT 122.750 10.325 125.850 11.325 ;
        RECT 128.975 11.300 134.200 11.325 ;
        RECT 128.975 10.350 134.220 11.300 ;
        RECT 128.975 10.325 134.200 10.350 ;
        RECT 121.285 8.325 122.375 9.325 ;
        RECT 121.960 6.125 122.330 8.325 ;
        RECT 122.750 6.125 123.120 10.325 ;
        RECT 125.130 10.205 125.580 10.325 ;
        RECT 129.025 10.295 130.025 10.325 ;
        RECT 133.695 9.950 134.200 10.325 ;
        RECT 134.625 10.280 135.625 11.370 ;
        RECT 136.585 11.325 136.955 17.350 ;
        RECT 135.950 10.325 136.955 11.325 ;
        RECT 133.695 9.455 134.735 9.950 ;
        RECT 135.045 9.050 135.620 10.280 ;
        RECT 133.200 8.675 134.255 9.050 ;
        RECT 134.675 8.675 135.620 9.050 ;
        RECT 117.450 6.080 118.450 6.125 ;
        RECT 131.015 5.285 132.155 5.315 ;
        RECT 133.200 5.285 134.200 8.675 ;
        RECT 135.955 7.125 136.955 10.325 ;
        RECT 134.755 6.125 136.955 7.125 ;
        RECT 137.375 11.370 137.745 17.350 ;
        RECT 141.575 16.925 142.575 16.955 ;
        RECT 141.575 15.925 144.345 16.925 ;
        RECT 141.575 15.895 142.575 15.925 ;
        RECT 138.600 12.825 139.600 15.275 ;
        RECT 140.075 12.825 141.020 13.350 ;
        RECT 141.300 12.825 142.300 15.275 ;
        RECT 142.775 12.825 143.720 13.350 ;
        RECT 139.095 11.700 140.135 12.175 ;
        RECT 137.375 11.325 138.375 11.370 ;
        RECT 139.095 11.325 139.600 11.700 ;
        RECT 140.445 11.325 141.020 12.825 ;
        RECT 141.795 11.700 142.835 12.175 ;
        RECT 141.795 11.325 142.300 11.700 ;
        RECT 143.145 11.325 143.720 12.825 ;
        RECT 144.685 11.325 145.055 17.350 ;
        RECT 145.475 11.325 145.845 17.350 ;
        RECT 147.385 11.325 147.755 17.350 ;
        RECT 137.375 11.300 139.600 11.325 ;
        RECT 137.375 10.355 139.620 11.300 ;
        RECT 137.375 10.325 139.600 10.355 ;
        RECT 139.980 10.325 142.300 11.325 ;
        RECT 142.725 10.325 145.055 11.325 ;
        RECT 145.430 10.325 146.520 11.325 ;
        RECT 146.750 10.325 147.755 11.325 ;
        RECT 137.375 10.280 138.375 10.325 ;
        RECT 137.375 6.125 137.745 10.280 ;
        RECT 139.095 9.950 139.600 10.325 ;
        RECT 139.095 9.455 140.135 9.950 ;
        RECT 140.445 9.050 141.020 10.325 ;
        RECT 141.795 9.950 142.300 10.325 ;
        RECT 141.795 9.455 142.835 9.950 ;
        RECT 143.145 9.050 143.720 10.325 ;
        RECT 138.600 8.675 139.655 9.050 ;
        RECT 140.075 8.675 141.020 9.050 ;
        RECT 141.300 8.675 142.355 9.050 ;
        RECT 142.775 8.675 143.720 9.050 ;
        RECT 138.600 7.800 139.600 8.675 ;
        RECT 141.300 7.800 142.300 8.675 ;
        RECT 138.600 6.800 142.300 7.800 ;
        RECT 142.875 7.125 143.875 7.170 ;
        RECT 144.055 7.125 145.055 10.325 ;
        RECT 138.600 5.285 139.600 6.800 ;
        RECT 142.875 6.125 145.055 7.125 ;
        RECT 145.475 6.125 145.845 10.325 ;
        RECT 146.755 9.325 147.755 10.325 ;
        RECT 148.175 11.325 148.545 17.350 ;
        RECT 150.555 11.875 151.005 12.515 ;
        RECT 150.275 11.325 151.275 11.875 ;
        RECT 148.175 10.325 151.275 11.325 ;
        RECT 146.710 8.325 147.800 9.325 ;
        RECT 147.385 6.125 147.755 8.325 ;
        RECT 148.175 6.125 148.545 10.325 ;
        RECT 150.555 10.205 151.005 10.325 ;
        RECT 142.875 6.080 143.875 6.125 ;
        RECT 1.850 5.275 14.575 5.285 ;
        RECT 15.350 5.275 19.390 5.285 ;
        RECT 19.590 5.275 40.000 5.285 ;
        RECT 40.775 5.275 44.815 5.285 ;
        RECT 45.015 5.275 65.425 5.285 ;
        RECT 66.200 5.275 70.240 5.285 ;
        RECT 70.440 5.275 90.850 5.285 ;
        RECT 91.625 5.275 95.665 5.285 ;
        RECT 95.865 5.275 116.275 5.285 ;
        RECT 117.050 5.275 121.090 5.285 ;
        RECT 121.290 5.275 141.700 5.285 ;
        RECT 142.475 5.275 146.515 5.285 ;
        RECT 146.715 5.275 151.360 5.285 ;
        RECT 1.850 4.175 151.360 5.275 ;
        RECT 1.850 4.170 19.390 4.175 ;
        RECT 19.590 4.170 44.815 4.175 ;
        RECT 45.015 4.170 70.240 4.175 ;
        RECT 70.440 4.170 95.665 4.175 ;
        RECT 95.865 4.170 121.090 4.175 ;
        RECT 121.290 4.170 146.515 4.175 ;
        RECT 146.715 4.170 151.360 4.175 ;
        RECT 3.890 4.140 5.030 4.170 ;
        RECT 29.315 4.140 30.455 4.170 ;
        RECT 54.740 4.140 55.880 4.170 ;
        RECT 80.165 4.140 81.305 4.170 ;
        RECT 105.590 4.140 106.730 4.170 ;
        RECT 131.015 4.140 132.155 4.170 ;
        RECT 19.370 3.225 21.325 3.245 ;
        RECT 44.795 3.225 46.750 3.245 ;
        RECT 70.220 3.225 72.175 3.245 ;
        RECT 95.645 3.225 97.600 3.245 ;
        RECT 121.070 3.225 123.025 3.245 ;
        RECT 146.495 3.225 148.450 3.245 ;
        RECT 9.550 3.200 10.550 3.225 ;
        RECT 15.750 3.200 16.750 3.225 ;
        RECT 17.650 3.200 18.650 3.225 ;
        RECT 9.530 2.250 10.570 3.200 ;
        RECT 15.730 2.250 16.770 3.200 ;
        RECT 17.630 2.250 18.670 3.200 ;
        RECT 9.550 2.225 10.550 2.250 ;
        RECT 15.750 2.225 16.750 2.250 ;
        RECT 17.650 2.225 18.650 2.250 ;
        RECT 19.365 2.225 21.350 3.225 ;
        RECT 34.975 3.200 35.975 3.225 ;
        RECT 41.175 3.200 42.175 3.225 ;
        RECT 43.075 3.200 44.075 3.225 ;
        RECT 34.955 2.250 35.995 3.200 ;
        RECT 41.155 2.250 42.195 3.200 ;
        RECT 43.055 2.250 44.095 3.200 ;
        RECT 34.975 2.225 35.975 2.250 ;
        RECT 41.175 2.225 42.175 2.250 ;
        RECT 43.075 2.225 44.075 2.250 ;
        RECT 44.790 2.225 46.775 3.225 ;
        RECT 60.400 3.200 61.400 3.225 ;
        RECT 66.600 3.200 67.600 3.225 ;
        RECT 68.500 3.200 69.500 3.225 ;
        RECT 60.380 2.250 61.420 3.200 ;
        RECT 66.580 2.250 67.620 3.200 ;
        RECT 68.480 2.250 69.520 3.200 ;
        RECT 60.400 2.225 61.400 2.250 ;
        RECT 66.600 2.225 67.600 2.250 ;
        RECT 68.500 2.225 69.500 2.250 ;
        RECT 70.215 2.225 72.200 3.225 ;
        RECT 85.825 3.200 86.825 3.225 ;
        RECT 92.025 3.200 93.025 3.225 ;
        RECT 93.925 3.200 94.925 3.225 ;
        RECT 85.805 2.250 86.845 3.200 ;
        RECT 92.005 2.250 93.045 3.200 ;
        RECT 93.905 2.250 94.945 3.200 ;
        RECT 85.825 2.225 86.825 2.250 ;
        RECT 92.025 2.225 93.025 2.250 ;
        RECT 93.925 2.225 94.925 2.250 ;
        RECT 95.640 2.225 97.625 3.225 ;
        RECT 111.250 3.200 112.250 3.225 ;
        RECT 117.450 3.200 118.450 3.225 ;
        RECT 119.350 3.200 120.350 3.225 ;
        RECT 111.230 2.250 112.270 3.200 ;
        RECT 117.430 2.250 118.470 3.200 ;
        RECT 119.330 2.250 120.370 3.200 ;
        RECT 111.250 2.225 112.250 2.250 ;
        RECT 117.450 2.225 118.450 2.250 ;
        RECT 119.350 2.225 120.350 2.250 ;
        RECT 121.065 2.225 123.050 3.225 ;
        RECT 136.675 3.200 137.675 3.225 ;
        RECT 142.875 3.200 143.875 3.225 ;
        RECT 144.775 3.200 145.775 3.225 ;
        RECT 136.655 2.250 137.695 3.200 ;
        RECT 142.855 2.250 143.895 3.200 ;
        RECT 144.755 2.250 145.795 3.200 ;
        RECT 136.675 2.225 137.675 2.250 ;
        RECT 142.875 2.225 143.875 2.250 ;
        RECT 144.775 2.225 145.775 2.250 ;
        RECT 146.490 2.225 148.475 3.225 ;
        RECT 19.370 2.205 21.325 2.225 ;
        RECT 44.795 2.205 46.750 2.225 ;
        RECT 70.220 2.205 72.175 2.225 ;
        RECT 95.645 2.205 97.600 2.225 ;
        RECT 121.070 2.205 123.025 2.225 ;
        RECT 146.495 2.205 148.450 2.225 ;
        RECT 48.680 0.950 49.580 0.995 ;
        RECT 156.435 0.950 157.285 0.970 ;
        RECT 48.680 0.050 157.310 0.950 ;
        RECT 48.680 0.005 49.580 0.050 ;
        RECT 156.435 0.030 157.285 0.050 ;
      LAYER met3 ;
        RECT 21.400 224.300 93.005 225.300 ;
        RECT 5.780 216.550 6.770 216.575 ;
        RECT 5.775 215.550 6.775 216.550 ;
        RECT 7.780 216.545 8.770 216.570 ;
        RECT 9.780 216.550 10.770 216.575 ;
        RECT 5.780 215.525 6.770 215.550 ;
        RECT 7.775 215.545 8.775 216.545 ;
        RECT 9.775 215.550 10.775 216.550 ;
        RECT 21.400 215.550 22.400 224.300 ;
        RECT 95.650 223.550 96.650 225.330 ;
        RECT 25.400 222.550 96.650 223.550 ;
        RECT 25.400 216.545 26.400 222.550 ;
        RECT 99.300 221.800 100.300 225.330 ;
        RECT 48.825 220.800 100.300 221.800 ;
        RECT 33.205 216.550 34.195 216.575 ;
        RECT 35.205 216.550 36.195 216.575 ;
        RECT 31.200 216.545 32.200 216.550 ;
        RECT 25.375 215.555 26.425 216.545 ;
        RECT 31.175 215.555 32.225 216.545 ;
        RECT 25.400 215.550 26.400 215.555 ;
        RECT 31.200 215.550 32.200 215.555 ;
        RECT 33.200 215.550 34.200 216.550 ;
        RECT 35.200 215.550 36.200 216.550 ;
        RECT 48.825 216.545 49.825 220.800 ;
        RECT 103.000 220.050 104.000 225.330 ;
        RECT 72.250 219.050 104.000 220.050 ;
        RECT 56.630 216.550 57.620 216.575 ;
        RECT 48.800 215.555 49.850 216.545 ;
        RECT 48.825 215.550 49.825 215.555 ;
        RECT 56.625 215.550 57.625 216.550 ;
        RECT 58.630 216.545 59.620 216.570 ;
        RECT 60.630 216.550 61.620 216.575 ;
        RECT 7.780 215.520 8.770 215.545 ;
        RECT 9.780 215.525 10.770 215.550 ;
        RECT 21.405 215.525 22.395 215.550 ;
        RECT 33.205 215.525 34.195 215.550 ;
        RECT 35.205 215.525 36.195 215.550 ;
        RECT 56.630 215.525 57.620 215.550 ;
        RECT 58.625 215.545 59.625 216.545 ;
        RECT 60.625 215.550 61.625 216.550 ;
        RECT 72.250 216.545 73.250 219.050 ;
        RECT 106.675 218.300 107.675 225.330 ;
        RECT 76.250 217.300 107.675 218.300 ;
        RECT 110.375 217.300 111.375 225.330 ;
        RECT 114.050 218.300 115.050 225.330 ;
        RECT 117.725 220.050 118.725 225.330 ;
        RECT 121.425 221.825 122.425 225.330 ;
        RECT 125.075 221.825 126.075 225.330 ;
        RECT 128.775 221.825 129.775 225.330 ;
        RECT 132.450 221.825 133.450 225.330 ;
        RECT 136.125 223.575 137.125 225.330 ;
        RECT 139.775 224.245 140.825 225.355 ;
        RECT 134.875 222.550 137.125 223.575 ;
        RECT 134.875 222.525 135.925 222.550 ;
        RECT 121.400 220.775 122.450 221.825 ;
        RECT 125.050 220.775 126.100 221.825 ;
        RECT 128.750 220.775 129.800 221.825 ;
        RECT 132.450 220.800 133.925 221.825 ;
        RECT 132.875 220.775 133.925 220.800 ;
        RECT 117.725 219.050 128.100 220.050 ;
        RECT 114.050 217.300 124.100 218.300 ;
        RECT 76.250 216.545 77.250 217.300 ;
        RECT 110.380 217.275 111.370 217.300 ;
        RECT 84.055 216.550 85.045 216.575 ;
        RECT 86.055 216.550 87.045 216.575 ;
        RECT 107.480 216.550 108.470 216.575 ;
        RECT 82.050 216.545 83.050 216.550 ;
        RECT 72.225 215.555 73.275 216.545 ;
        RECT 76.225 215.555 77.275 216.545 ;
        RECT 82.025 215.555 83.075 216.545 ;
        RECT 72.250 215.550 73.250 215.555 ;
        RECT 76.250 215.550 77.250 215.555 ;
        RECT 82.050 215.550 83.050 215.555 ;
        RECT 84.050 215.550 85.050 216.550 ;
        RECT 86.050 215.550 87.050 216.550 ;
        RECT 107.475 215.550 108.475 216.550 ;
        RECT 109.480 216.545 110.470 216.570 ;
        RECT 111.480 216.550 112.470 216.575 ;
        RECT 123.100 216.570 124.100 217.300 ;
        RECT 58.630 215.520 59.620 215.545 ;
        RECT 60.630 215.525 61.620 215.550 ;
        RECT 84.055 215.525 85.045 215.550 ;
        RECT 86.055 215.525 87.045 215.550 ;
        RECT 107.480 215.525 108.470 215.550 ;
        RECT 109.475 215.545 110.475 216.545 ;
        RECT 111.475 215.550 112.475 216.550 ;
        RECT 123.075 215.580 124.125 216.570 ;
        RECT 127.100 216.545 128.100 219.050 ;
        RECT 134.905 216.550 135.895 216.575 ;
        RECT 136.905 216.550 137.895 216.575 ;
        RECT 143.475 216.550 144.475 225.330 ;
        RECT 147.150 218.300 148.150 225.330 ;
        RECT 150.850 220.050 151.850 225.330 ;
        RECT 154.500 221.800 155.500 225.330 ;
        RECT 154.500 220.800 157.525 221.800 ;
        RECT 150.850 219.050 155.525 220.050 ;
        RECT 147.150 217.300 153.525 218.300 ;
        RECT 132.900 216.545 133.900 216.550 ;
        RECT 123.100 215.575 124.100 215.580 ;
        RECT 127.075 215.555 128.125 216.545 ;
        RECT 132.875 215.555 133.925 216.545 ;
        RECT 127.100 215.550 128.100 215.555 ;
        RECT 132.900 215.550 133.900 215.555 ;
        RECT 134.900 215.550 135.900 216.550 ;
        RECT 136.900 215.550 137.900 216.550 ;
        RECT 143.475 216.545 151.525 216.550 ;
        RECT 152.525 216.545 153.525 217.300 ;
        RECT 154.525 216.545 155.525 219.050 ;
        RECT 156.525 216.545 157.525 220.800 ;
        RECT 143.475 215.555 151.550 216.545 ;
        RECT 152.500 215.555 153.550 216.545 ;
        RECT 154.500 215.555 155.550 216.545 ;
        RECT 156.500 215.555 157.550 216.545 ;
        RECT 143.475 215.550 151.525 215.555 ;
        RECT 152.525 215.550 153.525 215.555 ;
        RECT 154.525 215.550 155.525 215.555 ;
        RECT 156.525 215.550 157.525 215.555 ;
        RECT 109.480 215.520 110.470 215.545 ;
        RECT 111.480 215.525 112.470 215.550 ;
        RECT 134.905 215.525 135.895 215.550 ;
        RECT 136.905 215.525 137.895 215.550 ;
        RECT 150.530 214.550 151.520 214.575 ;
        RECT 13.550 212.175 14.600 212.200 ;
        RECT 7.500 211.175 10.550 212.175 ;
        RECT 13.550 211.175 21.350 212.175 ;
        RECT 23.520 211.200 24.520 214.550 ;
        RECT 38.975 212.175 40.025 212.200 ;
        RECT 64.400 212.175 65.450 212.200 ;
        RECT 2.805 210.225 3.920 210.255 ;
        RECT 5.970 210.225 7.125 210.250 ;
        RECT 2.805 209.120 7.125 210.225 ;
        RECT 2.805 209.090 3.920 209.120 ;
        RECT 5.970 209.095 7.125 209.120 ;
        RECT 5.995 205.755 7.100 209.095 ;
        RECT 3.900 204.650 7.100 205.755 ;
        RECT 3.900 187.680 5.005 204.650 ;
        RECT 7.500 200.500 8.500 211.175 ;
        RECT 13.550 211.150 14.600 211.175 ;
        RECT 10.250 210.195 14.575 210.200 ;
        RECT 10.250 209.200 19.345 210.195 ;
        RECT 23.495 210.150 24.545 211.200 ;
        RECT 32.925 211.175 35.975 212.175 ;
        RECT 38.975 211.175 46.775 212.175 ;
        RECT 58.350 211.175 61.400 212.175 ;
        RECT 64.400 211.175 72.200 212.175 ;
        RECT 74.370 211.200 75.370 214.550 ;
        RECT 89.825 212.175 90.875 212.200 ;
        RECT 115.250 212.175 116.300 212.200 ;
        RECT 26.220 210.295 27.270 210.320 ;
        RECT 25.400 210.290 27.270 210.295 ;
        RECT 25.375 209.300 27.270 210.290 ;
        RECT 25.400 209.295 27.270 209.300 ;
        RECT 26.220 209.270 27.270 209.295 ;
        RECT 10.250 200.500 11.250 209.200 ;
        RECT 14.425 207.850 15.475 207.875 ;
        RECT 16.150 207.850 17.200 208.365 ;
        RECT 12.325 206.850 13.650 207.850 ;
        RECT 14.425 206.850 17.200 207.850 ;
        RECT 12.325 200.500 13.325 206.850 ;
        RECT 14.425 206.825 15.475 206.850 ;
        RECT 6.075 198.200 7.075 200.475 ;
        RECT 7.475 199.450 8.525 200.500 ;
        RECT 10.225 199.450 11.275 200.500 ;
        RECT 12.325 199.475 13.925 200.500 ;
        RECT 12.875 199.450 13.925 199.475 ;
        RECT 14.450 198.200 15.450 206.825 ;
        RECT 16.150 205.050 17.200 206.100 ;
        RECT 6.075 197.200 15.450 198.200 ;
        RECT 16.175 198.200 17.175 205.050 ;
        RECT 18.350 204.795 19.345 209.200 ;
        RECT 28.110 208.420 30.670 209.525 ;
        RECT 31.395 209.095 32.550 210.250 ;
        RECT 20.345 205.155 21.345 208.340 ;
        RECT 28.110 207.695 29.215 208.420 ;
        RECT 24.815 206.590 29.215 207.695 ;
        RECT 24.815 205.180 25.920 206.590 ;
        RECT 28.230 205.755 29.345 205.785 ;
        RECT 31.420 205.755 32.525 209.095 ;
        RECT 24.795 205.155 25.950 205.180 ;
        RECT 18.350 204.055 19.350 204.795 ;
        RECT 20.345 204.100 25.950 205.155 ;
        RECT 28.230 204.650 32.525 205.755 ;
        RECT 28.230 204.620 30.430 204.650 ;
        RECT 18.355 200.500 19.350 204.055 ;
        RECT 20.370 204.050 25.950 204.100 ;
        RECT 24.795 204.025 25.950 204.050 ;
        RECT 18.325 199.450 19.375 200.500 ;
        RECT 23.405 200.480 24.395 200.505 ;
        RECT 23.400 199.480 24.400 200.480 ;
        RECT 23.405 199.455 24.395 199.480 ;
        RECT 16.175 197.200 18.650 198.200 ;
        RECT 7.650 196.275 8.700 196.300 ;
        RECT 6.070 195.275 8.700 196.275 ;
        RECT 7.650 195.250 8.700 195.275 ;
        RECT 7.675 191.000 8.675 195.250 ;
        RECT 9.550 191.375 10.550 197.200 ;
        RECT 15.725 195.250 16.775 196.300 ;
        RECT 13.550 193.350 14.600 194.430 ;
        RECT 15.750 192.375 16.750 195.250 ;
        RECT 15.720 191.375 16.780 192.375 ;
        RECT 17.650 191.375 18.650 197.200 ;
        RECT 19.625 197.000 24.150 198.000 ;
        RECT 19.350 192.375 20.340 192.400 ;
        RECT 19.345 191.375 20.345 192.375 ;
        RECT 19.350 191.350 20.340 191.375 ;
        RECT 7.675 190.995 10.775 191.000 ;
        RECT 7.675 190.005 10.800 190.995 ;
        RECT 7.675 190.000 10.775 190.005 ;
        RECT 13.550 189.600 14.600 189.625 ;
        RECT 7.500 188.600 10.550 189.600 ;
        RECT 13.550 188.600 21.350 189.600 ;
        RECT 2.805 186.525 5.030 187.680 ;
        RECT 2.805 186.515 5.005 186.525 ;
        RECT 3.900 165.105 5.005 186.515 ;
        RECT 7.500 177.925 8.500 188.600 ;
        RECT 13.550 188.575 14.600 188.600 ;
        RECT 10.250 187.620 14.575 187.625 ;
        RECT 10.250 186.625 19.345 187.620 ;
        RECT 10.250 177.925 11.250 186.625 ;
        RECT 12.325 184.275 13.650 185.275 ;
        RECT 12.325 177.925 13.325 184.275 ;
        RECT 14.425 184.250 15.475 185.300 ;
        RECT 6.075 175.625 7.075 177.900 ;
        RECT 7.475 176.875 8.525 177.925 ;
        RECT 10.225 176.875 11.275 177.925 ;
        RECT 12.325 176.900 13.925 177.925 ;
        RECT 12.875 176.875 13.925 176.900 ;
        RECT 14.450 175.625 15.450 184.250 ;
        RECT 16.150 182.475 17.200 183.525 ;
        RECT 6.075 174.625 15.450 175.625 ;
        RECT 16.175 175.625 17.175 182.475 ;
        RECT 18.350 182.220 19.345 186.625 ;
        RECT 18.350 181.480 19.350 182.220 ;
        RECT 18.355 177.925 19.350 181.480 ;
        RECT 18.325 176.875 19.375 177.925 ;
        RECT 21.405 177.905 22.395 177.930 ;
        RECT 21.400 176.905 22.400 177.905 ;
        RECT 21.405 176.880 22.395 176.905 ;
        RECT 23.150 175.925 24.150 197.000 ;
        RECT 29.325 187.680 30.430 204.620 ;
        RECT 32.925 200.500 33.925 211.175 ;
        RECT 38.975 211.150 40.025 211.175 ;
        RECT 53.655 210.225 54.770 210.255 ;
        RECT 56.820 210.225 57.975 210.250 ;
        RECT 35.675 210.195 40.000 210.200 ;
        RECT 35.675 209.200 44.770 210.195 ;
        RECT 35.675 200.500 36.675 209.200 ;
        RECT 37.750 206.850 39.075 207.850 ;
        RECT 37.750 200.500 38.750 206.850 ;
        RECT 39.850 206.825 40.900 207.875 ;
        RECT 31.500 198.200 32.500 200.475 ;
        RECT 32.900 199.450 33.950 200.500 ;
        RECT 35.650 199.450 36.700 200.500 ;
        RECT 37.750 199.475 39.350 200.500 ;
        RECT 38.300 199.450 39.350 199.475 ;
        RECT 39.875 198.200 40.875 206.825 ;
        RECT 41.575 205.050 42.625 206.100 ;
        RECT 31.500 197.200 40.875 198.200 ;
        RECT 41.600 198.200 42.600 205.050 ;
        RECT 43.775 204.795 44.770 209.200 ;
        RECT 53.655 209.120 57.975 210.225 ;
        RECT 53.655 209.090 54.770 209.120 ;
        RECT 56.820 209.095 57.975 209.120 ;
        RECT 56.845 205.755 57.950 209.095 ;
        RECT 43.775 204.055 44.775 204.795 ;
        RECT 43.780 200.500 44.775 204.055 ;
        RECT 54.750 204.650 57.950 205.755 ;
        RECT 43.750 199.450 44.800 200.500 ;
        RECT 41.600 197.200 44.075 198.200 ;
        RECT 33.075 196.275 34.125 196.300 ;
        RECT 31.495 195.275 34.125 196.275 ;
        RECT 33.075 195.250 34.125 195.275 ;
        RECT 33.100 191.000 34.100 195.250 ;
        RECT 34.975 191.375 35.975 197.200 ;
        RECT 41.150 195.250 42.200 196.300 ;
        RECT 38.975 193.350 40.025 194.430 ;
        RECT 41.175 192.375 42.175 195.250 ;
        RECT 41.145 191.375 42.205 192.375 ;
        RECT 43.075 191.375 44.075 197.200 ;
        RECT 45.050 197.000 49.575 198.000 ;
        RECT 44.775 192.375 45.765 192.400 ;
        RECT 44.770 191.375 45.770 192.375 ;
        RECT 44.775 191.350 45.765 191.375 ;
        RECT 33.100 190.995 36.200 191.000 ;
        RECT 33.100 190.005 36.225 190.995 ;
        RECT 33.100 190.000 36.200 190.005 ;
        RECT 38.975 189.600 40.025 189.625 ;
        RECT 32.925 188.600 35.975 189.600 ;
        RECT 38.975 188.600 46.775 189.600 ;
        RECT 28.230 186.525 30.455 187.680 ;
        RECT 28.230 186.515 30.430 186.525 ;
        RECT 16.175 174.625 18.650 175.625 ;
        RECT 19.625 174.925 26.250 175.925 ;
        RECT 7.775 173.725 8.775 173.730 ;
        RECT 7.650 173.700 8.775 173.725 ;
        RECT 6.070 172.700 8.775 173.700 ;
        RECT 7.650 172.675 8.775 172.700 ;
        RECT 7.775 172.670 8.775 172.675 ;
        RECT 9.550 168.800 10.550 174.625 ;
        RECT 15.725 172.675 16.775 173.725 ;
        RECT 13.550 170.775 14.600 171.855 ;
        RECT 15.750 169.800 16.750 172.675 ;
        RECT 15.720 168.800 16.780 169.800 ;
        RECT 17.650 168.800 18.650 174.625 ;
        RECT 19.350 169.800 20.340 169.825 ;
        RECT 19.345 168.800 20.345 169.800 ;
        RECT 19.350 168.775 20.340 168.800 ;
        RECT 13.550 167.025 14.600 167.050 ;
        RECT 7.500 166.025 10.550 167.025 ;
        RECT 13.550 166.025 21.350 167.025 ;
        RECT 23.155 166.800 24.155 173.800 ;
        RECT 3.875 165.080 5.030 165.105 ;
        RECT 3.870 163.975 5.030 165.080 ;
        RECT 3.875 163.950 5.030 163.975 ;
        RECT 7.500 155.350 8.500 166.025 ;
        RECT 13.550 166.000 14.600 166.025 ;
        RECT 23.130 165.750 24.180 166.800 ;
        RECT 10.250 165.045 14.575 165.050 ;
        RECT 10.250 164.050 19.345 165.045 ;
        RECT 25.250 164.575 26.250 174.925 ;
        RECT 29.325 165.105 30.430 186.515 ;
        RECT 32.925 177.925 33.925 188.600 ;
        RECT 38.975 188.575 40.025 188.600 ;
        RECT 35.675 187.620 40.000 187.625 ;
        RECT 35.675 186.625 44.770 187.620 ;
        RECT 35.675 177.925 36.675 186.625 ;
        RECT 37.750 184.275 39.075 185.275 ;
        RECT 37.750 177.925 38.750 184.275 ;
        RECT 39.850 184.250 40.900 185.300 ;
        RECT 31.500 175.625 32.500 177.900 ;
        RECT 32.900 176.875 33.950 177.925 ;
        RECT 35.650 176.875 36.700 177.925 ;
        RECT 37.750 176.900 39.350 177.925 ;
        RECT 38.300 176.875 39.350 176.900 ;
        RECT 39.875 175.625 40.875 184.250 ;
        RECT 41.575 182.475 42.625 183.525 ;
        RECT 31.500 174.625 40.875 175.625 ;
        RECT 41.600 175.625 42.600 182.475 ;
        RECT 43.775 182.220 44.770 186.625 ;
        RECT 43.775 181.480 44.775 182.220 ;
        RECT 43.780 177.925 44.775 181.480 ;
        RECT 43.750 176.875 44.800 177.925 ;
        RECT 48.575 175.925 49.575 197.000 ;
        RECT 54.750 187.680 55.855 204.650 ;
        RECT 58.350 200.500 59.350 211.175 ;
        RECT 64.400 211.150 65.450 211.175 ;
        RECT 61.100 210.195 65.425 210.200 ;
        RECT 61.100 209.200 70.195 210.195 ;
        RECT 74.345 210.150 75.395 211.200 ;
        RECT 83.775 211.175 86.825 212.175 ;
        RECT 89.825 211.175 97.625 212.175 ;
        RECT 109.200 211.175 112.250 212.175 ;
        RECT 115.250 211.175 123.050 212.175 ;
        RECT 125.220 211.200 126.220 214.550 ;
        RECT 150.525 213.550 151.525 214.550 ;
        RECT 150.530 213.525 151.520 213.550 ;
        RECT 140.675 212.175 141.725 212.200 ;
        RECT 77.070 210.295 78.120 210.320 ;
        RECT 76.250 210.290 78.120 210.295 ;
        RECT 76.225 209.300 78.120 210.290 ;
        RECT 76.250 209.295 78.120 209.300 ;
        RECT 77.070 209.270 78.120 209.295 ;
        RECT 61.100 200.500 62.100 209.200 ;
        RECT 65.275 207.850 66.325 207.875 ;
        RECT 67.000 207.850 68.050 208.365 ;
        RECT 63.175 206.850 64.500 207.850 ;
        RECT 65.275 206.850 68.050 207.850 ;
        RECT 63.175 200.500 64.175 206.850 ;
        RECT 65.275 206.825 66.325 206.850 ;
        RECT 56.925 198.200 57.925 200.475 ;
        RECT 58.325 199.450 59.375 200.500 ;
        RECT 61.075 199.450 62.125 200.500 ;
        RECT 63.175 199.475 64.775 200.500 ;
        RECT 63.725 199.450 64.775 199.475 ;
        RECT 65.300 198.200 66.300 206.825 ;
        RECT 67.000 205.050 68.050 206.100 ;
        RECT 56.925 197.200 66.300 198.200 ;
        RECT 67.025 198.200 68.025 205.050 ;
        RECT 69.200 204.795 70.195 209.200 ;
        RECT 78.960 208.420 81.520 209.525 ;
        RECT 82.245 209.095 83.400 210.250 ;
        RECT 71.195 205.155 72.195 208.340 ;
        RECT 78.960 207.695 80.065 208.420 ;
        RECT 75.665 206.590 80.065 207.695 ;
        RECT 75.665 205.180 76.770 206.590 ;
        RECT 79.080 205.755 80.195 205.785 ;
        RECT 82.270 205.755 83.375 209.095 ;
        RECT 75.645 205.155 76.800 205.180 ;
        RECT 69.200 204.055 70.200 204.795 ;
        RECT 71.195 204.100 76.800 205.155 ;
        RECT 79.080 204.650 83.375 205.755 ;
        RECT 79.080 204.620 81.280 204.650 ;
        RECT 69.205 200.500 70.200 204.055 ;
        RECT 71.220 204.050 76.800 204.100 ;
        RECT 75.645 204.025 76.800 204.050 ;
        RECT 69.175 199.450 70.225 200.500 ;
        RECT 74.255 200.480 75.245 200.505 ;
        RECT 74.250 199.480 75.250 200.480 ;
        RECT 74.255 199.455 75.245 199.480 ;
        RECT 67.025 197.200 69.500 198.200 ;
        RECT 58.500 196.275 59.550 196.300 ;
        RECT 56.920 195.275 59.550 196.275 ;
        RECT 58.500 195.250 59.550 195.275 ;
        RECT 58.525 191.000 59.525 195.250 ;
        RECT 60.400 191.375 61.400 197.200 ;
        RECT 66.575 195.250 67.625 196.300 ;
        RECT 64.400 193.350 65.450 194.430 ;
        RECT 66.600 192.375 67.600 195.250 ;
        RECT 66.570 191.375 67.630 192.375 ;
        RECT 68.500 191.375 69.500 197.200 ;
        RECT 70.475 197.000 75.000 198.000 ;
        RECT 70.200 192.375 71.190 192.400 ;
        RECT 70.195 191.375 71.195 192.375 ;
        RECT 70.200 191.350 71.190 191.375 ;
        RECT 58.525 190.995 61.625 191.000 ;
        RECT 58.525 190.005 61.650 190.995 ;
        RECT 58.525 190.000 61.625 190.005 ;
        RECT 64.400 189.600 65.450 189.625 ;
        RECT 58.350 188.600 61.400 189.600 ;
        RECT 64.400 188.600 72.200 189.600 ;
        RECT 53.655 186.525 55.880 187.680 ;
        RECT 53.655 186.515 55.855 186.525 ;
        RECT 50.650 177.900 51.700 177.925 ;
        RECT 50.650 176.900 53.750 177.900 ;
        RECT 50.650 176.875 51.700 176.900 ;
        RECT 41.600 174.625 44.075 175.625 ;
        RECT 45.050 174.925 51.675 175.925 ;
        RECT 33.200 173.725 34.200 173.730 ;
        RECT 33.075 173.700 34.200 173.725 ;
        RECT 31.495 172.700 34.200 173.700 ;
        RECT 33.075 172.675 34.200 172.700 ;
        RECT 33.200 172.670 34.200 172.675 ;
        RECT 34.975 168.800 35.975 174.625 ;
        RECT 41.150 172.675 42.200 173.725 ;
        RECT 38.975 170.775 40.025 171.855 ;
        RECT 41.175 169.800 42.175 172.675 ;
        RECT 41.145 168.800 42.205 169.800 ;
        RECT 43.075 168.800 44.075 174.625 ;
        RECT 44.775 169.800 45.765 169.825 ;
        RECT 44.770 168.800 45.770 169.800 ;
        RECT 44.775 168.775 45.765 168.800 ;
        RECT 38.975 167.025 40.025 167.050 ;
        RECT 32.925 166.025 35.975 167.025 ;
        RECT 38.975 166.025 46.775 167.025 ;
        RECT 48.580 166.800 49.580 173.800 ;
        RECT 10.250 155.350 11.250 164.050 ;
        RECT 12.325 161.700 13.650 162.700 ;
        RECT 12.325 155.350 13.325 161.700 ;
        RECT 14.425 161.675 15.475 162.725 ;
        RECT 6.075 153.050 7.075 155.325 ;
        RECT 7.475 154.300 8.525 155.350 ;
        RECT 10.225 154.300 11.275 155.350 ;
        RECT 12.325 154.325 13.925 155.350 ;
        RECT 12.875 154.300 13.925 154.325 ;
        RECT 14.450 153.050 15.450 161.675 ;
        RECT 16.150 159.900 17.200 160.950 ;
        RECT 6.075 152.050 15.450 153.050 ;
        RECT 16.175 153.050 17.175 159.900 ;
        RECT 18.350 159.645 19.345 164.050 ;
        RECT 23.200 163.575 26.250 164.575 ;
        RECT 28.230 163.950 30.455 165.105 ;
        RECT 28.230 163.940 29.345 163.950 ;
        RECT 18.350 158.905 19.350 159.645 ;
        RECT 18.355 155.350 19.350 158.905 ;
        RECT 18.325 154.300 19.375 155.350 ;
        RECT 19.605 153.325 20.655 153.350 ;
        RECT 23.200 153.325 24.200 163.575 ;
        RECT 32.925 155.350 33.925 166.025 ;
        RECT 38.975 166.000 40.025 166.025 ;
        RECT 48.555 165.750 49.605 166.800 ;
        RECT 35.675 165.045 40.000 165.050 ;
        RECT 35.675 164.050 44.770 165.045 ;
        RECT 50.675 164.575 51.675 174.925 ;
        RECT 35.675 155.350 36.675 164.050 ;
        RECT 37.750 161.700 39.075 162.700 ;
        RECT 37.750 155.350 38.750 161.700 ;
        RECT 39.850 161.675 40.900 162.725 ;
        RECT 16.175 152.050 18.650 153.050 ;
        RECT 19.605 152.325 24.200 153.325 ;
        RECT 31.500 153.050 32.500 155.325 ;
        RECT 32.900 154.300 33.950 155.350 ;
        RECT 35.650 154.300 36.700 155.350 ;
        RECT 37.750 154.325 39.350 155.350 ;
        RECT 38.300 154.300 39.350 154.325 ;
        RECT 39.875 153.050 40.875 161.675 ;
        RECT 41.575 159.900 42.625 160.950 ;
        RECT 19.605 152.300 20.655 152.325 ;
        RECT 6.080 151.125 7.070 151.150 ;
        RECT 7.650 151.125 8.700 151.150 ;
        RECT 6.070 150.125 8.700 151.125 ;
        RECT 6.080 150.100 7.070 150.125 ;
        RECT 7.650 150.100 8.700 150.125 ;
        RECT 9.550 146.225 10.550 152.050 ;
        RECT 15.725 150.100 16.775 151.150 ;
        RECT 13.550 148.200 14.600 149.280 ;
        RECT 15.750 147.225 16.750 150.100 ;
        RECT 15.720 146.225 16.780 147.225 ;
        RECT 17.650 146.225 18.650 152.050 ;
        RECT 19.350 147.225 20.340 147.250 ;
        RECT 19.345 146.225 20.345 147.225 ;
        RECT 19.350 146.200 20.340 146.225 ;
        RECT 21.405 145.000 22.395 145.025 ;
        RECT 23.170 145.000 24.170 152.325 ;
        RECT 31.500 152.050 40.875 153.050 ;
        RECT 41.600 153.050 42.600 159.900 ;
        RECT 43.775 159.645 44.770 164.050 ;
        RECT 48.625 163.575 51.675 164.575 ;
        RECT 43.775 158.905 44.775 159.645 ;
        RECT 43.780 155.350 44.775 158.905 ;
        RECT 43.750 154.300 44.800 155.350 ;
        RECT 45.030 153.325 46.080 153.350 ;
        RECT 48.625 153.325 49.625 163.575 ;
        RECT 41.600 152.050 44.075 153.050 ;
        RECT 45.030 152.325 49.625 153.325 ;
        RECT 45.030 152.300 46.080 152.325 ;
        RECT 31.505 151.125 32.495 151.150 ;
        RECT 33.075 151.125 34.125 151.150 ;
        RECT 31.495 150.125 34.125 151.125 ;
        RECT 31.505 150.100 32.495 150.125 ;
        RECT 33.075 150.100 34.125 150.125 ;
        RECT 34.975 146.225 35.975 152.050 ;
        RECT 41.150 150.100 42.200 151.150 ;
        RECT 38.975 148.200 40.025 149.280 ;
        RECT 41.175 147.225 42.175 150.100 ;
        RECT 41.145 146.225 42.205 147.225 ;
        RECT 43.075 146.225 44.075 152.050 ;
        RECT 44.775 147.225 45.765 147.250 ;
        RECT 44.770 146.225 45.770 147.225 ;
        RECT 44.775 146.200 45.765 146.225 ;
        RECT 48.625 145.000 49.625 152.325 ;
        RECT 21.400 144.000 49.625 145.000 ;
        RECT 52.750 145.000 53.750 176.900 ;
        RECT 54.750 165.105 55.855 186.515 ;
        RECT 58.350 177.925 59.350 188.600 ;
        RECT 64.400 188.575 65.450 188.600 ;
        RECT 61.100 187.620 65.425 187.625 ;
        RECT 61.100 186.625 70.195 187.620 ;
        RECT 61.100 177.925 62.100 186.625 ;
        RECT 63.175 184.275 64.500 185.275 ;
        RECT 63.175 177.925 64.175 184.275 ;
        RECT 65.275 184.250 66.325 185.300 ;
        RECT 56.925 175.625 57.925 177.900 ;
        RECT 58.325 176.875 59.375 177.925 ;
        RECT 61.075 176.875 62.125 177.925 ;
        RECT 63.175 176.900 64.775 177.925 ;
        RECT 63.725 176.875 64.775 176.900 ;
        RECT 65.300 175.625 66.300 184.250 ;
        RECT 67.000 182.475 68.050 183.525 ;
        RECT 56.925 174.625 66.300 175.625 ;
        RECT 67.025 175.625 68.025 182.475 ;
        RECT 69.200 182.220 70.195 186.625 ;
        RECT 69.200 181.480 70.200 182.220 ;
        RECT 69.205 177.925 70.200 181.480 ;
        RECT 69.175 176.875 70.225 177.925 ;
        RECT 72.255 177.905 73.245 177.930 ;
        RECT 72.250 176.905 73.250 177.905 ;
        RECT 72.255 176.880 73.245 176.905 ;
        RECT 74.000 175.925 75.000 197.000 ;
        RECT 80.175 187.680 81.280 204.620 ;
        RECT 83.775 200.500 84.775 211.175 ;
        RECT 89.825 211.150 90.875 211.175 ;
        RECT 104.505 210.225 105.620 210.255 ;
        RECT 107.670 210.225 108.825 210.250 ;
        RECT 86.525 210.195 90.850 210.200 ;
        RECT 86.525 209.200 95.620 210.195 ;
        RECT 86.525 200.500 87.525 209.200 ;
        RECT 88.600 206.850 89.925 207.850 ;
        RECT 88.600 200.500 89.600 206.850 ;
        RECT 90.700 206.825 91.750 207.875 ;
        RECT 82.350 198.200 83.350 200.475 ;
        RECT 83.750 199.450 84.800 200.500 ;
        RECT 86.500 199.450 87.550 200.500 ;
        RECT 88.600 199.475 90.200 200.500 ;
        RECT 89.150 199.450 90.200 199.475 ;
        RECT 90.725 198.200 91.725 206.825 ;
        RECT 92.425 205.050 93.475 206.100 ;
        RECT 82.350 197.200 91.725 198.200 ;
        RECT 92.450 198.200 93.450 205.050 ;
        RECT 94.625 204.795 95.620 209.200 ;
        RECT 104.505 209.120 108.825 210.225 ;
        RECT 104.505 209.090 105.620 209.120 ;
        RECT 107.670 209.095 108.825 209.120 ;
        RECT 107.695 205.755 108.800 209.095 ;
        RECT 94.625 204.055 95.625 204.795 ;
        RECT 94.630 200.500 95.625 204.055 ;
        RECT 105.600 204.650 108.800 205.755 ;
        RECT 94.600 199.450 95.650 200.500 ;
        RECT 92.450 197.200 94.925 198.200 ;
        RECT 83.925 196.275 84.975 196.300 ;
        RECT 82.345 195.275 84.975 196.275 ;
        RECT 83.925 195.250 84.975 195.275 ;
        RECT 83.950 191.000 84.950 195.250 ;
        RECT 85.825 191.375 86.825 197.200 ;
        RECT 92.000 195.250 93.050 196.300 ;
        RECT 89.825 193.350 90.875 194.430 ;
        RECT 92.025 192.375 93.025 195.250 ;
        RECT 91.995 191.375 93.055 192.375 ;
        RECT 93.925 191.375 94.925 197.200 ;
        RECT 95.900 197.000 100.425 198.000 ;
        RECT 95.625 192.375 96.615 192.400 ;
        RECT 95.620 191.375 96.620 192.375 ;
        RECT 95.625 191.350 96.615 191.375 ;
        RECT 83.950 190.995 87.050 191.000 ;
        RECT 83.950 190.005 87.075 190.995 ;
        RECT 83.950 190.000 87.050 190.005 ;
        RECT 89.825 189.600 90.875 189.625 ;
        RECT 83.775 188.600 86.825 189.600 ;
        RECT 89.825 188.600 97.625 189.600 ;
        RECT 79.080 186.525 81.305 187.680 ;
        RECT 79.080 186.515 81.280 186.525 ;
        RECT 67.025 174.625 69.500 175.625 ;
        RECT 70.475 174.925 77.100 175.925 ;
        RECT 58.625 173.725 59.625 173.730 ;
        RECT 58.500 173.700 59.625 173.725 ;
        RECT 56.920 172.700 59.625 173.700 ;
        RECT 58.500 172.675 59.625 172.700 ;
        RECT 58.625 172.670 59.625 172.675 ;
        RECT 60.400 168.800 61.400 174.625 ;
        RECT 66.575 172.675 67.625 173.725 ;
        RECT 64.400 170.775 65.450 171.855 ;
        RECT 66.600 169.800 67.600 172.675 ;
        RECT 66.570 168.800 67.630 169.800 ;
        RECT 68.500 168.800 69.500 174.625 ;
        RECT 70.200 169.800 71.190 169.825 ;
        RECT 70.195 168.800 71.195 169.800 ;
        RECT 70.200 168.775 71.190 168.800 ;
        RECT 64.400 167.025 65.450 167.050 ;
        RECT 58.350 166.025 61.400 167.025 ;
        RECT 64.400 166.025 72.200 167.025 ;
        RECT 74.005 166.800 75.005 173.800 ;
        RECT 54.725 165.080 55.880 165.105 ;
        RECT 54.720 163.975 55.880 165.080 ;
        RECT 54.725 163.950 55.880 163.975 ;
        RECT 58.350 155.350 59.350 166.025 ;
        RECT 64.400 166.000 65.450 166.025 ;
        RECT 73.980 165.750 75.030 166.800 ;
        RECT 61.100 165.045 65.425 165.050 ;
        RECT 61.100 164.050 70.195 165.045 ;
        RECT 76.100 164.575 77.100 174.925 ;
        RECT 80.175 165.105 81.280 186.515 ;
        RECT 83.775 177.925 84.775 188.600 ;
        RECT 89.825 188.575 90.875 188.600 ;
        RECT 86.525 187.620 90.850 187.625 ;
        RECT 86.525 186.625 95.620 187.620 ;
        RECT 86.525 177.925 87.525 186.625 ;
        RECT 88.600 184.275 89.925 185.275 ;
        RECT 88.600 177.925 89.600 184.275 ;
        RECT 90.700 184.250 91.750 185.300 ;
        RECT 82.350 175.625 83.350 177.900 ;
        RECT 83.750 176.875 84.800 177.925 ;
        RECT 86.500 176.875 87.550 177.925 ;
        RECT 88.600 176.900 90.200 177.925 ;
        RECT 89.150 176.875 90.200 176.900 ;
        RECT 90.725 175.625 91.725 184.250 ;
        RECT 92.425 182.475 93.475 183.525 ;
        RECT 82.350 174.625 91.725 175.625 ;
        RECT 92.450 175.625 93.450 182.475 ;
        RECT 94.625 182.220 95.620 186.625 ;
        RECT 94.625 181.480 95.625 182.220 ;
        RECT 94.630 177.925 95.625 181.480 ;
        RECT 94.600 176.875 95.650 177.925 ;
        RECT 99.425 175.925 100.425 197.000 ;
        RECT 105.600 187.680 106.705 204.650 ;
        RECT 109.200 200.500 110.200 211.175 ;
        RECT 115.250 211.150 116.300 211.175 ;
        RECT 111.950 210.195 116.275 210.200 ;
        RECT 111.950 209.200 121.045 210.195 ;
        RECT 125.195 210.150 126.245 211.200 ;
        RECT 134.625 211.175 137.675 212.175 ;
        RECT 140.675 211.175 148.475 212.175 ;
        RECT 127.920 210.295 128.970 210.320 ;
        RECT 127.100 210.290 128.970 210.295 ;
        RECT 127.075 209.300 128.970 210.290 ;
        RECT 127.100 209.295 128.970 209.300 ;
        RECT 127.920 209.270 128.970 209.295 ;
        RECT 111.950 200.500 112.950 209.200 ;
        RECT 116.125 207.850 117.175 207.875 ;
        RECT 117.850 207.850 118.900 208.365 ;
        RECT 114.025 206.850 115.350 207.850 ;
        RECT 116.125 206.850 118.900 207.850 ;
        RECT 114.025 200.500 115.025 206.850 ;
        RECT 116.125 206.825 117.175 206.850 ;
        RECT 107.775 198.200 108.775 200.475 ;
        RECT 109.175 199.450 110.225 200.500 ;
        RECT 111.925 199.450 112.975 200.500 ;
        RECT 114.025 199.475 115.625 200.500 ;
        RECT 114.575 199.450 115.625 199.475 ;
        RECT 116.150 198.200 117.150 206.825 ;
        RECT 117.850 205.050 118.900 206.100 ;
        RECT 107.775 197.200 117.150 198.200 ;
        RECT 117.875 198.200 118.875 205.050 ;
        RECT 120.050 204.795 121.045 209.200 ;
        RECT 129.810 208.420 132.370 209.525 ;
        RECT 133.095 209.095 134.250 210.250 ;
        RECT 122.045 205.155 123.045 208.340 ;
        RECT 129.810 207.695 130.915 208.420 ;
        RECT 126.515 206.590 130.915 207.695 ;
        RECT 126.515 205.180 127.620 206.590 ;
        RECT 129.930 205.755 131.045 205.785 ;
        RECT 133.120 205.755 134.225 209.095 ;
        RECT 126.495 205.155 127.650 205.180 ;
        RECT 120.050 204.055 121.050 204.795 ;
        RECT 122.045 204.100 127.650 205.155 ;
        RECT 129.930 204.650 134.225 205.755 ;
        RECT 129.930 204.620 132.130 204.650 ;
        RECT 120.055 200.500 121.050 204.055 ;
        RECT 122.070 204.050 127.650 204.100 ;
        RECT 126.495 204.025 127.650 204.050 ;
        RECT 120.025 199.450 121.075 200.500 ;
        RECT 125.105 200.480 126.095 200.505 ;
        RECT 125.100 199.480 126.100 200.480 ;
        RECT 125.105 199.455 126.095 199.480 ;
        RECT 117.875 197.200 120.350 198.200 ;
        RECT 109.350 196.275 110.400 196.300 ;
        RECT 107.770 195.275 110.400 196.275 ;
        RECT 109.350 195.250 110.400 195.275 ;
        RECT 109.375 191.000 110.375 195.250 ;
        RECT 111.250 191.375 112.250 197.200 ;
        RECT 117.425 195.250 118.475 196.300 ;
        RECT 115.250 193.350 116.300 194.430 ;
        RECT 117.450 192.375 118.450 195.250 ;
        RECT 117.420 191.375 118.480 192.375 ;
        RECT 119.350 191.375 120.350 197.200 ;
        RECT 121.325 197.000 125.850 198.000 ;
        RECT 121.050 192.375 122.040 192.400 ;
        RECT 121.045 191.375 122.045 192.375 ;
        RECT 121.050 191.350 122.040 191.375 ;
        RECT 109.375 190.995 112.475 191.000 ;
        RECT 109.375 190.005 112.500 190.995 ;
        RECT 109.375 190.000 112.475 190.005 ;
        RECT 115.250 189.600 116.300 189.625 ;
        RECT 109.200 188.600 112.250 189.600 ;
        RECT 115.250 188.600 123.050 189.600 ;
        RECT 104.505 186.525 106.730 187.680 ;
        RECT 104.505 186.515 106.705 186.525 ;
        RECT 101.500 177.900 102.550 177.925 ;
        RECT 101.500 176.900 104.600 177.900 ;
        RECT 101.500 176.875 102.550 176.900 ;
        RECT 92.450 174.625 94.925 175.625 ;
        RECT 95.900 174.925 102.525 175.925 ;
        RECT 84.050 173.725 85.050 173.730 ;
        RECT 83.925 173.700 85.050 173.725 ;
        RECT 82.345 172.700 85.050 173.700 ;
        RECT 83.925 172.675 85.050 172.700 ;
        RECT 84.050 172.670 85.050 172.675 ;
        RECT 85.825 168.800 86.825 174.625 ;
        RECT 92.000 172.675 93.050 173.725 ;
        RECT 89.825 170.775 90.875 171.855 ;
        RECT 92.025 169.800 93.025 172.675 ;
        RECT 91.995 168.800 93.055 169.800 ;
        RECT 93.925 168.800 94.925 174.625 ;
        RECT 95.625 169.800 96.615 169.825 ;
        RECT 95.620 168.800 96.620 169.800 ;
        RECT 95.625 168.775 96.615 168.800 ;
        RECT 89.825 167.025 90.875 167.050 ;
        RECT 83.775 166.025 86.825 167.025 ;
        RECT 89.825 166.025 97.625 167.025 ;
        RECT 99.430 166.800 100.430 173.800 ;
        RECT 61.100 155.350 62.100 164.050 ;
        RECT 63.175 161.700 64.500 162.700 ;
        RECT 63.175 155.350 64.175 161.700 ;
        RECT 65.275 161.675 66.325 162.725 ;
        RECT 56.925 153.050 57.925 155.325 ;
        RECT 58.325 154.300 59.375 155.350 ;
        RECT 61.075 154.300 62.125 155.350 ;
        RECT 63.175 154.325 64.775 155.350 ;
        RECT 63.725 154.300 64.775 154.325 ;
        RECT 65.300 153.050 66.300 161.675 ;
        RECT 67.000 159.900 68.050 160.950 ;
        RECT 56.925 152.050 66.300 153.050 ;
        RECT 67.025 153.050 68.025 159.900 ;
        RECT 69.200 159.645 70.195 164.050 ;
        RECT 74.050 163.575 77.100 164.575 ;
        RECT 79.080 163.950 81.305 165.105 ;
        RECT 79.080 163.940 80.195 163.950 ;
        RECT 69.200 158.905 70.200 159.645 ;
        RECT 69.205 155.350 70.200 158.905 ;
        RECT 69.175 154.300 70.225 155.350 ;
        RECT 70.455 153.325 71.505 153.350 ;
        RECT 74.050 153.325 75.050 163.575 ;
        RECT 83.775 155.350 84.775 166.025 ;
        RECT 89.825 166.000 90.875 166.025 ;
        RECT 99.405 165.750 100.455 166.800 ;
        RECT 86.525 165.045 90.850 165.050 ;
        RECT 86.525 164.050 95.620 165.045 ;
        RECT 101.525 164.575 102.525 174.925 ;
        RECT 86.525 155.350 87.525 164.050 ;
        RECT 88.600 161.700 89.925 162.700 ;
        RECT 88.600 155.350 89.600 161.700 ;
        RECT 90.700 161.675 91.750 162.725 ;
        RECT 67.025 152.050 69.500 153.050 ;
        RECT 70.455 152.325 75.050 153.325 ;
        RECT 82.350 153.050 83.350 155.325 ;
        RECT 83.750 154.300 84.800 155.350 ;
        RECT 86.500 154.300 87.550 155.350 ;
        RECT 88.600 154.325 90.200 155.350 ;
        RECT 89.150 154.300 90.200 154.325 ;
        RECT 90.725 153.050 91.725 161.675 ;
        RECT 92.425 159.900 93.475 160.950 ;
        RECT 70.455 152.300 71.505 152.325 ;
        RECT 56.930 151.125 57.920 151.150 ;
        RECT 58.500 151.125 59.550 151.150 ;
        RECT 56.920 150.125 59.550 151.125 ;
        RECT 56.930 150.100 57.920 150.125 ;
        RECT 58.500 150.100 59.550 150.125 ;
        RECT 60.400 146.225 61.400 152.050 ;
        RECT 66.575 150.100 67.625 151.150 ;
        RECT 64.400 148.200 65.450 149.280 ;
        RECT 66.600 147.225 67.600 150.100 ;
        RECT 66.570 146.225 67.630 147.225 ;
        RECT 68.500 146.225 69.500 152.050 ;
        RECT 70.200 147.225 71.190 147.250 ;
        RECT 70.195 146.225 71.195 147.225 ;
        RECT 70.200 146.200 71.190 146.225 ;
        RECT 72.255 145.000 73.245 145.025 ;
        RECT 74.020 145.000 75.020 152.325 ;
        RECT 82.350 152.050 91.725 153.050 ;
        RECT 92.450 153.050 93.450 159.900 ;
        RECT 94.625 159.645 95.620 164.050 ;
        RECT 99.475 163.575 102.525 164.575 ;
        RECT 94.625 158.905 95.625 159.645 ;
        RECT 94.630 155.350 95.625 158.905 ;
        RECT 94.600 154.300 95.650 155.350 ;
        RECT 95.880 153.325 96.930 153.350 ;
        RECT 99.475 153.325 100.475 163.575 ;
        RECT 92.450 152.050 94.925 153.050 ;
        RECT 95.880 152.325 100.475 153.325 ;
        RECT 95.880 152.300 96.930 152.325 ;
        RECT 82.355 151.125 83.345 151.150 ;
        RECT 83.925 151.125 84.975 151.150 ;
        RECT 82.345 150.125 84.975 151.125 ;
        RECT 82.355 150.100 83.345 150.125 ;
        RECT 83.925 150.100 84.975 150.125 ;
        RECT 85.825 146.225 86.825 152.050 ;
        RECT 92.000 150.100 93.050 151.150 ;
        RECT 89.825 148.200 90.875 149.280 ;
        RECT 92.025 147.225 93.025 150.100 ;
        RECT 91.995 146.225 93.055 147.225 ;
        RECT 93.925 146.225 94.925 152.050 ;
        RECT 95.625 147.225 96.615 147.250 ;
        RECT 95.620 146.225 96.620 147.225 ;
        RECT 95.625 146.200 96.615 146.225 ;
        RECT 99.475 145.000 100.475 152.325 ;
        RECT 52.750 144.000 100.475 145.000 ;
        RECT 103.600 145.000 104.600 176.900 ;
        RECT 105.600 165.105 106.705 186.515 ;
        RECT 109.200 177.925 110.200 188.600 ;
        RECT 115.250 188.575 116.300 188.600 ;
        RECT 111.950 187.620 116.275 187.625 ;
        RECT 111.950 186.625 121.045 187.620 ;
        RECT 111.950 177.925 112.950 186.625 ;
        RECT 114.025 184.275 115.350 185.275 ;
        RECT 114.025 177.925 115.025 184.275 ;
        RECT 116.125 184.250 117.175 185.300 ;
        RECT 107.775 175.625 108.775 177.900 ;
        RECT 109.175 176.875 110.225 177.925 ;
        RECT 111.925 176.875 112.975 177.925 ;
        RECT 114.025 176.900 115.625 177.925 ;
        RECT 114.575 176.875 115.625 176.900 ;
        RECT 116.150 175.625 117.150 184.250 ;
        RECT 117.850 182.475 118.900 183.525 ;
        RECT 107.775 174.625 117.150 175.625 ;
        RECT 117.875 175.625 118.875 182.475 ;
        RECT 120.050 182.220 121.045 186.625 ;
        RECT 120.050 181.480 121.050 182.220 ;
        RECT 120.055 177.925 121.050 181.480 ;
        RECT 120.025 176.875 121.075 177.925 ;
        RECT 123.105 177.905 124.095 177.930 ;
        RECT 123.100 176.905 124.100 177.905 ;
        RECT 123.105 176.880 124.095 176.905 ;
        RECT 124.850 175.925 125.850 197.000 ;
        RECT 131.025 187.680 132.130 204.620 ;
        RECT 134.625 200.500 135.625 211.175 ;
        RECT 140.675 211.150 141.725 211.175 ;
        RECT 137.375 210.195 141.700 210.200 ;
        RECT 137.375 209.200 146.470 210.195 ;
        RECT 137.375 200.500 138.375 209.200 ;
        RECT 139.450 206.850 140.775 207.850 ;
        RECT 139.450 200.500 140.450 206.850 ;
        RECT 141.550 206.825 142.600 207.875 ;
        RECT 133.200 198.200 134.200 200.475 ;
        RECT 134.600 199.450 135.650 200.500 ;
        RECT 137.350 199.450 138.400 200.500 ;
        RECT 139.450 199.475 141.050 200.500 ;
        RECT 140.000 199.450 141.050 199.475 ;
        RECT 141.575 198.200 142.575 206.825 ;
        RECT 143.275 205.050 144.325 206.100 ;
        RECT 133.200 197.200 142.575 198.200 ;
        RECT 143.300 198.200 144.300 205.050 ;
        RECT 145.475 204.795 146.470 209.200 ;
        RECT 145.475 204.055 146.475 204.795 ;
        RECT 145.480 200.500 146.475 204.055 ;
        RECT 145.450 199.450 146.500 200.500 ;
        RECT 148.525 200.470 149.525 200.475 ;
        RECT 148.500 199.480 149.550 200.470 ;
        RECT 148.525 199.475 149.525 199.480 ;
        RECT 143.300 197.200 145.775 198.200 ;
        RECT 134.775 196.275 135.825 196.300 ;
        RECT 133.195 195.275 135.825 196.275 ;
        RECT 134.775 195.250 135.825 195.275 ;
        RECT 134.800 191.000 135.800 195.250 ;
        RECT 136.675 191.375 137.675 197.200 ;
        RECT 142.850 195.250 143.900 196.300 ;
        RECT 140.675 193.350 141.725 194.430 ;
        RECT 142.875 192.375 143.875 195.250 ;
        RECT 142.845 191.375 143.905 192.375 ;
        RECT 144.775 191.375 145.775 197.200 ;
        RECT 146.750 197.000 151.275 198.000 ;
        RECT 146.475 192.375 147.465 192.400 ;
        RECT 146.470 191.375 147.470 192.375 ;
        RECT 146.475 191.350 147.465 191.375 ;
        RECT 134.800 190.995 137.900 191.000 ;
        RECT 134.800 190.005 137.925 190.995 ;
        RECT 134.800 190.000 137.900 190.005 ;
        RECT 140.675 189.600 141.725 189.625 ;
        RECT 134.625 188.600 137.675 189.600 ;
        RECT 140.675 188.600 148.475 189.600 ;
        RECT 129.930 186.525 132.155 187.680 ;
        RECT 129.930 186.515 132.130 186.525 ;
        RECT 117.875 174.625 120.350 175.625 ;
        RECT 121.325 174.925 127.950 175.925 ;
        RECT 109.475 173.725 110.475 173.730 ;
        RECT 109.350 173.700 110.475 173.725 ;
        RECT 107.770 172.700 110.475 173.700 ;
        RECT 109.350 172.675 110.475 172.700 ;
        RECT 109.475 172.670 110.475 172.675 ;
        RECT 111.250 168.800 112.250 174.625 ;
        RECT 117.425 172.675 118.475 173.725 ;
        RECT 115.250 170.775 116.300 171.855 ;
        RECT 117.450 169.800 118.450 172.675 ;
        RECT 117.420 168.800 118.480 169.800 ;
        RECT 119.350 168.800 120.350 174.625 ;
        RECT 121.050 169.800 122.040 169.825 ;
        RECT 121.045 168.800 122.045 169.800 ;
        RECT 121.050 168.775 122.040 168.800 ;
        RECT 115.250 167.025 116.300 167.050 ;
        RECT 109.200 166.025 112.250 167.025 ;
        RECT 115.250 166.025 123.050 167.025 ;
        RECT 124.855 166.800 125.855 173.800 ;
        RECT 105.575 165.080 106.730 165.105 ;
        RECT 105.570 163.975 106.730 165.080 ;
        RECT 105.575 163.950 106.730 163.975 ;
        RECT 109.200 155.350 110.200 166.025 ;
        RECT 115.250 166.000 116.300 166.025 ;
        RECT 124.830 165.750 125.880 166.800 ;
        RECT 111.950 165.045 116.275 165.050 ;
        RECT 111.950 164.050 121.045 165.045 ;
        RECT 126.950 164.575 127.950 174.925 ;
        RECT 131.025 165.105 132.130 186.515 ;
        RECT 134.625 177.925 135.625 188.600 ;
        RECT 140.675 188.575 141.725 188.600 ;
        RECT 137.375 187.620 141.700 187.625 ;
        RECT 137.375 186.625 146.470 187.620 ;
        RECT 137.375 177.925 138.375 186.625 ;
        RECT 139.450 184.275 140.775 185.275 ;
        RECT 139.450 177.925 140.450 184.275 ;
        RECT 141.550 184.250 142.600 185.300 ;
        RECT 133.200 175.625 134.200 177.900 ;
        RECT 134.600 176.875 135.650 177.925 ;
        RECT 137.350 176.875 138.400 177.925 ;
        RECT 139.450 176.900 141.050 177.925 ;
        RECT 140.000 176.875 141.050 176.900 ;
        RECT 141.575 175.625 142.575 184.250 ;
        RECT 143.275 182.475 144.325 183.525 ;
        RECT 133.200 174.625 142.575 175.625 ;
        RECT 143.300 175.625 144.300 182.475 ;
        RECT 145.475 182.220 146.470 186.625 ;
        RECT 145.475 181.480 146.475 182.220 ;
        RECT 145.480 177.925 146.475 181.480 ;
        RECT 145.450 176.875 146.500 177.925 ;
        RECT 150.275 175.925 151.275 197.000 ;
        RECT 156.500 176.875 157.550 177.955 ;
        RECT 143.300 174.625 145.775 175.625 ;
        RECT 146.750 174.925 153.375 175.925 ;
        RECT 134.900 173.725 135.900 173.730 ;
        RECT 134.775 173.700 135.900 173.725 ;
        RECT 133.195 172.700 135.900 173.700 ;
        RECT 134.775 172.675 135.900 172.700 ;
        RECT 134.900 172.670 135.900 172.675 ;
        RECT 136.675 168.800 137.675 174.625 ;
        RECT 142.850 172.675 143.900 173.725 ;
        RECT 140.675 170.775 141.725 171.855 ;
        RECT 142.875 169.800 143.875 172.675 ;
        RECT 142.845 168.800 143.905 169.800 ;
        RECT 144.775 168.800 145.775 174.625 ;
        RECT 146.475 169.800 147.465 169.825 ;
        RECT 146.470 168.800 147.470 169.800 ;
        RECT 146.475 168.775 147.465 168.800 ;
        RECT 140.675 167.025 141.725 167.050 ;
        RECT 134.625 166.025 137.675 167.025 ;
        RECT 140.675 166.025 148.475 167.025 ;
        RECT 150.280 166.800 151.280 173.800 ;
        RECT 111.950 155.350 112.950 164.050 ;
        RECT 114.025 161.700 115.350 162.700 ;
        RECT 114.025 155.350 115.025 161.700 ;
        RECT 116.125 161.675 117.175 162.725 ;
        RECT 107.775 153.050 108.775 155.325 ;
        RECT 109.175 154.300 110.225 155.350 ;
        RECT 111.925 154.300 112.975 155.350 ;
        RECT 114.025 154.325 115.625 155.350 ;
        RECT 114.575 154.300 115.625 154.325 ;
        RECT 116.150 153.050 117.150 161.675 ;
        RECT 117.850 159.900 118.900 160.950 ;
        RECT 107.775 152.050 117.150 153.050 ;
        RECT 117.875 153.050 118.875 159.900 ;
        RECT 120.050 159.645 121.045 164.050 ;
        RECT 124.900 163.575 127.950 164.575 ;
        RECT 129.930 163.950 132.155 165.105 ;
        RECT 129.930 163.940 131.045 163.950 ;
        RECT 120.050 158.905 121.050 159.645 ;
        RECT 120.055 155.350 121.050 158.905 ;
        RECT 120.025 154.300 121.075 155.350 ;
        RECT 121.305 153.325 122.355 153.350 ;
        RECT 124.900 153.325 125.900 163.575 ;
        RECT 134.625 155.350 135.625 166.025 ;
        RECT 140.675 166.000 141.725 166.025 ;
        RECT 150.255 165.750 151.305 166.800 ;
        RECT 137.375 165.045 141.700 165.050 ;
        RECT 137.375 164.050 146.470 165.045 ;
        RECT 152.375 164.575 153.375 174.925 ;
        RECT 137.375 155.350 138.375 164.050 ;
        RECT 139.450 161.700 140.775 162.700 ;
        RECT 139.450 155.350 140.450 161.700 ;
        RECT 141.550 161.675 142.600 162.725 ;
        RECT 117.875 152.050 120.350 153.050 ;
        RECT 121.305 152.325 125.900 153.325 ;
        RECT 133.200 153.050 134.200 155.325 ;
        RECT 134.600 154.300 135.650 155.350 ;
        RECT 137.350 154.300 138.400 155.350 ;
        RECT 139.450 154.325 141.050 155.350 ;
        RECT 140.000 154.300 141.050 154.325 ;
        RECT 141.575 153.050 142.575 161.675 ;
        RECT 143.275 159.900 144.325 160.950 ;
        RECT 121.305 152.300 122.355 152.325 ;
        RECT 107.780 151.125 108.770 151.150 ;
        RECT 109.350 151.125 110.400 151.150 ;
        RECT 107.770 150.125 110.400 151.125 ;
        RECT 107.780 150.100 108.770 150.125 ;
        RECT 109.350 150.100 110.400 150.125 ;
        RECT 111.250 146.225 112.250 152.050 ;
        RECT 117.425 150.100 118.475 151.150 ;
        RECT 115.250 148.200 116.300 149.280 ;
        RECT 117.450 147.225 118.450 150.100 ;
        RECT 117.420 146.225 118.480 147.225 ;
        RECT 119.350 146.225 120.350 152.050 ;
        RECT 121.050 147.225 122.040 147.250 ;
        RECT 121.045 146.225 122.045 147.225 ;
        RECT 121.050 146.200 122.040 146.225 ;
        RECT 123.105 145.000 124.095 145.025 ;
        RECT 124.870 145.000 125.870 152.325 ;
        RECT 133.200 152.050 142.575 153.050 ;
        RECT 143.300 153.050 144.300 159.900 ;
        RECT 145.475 159.645 146.470 164.050 ;
        RECT 150.325 163.575 153.375 164.575 ;
        RECT 145.475 158.905 146.475 159.645 ;
        RECT 145.480 155.350 146.475 158.905 ;
        RECT 145.450 154.300 146.500 155.350 ;
        RECT 146.730 153.325 147.780 153.350 ;
        RECT 150.325 153.325 151.325 163.575 ;
        RECT 143.300 152.050 145.775 153.050 ;
        RECT 146.730 152.325 151.325 153.325 ;
        RECT 146.730 152.300 147.780 152.325 ;
        RECT 133.205 151.125 134.195 151.150 ;
        RECT 134.775 151.125 135.825 151.150 ;
        RECT 133.195 150.125 135.825 151.125 ;
        RECT 133.205 150.100 134.195 150.125 ;
        RECT 134.775 150.100 135.825 150.125 ;
        RECT 136.675 146.225 137.675 152.050 ;
        RECT 142.850 150.100 143.900 151.150 ;
        RECT 140.675 148.200 141.725 149.280 ;
        RECT 142.875 147.225 143.875 150.100 ;
        RECT 142.845 146.225 143.905 147.225 ;
        RECT 144.775 146.225 145.775 152.050 ;
        RECT 146.475 147.225 147.465 147.250 ;
        RECT 146.470 146.225 147.470 147.225 ;
        RECT 146.475 146.200 147.465 146.225 ;
        RECT 150.325 145.000 151.325 152.325 ;
        RECT 103.600 144.000 151.325 145.000 ;
        RECT 21.405 143.975 22.395 144.000 ;
        RECT 72.255 143.975 73.245 144.000 ;
        RECT 123.105 143.975 124.095 144.000 ;
        RECT 99.680 142.550 100.670 142.575 ;
        RECT 13.550 140.175 14.600 140.200 ;
        RECT 7.500 139.175 10.550 140.175 ;
        RECT 13.550 139.175 21.350 140.175 ;
        RECT 23.520 139.200 24.520 142.550 ;
        RECT 38.975 140.175 40.025 140.200 ;
        RECT 64.400 140.175 65.450 140.200 ;
        RECT 2.805 138.225 3.920 138.255 ;
        RECT 5.970 138.225 7.125 138.250 ;
        RECT 2.805 137.120 7.125 138.225 ;
        RECT 2.805 137.090 3.920 137.120 ;
        RECT 5.970 137.095 7.125 137.120 ;
        RECT 5.995 133.755 7.100 137.095 ;
        RECT 3.900 132.650 7.100 133.755 ;
        RECT 3.900 115.680 5.005 132.650 ;
        RECT 7.500 128.500 8.500 139.175 ;
        RECT 13.550 139.150 14.600 139.175 ;
        RECT 10.250 138.195 14.575 138.200 ;
        RECT 10.250 137.200 19.345 138.195 ;
        RECT 23.495 138.150 24.545 139.200 ;
        RECT 32.925 139.175 35.975 140.175 ;
        RECT 38.975 139.175 46.775 140.175 ;
        RECT 58.350 139.175 61.400 140.175 ;
        RECT 64.400 139.175 72.200 140.175 ;
        RECT 74.370 139.200 75.370 142.550 ;
        RECT 99.675 141.550 100.675 142.550 ;
        RECT 99.680 141.525 100.670 141.550 ;
        RECT 89.825 140.175 90.875 140.200 ;
        RECT 115.250 140.175 116.300 140.200 ;
        RECT 26.220 138.295 27.270 138.320 ;
        RECT 25.400 138.290 27.270 138.295 ;
        RECT 25.375 137.300 27.270 138.290 ;
        RECT 25.400 137.295 27.270 137.300 ;
        RECT 26.220 137.270 27.270 137.295 ;
        RECT 10.250 128.500 11.250 137.200 ;
        RECT 14.425 135.850 15.475 135.875 ;
        RECT 16.150 135.850 17.200 136.365 ;
        RECT 12.325 134.850 13.650 135.850 ;
        RECT 14.425 134.850 17.200 135.850 ;
        RECT 12.325 128.500 13.325 134.850 ;
        RECT 14.425 134.825 15.475 134.850 ;
        RECT 6.075 126.200 7.075 128.475 ;
        RECT 7.475 127.450 8.525 128.500 ;
        RECT 10.225 127.450 11.275 128.500 ;
        RECT 12.325 127.475 13.925 128.500 ;
        RECT 12.875 127.450 13.925 127.475 ;
        RECT 14.450 126.200 15.450 134.825 ;
        RECT 16.150 133.050 17.200 134.100 ;
        RECT 6.075 125.200 15.450 126.200 ;
        RECT 16.175 126.200 17.175 133.050 ;
        RECT 18.350 132.795 19.345 137.200 ;
        RECT 28.110 136.420 30.670 137.525 ;
        RECT 31.395 137.095 32.550 138.250 ;
        RECT 20.345 133.155 21.345 136.340 ;
        RECT 28.110 135.695 29.215 136.420 ;
        RECT 24.815 134.590 29.215 135.695 ;
        RECT 24.815 133.180 25.920 134.590 ;
        RECT 28.230 133.755 29.345 133.785 ;
        RECT 31.420 133.755 32.525 137.095 ;
        RECT 24.795 133.155 25.950 133.180 ;
        RECT 18.350 132.055 19.350 132.795 ;
        RECT 20.345 132.100 25.950 133.155 ;
        RECT 28.230 132.650 32.525 133.755 ;
        RECT 28.230 132.620 30.430 132.650 ;
        RECT 18.355 128.500 19.350 132.055 ;
        RECT 20.370 132.050 25.950 132.100 ;
        RECT 24.795 132.025 25.950 132.050 ;
        RECT 18.325 127.450 19.375 128.500 ;
        RECT 23.405 128.480 24.395 128.505 ;
        RECT 23.400 127.480 24.400 128.480 ;
        RECT 23.405 127.455 24.395 127.480 ;
        RECT 16.175 125.200 18.650 126.200 ;
        RECT 7.650 124.275 8.700 124.300 ;
        RECT 6.070 123.275 8.700 124.275 ;
        RECT 7.650 123.250 8.700 123.275 ;
        RECT 7.675 119.000 8.675 123.250 ;
        RECT 9.550 119.375 10.550 125.200 ;
        RECT 15.725 123.250 16.775 124.300 ;
        RECT 13.550 121.350 14.600 122.430 ;
        RECT 15.750 120.375 16.750 123.250 ;
        RECT 15.720 119.375 16.780 120.375 ;
        RECT 17.650 119.375 18.650 125.200 ;
        RECT 19.625 125.000 24.150 126.000 ;
        RECT 19.350 120.375 20.340 120.400 ;
        RECT 19.345 119.375 20.345 120.375 ;
        RECT 19.350 119.350 20.340 119.375 ;
        RECT 7.675 118.995 10.775 119.000 ;
        RECT 7.675 118.005 10.800 118.995 ;
        RECT 7.675 118.000 10.775 118.005 ;
        RECT 13.550 117.600 14.600 117.625 ;
        RECT 7.500 116.600 10.550 117.600 ;
        RECT 13.550 116.600 21.350 117.600 ;
        RECT 2.805 114.525 5.030 115.680 ;
        RECT 2.805 114.515 5.005 114.525 ;
        RECT 3.900 93.105 5.005 114.515 ;
        RECT 7.500 105.925 8.500 116.600 ;
        RECT 13.550 116.575 14.600 116.600 ;
        RECT 10.250 115.620 14.575 115.625 ;
        RECT 10.250 114.625 19.345 115.620 ;
        RECT 10.250 105.925 11.250 114.625 ;
        RECT 12.325 112.275 13.650 113.275 ;
        RECT 12.325 105.925 13.325 112.275 ;
        RECT 14.425 112.250 15.475 113.300 ;
        RECT 6.075 103.625 7.075 105.900 ;
        RECT 7.475 104.875 8.525 105.925 ;
        RECT 10.225 104.875 11.275 105.925 ;
        RECT 12.325 104.900 13.925 105.925 ;
        RECT 12.875 104.875 13.925 104.900 ;
        RECT 14.450 103.625 15.450 112.250 ;
        RECT 16.150 110.475 17.200 111.525 ;
        RECT 6.075 102.625 15.450 103.625 ;
        RECT 16.175 103.625 17.175 110.475 ;
        RECT 18.350 110.220 19.345 114.625 ;
        RECT 18.350 109.480 19.350 110.220 ;
        RECT 18.355 105.925 19.350 109.480 ;
        RECT 18.325 104.875 19.375 105.925 ;
        RECT 21.405 105.905 22.395 105.930 ;
        RECT 21.400 104.905 22.400 105.905 ;
        RECT 21.405 104.880 22.395 104.905 ;
        RECT 23.150 103.925 24.150 125.000 ;
        RECT 29.325 115.680 30.430 132.620 ;
        RECT 32.925 128.500 33.925 139.175 ;
        RECT 38.975 139.150 40.025 139.175 ;
        RECT 53.655 138.225 54.770 138.255 ;
        RECT 56.820 138.225 57.975 138.250 ;
        RECT 35.675 138.195 40.000 138.200 ;
        RECT 35.675 137.200 44.770 138.195 ;
        RECT 35.675 128.500 36.675 137.200 ;
        RECT 37.750 134.850 39.075 135.850 ;
        RECT 37.750 128.500 38.750 134.850 ;
        RECT 39.850 134.825 40.900 135.875 ;
        RECT 31.500 126.200 32.500 128.475 ;
        RECT 32.900 127.450 33.950 128.500 ;
        RECT 35.650 127.450 36.700 128.500 ;
        RECT 37.750 127.475 39.350 128.500 ;
        RECT 38.300 127.450 39.350 127.475 ;
        RECT 39.875 126.200 40.875 134.825 ;
        RECT 41.575 133.050 42.625 134.100 ;
        RECT 31.500 125.200 40.875 126.200 ;
        RECT 41.600 126.200 42.600 133.050 ;
        RECT 43.775 132.795 44.770 137.200 ;
        RECT 53.655 137.120 57.975 138.225 ;
        RECT 53.655 137.090 54.770 137.120 ;
        RECT 56.820 137.095 57.975 137.120 ;
        RECT 56.845 133.755 57.950 137.095 ;
        RECT 43.775 132.055 44.775 132.795 ;
        RECT 43.780 128.500 44.775 132.055 ;
        RECT 54.750 132.650 57.950 133.755 ;
        RECT 43.750 127.450 44.800 128.500 ;
        RECT 41.600 125.200 44.075 126.200 ;
        RECT 33.075 124.275 34.125 124.300 ;
        RECT 31.495 123.275 34.125 124.275 ;
        RECT 33.075 123.250 34.125 123.275 ;
        RECT 33.100 119.000 34.100 123.250 ;
        RECT 34.975 119.375 35.975 125.200 ;
        RECT 41.150 123.250 42.200 124.300 ;
        RECT 38.975 121.350 40.025 122.430 ;
        RECT 41.175 120.375 42.175 123.250 ;
        RECT 41.145 119.375 42.205 120.375 ;
        RECT 43.075 119.375 44.075 125.200 ;
        RECT 45.050 125.000 49.575 126.000 ;
        RECT 44.775 120.375 45.765 120.400 ;
        RECT 44.770 119.375 45.770 120.375 ;
        RECT 44.775 119.350 45.765 119.375 ;
        RECT 33.100 118.995 36.200 119.000 ;
        RECT 33.100 118.005 36.225 118.995 ;
        RECT 33.100 118.000 36.200 118.005 ;
        RECT 38.975 117.600 40.025 117.625 ;
        RECT 32.925 116.600 35.975 117.600 ;
        RECT 38.975 116.600 46.775 117.600 ;
        RECT 28.230 114.525 30.455 115.680 ;
        RECT 28.230 114.515 30.430 114.525 ;
        RECT 16.175 102.625 18.650 103.625 ;
        RECT 19.625 102.925 26.250 103.925 ;
        RECT 7.775 101.725 8.775 101.730 ;
        RECT 7.650 101.700 8.775 101.725 ;
        RECT 6.070 100.700 8.775 101.700 ;
        RECT 7.650 100.675 8.775 100.700 ;
        RECT 7.775 100.670 8.775 100.675 ;
        RECT 9.550 96.800 10.550 102.625 ;
        RECT 15.725 100.675 16.775 101.725 ;
        RECT 13.550 98.775 14.600 99.855 ;
        RECT 15.750 97.800 16.750 100.675 ;
        RECT 15.720 96.800 16.780 97.800 ;
        RECT 17.650 96.800 18.650 102.625 ;
        RECT 19.350 97.800 20.340 97.825 ;
        RECT 19.345 96.800 20.345 97.800 ;
        RECT 19.350 96.775 20.340 96.800 ;
        RECT 13.550 95.025 14.600 95.050 ;
        RECT 7.500 94.025 10.550 95.025 ;
        RECT 13.550 94.025 21.350 95.025 ;
        RECT 23.155 94.800 24.155 101.800 ;
        RECT 3.875 93.080 5.030 93.105 ;
        RECT 3.870 91.975 5.030 93.080 ;
        RECT 3.875 91.950 5.030 91.975 ;
        RECT 7.500 83.350 8.500 94.025 ;
        RECT 13.550 94.000 14.600 94.025 ;
        RECT 23.130 93.750 24.180 94.800 ;
        RECT 10.250 93.045 14.575 93.050 ;
        RECT 10.250 92.050 19.345 93.045 ;
        RECT 25.250 92.575 26.250 102.925 ;
        RECT 29.325 93.105 30.430 114.515 ;
        RECT 32.925 105.925 33.925 116.600 ;
        RECT 38.975 116.575 40.025 116.600 ;
        RECT 35.675 115.620 40.000 115.625 ;
        RECT 35.675 114.625 44.770 115.620 ;
        RECT 35.675 105.925 36.675 114.625 ;
        RECT 37.750 112.275 39.075 113.275 ;
        RECT 37.750 105.925 38.750 112.275 ;
        RECT 39.850 112.250 40.900 113.300 ;
        RECT 31.500 103.625 32.500 105.900 ;
        RECT 32.900 104.875 33.950 105.925 ;
        RECT 35.650 104.875 36.700 105.925 ;
        RECT 37.750 104.900 39.350 105.925 ;
        RECT 38.300 104.875 39.350 104.900 ;
        RECT 39.875 103.625 40.875 112.250 ;
        RECT 41.575 110.475 42.625 111.525 ;
        RECT 31.500 102.625 40.875 103.625 ;
        RECT 41.600 103.625 42.600 110.475 ;
        RECT 43.775 110.220 44.770 114.625 ;
        RECT 43.775 109.480 44.775 110.220 ;
        RECT 43.780 105.925 44.775 109.480 ;
        RECT 43.750 104.875 44.800 105.925 ;
        RECT 48.575 103.925 49.575 125.000 ;
        RECT 54.750 115.680 55.855 132.650 ;
        RECT 58.350 128.500 59.350 139.175 ;
        RECT 64.400 139.150 65.450 139.175 ;
        RECT 61.100 138.195 65.425 138.200 ;
        RECT 61.100 137.200 70.195 138.195 ;
        RECT 74.345 138.150 75.395 139.200 ;
        RECT 83.775 139.175 86.825 140.175 ;
        RECT 89.825 139.175 97.625 140.175 ;
        RECT 109.200 139.175 112.250 140.175 ;
        RECT 115.250 139.175 123.050 140.175 ;
        RECT 125.220 139.200 126.220 142.550 ;
        RECT 140.675 140.175 141.725 140.200 ;
        RECT 77.070 138.295 78.120 138.320 ;
        RECT 76.250 138.290 78.120 138.295 ;
        RECT 76.225 137.300 78.120 138.290 ;
        RECT 76.250 137.295 78.120 137.300 ;
        RECT 77.070 137.270 78.120 137.295 ;
        RECT 61.100 128.500 62.100 137.200 ;
        RECT 65.275 135.850 66.325 135.875 ;
        RECT 67.000 135.850 68.050 136.365 ;
        RECT 63.175 134.850 64.500 135.850 ;
        RECT 65.275 134.850 68.050 135.850 ;
        RECT 63.175 128.500 64.175 134.850 ;
        RECT 65.275 134.825 66.325 134.850 ;
        RECT 56.925 126.200 57.925 128.475 ;
        RECT 58.325 127.450 59.375 128.500 ;
        RECT 61.075 127.450 62.125 128.500 ;
        RECT 63.175 127.475 64.775 128.500 ;
        RECT 63.725 127.450 64.775 127.475 ;
        RECT 65.300 126.200 66.300 134.825 ;
        RECT 67.000 133.050 68.050 134.100 ;
        RECT 56.925 125.200 66.300 126.200 ;
        RECT 67.025 126.200 68.025 133.050 ;
        RECT 69.200 132.795 70.195 137.200 ;
        RECT 78.960 136.420 81.520 137.525 ;
        RECT 82.245 137.095 83.400 138.250 ;
        RECT 71.195 133.155 72.195 136.340 ;
        RECT 78.960 135.695 80.065 136.420 ;
        RECT 75.665 134.590 80.065 135.695 ;
        RECT 75.665 133.180 76.770 134.590 ;
        RECT 79.080 133.755 80.195 133.785 ;
        RECT 82.270 133.755 83.375 137.095 ;
        RECT 75.645 133.155 76.800 133.180 ;
        RECT 69.200 132.055 70.200 132.795 ;
        RECT 71.195 132.100 76.800 133.155 ;
        RECT 79.080 132.650 83.375 133.755 ;
        RECT 79.080 132.620 81.280 132.650 ;
        RECT 69.205 128.500 70.200 132.055 ;
        RECT 71.220 132.050 76.800 132.100 ;
        RECT 75.645 132.025 76.800 132.050 ;
        RECT 69.175 127.450 70.225 128.500 ;
        RECT 74.255 128.480 75.245 128.505 ;
        RECT 74.250 127.480 75.250 128.480 ;
        RECT 74.255 127.455 75.245 127.480 ;
        RECT 67.025 125.200 69.500 126.200 ;
        RECT 58.500 124.275 59.550 124.300 ;
        RECT 56.920 123.275 59.550 124.275 ;
        RECT 58.500 123.250 59.550 123.275 ;
        RECT 58.525 119.000 59.525 123.250 ;
        RECT 60.400 119.375 61.400 125.200 ;
        RECT 66.575 123.250 67.625 124.300 ;
        RECT 64.400 121.350 65.450 122.430 ;
        RECT 66.600 120.375 67.600 123.250 ;
        RECT 66.570 119.375 67.630 120.375 ;
        RECT 68.500 119.375 69.500 125.200 ;
        RECT 70.475 125.000 75.000 126.000 ;
        RECT 70.200 120.375 71.190 120.400 ;
        RECT 70.195 119.375 71.195 120.375 ;
        RECT 70.200 119.350 71.190 119.375 ;
        RECT 58.525 118.995 61.625 119.000 ;
        RECT 58.525 118.005 61.650 118.995 ;
        RECT 58.525 118.000 61.625 118.005 ;
        RECT 64.400 117.600 65.450 117.625 ;
        RECT 58.350 116.600 61.400 117.600 ;
        RECT 64.400 116.600 72.200 117.600 ;
        RECT 53.655 114.525 55.880 115.680 ;
        RECT 53.655 114.515 55.855 114.525 ;
        RECT 50.650 105.900 51.700 105.925 ;
        RECT 50.650 104.900 53.750 105.900 ;
        RECT 50.650 104.875 51.700 104.900 ;
        RECT 41.600 102.625 44.075 103.625 ;
        RECT 45.050 102.925 51.675 103.925 ;
        RECT 33.200 101.725 34.200 101.730 ;
        RECT 33.075 101.700 34.200 101.725 ;
        RECT 31.495 100.700 34.200 101.700 ;
        RECT 33.075 100.675 34.200 100.700 ;
        RECT 33.200 100.670 34.200 100.675 ;
        RECT 34.975 96.800 35.975 102.625 ;
        RECT 41.150 100.675 42.200 101.725 ;
        RECT 38.975 98.775 40.025 99.855 ;
        RECT 41.175 97.800 42.175 100.675 ;
        RECT 41.145 96.800 42.205 97.800 ;
        RECT 43.075 96.800 44.075 102.625 ;
        RECT 44.775 97.800 45.765 97.825 ;
        RECT 44.770 96.800 45.770 97.800 ;
        RECT 44.775 96.775 45.765 96.800 ;
        RECT 38.975 95.025 40.025 95.050 ;
        RECT 32.925 94.025 35.975 95.025 ;
        RECT 38.975 94.025 46.775 95.025 ;
        RECT 48.580 94.800 49.580 101.800 ;
        RECT 10.250 83.350 11.250 92.050 ;
        RECT 12.325 89.700 13.650 90.700 ;
        RECT 12.325 83.350 13.325 89.700 ;
        RECT 14.425 89.675 15.475 90.725 ;
        RECT 6.075 81.050 7.075 83.325 ;
        RECT 7.475 82.300 8.525 83.350 ;
        RECT 10.225 82.300 11.275 83.350 ;
        RECT 12.325 82.325 13.925 83.350 ;
        RECT 12.875 82.300 13.925 82.325 ;
        RECT 14.450 81.050 15.450 89.675 ;
        RECT 16.150 87.900 17.200 88.950 ;
        RECT 6.075 80.050 15.450 81.050 ;
        RECT 16.175 81.050 17.175 87.900 ;
        RECT 18.350 87.645 19.345 92.050 ;
        RECT 23.200 91.575 26.250 92.575 ;
        RECT 28.230 91.950 30.455 93.105 ;
        RECT 28.230 91.940 29.345 91.950 ;
        RECT 18.350 86.905 19.350 87.645 ;
        RECT 18.355 83.350 19.350 86.905 ;
        RECT 18.325 82.300 19.375 83.350 ;
        RECT 19.605 81.325 20.655 81.350 ;
        RECT 23.200 81.325 24.200 91.575 ;
        RECT 32.925 83.350 33.925 94.025 ;
        RECT 38.975 94.000 40.025 94.025 ;
        RECT 48.555 93.750 49.605 94.800 ;
        RECT 35.675 93.045 40.000 93.050 ;
        RECT 35.675 92.050 44.770 93.045 ;
        RECT 50.675 92.575 51.675 102.925 ;
        RECT 35.675 83.350 36.675 92.050 ;
        RECT 37.750 89.700 39.075 90.700 ;
        RECT 37.750 83.350 38.750 89.700 ;
        RECT 39.850 89.675 40.900 90.725 ;
        RECT 16.175 80.050 18.650 81.050 ;
        RECT 19.605 80.325 24.200 81.325 ;
        RECT 31.500 81.050 32.500 83.325 ;
        RECT 32.900 82.300 33.950 83.350 ;
        RECT 35.650 82.300 36.700 83.350 ;
        RECT 37.750 82.325 39.350 83.350 ;
        RECT 38.300 82.300 39.350 82.325 ;
        RECT 39.875 81.050 40.875 89.675 ;
        RECT 41.575 87.900 42.625 88.950 ;
        RECT 19.605 80.300 20.655 80.325 ;
        RECT 6.080 79.125 7.070 79.150 ;
        RECT 7.650 79.125 8.700 79.150 ;
        RECT 6.070 78.125 8.700 79.125 ;
        RECT 6.080 78.100 7.070 78.125 ;
        RECT 7.650 78.100 8.700 78.125 ;
        RECT 9.550 74.225 10.550 80.050 ;
        RECT 15.725 78.100 16.775 79.150 ;
        RECT 13.550 76.200 14.600 77.280 ;
        RECT 15.750 75.225 16.750 78.100 ;
        RECT 15.720 74.225 16.780 75.225 ;
        RECT 17.650 74.225 18.650 80.050 ;
        RECT 19.350 75.225 20.340 75.250 ;
        RECT 19.345 74.225 20.345 75.225 ;
        RECT 19.350 74.200 20.340 74.225 ;
        RECT 21.405 73.000 22.395 73.025 ;
        RECT 23.170 73.000 24.170 80.325 ;
        RECT 31.500 80.050 40.875 81.050 ;
        RECT 41.600 81.050 42.600 87.900 ;
        RECT 43.775 87.645 44.770 92.050 ;
        RECT 48.625 91.575 51.675 92.575 ;
        RECT 43.775 86.905 44.775 87.645 ;
        RECT 43.780 83.350 44.775 86.905 ;
        RECT 43.750 82.300 44.800 83.350 ;
        RECT 45.030 81.325 46.080 81.350 ;
        RECT 48.625 81.325 49.625 91.575 ;
        RECT 41.600 80.050 44.075 81.050 ;
        RECT 45.030 80.325 49.625 81.325 ;
        RECT 45.030 80.300 46.080 80.325 ;
        RECT 31.505 79.125 32.495 79.150 ;
        RECT 33.075 79.125 34.125 79.150 ;
        RECT 31.495 78.125 34.125 79.125 ;
        RECT 31.505 78.100 32.495 78.125 ;
        RECT 33.075 78.100 34.125 78.125 ;
        RECT 34.975 74.225 35.975 80.050 ;
        RECT 41.150 78.100 42.200 79.150 ;
        RECT 38.975 76.200 40.025 77.280 ;
        RECT 41.175 75.225 42.175 78.100 ;
        RECT 41.145 74.225 42.205 75.225 ;
        RECT 43.075 74.225 44.075 80.050 ;
        RECT 44.775 75.225 45.765 75.250 ;
        RECT 44.770 74.225 45.770 75.225 ;
        RECT 44.775 74.200 45.765 74.225 ;
        RECT 48.625 73.000 49.625 80.325 ;
        RECT 21.400 72.000 49.625 73.000 ;
        RECT 52.750 73.000 53.750 104.900 ;
        RECT 54.750 93.105 55.855 114.515 ;
        RECT 58.350 105.925 59.350 116.600 ;
        RECT 64.400 116.575 65.450 116.600 ;
        RECT 61.100 115.620 65.425 115.625 ;
        RECT 61.100 114.625 70.195 115.620 ;
        RECT 61.100 105.925 62.100 114.625 ;
        RECT 63.175 112.275 64.500 113.275 ;
        RECT 63.175 105.925 64.175 112.275 ;
        RECT 65.275 112.250 66.325 113.300 ;
        RECT 56.925 103.625 57.925 105.900 ;
        RECT 58.325 104.875 59.375 105.925 ;
        RECT 61.075 104.875 62.125 105.925 ;
        RECT 63.175 104.900 64.775 105.925 ;
        RECT 63.725 104.875 64.775 104.900 ;
        RECT 65.300 103.625 66.300 112.250 ;
        RECT 67.000 110.475 68.050 111.525 ;
        RECT 56.925 102.625 66.300 103.625 ;
        RECT 67.025 103.625 68.025 110.475 ;
        RECT 69.200 110.220 70.195 114.625 ;
        RECT 69.200 109.480 70.200 110.220 ;
        RECT 69.205 105.925 70.200 109.480 ;
        RECT 69.175 104.875 70.225 105.925 ;
        RECT 72.255 105.905 73.245 105.930 ;
        RECT 72.250 104.905 73.250 105.905 ;
        RECT 72.255 104.880 73.245 104.905 ;
        RECT 74.000 103.925 75.000 125.000 ;
        RECT 80.175 115.680 81.280 132.620 ;
        RECT 83.775 128.500 84.775 139.175 ;
        RECT 89.825 139.150 90.875 139.175 ;
        RECT 104.505 138.225 105.620 138.255 ;
        RECT 107.670 138.225 108.825 138.250 ;
        RECT 86.525 138.195 90.850 138.200 ;
        RECT 86.525 137.200 95.620 138.195 ;
        RECT 86.525 128.500 87.525 137.200 ;
        RECT 88.600 134.850 89.925 135.850 ;
        RECT 88.600 128.500 89.600 134.850 ;
        RECT 90.700 134.825 91.750 135.875 ;
        RECT 82.350 126.200 83.350 128.475 ;
        RECT 83.750 127.450 84.800 128.500 ;
        RECT 86.500 127.450 87.550 128.500 ;
        RECT 88.600 127.475 90.200 128.500 ;
        RECT 89.150 127.450 90.200 127.475 ;
        RECT 90.725 126.200 91.725 134.825 ;
        RECT 92.425 133.050 93.475 134.100 ;
        RECT 82.350 125.200 91.725 126.200 ;
        RECT 92.450 126.200 93.450 133.050 ;
        RECT 94.625 132.795 95.620 137.200 ;
        RECT 104.505 137.120 108.825 138.225 ;
        RECT 104.505 137.090 105.620 137.120 ;
        RECT 107.670 137.095 108.825 137.120 ;
        RECT 107.695 133.755 108.800 137.095 ;
        RECT 94.625 132.055 95.625 132.795 ;
        RECT 94.630 128.500 95.625 132.055 ;
        RECT 105.600 132.650 108.800 133.755 ;
        RECT 94.600 127.450 95.650 128.500 ;
        RECT 97.675 128.470 98.675 128.475 ;
        RECT 97.650 127.480 98.700 128.470 ;
        RECT 97.675 127.475 98.675 127.480 ;
        RECT 92.450 125.200 94.925 126.200 ;
        RECT 83.925 124.275 84.975 124.300 ;
        RECT 82.345 123.275 84.975 124.275 ;
        RECT 83.925 123.250 84.975 123.275 ;
        RECT 83.950 119.000 84.950 123.250 ;
        RECT 85.825 119.375 86.825 125.200 ;
        RECT 92.000 123.250 93.050 124.300 ;
        RECT 89.825 121.350 90.875 122.430 ;
        RECT 92.025 120.375 93.025 123.250 ;
        RECT 91.995 119.375 93.055 120.375 ;
        RECT 93.925 119.375 94.925 125.200 ;
        RECT 95.900 125.000 100.425 126.000 ;
        RECT 95.625 120.375 96.615 120.400 ;
        RECT 95.620 119.375 96.620 120.375 ;
        RECT 95.625 119.350 96.615 119.375 ;
        RECT 83.950 118.995 87.050 119.000 ;
        RECT 83.950 118.005 87.075 118.995 ;
        RECT 83.950 118.000 87.050 118.005 ;
        RECT 89.825 117.600 90.875 117.625 ;
        RECT 83.775 116.600 86.825 117.600 ;
        RECT 89.825 116.600 97.625 117.600 ;
        RECT 79.080 114.525 81.305 115.680 ;
        RECT 79.080 114.515 81.280 114.525 ;
        RECT 67.025 102.625 69.500 103.625 ;
        RECT 70.475 102.925 77.100 103.925 ;
        RECT 58.625 101.725 59.625 101.730 ;
        RECT 58.500 101.700 59.625 101.725 ;
        RECT 56.920 100.700 59.625 101.700 ;
        RECT 58.500 100.675 59.625 100.700 ;
        RECT 58.625 100.670 59.625 100.675 ;
        RECT 60.400 96.800 61.400 102.625 ;
        RECT 66.575 100.675 67.625 101.725 ;
        RECT 64.400 98.775 65.450 99.855 ;
        RECT 66.600 97.800 67.600 100.675 ;
        RECT 66.570 96.800 67.630 97.800 ;
        RECT 68.500 96.800 69.500 102.625 ;
        RECT 70.200 97.800 71.190 97.825 ;
        RECT 70.195 96.800 71.195 97.800 ;
        RECT 70.200 96.775 71.190 96.800 ;
        RECT 64.400 95.025 65.450 95.050 ;
        RECT 58.350 94.025 61.400 95.025 ;
        RECT 64.400 94.025 72.200 95.025 ;
        RECT 74.005 94.800 75.005 101.800 ;
        RECT 54.725 93.080 55.880 93.105 ;
        RECT 54.720 91.975 55.880 93.080 ;
        RECT 54.725 91.950 55.880 91.975 ;
        RECT 58.350 83.350 59.350 94.025 ;
        RECT 64.400 94.000 65.450 94.025 ;
        RECT 73.980 93.750 75.030 94.800 ;
        RECT 61.100 93.045 65.425 93.050 ;
        RECT 61.100 92.050 70.195 93.045 ;
        RECT 76.100 92.575 77.100 102.925 ;
        RECT 80.175 93.105 81.280 114.515 ;
        RECT 83.775 105.925 84.775 116.600 ;
        RECT 89.825 116.575 90.875 116.600 ;
        RECT 86.525 115.620 90.850 115.625 ;
        RECT 86.525 114.625 95.620 115.620 ;
        RECT 86.525 105.925 87.525 114.625 ;
        RECT 88.600 112.275 89.925 113.275 ;
        RECT 88.600 105.925 89.600 112.275 ;
        RECT 90.700 112.250 91.750 113.300 ;
        RECT 82.350 103.625 83.350 105.900 ;
        RECT 83.750 104.875 84.800 105.925 ;
        RECT 86.500 104.875 87.550 105.925 ;
        RECT 88.600 104.900 90.200 105.925 ;
        RECT 89.150 104.875 90.200 104.900 ;
        RECT 90.725 103.625 91.725 112.250 ;
        RECT 92.425 110.475 93.475 111.525 ;
        RECT 82.350 102.625 91.725 103.625 ;
        RECT 92.450 103.625 93.450 110.475 ;
        RECT 94.625 110.220 95.620 114.625 ;
        RECT 94.625 109.480 95.625 110.220 ;
        RECT 94.630 105.925 95.625 109.480 ;
        RECT 94.600 104.875 95.650 105.925 ;
        RECT 99.425 103.925 100.425 125.000 ;
        RECT 105.600 115.680 106.705 132.650 ;
        RECT 109.200 128.500 110.200 139.175 ;
        RECT 115.250 139.150 116.300 139.175 ;
        RECT 111.950 138.195 116.275 138.200 ;
        RECT 111.950 137.200 121.045 138.195 ;
        RECT 125.195 138.150 126.245 139.200 ;
        RECT 134.625 139.175 137.675 140.175 ;
        RECT 140.675 139.175 148.475 140.175 ;
        RECT 127.920 138.295 128.970 138.320 ;
        RECT 127.100 138.290 128.970 138.295 ;
        RECT 127.075 137.300 128.970 138.290 ;
        RECT 127.100 137.295 128.970 137.300 ;
        RECT 127.920 137.270 128.970 137.295 ;
        RECT 111.950 128.500 112.950 137.200 ;
        RECT 116.125 135.850 117.175 135.875 ;
        RECT 117.850 135.850 118.900 136.365 ;
        RECT 114.025 134.850 115.350 135.850 ;
        RECT 116.125 134.850 118.900 135.850 ;
        RECT 114.025 128.500 115.025 134.850 ;
        RECT 116.125 134.825 117.175 134.850 ;
        RECT 107.775 126.200 108.775 128.475 ;
        RECT 109.175 127.450 110.225 128.500 ;
        RECT 111.925 127.450 112.975 128.500 ;
        RECT 114.025 127.475 115.625 128.500 ;
        RECT 114.575 127.450 115.625 127.475 ;
        RECT 116.150 126.200 117.150 134.825 ;
        RECT 117.850 133.050 118.900 134.100 ;
        RECT 107.775 125.200 117.150 126.200 ;
        RECT 117.875 126.200 118.875 133.050 ;
        RECT 120.050 132.795 121.045 137.200 ;
        RECT 129.810 136.420 132.370 137.525 ;
        RECT 133.095 137.095 134.250 138.250 ;
        RECT 122.045 133.155 123.045 136.340 ;
        RECT 129.810 135.695 130.915 136.420 ;
        RECT 126.515 134.590 130.915 135.695 ;
        RECT 126.515 133.180 127.620 134.590 ;
        RECT 129.930 133.755 131.045 133.785 ;
        RECT 133.120 133.755 134.225 137.095 ;
        RECT 126.495 133.155 127.650 133.180 ;
        RECT 120.050 132.055 121.050 132.795 ;
        RECT 122.045 132.100 127.650 133.155 ;
        RECT 129.930 132.650 134.225 133.755 ;
        RECT 129.930 132.620 132.130 132.650 ;
        RECT 120.055 128.500 121.050 132.055 ;
        RECT 122.070 132.050 127.650 132.100 ;
        RECT 126.495 132.025 127.650 132.050 ;
        RECT 120.025 127.450 121.075 128.500 ;
        RECT 125.105 128.480 126.095 128.505 ;
        RECT 125.100 127.480 126.100 128.480 ;
        RECT 125.105 127.455 126.095 127.480 ;
        RECT 117.875 125.200 120.350 126.200 ;
        RECT 109.350 124.275 110.400 124.300 ;
        RECT 107.770 123.275 110.400 124.275 ;
        RECT 109.350 123.250 110.400 123.275 ;
        RECT 109.375 119.000 110.375 123.250 ;
        RECT 111.250 119.375 112.250 125.200 ;
        RECT 117.425 123.250 118.475 124.300 ;
        RECT 115.250 121.350 116.300 122.430 ;
        RECT 117.450 120.375 118.450 123.250 ;
        RECT 117.420 119.375 118.480 120.375 ;
        RECT 119.350 119.375 120.350 125.200 ;
        RECT 121.325 125.000 125.850 126.000 ;
        RECT 121.050 120.375 122.040 120.400 ;
        RECT 121.045 119.375 122.045 120.375 ;
        RECT 121.050 119.350 122.040 119.375 ;
        RECT 109.375 118.995 112.475 119.000 ;
        RECT 109.375 118.005 112.500 118.995 ;
        RECT 109.375 118.000 112.475 118.005 ;
        RECT 115.250 117.600 116.300 117.625 ;
        RECT 109.200 116.600 112.250 117.600 ;
        RECT 115.250 116.600 123.050 117.600 ;
        RECT 104.505 114.525 106.730 115.680 ;
        RECT 104.505 114.515 106.705 114.525 ;
        RECT 101.500 105.900 102.550 105.925 ;
        RECT 101.500 104.900 104.600 105.900 ;
        RECT 101.500 104.875 102.550 104.900 ;
        RECT 92.450 102.625 94.925 103.625 ;
        RECT 95.900 102.925 102.525 103.925 ;
        RECT 84.050 101.725 85.050 101.730 ;
        RECT 83.925 101.700 85.050 101.725 ;
        RECT 82.345 100.700 85.050 101.700 ;
        RECT 83.925 100.675 85.050 100.700 ;
        RECT 84.050 100.670 85.050 100.675 ;
        RECT 85.825 96.800 86.825 102.625 ;
        RECT 92.000 100.675 93.050 101.725 ;
        RECT 89.825 98.775 90.875 99.855 ;
        RECT 92.025 97.800 93.025 100.675 ;
        RECT 91.995 96.800 93.055 97.800 ;
        RECT 93.925 96.800 94.925 102.625 ;
        RECT 95.625 97.800 96.615 97.825 ;
        RECT 95.620 96.800 96.620 97.800 ;
        RECT 95.625 96.775 96.615 96.800 ;
        RECT 89.825 95.025 90.875 95.050 ;
        RECT 83.775 94.025 86.825 95.025 ;
        RECT 89.825 94.025 97.625 95.025 ;
        RECT 99.430 94.800 100.430 101.800 ;
        RECT 61.100 83.350 62.100 92.050 ;
        RECT 63.175 89.700 64.500 90.700 ;
        RECT 63.175 83.350 64.175 89.700 ;
        RECT 65.275 89.675 66.325 90.725 ;
        RECT 56.925 81.050 57.925 83.325 ;
        RECT 58.325 82.300 59.375 83.350 ;
        RECT 61.075 82.300 62.125 83.350 ;
        RECT 63.175 82.325 64.775 83.350 ;
        RECT 63.725 82.300 64.775 82.325 ;
        RECT 65.300 81.050 66.300 89.675 ;
        RECT 67.000 87.900 68.050 88.950 ;
        RECT 56.925 80.050 66.300 81.050 ;
        RECT 67.025 81.050 68.025 87.900 ;
        RECT 69.200 87.645 70.195 92.050 ;
        RECT 74.050 91.575 77.100 92.575 ;
        RECT 79.080 91.950 81.305 93.105 ;
        RECT 79.080 91.940 80.195 91.950 ;
        RECT 69.200 86.905 70.200 87.645 ;
        RECT 69.205 83.350 70.200 86.905 ;
        RECT 69.175 82.300 70.225 83.350 ;
        RECT 70.455 81.325 71.505 81.350 ;
        RECT 74.050 81.325 75.050 91.575 ;
        RECT 83.775 83.350 84.775 94.025 ;
        RECT 89.825 94.000 90.875 94.025 ;
        RECT 99.405 93.750 100.455 94.800 ;
        RECT 86.525 93.045 90.850 93.050 ;
        RECT 86.525 92.050 95.620 93.045 ;
        RECT 101.525 92.575 102.525 102.925 ;
        RECT 86.525 83.350 87.525 92.050 ;
        RECT 88.600 89.700 89.925 90.700 ;
        RECT 88.600 83.350 89.600 89.700 ;
        RECT 90.700 89.675 91.750 90.725 ;
        RECT 67.025 80.050 69.500 81.050 ;
        RECT 70.455 80.325 75.050 81.325 ;
        RECT 82.350 81.050 83.350 83.325 ;
        RECT 83.750 82.300 84.800 83.350 ;
        RECT 86.500 82.300 87.550 83.350 ;
        RECT 88.600 82.325 90.200 83.350 ;
        RECT 89.150 82.300 90.200 82.325 ;
        RECT 90.725 81.050 91.725 89.675 ;
        RECT 92.425 87.900 93.475 88.950 ;
        RECT 70.455 80.300 71.505 80.325 ;
        RECT 56.930 79.125 57.920 79.150 ;
        RECT 58.500 79.125 59.550 79.150 ;
        RECT 56.920 78.125 59.550 79.125 ;
        RECT 56.930 78.100 57.920 78.125 ;
        RECT 58.500 78.100 59.550 78.125 ;
        RECT 60.400 74.225 61.400 80.050 ;
        RECT 66.575 78.100 67.625 79.150 ;
        RECT 64.400 76.200 65.450 77.280 ;
        RECT 66.600 75.225 67.600 78.100 ;
        RECT 66.570 74.225 67.630 75.225 ;
        RECT 68.500 74.225 69.500 80.050 ;
        RECT 70.200 75.225 71.190 75.250 ;
        RECT 70.195 74.225 71.195 75.225 ;
        RECT 70.200 74.200 71.190 74.225 ;
        RECT 72.255 73.000 73.245 73.025 ;
        RECT 74.020 73.000 75.020 80.325 ;
        RECT 82.350 80.050 91.725 81.050 ;
        RECT 92.450 81.050 93.450 87.900 ;
        RECT 94.625 87.645 95.620 92.050 ;
        RECT 99.475 91.575 102.525 92.575 ;
        RECT 94.625 86.905 95.625 87.645 ;
        RECT 94.630 83.350 95.625 86.905 ;
        RECT 94.600 82.300 95.650 83.350 ;
        RECT 95.880 81.325 96.930 81.350 ;
        RECT 99.475 81.325 100.475 91.575 ;
        RECT 92.450 80.050 94.925 81.050 ;
        RECT 95.880 80.325 100.475 81.325 ;
        RECT 95.880 80.300 96.930 80.325 ;
        RECT 82.355 79.125 83.345 79.150 ;
        RECT 83.925 79.125 84.975 79.150 ;
        RECT 82.345 78.125 84.975 79.125 ;
        RECT 82.355 78.100 83.345 78.125 ;
        RECT 83.925 78.100 84.975 78.125 ;
        RECT 85.825 74.225 86.825 80.050 ;
        RECT 92.000 78.100 93.050 79.150 ;
        RECT 89.825 76.200 90.875 77.280 ;
        RECT 92.025 75.225 93.025 78.100 ;
        RECT 91.995 74.225 93.055 75.225 ;
        RECT 93.925 74.225 94.925 80.050 ;
        RECT 95.625 75.225 96.615 75.250 ;
        RECT 95.620 74.225 96.620 75.225 ;
        RECT 95.625 74.200 96.615 74.225 ;
        RECT 99.475 73.000 100.475 80.325 ;
        RECT 52.750 72.000 100.475 73.000 ;
        RECT 103.600 73.000 104.600 104.900 ;
        RECT 105.600 93.105 106.705 114.515 ;
        RECT 109.200 105.925 110.200 116.600 ;
        RECT 115.250 116.575 116.300 116.600 ;
        RECT 111.950 115.620 116.275 115.625 ;
        RECT 111.950 114.625 121.045 115.620 ;
        RECT 111.950 105.925 112.950 114.625 ;
        RECT 114.025 112.275 115.350 113.275 ;
        RECT 114.025 105.925 115.025 112.275 ;
        RECT 116.125 112.250 117.175 113.300 ;
        RECT 107.775 103.625 108.775 105.900 ;
        RECT 109.175 104.875 110.225 105.925 ;
        RECT 111.925 104.875 112.975 105.925 ;
        RECT 114.025 104.900 115.625 105.925 ;
        RECT 114.575 104.875 115.625 104.900 ;
        RECT 116.150 103.625 117.150 112.250 ;
        RECT 117.850 110.475 118.900 111.525 ;
        RECT 107.775 102.625 117.150 103.625 ;
        RECT 117.875 103.625 118.875 110.475 ;
        RECT 120.050 110.220 121.045 114.625 ;
        RECT 120.050 109.480 121.050 110.220 ;
        RECT 120.055 105.925 121.050 109.480 ;
        RECT 120.025 104.875 121.075 105.925 ;
        RECT 123.105 105.905 124.095 105.930 ;
        RECT 123.100 104.905 124.100 105.905 ;
        RECT 123.105 104.880 124.095 104.905 ;
        RECT 124.850 103.925 125.850 125.000 ;
        RECT 131.025 115.680 132.130 132.620 ;
        RECT 134.625 128.500 135.625 139.175 ;
        RECT 140.675 139.150 141.725 139.175 ;
        RECT 137.375 138.195 141.700 138.200 ;
        RECT 137.375 137.200 146.470 138.195 ;
        RECT 137.375 128.500 138.375 137.200 ;
        RECT 139.450 134.850 140.775 135.850 ;
        RECT 139.450 128.500 140.450 134.850 ;
        RECT 141.550 134.825 142.600 135.875 ;
        RECT 133.200 126.200 134.200 128.475 ;
        RECT 134.600 127.450 135.650 128.500 ;
        RECT 137.350 127.450 138.400 128.500 ;
        RECT 139.450 127.475 141.050 128.500 ;
        RECT 140.000 127.450 141.050 127.475 ;
        RECT 141.575 126.200 142.575 134.825 ;
        RECT 143.275 133.050 144.325 134.100 ;
        RECT 133.200 125.200 142.575 126.200 ;
        RECT 143.300 126.200 144.300 133.050 ;
        RECT 145.475 132.795 146.470 137.200 ;
        RECT 145.475 132.055 146.475 132.795 ;
        RECT 145.480 128.500 146.475 132.055 ;
        RECT 145.450 127.450 146.500 128.500 ;
        RECT 143.300 125.200 145.775 126.200 ;
        RECT 134.775 124.275 135.825 124.300 ;
        RECT 133.195 123.275 135.825 124.275 ;
        RECT 134.775 123.250 135.825 123.275 ;
        RECT 134.800 119.000 135.800 123.250 ;
        RECT 136.675 119.375 137.675 125.200 ;
        RECT 142.850 123.250 143.900 124.300 ;
        RECT 140.675 121.350 141.725 122.430 ;
        RECT 142.875 120.375 143.875 123.250 ;
        RECT 142.845 119.375 143.905 120.375 ;
        RECT 144.775 119.375 145.775 125.200 ;
        RECT 146.750 125.000 151.275 126.000 ;
        RECT 146.475 120.375 147.465 120.400 ;
        RECT 146.470 119.375 147.470 120.375 ;
        RECT 146.475 119.350 147.465 119.375 ;
        RECT 134.800 118.995 137.900 119.000 ;
        RECT 134.800 118.005 137.925 118.995 ;
        RECT 134.800 118.000 137.900 118.005 ;
        RECT 140.675 117.600 141.725 117.625 ;
        RECT 134.625 116.600 137.675 117.600 ;
        RECT 140.675 116.600 148.475 117.600 ;
        RECT 129.930 114.525 132.155 115.680 ;
        RECT 129.930 114.515 132.130 114.525 ;
        RECT 117.875 102.625 120.350 103.625 ;
        RECT 121.325 102.925 127.950 103.925 ;
        RECT 109.475 101.725 110.475 101.730 ;
        RECT 109.350 101.700 110.475 101.725 ;
        RECT 107.770 100.700 110.475 101.700 ;
        RECT 109.350 100.675 110.475 100.700 ;
        RECT 109.475 100.670 110.475 100.675 ;
        RECT 111.250 96.800 112.250 102.625 ;
        RECT 117.425 100.675 118.475 101.725 ;
        RECT 115.250 98.775 116.300 99.855 ;
        RECT 117.450 97.800 118.450 100.675 ;
        RECT 117.420 96.800 118.480 97.800 ;
        RECT 119.350 96.800 120.350 102.625 ;
        RECT 121.050 97.800 122.040 97.825 ;
        RECT 121.045 96.800 122.045 97.800 ;
        RECT 121.050 96.775 122.040 96.800 ;
        RECT 115.250 95.025 116.300 95.050 ;
        RECT 109.200 94.025 112.250 95.025 ;
        RECT 115.250 94.025 123.050 95.025 ;
        RECT 124.855 94.800 125.855 101.800 ;
        RECT 105.575 93.080 106.730 93.105 ;
        RECT 105.570 91.975 106.730 93.080 ;
        RECT 105.575 91.950 106.730 91.975 ;
        RECT 109.200 83.350 110.200 94.025 ;
        RECT 115.250 94.000 116.300 94.025 ;
        RECT 124.830 93.750 125.880 94.800 ;
        RECT 111.950 93.045 116.275 93.050 ;
        RECT 111.950 92.050 121.045 93.045 ;
        RECT 126.950 92.575 127.950 102.925 ;
        RECT 131.025 93.105 132.130 114.515 ;
        RECT 134.625 105.925 135.625 116.600 ;
        RECT 140.675 116.575 141.725 116.600 ;
        RECT 137.375 115.620 141.700 115.625 ;
        RECT 137.375 114.625 146.470 115.620 ;
        RECT 137.375 105.925 138.375 114.625 ;
        RECT 139.450 112.275 140.775 113.275 ;
        RECT 139.450 105.925 140.450 112.275 ;
        RECT 141.550 112.250 142.600 113.300 ;
        RECT 133.200 103.625 134.200 105.900 ;
        RECT 134.600 104.875 135.650 105.925 ;
        RECT 137.350 104.875 138.400 105.925 ;
        RECT 139.450 104.900 141.050 105.925 ;
        RECT 140.000 104.875 141.050 104.900 ;
        RECT 141.575 103.625 142.575 112.250 ;
        RECT 143.275 110.475 144.325 111.525 ;
        RECT 133.200 102.625 142.575 103.625 ;
        RECT 143.300 103.625 144.300 110.475 ;
        RECT 145.475 110.220 146.470 114.625 ;
        RECT 145.475 109.480 146.475 110.220 ;
        RECT 145.480 105.925 146.475 109.480 ;
        RECT 145.450 104.875 146.500 105.925 ;
        RECT 150.275 103.925 151.275 125.000 ;
        RECT 154.500 104.875 155.550 105.955 ;
        RECT 143.300 102.625 145.775 103.625 ;
        RECT 146.750 102.925 153.375 103.925 ;
        RECT 134.900 101.725 135.900 101.730 ;
        RECT 134.775 101.700 135.900 101.725 ;
        RECT 133.195 100.700 135.900 101.700 ;
        RECT 134.775 100.675 135.900 100.700 ;
        RECT 134.900 100.670 135.900 100.675 ;
        RECT 136.675 96.800 137.675 102.625 ;
        RECT 142.850 100.675 143.900 101.725 ;
        RECT 140.675 98.775 141.725 99.855 ;
        RECT 142.875 97.800 143.875 100.675 ;
        RECT 142.845 96.800 143.905 97.800 ;
        RECT 144.775 96.800 145.775 102.625 ;
        RECT 146.475 97.800 147.465 97.825 ;
        RECT 146.470 96.800 147.470 97.800 ;
        RECT 146.475 96.775 147.465 96.800 ;
        RECT 140.675 95.025 141.725 95.050 ;
        RECT 134.625 94.025 137.675 95.025 ;
        RECT 140.675 94.025 148.475 95.025 ;
        RECT 150.280 94.800 151.280 101.800 ;
        RECT 111.950 83.350 112.950 92.050 ;
        RECT 114.025 89.700 115.350 90.700 ;
        RECT 114.025 83.350 115.025 89.700 ;
        RECT 116.125 89.675 117.175 90.725 ;
        RECT 107.775 81.050 108.775 83.325 ;
        RECT 109.175 82.300 110.225 83.350 ;
        RECT 111.925 82.300 112.975 83.350 ;
        RECT 114.025 82.325 115.625 83.350 ;
        RECT 114.575 82.300 115.625 82.325 ;
        RECT 116.150 81.050 117.150 89.675 ;
        RECT 117.850 87.900 118.900 88.950 ;
        RECT 107.775 80.050 117.150 81.050 ;
        RECT 117.875 81.050 118.875 87.900 ;
        RECT 120.050 87.645 121.045 92.050 ;
        RECT 124.900 91.575 127.950 92.575 ;
        RECT 129.930 91.950 132.155 93.105 ;
        RECT 129.930 91.940 131.045 91.950 ;
        RECT 120.050 86.905 121.050 87.645 ;
        RECT 120.055 83.350 121.050 86.905 ;
        RECT 120.025 82.300 121.075 83.350 ;
        RECT 121.305 81.325 122.355 81.350 ;
        RECT 124.900 81.325 125.900 91.575 ;
        RECT 134.625 83.350 135.625 94.025 ;
        RECT 140.675 94.000 141.725 94.025 ;
        RECT 150.255 93.750 151.305 94.800 ;
        RECT 137.375 93.045 141.700 93.050 ;
        RECT 137.375 92.050 146.470 93.045 ;
        RECT 152.375 92.575 153.375 102.925 ;
        RECT 137.375 83.350 138.375 92.050 ;
        RECT 139.450 89.700 140.775 90.700 ;
        RECT 139.450 83.350 140.450 89.700 ;
        RECT 141.550 89.675 142.600 90.725 ;
        RECT 117.875 80.050 120.350 81.050 ;
        RECT 121.305 80.325 125.900 81.325 ;
        RECT 133.200 81.050 134.200 83.325 ;
        RECT 134.600 82.300 135.650 83.350 ;
        RECT 137.350 82.300 138.400 83.350 ;
        RECT 139.450 82.325 141.050 83.350 ;
        RECT 140.000 82.300 141.050 82.325 ;
        RECT 141.575 81.050 142.575 89.675 ;
        RECT 143.275 87.900 144.325 88.950 ;
        RECT 121.305 80.300 122.355 80.325 ;
        RECT 107.780 79.125 108.770 79.150 ;
        RECT 109.350 79.125 110.400 79.150 ;
        RECT 107.770 78.125 110.400 79.125 ;
        RECT 107.780 78.100 108.770 78.125 ;
        RECT 109.350 78.100 110.400 78.125 ;
        RECT 111.250 74.225 112.250 80.050 ;
        RECT 117.425 78.100 118.475 79.150 ;
        RECT 115.250 76.200 116.300 77.280 ;
        RECT 117.450 75.225 118.450 78.100 ;
        RECT 117.420 74.225 118.480 75.225 ;
        RECT 119.350 74.225 120.350 80.050 ;
        RECT 121.050 75.225 122.040 75.250 ;
        RECT 121.045 74.225 122.045 75.225 ;
        RECT 121.050 74.200 122.040 74.225 ;
        RECT 123.105 73.000 124.095 73.025 ;
        RECT 124.870 73.000 125.870 80.325 ;
        RECT 133.200 80.050 142.575 81.050 ;
        RECT 143.300 81.050 144.300 87.900 ;
        RECT 145.475 87.645 146.470 92.050 ;
        RECT 150.325 91.575 153.375 92.575 ;
        RECT 145.475 86.905 146.475 87.645 ;
        RECT 145.480 83.350 146.475 86.905 ;
        RECT 145.450 82.300 146.500 83.350 ;
        RECT 146.730 81.325 147.780 81.350 ;
        RECT 150.325 81.325 151.325 91.575 ;
        RECT 143.300 80.050 145.775 81.050 ;
        RECT 146.730 80.325 151.325 81.325 ;
        RECT 146.730 80.300 147.780 80.325 ;
        RECT 133.205 79.125 134.195 79.150 ;
        RECT 134.775 79.125 135.825 79.150 ;
        RECT 133.195 78.125 135.825 79.125 ;
        RECT 133.205 78.100 134.195 78.125 ;
        RECT 134.775 78.100 135.825 78.125 ;
        RECT 136.675 74.225 137.675 80.050 ;
        RECT 142.850 78.100 143.900 79.150 ;
        RECT 140.675 76.200 141.725 77.280 ;
        RECT 142.875 75.225 143.875 78.100 ;
        RECT 142.845 74.225 143.905 75.225 ;
        RECT 144.775 74.225 145.775 80.050 ;
        RECT 146.475 75.225 147.465 75.250 ;
        RECT 146.470 74.225 147.470 75.225 ;
        RECT 146.475 74.200 147.465 74.225 ;
        RECT 150.325 73.000 151.325 80.325 ;
        RECT 103.600 72.000 151.325 73.000 ;
        RECT 21.405 71.975 22.395 72.000 ;
        RECT 72.255 71.975 73.245 72.000 ;
        RECT 123.105 71.975 124.095 72.000 ;
        RECT 48.830 70.550 49.820 70.575 ;
        RECT 13.550 68.175 14.600 68.200 ;
        RECT 7.500 67.175 10.550 68.175 ;
        RECT 13.550 67.175 21.350 68.175 ;
        RECT 23.520 67.200 24.520 70.550 ;
        RECT 48.825 69.550 49.825 70.550 ;
        RECT 48.830 69.525 49.820 69.550 ;
        RECT 38.975 68.175 40.025 68.200 ;
        RECT 64.400 68.175 65.450 68.200 ;
        RECT 2.805 66.225 3.920 66.255 ;
        RECT 5.970 66.225 7.125 66.250 ;
        RECT 2.805 65.120 7.125 66.225 ;
        RECT 2.805 65.090 3.920 65.120 ;
        RECT 5.970 65.095 7.125 65.120 ;
        RECT 5.995 61.755 7.100 65.095 ;
        RECT 3.900 60.650 7.100 61.755 ;
        RECT 3.900 43.680 5.005 60.650 ;
        RECT 7.500 56.500 8.500 67.175 ;
        RECT 13.550 67.150 14.600 67.175 ;
        RECT 10.250 66.195 14.575 66.200 ;
        RECT 10.250 65.200 19.345 66.195 ;
        RECT 23.495 66.150 24.545 67.200 ;
        RECT 32.925 67.175 35.975 68.175 ;
        RECT 38.975 67.175 46.775 68.175 ;
        RECT 58.350 67.175 61.400 68.175 ;
        RECT 64.400 67.175 72.200 68.175 ;
        RECT 74.370 67.200 75.370 70.550 ;
        RECT 89.825 68.175 90.875 68.200 ;
        RECT 115.250 68.175 116.300 68.200 ;
        RECT 26.220 66.295 27.270 66.320 ;
        RECT 25.400 66.290 27.270 66.295 ;
        RECT 25.375 65.300 27.270 66.290 ;
        RECT 25.400 65.295 27.270 65.300 ;
        RECT 26.220 65.270 27.270 65.295 ;
        RECT 10.250 56.500 11.250 65.200 ;
        RECT 14.425 63.850 15.475 63.875 ;
        RECT 16.150 63.850 17.200 64.365 ;
        RECT 12.325 62.850 13.650 63.850 ;
        RECT 14.425 62.850 17.200 63.850 ;
        RECT 12.325 56.500 13.325 62.850 ;
        RECT 14.425 62.825 15.475 62.850 ;
        RECT 6.075 54.200 7.075 56.475 ;
        RECT 7.475 55.450 8.525 56.500 ;
        RECT 10.225 55.450 11.275 56.500 ;
        RECT 12.325 55.475 13.925 56.500 ;
        RECT 12.875 55.450 13.925 55.475 ;
        RECT 14.450 54.200 15.450 62.825 ;
        RECT 16.150 61.050 17.200 62.100 ;
        RECT 6.075 53.200 15.450 54.200 ;
        RECT 16.175 54.200 17.175 61.050 ;
        RECT 18.350 60.795 19.345 65.200 ;
        RECT 28.110 64.420 30.670 65.525 ;
        RECT 31.395 65.095 32.550 66.250 ;
        RECT 20.345 61.155 21.345 64.340 ;
        RECT 28.110 63.695 29.215 64.420 ;
        RECT 24.815 62.590 29.215 63.695 ;
        RECT 24.815 61.180 25.920 62.590 ;
        RECT 28.230 61.755 29.345 61.785 ;
        RECT 31.420 61.755 32.525 65.095 ;
        RECT 24.795 61.155 25.950 61.180 ;
        RECT 18.350 60.055 19.350 60.795 ;
        RECT 20.345 60.100 25.950 61.155 ;
        RECT 28.230 60.650 32.525 61.755 ;
        RECT 28.230 60.620 30.430 60.650 ;
        RECT 18.355 56.500 19.350 60.055 ;
        RECT 20.370 60.050 25.950 60.100 ;
        RECT 24.795 60.025 25.950 60.050 ;
        RECT 18.325 55.450 19.375 56.500 ;
        RECT 23.405 56.480 24.395 56.505 ;
        RECT 23.400 55.480 24.400 56.480 ;
        RECT 23.405 55.455 24.395 55.480 ;
        RECT 16.175 53.200 18.650 54.200 ;
        RECT 7.650 52.275 8.700 52.300 ;
        RECT 6.070 51.275 8.700 52.275 ;
        RECT 7.650 51.250 8.700 51.275 ;
        RECT 7.675 47.000 8.675 51.250 ;
        RECT 9.550 47.375 10.550 53.200 ;
        RECT 15.725 51.250 16.775 52.300 ;
        RECT 13.550 49.350 14.600 50.430 ;
        RECT 15.750 48.375 16.750 51.250 ;
        RECT 15.720 47.375 16.780 48.375 ;
        RECT 17.650 47.375 18.650 53.200 ;
        RECT 19.625 53.000 24.150 54.000 ;
        RECT 19.350 48.375 20.340 48.400 ;
        RECT 19.345 47.375 20.345 48.375 ;
        RECT 19.350 47.350 20.340 47.375 ;
        RECT 7.675 46.995 10.775 47.000 ;
        RECT 7.675 46.005 10.800 46.995 ;
        RECT 7.675 46.000 10.775 46.005 ;
        RECT 13.550 45.600 14.600 45.625 ;
        RECT 7.500 44.600 10.550 45.600 ;
        RECT 13.550 44.600 21.350 45.600 ;
        RECT 2.805 42.525 5.030 43.680 ;
        RECT 2.805 42.515 5.005 42.525 ;
        RECT 3.900 21.105 5.005 42.515 ;
        RECT 7.500 33.925 8.500 44.600 ;
        RECT 13.550 44.575 14.600 44.600 ;
        RECT 10.250 43.620 14.575 43.625 ;
        RECT 10.250 42.625 19.345 43.620 ;
        RECT 10.250 33.925 11.250 42.625 ;
        RECT 12.325 40.275 13.650 41.275 ;
        RECT 12.325 33.925 13.325 40.275 ;
        RECT 14.425 40.250 15.475 41.300 ;
        RECT 6.075 31.625 7.075 33.900 ;
        RECT 7.475 32.875 8.525 33.925 ;
        RECT 10.225 32.875 11.275 33.925 ;
        RECT 12.325 32.900 13.925 33.925 ;
        RECT 12.875 32.875 13.925 32.900 ;
        RECT 14.450 31.625 15.450 40.250 ;
        RECT 16.150 38.475 17.200 39.525 ;
        RECT 6.075 30.625 15.450 31.625 ;
        RECT 16.175 31.625 17.175 38.475 ;
        RECT 18.350 38.220 19.345 42.625 ;
        RECT 18.350 37.480 19.350 38.220 ;
        RECT 18.355 33.925 19.350 37.480 ;
        RECT 18.325 32.875 19.375 33.925 ;
        RECT 21.405 33.905 22.395 33.930 ;
        RECT 21.400 32.905 22.400 33.905 ;
        RECT 21.405 32.880 22.395 32.905 ;
        RECT 23.150 31.925 24.150 53.000 ;
        RECT 29.325 43.680 30.430 60.620 ;
        RECT 32.925 56.500 33.925 67.175 ;
        RECT 38.975 67.150 40.025 67.175 ;
        RECT 53.655 66.225 54.770 66.255 ;
        RECT 56.820 66.225 57.975 66.250 ;
        RECT 35.675 66.195 40.000 66.200 ;
        RECT 35.675 65.200 44.770 66.195 ;
        RECT 35.675 56.500 36.675 65.200 ;
        RECT 37.750 62.850 39.075 63.850 ;
        RECT 37.750 56.500 38.750 62.850 ;
        RECT 39.850 62.825 40.900 63.875 ;
        RECT 31.500 54.200 32.500 56.475 ;
        RECT 32.900 55.450 33.950 56.500 ;
        RECT 35.650 55.450 36.700 56.500 ;
        RECT 37.750 55.475 39.350 56.500 ;
        RECT 38.300 55.450 39.350 55.475 ;
        RECT 39.875 54.200 40.875 62.825 ;
        RECT 41.575 61.050 42.625 62.100 ;
        RECT 31.500 53.200 40.875 54.200 ;
        RECT 41.600 54.200 42.600 61.050 ;
        RECT 43.775 60.795 44.770 65.200 ;
        RECT 53.655 65.120 57.975 66.225 ;
        RECT 53.655 65.090 54.770 65.120 ;
        RECT 56.820 65.095 57.975 65.120 ;
        RECT 56.845 61.755 57.950 65.095 ;
        RECT 43.775 60.055 44.775 60.795 ;
        RECT 43.780 56.500 44.775 60.055 ;
        RECT 54.750 60.650 57.950 61.755 ;
        RECT 43.750 55.450 44.800 56.500 ;
        RECT 46.825 56.470 47.825 56.475 ;
        RECT 46.800 55.480 47.850 56.470 ;
        RECT 46.825 55.475 47.825 55.480 ;
        RECT 41.600 53.200 44.075 54.200 ;
        RECT 33.075 52.275 34.125 52.300 ;
        RECT 31.495 51.275 34.125 52.275 ;
        RECT 33.075 51.250 34.125 51.275 ;
        RECT 33.100 47.000 34.100 51.250 ;
        RECT 34.975 47.375 35.975 53.200 ;
        RECT 41.150 51.250 42.200 52.300 ;
        RECT 38.975 49.350 40.025 50.430 ;
        RECT 41.175 48.375 42.175 51.250 ;
        RECT 41.145 47.375 42.205 48.375 ;
        RECT 43.075 47.375 44.075 53.200 ;
        RECT 45.050 53.000 49.575 54.000 ;
        RECT 44.775 48.375 45.765 48.400 ;
        RECT 44.770 47.375 45.770 48.375 ;
        RECT 44.775 47.350 45.765 47.375 ;
        RECT 33.100 46.995 36.200 47.000 ;
        RECT 33.100 46.005 36.225 46.995 ;
        RECT 33.100 46.000 36.200 46.005 ;
        RECT 38.975 45.600 40.025 45.625 ;
        RECT 32.925 44.600 35.975 45.600 ;
        RECT 38.975 44.600 46.775 45.600 ;
        RECT 28.230 42.525 30.455 43.680 ;
        RECT 28.230 42.515 30.430 42.525 ;
        RECT 16.175 30.625 18.650 31.625 ;
        RECT 19.625 30.925 26.250 31.925 ;
        RECT 7.775 29.725 8.775 29.730 ;
        RECT 7.650 29.700 8.775 29.725 ;
        RECT 6.070 28.700 8.775 29.700 ;
        RECT 7.650 28.675 8.775 28.700 ;
        RECT 7.775 28.670 8.775 28.675 ;
        RECT 9.550 24.800 10.550 30.625 ;
        RECT 15.725 28.675 16.775 29.725 ;
        RECT 13.550 26.775 14.600 27.855 ;
        RECT 15.750 25.800 16.750 28.675 ;
        RECT 15.720 24.800 16.780 25.800 ;
        RECT 17.650 24.800 18.650 30.625 ;
        RECT 19.350 25.800 20.340 25.825 ;
        RECT 19.345 24.800 20.345 25.800 ;
        RECT 19.350 24.775 20.340 24.800 ;
        RECT 13.550 23.025 14.600 23.050 ;
        RECT 7.500 22.025 10.550 23.025 ;
        RECT 13.550 22.025 21.350 23.025 ;
        RECT 23.155 22.800 24.155 29.800 ;
        RECT 3.875 21.080 5.030 21.105 ;
        RECT 3.870 19.975 5.030 21.080 ;
        RECT 3.875 19.950 5.030 19.975 ;
        RECT 7.500 11.350 8.500 22.025 ;
        RECT 13.550 22.000 14.600 22.025 ;
        RECT 23.130 21.750 24.180 22.800 ;
        RECT 10.250 21.045 14.575 21.050 ;
        RECT 10.250 20.050 19.345 21.045 ;
        RECT 25.250 20.575 26.250 30.925 ;
        RECT 29.325 21.105 30.430 42.515 ;
        RECT 32.925 33.925 33.925 44.600 ;
        RECT 38.975 44.575 40.025 44.600 ;
        RECT 35.675 43.620 40.000 43.625 ;
        RECT 35.675 42.625 44.770 43.620 ;
        RECT 35.675 33.925 36.675 42.625 ;
        RECT 37.750 40.275 39.075 41.275 ;
        RECT 37.750 33.925 38.750 40.275 ;
        RECT 39.850 40.250 40.900 41.300 ;
        RECT 31.500 31.625 32.500 33.900 ;
        RECT 32.900 32.875 33.950 33.925 ;
        RECT 35.650 32.875 36.700 33.925 ;
        RECT 37.750 32.900 39.350 33.925 ;
        RECT 38.300 32.875 39.350 32.900 ;
        RECT 39.875 31.625 40.875 40.250 ;
        RECT 41.575 38.475 42.625 39.525 ;
        RECT 31.500 30.625 40.875 31.625 ;
        RECT 41.600 31.625 42.600 38.475 ;
        RECT 43.775 38.220 44.770 42.625 ;
        RECT 43.775 37.480 44.775 38.220 ;
        RECT 43.780 33.925 44.775 37.480 ;
        RECT 43.750 32.875 44.800 33.925 ;
        RECT 48.575 31.925 49.575 53.000 ;
        RECT 54.750 43.680 55.855 60.650 ;
        RECT 58.350 56.500 59.350 67.175 ;
        RECT 64.400 67.150 65.450 67.175 ;
        RECT 61.100 66.195 65.425 66.200 ;
        RECT 61.100 65.200 70.195 66.195 ;
        RECT 74.345 66.150 75.395 67.200 ;
        RECT 83.775 67.175 86.825 68.175 ;
        RECT 89.825 67.175 97.625 68.175 ;
        RECT 109.200 67.175 112.250 68.175 ;
        RECT 115.250 67.175 123.050 68.175 ;
        RECT 125.220 67.200 126.220 70.550 ;
        RECT 140.675 68.175 141.725 68.200 ;
        RECT 77.070 66.295 78.120 66.320 ;
        RECT 76.250 66.290 78.120 66.295 ;
        RECT 76.225 65.300 78.120 66.290 ;
        RECT 76.250 65.295 78.120 65.300 ;
        RECT 77.070 65.270 78.120 65.295 ;
        RECT 61.100 56.500 62.100 65.200 ;
        RECT 65.275 63.850 66.325 63.875 ;
        RECT 67.000 63.850 68.050 64.365 ;
        RECT 63.175 62.850 64.500 63.850 ;
        RECT 65.275 62.850 68.050 63.850 ;
        RECT 63.175 56.500 64.175 62.850 ;
        RECT 65.275 62.825 66.325 62.850 ;
        RECT 56.925 54.200 57.925 56.475 ;
        RECT 58.325 55.450 59.375 56.500 ;
        RECT 61.075 55.450 62.125 56.500 ;
        RECT 63.175 55.475 64.775 56.500 ;
        RECT 63.725 55.450 64.775 55.475 ;
        RECT 65.300 54.200 66.300 62.825 ;
        RECT 67.000 61.050 68.050 62.100 ;
        RECT 56.925 53.200 66.300 54.200 ;
        RECT 67.025 54.200 68.025 61.050 ;
        RECT 69.200 60.795 70.195 65.200 ;
        RECT 78.960 64.420 81.520 65.525 ;
        RECT 82.245 65.095 83.400 66.250 ;
        RECT 71.195 61.155 72.195 64.340 ;
        RECT 78.960 63.695 80.065 64.420 ;
        RECT 75.665 62.590 80.065 63.695 ;
        RECT 75.665 61.180 76.770 62.590 ;
        RECT 79.080 61.755 80.195 61.785 ;
        RECT 82.270 61.755 83.375 65.095 ;
        RECT 75.645 61.155 76.800 61.180 ;
        RECT 69.200 60.055 70.200 60.795 ;
        RECT 71.195 60.100 76.800 61.155 ;
        RECT 79.080 60.650 83.375 61.755 ;
        RECT 79.080 60.620 81.280 60.650 ;
        RECT 69.205 56.500 70.200 60.055 ;
        RECT 71.220 60.050 76.800 60.100 ;
        RECT 75.645 60.025 76.800 60.050 ;
        RECT 69.175 55.450 70.225 56.500 ;
        RECT 74.255 56.480 75.245 56.505 ;
        RECT 74.250 55.480 75.250 56.480 ;
        RECT 74.255 55.455 75.245 55.480 ;
        RECT 67.025 53.200 69.500 54.200 ;
        RECT 58.500 52.275 59.550 52.300 ;
        RECT 56.920 51.275 59.550 52.275 ;
        RECT 58.500 51.250 59.550 51.275 ;
        RECT 58.525 47.000 59.525 51.250 ;
        RECT 60.400 47.375 61.400 53.200 ;
        RECT 66.575 51.250 67.625 52.300 ;
        RECT 64.400 49.350 65.450 50.430 ;
        RECT 66.600 48.375 67.600 51.250 ;
        RECT 66.570 47.375 67.630 48.375 ;
        RECT 68.500 47.375 69.500 53.200 ;
        RECT 70.475 53.000 75.000 54.000 ;
        RECT 70.200 48.375 71.190 48.400 ;
        RECT 70.195 47.375 71.195 48.375 ;
        RECT 70.200 47.350 71.190 47.375 ;
        RECT 58.525 46.995 61.625 47.000 ;
        RECT 58.525 46.005 61.650 46.995 ;
        RECT 58.525 46.000 61.625 46.005 ;
        RECT 64.400 45.600 65.450 45.625 ;
        RECT 58.350 44.600 61.400 45.600 ;
        RECT 64.400 44.600 72.200 45.600 ;
        RECT 53.655 42.525 55.880 43.680 ;
        RECT 53.655 42.515 55.855 42.525 ;
        RECT 50.650 33.900 51.700 33.925 ;
        RECT 50.650 32.900 53.750 33.900 ;
        RECT 50.650 32.875 51.700 32.900 ;
        RECT 41.600 30.625 44.075 31.625 ;
        RECT 45.050 30.925 51.675 31.925 ;
        RECT 33.200 29.725 34.200 29.730 ;
        RECT 33.075 29.700 34.200 29.725 ;
        RECT 31.495 28.700 34.200 29.700 ;
        RECT 33.075 28.675 34.200 28.700 ;
        RECT 33.200 28.670 34.200 28.675 ;
        RECT 34.975 24.800 35.975 30.625 ;
        RECT 41.150 28.675 42.200 29.725 ;
        RECT 38.975 26.775 40.025 27.855 ;
        RECT 41.175 25.800 42.175 28.675 ;
        RECT 41.145 24.800 42.205 25.800 ;
        RECT 43.075 24.800 44.075 30.625 ;
        RECT 44.775 25.800 45.765 25.825 ;
        RECT 44.770 24.800 45.770 25.800 ;
        RECT 44.775 24.775 45.765 24.800 ;
        RECT 38.975 23.025 40.025 23.050 ;
        RECT 32.925 22.025 35.975 23.025 ;
        RECT 38.975 22.025 46.775 23.025 ;
        RECT 48.580 22.800 49.580 29.800 ;
        RECT 10.250 11.350 11.250 20.050 ;
        RECT 12.325 17.700 13.650 18.700 ;
        RECT 12.325 11.350 13.325 17.700 ;
        RECT 14.425 17.675 15.475 18.725 ;
        RECT 6.075 9.050 7.075 11.325 ;
        RECT 7.475 10.300 8.525 11.350 ;
        RECT 10.225 10.300 11.275 11.350 ;
        RECT 12.325 10.325 13.925 11.350 ;
        RECT 12.875 10.300 13.925 10.325 ;
        RECT 14.450 9.050 15.450 17.675 ;
        RECT 16.150 15.900 17.200 16.950 ;
        RECT 6.075 8.050 15.450 9.050 ;
        RECT 16.175 9.050 17.175 15.900 ;
        RECT 18.350 15.645 19.345 20.050 ;
        RECT 23.200 19.575 26.250 20.575 ;
        RECT 28.230 19.950 30.455 21.105 ;
        RECT 28.230 19.940 29.345 19.950 ;
        RECT 18.350 14.905 19.350 15.645 ;
        RECT 18.355 11.350 19.350 14.905 ;
        RECT 18.325 10.300 19.375 11.350 ;
        RECT 19.605 9.325 20.655 9.350 ;
        RECT 23.200 9.325 24.200 19.575 ;
        RECT 32.925 11.350 33.925 22.025 ;
        RECT 38.975 22.000 40.025 22.025 ;
        RECT 48.555 21.750 49.605 22.800 ;
        RECT 35.675 21.045 40.000 21.050 ;
        RECT 35.675 20.050 44.770 21.045 ;
        RECT 50.675 20.575 51.675 30.925 ;
        RECT 35.675 11.350 36.675 20.050 ;
        RECT 37.750 17.700 39.075 18.700 ;
        RECT 37.750 11.350 38.750 17.700 ;
        RECT 39.850 17.675 40.900 18.725 ;
        RECT 16.175 8.050 18.650 9.050 ;
        RECT 19.605 8.325 24.200 9.325 ;
        RECT 31.500 9.050 32.500 11.325 ;
        RECT 32.900 10.300 33.950 11.350 ;
        RECT 35.650 10.300 36.700 11.350 ;
        RECT 37.750 10.325 39.350 11.350 ;
        RECT 38.300 10.300 39.350 10.325 ;
        RECT 39.875 9.050 40.875 17.675 ;
        RECT 41.575 15.900 42.625 16.950 ;
        RECT 19.605 8.300 20.655 8.325 ;
        RECT 6.080 7.125 7.070 7.150 ;
        RECT 7.650 7.125 8.700 7.150 ;
        RECT 6.070 6.125 8.700 7.125 ;
        RECT 6.080 6.100 7.070 6.125 ;
        RECT 7.650 6.100 8.700 6.125 ;
        RECT 9.550 2.225 10.550 8.050 ;
        RECT 15.725 6.100 16.775 7.150 ;
        RECT 13.550 4.200 14.600 5.280 ;
        RECT 15.750 3.225 16.750 6.100 ;
        RECT 15.720 2.225 16.780 3.225 ;
        RECT 17.650 2.225 18.650 8.050 ;
        RECT 19.350 3.225 20.340 3.250 ;
        RECT 19.345 2.225 20.345 3.225 ;
        RECT 19.350 2.200 20.340 2.225 ;
        RECT 23.170 1.000 24.170 8.325 ;
        RECT 31.500 8.050 40.875 9.050 ;
        RECT 41.600 9.050 42.600 15.900 ;
        RECT 43.775 15.645 44.770 20.050 ;
        RECT 48.625 19.575 51.675 20.575 ;
        RECT 43.775 14.905 44.775 15.645 ;
        RECT 43.780 11.350 44.775 14.905 ;
        RECT 43.750 10.300 44.800 11.350 ;
        RECT 45.030 9.325 46.080 9.350 ;
        RECT 48.625 9.325 49.625 19.575 ;
        RECT 41.600 8.050 44.075 9.050 ;
        RECT 45.030 8.325 49.625 9.325 ;
        RECT 45.030 8.300 46.080 8.325 ;
        RECT 31.505 7.125 32.495 7.150 ;
        RECT 33.075 7.125 34.125 7.150 ;
        RECT 31.495 6.125 34.125 7.125 ;
        RECT 31.505 6.100 32.495 6.125 ;
        RECT 33.075 6.100 34.125 6.125 ;
        RECT 34.975 2.225 35.975 8.050 ;
        RECT 41.150 6.100 42.200 7.150 ;
        RECT 38.975 4.200 40.025 5.280 ;
        RECT 41.175 3.225 42.175 6.100 ;
        RECT 41.145 2.225 42.205 3.225 ;
        RECT 43.075 2.225 44.075 8.050 ;
        RECT 44.775 3.225 45.765 3.250 ;
        RECT 44.770 2.225 45.770 3.225 ;
        RECT 44.775 2.200 45.765 2.225 ;
        RECT 48.625 1.000 49.625 8.325 ;
        RECT 23.170 0.000 49.625 1.000 ;
        RECT 52.750 1.000 53.750 32.900 ;
        RECT 54.750 21.105 55.855 42.515 ;
        RECT 58.350 33.925 59.350 44.600 ;
        RECT 64.400 44.575 65.450 44.600 ;
        RECT 61.100 43.620 65.425 43.625 ;
        RECT 61.100 42.625 70.195 43.620 ;
        RECT 61.100 33.925 62.100 42.625 ;
        RECT 63.175 40.275 64.500 41.275 ;
        RECT 63.175 33.925 64.175 40.275 ;
        RECT 65.275 40.250 66.325 41.300 ;
        RECT 56.925 31.625 57.925 33.900 ;
        RECT 58.325 32.875 59.375 33.925 ;
        RECT 61.075 32.875 62.125 33.925 ;
        RECT 63.175 32.900 64.775 33.925 ;
        RECT 63.725 32.875 64.775 32.900 ;
        RECT 65.300 31.625 66.300 40.250 ;
        RECT 67.000 38.475 68.050 39.525 ;
        RECT 56.925 30.625 66.300 31.625 ;
        RECT 67.025 31.625 68.025 38.475 ;
        RECT 69.200 38.220 70.195 42.625 ;
        RECT 69.200 37.480 70.200 38.220 ;
        RECT 69.205 33.925 70.200 37.480 ;
        RECT 69.175 32.875 70.225 33.925 ;
        RECT 72.255 33.905 73.245 33.930 ;
        RECT 72.250 32.905 73.250 33.905 ;
        RECT 72.255 32.880 73.245 32.905 ;
        RECT 74.000 31.925 75.000 53.000 ;
        RECT 80.175 43.680 81.280 60.620 ;
        RECT 83.775 56.500 84.775 67.175 ;
        RECT 89.825 67.150 90.875 67.175 ;
        RECT 104.505 66.225 105.620 66.255 ;
        RECT 107.670 66.225 108.825 66.250 ;
        RECT 86.525 66.195 90.850 66.200 ;
        RECT 86.525 65.200 95.620 66.195 ;
        RECT 86.525 56.500 87.525 65.200 ;
        RECT 88.600 62.850 89.925 63.850 ;
        RECT 88.600 56.500 89.600 62.850 ;
        RECT 90.700 62.825 91.750 63.875 ;
        RECT 82.350 54.200 83.350 56.475 ;
        RECT 83.750 55.450 84.800 56.500 ;
        RECT 86.500 55.450 87.550 56.500 ;
        RECT 88.600 55.475 90.200 56.500 ;
        RECT 89.150 55.450 90.200 55.475 ;
        RECT 90.725 54.200 91.725 62.825 ;
        RECT 92.425 61.050 93.475 62.100 ;
        RECT 82.350 53.200 91.725 54.200 ;
        RECT 92.450 54.200 93.450 61.050 ;
        RECT 94.625 60.795 95.620 65.200 ;
        RECT 104.505 65.120 108.825 66.225 ;
        RECT 104.505 65.090 105.620 65.120 ;
        RECT 107.670 65.095 108.825 65.120 ;
        RECT 107.695 61.755 108.800 65.095 ;
        RECT 94.625 60.055 95.625 60.795 ;
        RECT 94.630 56.500 95.625 60.055 ;
        RECT 105.600 60.650 108.800 61.755 ;
        RECT 94.600 55.450 95.650 56.500 ;
        RECT 92.450 53.200 94.925 54.200 ;
        RECT 83.925 52.275 84.975 52.300 ;
        RECT 82.345 51.275 84.975 52.275 ;
        RECT 83.925 51.250 84.975 51.275 ;
        RECT 83.950 47.000 84.950 51.250 ;
        RECT 85.825 47.375 86.825 53.200 ;
        RECT 92.000 51.250 93.050 52.300 ;
        RECT 89.825 49.350 90.875 50.430 ;
        RECT 92.025 48.375 93.025 51.250 ;
        RECT 91.995 47.375 93.055 48.375 ;
        RECT 93.925 47.375 94.925 53.200 ;
        RECT 95.900 53.000 100.425 54.000 ;
        RECT 95.625 48.375 96.615 48.400 ;
        RECT 95.620 47.375 96.620 48.375 ;
        RECT 95.625 47.350 96.615 47.375 ;
        RECT 83.950 46.995 87.050 47.000 ;
        RECT 83.950 46.005 87.075 46.995 ;
        RECT 83.950 46.000 87.050 46.005 ;
        RECT 89.825 45.600 90.875 45.625 ;
        RECT 83.775 44.600 86.825 45.600 ;
        RECT 89.825 44.600 97.625 45.600 ;
        RECT 79.080 42.525 81.305 43.680 ;
        RECT 79.080 42.515 81.280 42.525 ;
        RECT 67.025 30.625 69.500 31.625 ;
        RECT 70.475 30.925 77.100 31.925 ;
        RECT 58.625 29.725 59.625 29.730 ;
        RECT 58.500 29.700 59.625 29.725 ;
        RECT 56.920 28.700 59.625 29.700 ;
        RECT 58.500 28.675 59.625 28.700 ;
        RECT 58.625 28.670 59.625 28.675 ;
        RECT 60.400 24.800 61.400 30.625 ;
        RECT 66.575 28.675 67.625 29.725 ;
        RECT 64.400 26.775 65.450 27.855 ;
        RECT 66.600 25.800 67.600 28.675 ;
        RECT 66.570 24.800 67.630 25.800 ;
        RECT 68.500 24.800 69.500 30.625 ;
        RECT 70.200 25.800 71.190 25.825 ;
        RECT 70.195 24.800 71.195 25.800 ;
        RECT 70.200 24.775 71.190 24.800 ;
        RECT 64.400 23.025 65.450 23.050 ;
        RECT 58.350 22.025 61.400 23.025 ;
        RECT 64.400 22.025 72.200 23.025 ;
        RECT 74.005 22.800 75.005 29.800 ;
        RECT 54.725 21.080 55.880 21.105 ;
        RECT 54.720 19.975 55.880 21.080 ;
        RECT 54.725 19.950 55.880 19.975 ;
        RECT 58.350 11.350 59.350 22.025 ;
        RECT 64.400 22.000 65.450 22.025 ;
        RECT 73.980 21.750 75.030 22.800 ;
        RECT 61.100 21.045 65.425 21.050 ;
        RECT 61.100 20.050 70.195 21.045 ;
        RECT 76.100 20.575 77.100 30.925 ;
        RECT 80.175 21.105 81.280 42.515 ;
        RECT 83.775 33.925 84.775 44.600 ;
        RECT 89.825 44.575 90.875 44.600 ;
        RECT 86.525 43.620 90.850 43.625 ;
        RECT 86.525 42.625 95.620 43.620 ;
        RECT 86.525 33.925 87.525 42.625 ;
        RECT 88.600 40.275 89.925 41.275 ;
        RECT 88.600 33.925 89.600 40.275 ;
        RECT 90.700 40.250 91.750 41.300 ;
        RECT 82.350 31.625 83.350 33.900 ;
        RECT 83.750 32.875 84.800 33.925 ;
        RECT 86.500 32.875 87.550 33.925 ;
        RECT 88.600 32.900 90.200 33.925 ;
        RECT 89.150 32.875 90.200 32.900 ;
        RECT 90.725 31.625 91.725 40.250 ;
        RECT 92.425 38.475 93.475 39.525 ;
        RECT 82.350 30.625 91.725 31.625 ;
        RECT 92.450 31.625 93.450 38.475 ;
        RECT 94.625 38.220 95.620 42.625 ;
        RECT 94.625 37.480 95.625 38.220 ;
        RECT 94.630 33.925 95.625 37.480 ;
        RECT 94.600 32.875 95.650 33.925 ;
        RECT 99.425 31.925 100.425 53.000 ;
        RECT 105.600 43.680 106.705 60.650 ;
        RECT 109.200 56.500 110.200 67.175 ;
        RECT 115.250 67.150 116.300 67.175 ;
        RECT 111.950 66.195 116.275 66.200 ;
        RECT 111.950 65.200 121.045 66.195 ;
        RECT 125.195 66.150 126.245 67.200 ;
        RECT 134.625 67.175 137.675 68.175 ;
        RECT 140.675 67.175 148.475 68.175 ;
        RECT 127.920 66.295 128.970 66.320 ;
        RECT 127.100 66.290 128.970 66.295 ;
        RECT 127.075 65.300 128.970 66.290 ;
        RECT 127.100 65.295 128.970 65.300 ;
        RECT 127.920 65.270 128.970 65.295 ;
        RECT 111.950 56.500 112.950 65.200 ;
        RECT 116.125 63.850 117.175 63.875 ;
        RECT 117.850 63.850 118.900 64.365 ;
        RECT 114.025 62.850 115.350 63.850 ;
        RECT 116.125 62.850 118.900 63.850 ;
        RECT 114.025 56.500 115.025 62.850 ;
        RECT 116.125 62.825 117.175 62.850 ;
        RECT 107.775 54.200 108.775 56.475 ;
        RECT 109.175 55.450 110.225 56.500 ;
        RECT 111.925 55.450 112.975 56.500 ;
        RECT 114.025 55.475 115.625 56.500 ;
        RECT 114.575 55.450 115.625 55.475 ;
        RECT 116.150 54.200 117.150 62.825 ;
        RECT 117.850 61.050 118.900 62.100 ;
        RECT 107.775 53.200 117.150 54.200 ;
        RECT 117.875 54.200 118.875 61.050 ;
        RECT 120.050 60.795 121.045 65.200 ;
        RECT 129.810 64.420 132.370 65.525 ;
        RECT 133.095 65.095 134.250 66.250 ;
        RECT 122.045 61.155 123.045 64.340 ;
        RECT 129.810 63.695 130.915 64.420 ;
        RECT 126.515 62.590 130.915 63.695 ;
        RECT 126.515 61.180 127.620 62.590 ;
        RECT 129.930 61.755 131.045 61.785 ;
        RECT 133.120 61.755 134.225 65.095 ;
        RECT 126.495 61.155 127.650 61.180 ;
        RECT 120.050 60.055 121.050 60.795 ;
        RECT 122.045 60.100 127.650 61.155 ;
        RECT 129.930 60.650 134.225 61.755 ;
        RECT 129.930 60.620 132.130 60.650 ;
        RECT 120.055 56.500 121.050 60.055 ;
        RECT 122.070 60.050 127.650 60.100 ;
        RECT 126.495 60.025 127.650 60.050 ;
        RECT 120.025 55.450 121.075 56.500 ;
        RECT 125.105 56.480 126.095 56.505 ;
        RECT 125.100 55.480 126.100 56.480 ;
        RECT 125.105 55.455 126.095 55.480 ;
        RECT 117.875 53.200 120.350 54.200 ;
        RECT 109.350 52.275 110.400 52.300 ;
        RECT 107.770 51.275 110.400 52.275 ;
        RECT 109.350 51.250 110.400 51.275 ;
        RECT 109.375 47.000 110.375 51.250 ;
        RECT 111.250 47.375 112.250 53.200 ;
        RECT 117.425 51.250 118.475 52.300 ;
        RECT 115.250 49.350 116.300 50.430 ;
        RECT 117.450 48.375 118.450 51.250 ;
        RECT 117.420 47.375 118.480 48.375 ;
        RECT 119.350 47.375 120.350 53.200 ;
        RECT 121.325 53.000 125.850 54.000 ;
        RECT 121.050 48.375 122.040 48.400 ;
        RECT 121.045 47.375 122.045 48.375 ;
        RECT 121.050 47.350 122.040 47.375 ;
        RECT 109.375 46.995 112.475 47.000 ;
        RECT 109.375 46.005 112.500 46.995 ;
        RECT 109.375 46.000 112.475 46.005 ;
        RECT 115.250 45.600 116.300 45.625 ;
        RECT 109.200 44.600 112.250 45.600 ;
        RECT 115.250 44.600 123.050 45.600 ;
        RECT 104.505 42.525 106.730 43.680 ;
        RECT 104.505 42.515 106.705 42.525 ;
        RECT 101.500 33.900 102.550 33.925 ;
        RECT 101.500 32.900 104.600 33.900 ;
        RECT 101.500 32.875 102.550 32.900 ;
        RECT 92.450 30.625 94.925 31.625 ;
        RECT 95.900 30.925 102.525 31.925 ;
        RECT 84.050 29.725 85.050 29.730 ;
        RECT 83.925 29.700 85.050 29.725 ;
        RECT 82.345 28.700 85.050 29.700 ;
        RECT 83.925 28.675 85.050 28.700 ;
        RECT 84.050 28.670 85.050 28.675 ;
        RECT 85.825 24.800 86.825 30.625 ;
        RECT 92.000 28.675 93.050 29.725 ;
        RECT 89.825 26.775 90.875 27.855 ;
        RECT 92.025 25.800 93.025 28.675 ;
        RECT 91.995 24.800 93.055 25.800 ;
        RECT 93.925 24.800 94.925 30.625 ;
        RECT 95.625 25.800 96.615 25.825 ;
        RECT 95.620 24.800 96.620 25.800 ;
        RECT 95.625 24.775 96.615 24.800 ;
        RECT 89.825 23.025 90.875 23.050 ;
        RECT 83.775 22.025 86.825 23.025 ;
        RECT 89.825 22.025 97.625 23.025 ;
        RECT 99.430 22.800 100.430 29.800 ;
        RECT 61.100 11.350 62.100 20.050 ;
        RECT 63.175 17.700 64.500 18.700 ;
        RECT 63.175 11.350 64.175 17.700 ;
        RECT 65.275 17.675 66.325 18.725 ;
        RECT 56.925 9.050 57.925 11.325 ;
        RECT 58.325 10.300 59.375 11.350 ;
        RECT 61.075 10.300 62.125 11.350 ;
        RECT 63.175 10.325 64.775 11.350 ;
        RECT 63.725 10.300 64.775 10.325 ;
        RECT 65.300 9.050 66.300 17.675 ;
        RECT 67.000 15.900 68.050 16.950 ;
        RECT 56.925 8.050 66.300 9.050 ;
        RECT 67.025 9.050 68.025 15.900 ;
        RECT 69.200 15.645 70.195 20.050 ;
        RECT 74.050 19.575 77.100 20.575 ;
        RECT 79.080 19.950 81.305 21.105 ;
        RECT 79.080 19.940 80.195 19.950 ;
        RECT 69.200 14.905 70.200 15.645 ;
        RECT 69.205 11.350 70.200 14.905 ;
        RECT 69.175 10.300 70.225 11.350 ;
        RECT 70.455 9.325 71.505 9.350 ;
        RECT 74.050 9.325 75.050 19.575 ;
        RECT 83.775 11.350 84.775 22.025 ;
        RECT 89.825 22.000 90.875 22.025 ;
        RECT 99.405 21.750 100.455 22.800 ;
        RECT 86.525 21.045 90.850 21.050 ;
        RECT 86.525 20.050 95.620 21.045 ;
        RECT 101.525 20.575 102.525 30.925 ;
        RECT 86.525 11.350 87.525 20.050 ;
        RECT 88.600 17.700 89.925 18.700 ;
        RECT 88.600 11.350 89.600 17.700 ;
        RECT 90.700 17.675 91.750 18.725 ;
        RECT 67.025 8.050 69.500 9.050 ;
        RECT 70.455 8.325 75.050 9.325 ;
        RECT 82.350 9.050 83.350 11.325 ;
        RECT 83.750 10.300 84.800 11.350 ;
        RECT 86.500 10.300 87.550 11.350 ;
        RECT 88.600 10.325 90.200 11.350 ;
        RECT 89.150 10.300 90.200 10.325 ;
        RECT 90.725 9.050 91.725 17.675 ;
        RECT 92.425 15.900 93.475 16.950 ;
        RECT 70.455 8.300 71.505 8.325 ;
        RECT 56.930 7.125 57.920 7.150 ;
        RECT 58.500 7.125 59.550 7.150 ;
        RECT 56.920 6.125 59.550 7.125 ;
        RECT 56.930 6.100 57.920 6.125 ;
        RECT 58.500 6.100 59.550 6.125 ;
        RECT 60.400 2.225 61.400 8.050 ;
        RECT 66.575 6.100 67.625 7.150 ;
        RECT 64.400 4.200 65.450 5.280 ;
        RECT 66.600 3.225 67.600 6.100 ;
        RECT 66.570 2.225 67.630 3.225 ;
        RECT 68.500 2.225 69.500 8.050 ;
        RECT 70.200 3.225 71.190 3.250 ;
        RECT 70.195 2.225 71.195 3.225 ;
        RECT 70.200 2.200 71.190 2.225 ;
        RECT 74.020 1.000 75.020 8.325 ;
        RECT 82.350 8.050 91.725 9.050 ;
        RECT 92.450 9.050 93.450 15.900 ;
        RECT 94.625 15.645 95.620 20.050 ;
        RECT 99.475 19.575 102.525 20.575 ;
        RECT 94.625 14.905 95.625 15.645 ;
        RECT 94.630 11.350 95.625 14.905 ;
        RECT 94.600 10.300 95.650 11.350 ;
        RECT 95.880 9.325 96.930 9.350 ;
        RECT 99.475 9.325 100.475 19.575 ;
        RECT 92.450 8.050 94.925 9.050 ;
        RECT 95.880 8.325 100.475 9.325 ;
        RECT 95.880 8.300 96.930 8.325 ;
        RECT 82.355 7.125 83.345 7.150 ;
        RECT 83.925 7.125 84.975 7.150 ;
        RECT 82.345 6.125 84.975 7.125 ;
        RECT 82.355 6.100 83.345 6.125 ;
        RECT 83.925 6.100 84.975 6.125 ;
        RECT 85.825 2.225 86.825 8.050 ;
        RECT 92.000 6.100 93.050 7.150 ;
        RECT 89.825 4.200 90.875 5.280 ;
        RECT 92.025 3.225 93.025 6.100 ;
        RECT 91.995 2.225 93.055 3.225 ;
        RECT 93.925 2.225 94.925 8.050 ;
        RECT 95.625 3.225 96.615 3.250 ;
        RECT 95.620 2.225 96.620 3.225 ;
        RECT 95.625 2.200 96.615 2.225 ;
        RECT 99.475 1.000 100.475 8.325 ;
        RECT 52.750 0.000 100.475 1.000 ;
        RECT 103.600 1.000 104.600 32.900 ;
        RECT 105.600 21.105 106.705 42.515 ;
        RECT 109.200 33.925 110.200 44.600 ;
        RECT 115.250 44.575 116.300 44.600 ;
        RECT 111.950 43.620 116.275 43.625 ;
        RECT 111.950 42.625 121.045 43.620 ;
        RECT 111.950 33.925 112.950 42.625 ;
        RECT 114.025 40.275 115.350 41.275 ;
        RECT 114.025 33.925 115.025 40.275 ;
        RECT 116.125 40.250 117.175 41.300 ;
        RECT 107.775 31.625 108.775 33.900 ;
        RECT 109.175 32.875 110.225 33.925 ;
        RECT 111.925 32.875 112.975 33.925 ;
        RECT 114.025 32.900 115.625 33.925 ;
        RECT 114.575 32.875 115.625 32.900 ;
        RECT 116.150 31.625 117.150 40.250 ;
        RECT 117.850 38.475 118.900 39.525 ;
        RECT 107.775 30.625 117.150 31.625 ;
        RECT 117.875 31.625 118.875 38.475 ;
        RECT 120.050 38.220 121.045 42.625 ;
        RECT 120.050 37.480 121.050 38.220 ;
        RECT 120.055 33.925 121.050 37.480 ;
        RECT 120.025 32.875 121.075 33.925 ;
        RECT 123.105 33.905 124.095 33.930 ;
        RECT 123.100 32.905 124.100 33.905 ;
        RECT 123.105 32.880 124.095 32.905 ;
        RECT 124.850 31.925 125.850 53.000 ;
        RECT 131.025 43.680 132.130 60.620 ;
        RECT 134.625 56.500 135.625 67.175 ;
        RECT 140.675 67.150 141.725 67.175 ;
        RECT 137.375 66.195 141.700 66.200 ;
        RECT 137.375 65.200 146.470 66.195 ;
        RECT 137.375 56.500 138.375 65.200 ;
        RECT 139.450 62.850 140.775 63.850 ;
        RECT 139.450 56.500 140.450 62.850 ;
        RECT 141.550 62.825 142.600 63.875 ;
        RECT 133.200 54.200 134.200 56.475 ;
        RECT 134.600 55.450 135.650 56.500 ;
        RECT 137.350 55.450 138.400 56.500 ;
        RECT 139.450 55.475 141.050 56.500 ;
        RECT 140.000 55.450 141.050 55.475 ;
        RECT 141.575 54.200 142.575 62.825 ;
        RECT 143.275 61.050 144.325 62.100 ;
        RECT 133.200 53.200 142.575 54.200 ;
        RECT 143.300 54.200 144.300 61.050 ;
        RECT 145.475 60.795 146.470 65.200 ;
        RECT 145.475 60.055 146.475 60.795 ;
        RECT 145.480 56.500 146.475 60.055 ;
        RECT 145.450 55.450 146.500 56.500 ;
        RECT 143.300 53.200 145.775 54.200 ;
        RECT 134.775 52.275 135.825 52.300 ;
        RECT 133.195 51.275 135.825 52.275 ;
        RECT 134.775 51.250 135.825 51.275 ;
        RECT 134.800 47.000 135.800 51.250 ;
        RECT 136.675 47.375 137.675 53.200 ;
        RECT 142.850 51.250 143.900 52.300 ;
        RECT 140.675 49.350 141.725 50.430 ;
        RECT 142.875 48.375 143.875 51.250 ;
        RECT 142.845 47.375 143.905 48.375 ;
        RECT 144.775 47.375 145.775 53.200 ;
        RECT 146.750 53.000 151.275 54.000 ;
        RECT 146.475 48.375 147.465 48.400 ;
        RECT 146.470 47.375 147.470 48.375 ;
        RECT 146.475 47.350 147.465 47.375 ;
        RECT 134.800 46.995 137.900 47.000 ;
        RECT 134.800 46.005 137.925 46.995 ;
        RECT 134.800 46.000 137.900 46.005 ;
        RECT 140.675 45.600 141.725 45.625 ;
        RECT 134.625 44.600 137.675 45.600 ;
        RECT 140.675 44.600 148.475 45.600 ;
        RECT 129.930 42.525 132.155 43.680 ;
        RECT 129.930 42.515 132.130 42.525 ;
        RECT 117.875 30.625 120.350 31.625 ;
        RECT 121.325 30.925 127.950 31.925 ;
        RECT 109.475 29.725 110.475 29.730 ;
        RECT 109.350 29.700 110.475 29.725 ;
        RECT 107.770 28.700 110.475 29.700 ;
        RECT 109.350 28.675 110.475 28.700 ;
        RECT 109.475 28.670 110.475 28.675 ;
        RECT 111.250 24.800 112.250 30.625 ;
        RECT 117.425 28.675 118.475 29.725 ;
        RECT 115.250 26.775 116.300 27.855 ;
        RECT 117.450 25.800 118.450 28.675 ;
        RECT 117.420 24.800 118.480 25.800 ;
        RECT 119.350 24.800 120.350 30.625 ;
        RECT 121.050 25.800 122.040 25.825 ;
        RECT 121.045 24.800 122.045 25.800 ;
        RECT 121.050 24.775 122.040 24.800 ;
        RECT 115.250 23.025 116.300 23.050 ;
        RECT 109.200 22.025 112.250 23.025 ;
        RECT 115.250 22.025 123.050 23.025 ;
        RECT 124.855 22.800 125.855 29.800 ;
        RECT 105.575 21.080 106.730 21.105 ;
        RECT 105.570 19.975 106.730 21.080 ;
        RECT 105.575 19.950 106.730 19.975 ;
        RECT 109.200 11.350 110.200 22.025 ;
        RECT 115.250 22.000 116.300 22.025 ;
        RECT 124.830 21.750 125.880 22.800 ;
        RECT 111.950 21.045 116.275 21.050 ;
        RECT 111.950 20.050 121.045 21.045 ;
        RECT 126.950 20.575 127.950 30.925 ;
        RECT 131.025 21.105 132.130 42.515 ;
        RECT 134.625 33.925 135.625 44.600 ;
        RECT 140.675 44.575 141.725 44.600 ;
        RECT 137.375 43.620 141.700 43.625 ;
        RECT 137.375 42.625 146.470 43.620 ;
        RECT 137.375 33.925 138.375 42.625 ;
        RECT 139.450 40.275 140.775 41.275 ;
        RECT 139.450 33.925 140.450 40.275 ;
        RECT 141.550 40.250 142.600 41.300 ;
        RECT 133.200 31.625 134.200 33.900 ;
        RECT 134.600 32.875 135.650 33.925 ;
        RECT 137.350 32.875 138.400 33.925 ;
        RECT 139.450 32.900 141.050 33.925 ;
        RECT 140.000 32.875 141.050 32.900 ;
        RECT 141.575 31.625 142.575 40.250 ;
        RECT 143.275 38.475 144.325 39.525 ;
        RECT 133.200 30.625 142.575 31.625 ;
        RECT 143.300 31.625 144.300 38.475 ;
        RECT 145.475 38.220 146.470 42.625 ;
        RECT 145.475 37.480 146.475 38.220 ;
        RECT 145.480 33.925 146.475 37.480 ;
        RECT 145.450 32.875 146.500 33.925 ;
        RECT 150.275 31.925 151.275 53.000 ;
        RECT 152.500 32.875 153.550 33.955 ;
        RECT 143.300 30.625 145.775 31.625 ;
        RECT 146.750 30.925 153.375 31.925 ;
        RECT 134.900 29.725 135.900 29.730 ;
        RECT 134.775 29.700 135.900 29.725 ;
        RECT 133.195 28.700 135.900 29.700 ;
        RECT 134.775 28.675 135.900 28.700 ;
        RECT 134.900 28.670 135.900 28.675 ;
        RECT 136.675 24.800 137.675 30.625 ;
        RECT 142.850 28.675 143.900 29.725 ;
        RECT 140.675 26.775 141.725 27.855 ;
        RECT 142.875 25.800 143.875 28.675 ;
        RECT 142.845 24.800 143.905 25.800 ;
        RECT 144.775 24.800 145.775 30.625 ;
        RECT 146.475 25.800 147.465 25.825 ;
        RECT 146.470 24.800 147.470 25.800 ;
        RECT 146.475 24.775 147.465 24.800 ;
        RECT 140.675 23.025 141.725 23.050 ;
        RECT 134.625 22.025 137.675 23.025 ;
        RECT 140.675 22.025 148.475 23.025 ;
        RECT 150.280 22.800 151.280 29.800 ;
        RECT 111.950 11.350 112.950 20.050 ;
        RECT 114.025 17.700 115.350 18.700 ;
        RECT 114.025 11.350 115.025 17.700 ;
        RECT 116.125 17.675 117.175 18.725 ;
        RECT 107.775 9.050 108.775 11.325 ;
        RECT 109.175 10.300 110.225 11.350 ;
        RECT 111.925 10.300 112.975 11.350 ;
        RECT 114.025 10.325 115.625 11.350 ;
        RECT 114.575 10.300 115.625 10.325 ;
        RECT 116.150 9.050 117.150 17.675 ;
        RECT 117.850 15.900 118.900 16.950 ;
        RECT 107.775 8.050 117.150 9.050 ;
        RECT 117.875 9.050 118.875 15.900 ;
        RECT 120.050 15.645 121.045 20.050 ;
        RECT 124.900 19.575 127.950 20.575 ;
        RECT 129.930 19.950 132.155 21.105 ;
        RECT 129.930 19.940 131.045 19.950 ;
        RECT 120.050 14.905 121.050 15.645 ;
        RECT 120.055 11.350 121.050 14.905 ;
        RECT 120.025 10.300 121.075 11.350 ;
        RECT 121.305 9.325 122.355 9.350 ;
        RECT 124.900 9.325 125.900 19.575 ;
        RECT 134.625 11.350 135.625 22.025 ;
        RECT 140.675 22.000 141.725 22.025 ;
        RECT 150.255 21.750 151.305 22.800 ;
        RECT 137.375 21.045 141.700 21.050 ;
        RECT 137.375 20.050 146.470 21.045 ;
        RECT 152.375 20.575 153.375 30.925 ;
        RECT 137.375 11.350 138.375 20.050 ;
        RECT 139.450 17.700 140.775 18.700 ;
        RECT 139.450 11.350 140.450 17.700 ;
        RECT 141.550 17.675 142.600 18.725 ;
        RECT 117.875 8.050 120.350 9.050 ;
        RECT 121.305 8.325 125.900 9.325 ;
        RECT 133.200 9.050 134.200 11.325 ;
        RECT 134.600 10.300 135.650 11.350 ;
        RECT 137.350 10.300 138.400 11.350 ;
        RECT 139.450 10.325 141.050 11.350 ;
        RECT 140.000 10.300 141.050 10.325 ;
        RECT 141.575 9.050 142.575 17.675 ;
        RECT 143.275 15.900 144.325 16.950 ;
        RECT 121.305 8.300 122.355 8.325 ;
        RECT 107.780 7.125 108.770 7.150 ;
        RECT 109.350 7.125 110.400 7.150 ;
        RECT 107.770 6.125 110.400 7.125 ;
        RECT 107.780 6.100 108.770 6.125 ;
        RECT 109.350 6.100 110.400 6.125 ;
        RECT 111.250 2.225 112.250 8.050 ;
        RECT 117.425 6.100 118.475 7.150 ;
        RECT 115.250 4.200 116.300 5.280 ;
        RECT 117.450 3.225 118.450 6.100 ;
        RECT 117.420 2.225 118.480 3.225 ;
        RECT 119.350 2.225 120.350 8.050 ;
        RECT 121.050 3.225 122.040 3.250 ;
        RECT 121.045 2.225 122.045 3.225 ;
        RECT 121.050 2.200 122.040 2.225 ;
        RECT 124.870 1.000 125.870 8.325 ;
        RECT 133.200 8.050 142.575 9.050 ;
        RECT 143.300 9.050 144.300 15.900 ;
        RECT 145.475 15.645 146.470 20.050 ;
        RECT 150.325 19.575 153.375 20.575 ;
        RECT 145.475 14.905 146.475 15.645 ;
        RECT 145.480 11.350 146.475 14.905 ;
        RECT 145.450 10.300 146.500 11.350 ;
        RECT 146.730 9.325 147.780 9.350 ;
        RECT 150.325 9.325 151.325 19.575 ;
        RECT 143.300 8.050 145.775 9.050 ;
        RECT 146.730 8.325 151.325 9.325 ;
        RECT 146.730 8.300 147.780 8.325 ;
        RECT 133.205 7.125 134.195 7.150 ;
        RECT 134.775 7.125 135.825 7.150 ;
        RECT 133.195 6.125 135.825 7.125 ;
        RECT 133.205 6.100 134.195 6.125 ;
        RECT 134.775 6.100 135.825 6.125 ;
        RECT 136.675 2.225 137.675 8.050 ;
        RECT 142.850 6.100 143.900 7.150 ;
        RECT 140.675 4.200 141.725 5.280 ;
        RECT 142.875 3.225 143.875 6.100 ;
        RECT 142.845 2.225 143.905 3.225 ;
        RECT 144.775 2.225 145.775 8.050 ;
        RECT 146.475 3.225 147.465 3.250 ;
        RECT 146.470 2.225 147.470 3.225 ;
        RECT 146.475 2.200 147.465 2.225 ;
        RECT 150.325 1.000 151.325 8.325 ;
        RECT 103.600 0.000 151.325 1.000 ;
        RECT 156.415 0.950 157.305 0.975 ;
        RECT 156.410 0.050 157.310 0.950 ;
        RECT 156.415 0.025 157.305 0.050 ;
      LAYER met4 ;
        RECT 91.970 224.760 92.310 225.305 ;
        RECT 92.610 224.760 92.980 225.305 ;
        RECT 91.970 224.295 92.980 224.760 ;
        RECT 95.645 224.760 95.990 225.305 ;
        RECT 96.290 224.760 96.655 225.305 ;
        RECT 95.645 224.295 96.655 224.760 ;
        RECT 99.295 224.760 99.670 225.305 ;
        RECT 99.970 224.760 100.305 225.305 ;
        RECT 99.295 224.295 100.305 224.760 ;
        RECT 102.995 224.760 103.350 225.305 ;
        RECT 103.650 224.760 104.005 225.305 ;
        RECT 102.995 224.295 104.005 224.760 ;
        RECT 106.670 224.760 107.030 225.305 ;
        RECT 107.330 224.760 107.680 225.305 ;
        RECT 106.670 224.295 107.680 224.760 ;
        RECT 110.370 224.760 110.710 225.305 ;
        RECT 111.010 224.760 111.380 225.305 ;
        RECT 110.370 224.295 111.380 224.760 ;
        RECT 114.045 224.760 114.390 225.305 ;
        RECT 114.690 224.760 115.055 225.305 ;
        RECT 114.045 224.295 115.055 224.760 ;
        RECT 117.720 224.760 118.070 225.305 ;
        RECT 118.370 224.760 118.730 225.305 ;
        RECT 117.720 224.295 118.730 224.760 ;
        RECT 121.420 224.760 121.750 225.305 ;
        RECT 122.050 224.760 122.430 225.305 ;
        RECT 121.420 224.295 122.430 224.760 ;
        RECT 125.070 224.760 125.430 225.305 ;
        RECT 125.730 224.760 126.080 225.305 ;
        RECT 125.070 224.295 126.080 224.760 ;
        RECT 128.770 224.760 129.110 225.305 ;
        RECT 129.410 224.760 129.780 225.305 ;
        RECT 128.770 224.295 129.780 224.760 ;
        RECT 132.445 224.760 132.790 225.305 ;
        RECT 133.090 224.760 133.455 225.305 ;
        RECT 132.445 224.295 133.455 224.760 ;
        RECT 136.120 224.760 136.470 225.305 ;
        RECT 136.770 224.760 137.130 225.305 ;
        RECT 136.120 224.295 137.130 224.760 ;
        RECT 139.770 224.760 140.150 225.330 ;
        RECT 140.450 224.760 140.830 225.330 ;
        RECT 139.770 224.270 140.830 224.760 ;
        RECT 143.470 224.760 143.830 225.305 ;
        RECT 144.130 224.760 144.480 225.305 ;
        RECT 143.470 224.295 144.480 224.760 ;
        RECT 147.145 224.760 147.510 225.305 ;
        RECT 147.810 224.760 148.155 225.305 ;
        RECT 147.145 224.295 148.155 224.760 ;
        RECT 150.845 224.760 151.190 225.305 ;
        RECT 151.490 224.760 151.855 225.305 ;
        RECT 150.845 224.295 151.855 224.760 ;
        RECT 154.495 224.760 154.870 225.305 ;
        RECT 155.170 224.760 155.505 225.305 ;
        RECT 154.495 224.295 155.505 224.760 ;
        RECT 13.275 216.550 14.875 221.975 ;
        RECT 99.675 217.300 111.375 218.300 ;
        RECT 4.175 163.970 4.960 165.085 ;
        RECT 5.775 151.125 6.775 216.550 ;
        RECT 7.775 173.705 8.775 216.545 ;
        RECT 7.770 172.695 8.780 173.705 ;
        RECT 5.775 150.125 7.105 151.125 ;
        RECT 4.175 91.970 4.960 93.085 ;
        RECT 5.775 79.125 6.775 150.125 ;
        RECT 7.775 101.705 8.775 172.695 ;
        RECT 7.770 100.695 8.780 101.705 ;
        RECT 5.775 78.125 7.105 79.125 ;
        RECT 4.175 19.970 4.960 21.085 ;
        RECT 5.775 7.125 6.775 78.125 ;
        RECT 7.775 29.705 8.775 100.695 ;
        RECT 7.770 28.695 8.780 29.705 ;
        RECT 5.775 6.125 7.105 7.125 ;
        RECT 5.775 1.535 6.775 6.125 ;
        RECT 7.775 1.535 8.775 28.695 ;
        RECT 9.775 1.535 10.775 216.550 ;
        RECT 15.745 192.375 16.755 192.380 ;
        RECT 15.745 191.375 20.345 192.375 ;
        RECT 15.745 191.370 16.755 191.375 ;
        RECT 15.745 169.800 16.755 169.805 ;
        RECT 15.745 168.800 20.345 169.800 ;
        RECT 15.745 168.795 16.755 168.800 ;
        RECT 21.400 147.850 22.400 216.550 ;
        RECT 15.745 147.225 16.755 147.230 ;
        RECT 15.745 146.225 20.345 147.225 ;
        RECT 15.745 146.220 16.755 146.225 ;
        RECT 15.745 120.375 16.755 120.380 ;
        RECT 15.745 119.375 20.345 120.375 ;
        RECT 15.745 119.370 16.755 119.375 ;
        RECT 15.745 97.800 16.755 97.805 ;
        RECT 15.745 96.800 20.345 97.800 ;
        RECT 15.745 96.795 16.755 96.800 ;
        RECT 21.400 75.850 22.400 145.000 ;
        RECT 15.745 75.225 16.755 75.230 ;
        RECT 15.745 74.225 20.345 75.225 ;
        RECT 15.745 74.220 16.755 74.225 ;
        RECT 15.745 48.375 16.755 48.380 ;
        RECT 15.745 47.375 20.345 48.375 ;
        RECT 15.745 47.370 16.755 47.375 ;
        RECT 15.745 25.800 16.755 25.805 ;
        RECT 15.745 24.800 20.345 25.800 ;
        RECT 15.745 24.795 16.755 24.800 ;
        RECT 15.745 3.225 16.755 3.230 ;
        RECT 15.745 2.225 20.345 3.225 ;
        RECT 15.745 2.220 16.755 2.225 ;
        RECT 21.400 1.540 22.400 73.000 ;
        RECT 23.400 1.540 24.400 214.550 ;
        RECT 25.400 1.540 26.400 216.550 ;
        RECT 31.200 151.125 32.200 216.550 ;
        RECT 33.200 173.705 34.200 216.550 ;
        RECT 33.195 172.695 34.205 173.705 ;
        RECT 31.200 150.125 32.530 151.125 ;
        RECT 31.200 79.125 32.200 150.125 ;
        RECT 33.200 101.705 34.200 172.695 ;
        RECT 33.195 100.695 34.205 101.705 ;
        RECT 31.200 78.125 32.530 79.125 ;
        RECT 31.200 7.125 32.200 78.125 ;
        RECT 33.200 29.705 34.200 100.695 ;
        RECT 33.195 28.695 34.205 29.705 ;
        RECT 31.200 6.125 32.530 7.125 ;
        RECT 31.200 1.535 32.200 6.125 ;
        RECT 33.200 1.535 34.200 28.695 ;
        RECT 35.200 1.535 36.200 216.550 ;
        RECT 41.170 192.375 42.180 192.380 ;
        RECT 41.170 191.375 45.770 192.375 ;
        RECT 41.170 191.370 42.180 191.375 ;
        RECT 41.170 169.800 42.180 169.805 ;
        RECT 41.170 168.800 45.770 169.800 ;
        RECT 41.170 168.795 42.180 168.800 ;
        RECT 41.170 147.225 42.180 147.230 ;
        RECT 41.170 146.225 45.770 147.225 ;
        RECT 41.170 146.220 42.180 146.225 ;
        RECT 41.170 120.375 42.180 120.380 ;
        RECT 41.170 119.375 45.770 120.375 ;
        RECT 41.170 119.370 42.180 119.375 ;
        RECT 41.170 97.800 42.180 97.805 ;
        RECT 41.170 96.800 45.770 97.800 ;
        RECT 41.170 96.795 42.180 96.800 ;
        RECT 41.170 75.225 42.180 75.230 ;
        RECT 41.170 74.225 45.770 75.225 ;
        RECT 41.170 74.220 42.180 74.225 ;
        RECT 41.170 48.375 42.180 48.380 ;
        RECT 41.170 47.375 45.770 48.375 ;
        RECT 41.170 47.370 42.180 47.375 ;
        RECT 41.170 25.800 42.180 25.805 ;
        RECT 41.170 24.800 45.770 25.800 ;
        RECT 41.170 24.795 42.180 24.800 ;
        RECT 41.170 3.225 42.180 3.230 ;
        RECT 41.170 2.225 45.770 3.225 ;
        RECT 41.170 2.220 42.180 2.225 ;
        RECT 46.825 1.540 47.825 214.550 ;
        RECT 48.825 1.540 49.825 216.550 ;
        RECT 55.025 163.970 55.810 165.085 ;
        RECT 56.625 151.125 57.625 216.550 ;
        RECT 58.625 173.705 59.625 216.545 ;
        RECT 58.620 172.695 59.630 173.705 ;
        RECT 56.625 150.125 57.955 151.125 ;
        RECT 55.025 91.970 55.810 93.085 ;
        RECT 56.625 79.125 57.625 150.125 ;
        RECT 58.625 101.705 59.625 172.695 ;
        RECT 58.620 100.695 59.630 101.705 ;
        RECT 56.625 78.125 57.955 79.125 ;
        RECT 55.025 19.970 55.810 21.085 ;
        RECT 56.625 7.125 57.625 78.125 ;
        RECT 58.625 29.705 59.625 100.695 ;
        RECT 58.620 28.695 59.630 29.705 ;
        RECT 56.625 6.125 57.955 7.125 ;
        RECT 56.625 1.535 57.625 6.125 ;
        RECT 58.625 1.535 59.625 28.695 ;
        RECT 60.625 1.535 61.625 216.550 ;
        RECT 66.595 192.375 67.605 192.380 ;
        RECT 66.595 191.375 71.195 192.375 ;
        RECT 66.595 191.370 67.605 191.375 ;
        RECT 66.595 169.800 67.605 169.805 ;
        RECT 66.595 168.800 71.195 169.800 ;
        RECT 66.595 168.795 67.605 168.800 ;
        RECT 72.250 147.850 73.250 216.550 ;
        RECT 66.595 147.225 67.605 147.230 ;
        RECT 66.595 146.225 71.195 147.225 ;
        RECT 66.595 146.220 67.605 146.225 ;
        RECT 66.595 120.375 67.605 120.380 ;
        RECT 66.595 119.375 71.195 120.375 ;
        RECT 66.595 119.370 67.605 119.375 ;
        RECT 66.595 97.800 67.605 97.805 ;
        RECT 66.595 96.800 71.195 97.800 ;
        RECT 66.595 96.795 67.605 96.800 ;
        RECT 72.250 75.850 73.250 145.000 ;
        RECT 66.595 75.225 67.605 75.230 ;
        RECT 66.595 74.225 71.195 75.225 ;
        RECT 66.595 74.220 67.605 74.225 ;
        RECT 66.595 48.375 67.605 48.380 ;
        RECT 66.595 47.375 71.195 48.375 ;
        RECT 66.595 47.370 67.605 47.375 ;
        RECT 66.595 25.800 67.605 25.805 ;
        RECT 66.595 24.800 71.195 25.800 ;
        RECT 66.595 24.795 67.605 24.800 ;
        RECT 66.595 3.225 67.605 3.230 ;
        RECT 66.595 2.225 71.195 3.225 ;
        RECT 66.595 2.220 67.605 2.225 ;
        RECT 72.250 1.540 73.250 73.000 ;
        RECT 74.250 1.540 75.250 214.550 ;
        RECT 76.250 1.540 77.250 216.550 ;
        RECT 82.050 151.125 83.050 216.550 ;
        RECT 84.050 173.705 85.050 216.550 ;
        RECT 84.045 172.695 85.055 173.705 ;
        RECT 82.050 150.125 83.380 151.125 ;
        RECT 82.050 79.125 83.050 150.125 ;
        RECT 84.050 101.705 85.050 172.695 ;
        RECT 84.045 100.695 85.055 101.705 ;
        RECT 82.050 78.125 83.380 79.125 ;
        RECT 82.050 7.125 83.050 78.125 ;
        RECT 84.050 29.705 85.050 100.695 ;
        RECT 84.045 28.695 85.055 29.705 ;
        RECT 82.050 6.125 83.380 7.125 ;
        RECT 82.050 1.535 83.050 6.125 ;
        RECT 84.050 1.535 85.050 28.695 ;
        RECT 86.050 1.535 87.050 216.550 ;
        RECT 92.020 192.375 93.030 192.380 ;
        RECT 92.020 191.375 96.620 192.375 ;
        RECT 92.020 191.370 93.030 191.375 ;
        RECT 92.020 169.800 93.030 169.805 ;
        RECT 92.020 168.800 96.620 169.800 ;
        RECT 92.020 168.795 93.030 168.800 ;
        RECT 92.020 147.225 93.030 147.230 ;
        RECT 92.020 146.225 96.620 147.225 ;
        RECT 92.020 146.220 93.030 146.225 ;
        RECT 92.020 120.375 93.030 120.380 ;
        RECT 92.020 119.375 96.620 120.375 ;
        RECT 92.020 119.370 93.030 119.375 ;
        RECT 92.020 97.800 93.030 97.805 ;
        RECT 92.020 96.800 96.620 97.800 ;
        RECT 92.020 96.795 93.030 96.800 ;
        RECT 92.020 75.225 93.030 75.230 ;
        RECT 92.020 74.225 96.620 75.225 ;
        RECT 92.020 74.220 93.030 74.225 ;
        RECT 92.020 48.375 93.030 48.380 ;
        RECT 92.020 47.375 96.620 48.375 ;
        RECT 92.020 47.370 93.030 47.375 ;
        RECT 92.020 25.800 93.030 25.805 ;
        RECT 92.020 24.800 96.620 25.800 ;
        RECT 92.020 24.795 93.030 24.800 ;
        RECT 92.020 3.225 93.030 3.230 ;
        RECT 92.020 2.225 96.620 3.225 ;
        RECT 92.020 2.220 93.030 2.225 ;
        RECT 97.675 1.540 98.675 214.550 ;
        RECT 99.675 1.540 100.675 217.300 ;
        RECT 105.875 163.970 106.660 165.085 ;
        RECT 107.475 151.125 108.475 216.550 ;
        RECT 109.475 173.705 110.475 216.545 ;
        RECT 109.470 172.695 110.480 173.705 ;
        RECT 107.475 150.125 108.805 151.125 ;
        RECT 105.875 91.970 106.660 93.085 ;
        RECT 107.475 79.125 108.475 150.125 ;
        RECT 109.475 101.705 110.475 172.695 ;
        RECT 109.470 100.695 110.480 101.705 ;
        RECT 107.475 78.125 108.805 79.125 ;
        RECT 105.875 19.970 106.660 21.085 ;
        RECT 107.475 7.125 108.475 78.125 ;
        RECT 109.475 29.705 110.475 100.695 ;
        RECT 109.470 28.695 110.480 29.705 ;
        RECT 107.475 6.125 108.805 7.125 ;
        RECT 107.475 1.535 108.475 6.125 ;
        RECT 109.475 1.535 110.475 28.695 ;
        RECT 111.475 1.535 112.475 216.550 ;
        RECT 117.445 192.375 118.455 192.380 ;
        RECT 117.445 191.375 122.045 192.375 ;
        RECT 117.445 191.370 118.455 191.375 ;
        RECT 117.445 169.800 118.455 169.805 ;
        RECT 117.445 168.800 122.045 169.800 ;
        RECT 117.445 168.795 118.455 168.800 ;
        RECT 123.100 147.850 124.100 216.575 ;
        RECT 117.445 147.225 118.455 147.230 ;
        RECT 117.445 146.225 122.045 147.225 ;
        RECT 117.445 146.220 118.455 146.225 ;
        RECT 117.445 120.375 118.455 120.380 ;
        RECT 117.445 119.375 122.045 120.375 ;
        RECT 117.445 119.370 118.455 119.375 ;
        RECT 117.445 97.800 118.455 97.805 ;
        RECT 117.445 96.800 122.045 97.800 ;
        RECT 117.445 96.795 118.455 96.800 ;
        RECT 123.100 75.850 124.100 145.000 ;
        RECT 117.445 75.225 118.455 75.230 ;
        RECT 117.445 74.225 122.045 75.225 ;
        RECT 117.445 74.220 118.455 74.225 ;
        RECT 117.445 48.375 118.455 48.380 ;
        RECT 117.445 47.375 122.045 48.375 ;
        RECT 117.445 47.370 118.455 47.375 ;
        RECT 117.445 25.800 118.455 25.805 ;
        RECT 117.445 24.800 122.045 25.800 ;
        RECT 117.445 24.795 118.455 24.800 ;
        RECT 117.445 3.225 118.455 3.230 ;
        RECT 117.445 2.225 122.045 3.225 ;
        RECT 117.445 2.220 118.455 2.225 ;
        RECT 123.100 1.540 124.100 73.000 ;
        RECT 125.100 1.540 126.100 214.550 ;
        RECT 127.100 1.540 128.100 216.550 ;
        RECT 132.900 151.125 133.900 216.550 ;
        RECT 134.900 173.705 135.900 216.550 ;
        RECT 134.895 172.695 135.905 173.705 ;
        RECT 132.900 150.125 134.230 151.125 ;
        RECT 132.900 79.125 133.900 150.125 ;
        RECT 134.900 101.705 135.900 172.695 ;
        RECT 134.895 100.695 135.905 101.705 ;
        RECT 132.900 78.125 134.230 79.125 ;
        RECT 132.900 7.125 133.900 78.125 ;
        RECT 134.900 29.705 135.900 100.695 ;
        RECT 134.895 28.695 135.905 29.705 ;
        RECT 132.900 6.125 134.230 7.125 ;
        RECT 132.900 1.535 133.900 6.125 ;
        RECT 134.900 1.535 135.900 28.695 ;
        RECT 136.900 1.535 137.900 216.550 ;
        RECT 142.870 192.375 143.880 192.380 ;
        RECT 142.870 191.375 147.470 192.375 ;
        RECT 142.870 191.370 143.880 191.375 ;
        RECT 142.870 169.800 143.880 169.805 ;
        RECT 142.870 168.800 147.470 169.800 ;
        RECT 142.870 168.795 143.880 168.800 ;
        RECT 142.870 147.225 143.880 147.230 ;
        RECT 142.870 146.225 147.470 147.225 ;
        RECT 142.870 146.220 143.880 146.225 ;
        RECT 142.870 120.375 143.880 120.380 ;
        RECT 142.870 119.375 147.470 120.375 ;
        RECT 142.870 119.370 143.880 119.375 ;
        RECT 142.870 97.800 143.880 97.805 ;
        RECT 142.870 96.800 147.470 97.800 ;
        RECT 142.870 96.795 143.880 96.800 ;
        RECT 142.870 75.225 143.880 75.230 ;
        RECT 142.870 74.225 147.470 75.225 ;
        RECT 142.870 74.220 143.880 74.225 ;
        RECT 142.870 48.375 143.880 48.380 ;
        RECT 142.870 47.375 147.470 48.375 ;
        RECT 142.870 47.370 143.880 47.375 ;
        RECT 142.870 25.800 143.880 25.805 ;
        RECT 142.870 24.800 147.470 25.800 ;
        RECT 142.870 24.795 143.880 24.800 ;
        RECT 142.870 3.225 143.880 3.230 ;
        RECT 142.870 2.225 147.470 3.225 ;
        RECT 142.870 2.220 143.880 2.225 ;
        RECT 148.525 1.540 149.525 214.550 ;
        RECT 150.525 1.540 151.525 216.550 ;
        RECT 152.525 33.930 153.525 216.550 ;
        RECT 154.525 105.930 155.525 216.550 ;
        RECT 156.525 177.930 157.525 216.550 ;
        RECT 156.495 176.920 157.555 177.930 ;
        RECT 154.495 104.920 155.555 105.930 ;
        RECT 152.495 32.920 153.555 33.930 ;
        RECT 152.525 1.540 153.525 32.920 ;
        RECT 154.525 1.535 155.525 104.920 ;
        RECT 156.525 1.535 157.525 176.920 ;
  END
END tt_um_htfab_fprn
END LIBRARY

