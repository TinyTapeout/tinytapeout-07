MACRO tt_um_brucemack_sb_mixer
  CLASS BLOCK ;
  FOREIGN tt_um_brucemack_sb_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 40.000000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.450000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.450000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 22.813499 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 129.470 20.700 135.980 23.050 ;
        RECT 138.050 22.480 145.150 25.000 ;
        RECT 137.790 21.380 145.150 22.480 ;
        RECT 137.800 21.360 145.150 21.380 ;
        RECT 138.050 18.750 145.150 21.360 ;
      LAYER nwell ;
        RECT 136.890 13.830 138.495 16.430 ;
      LAYER pwell ;
        RECT 138.785 15.175 139.695 16.000 ;
        RECT 138.785 15.070 139.885 15.175 ;
        RECT 139.715 15.005 139.885 15.070 ;
      LAYER nwell ;
        RECT 141.190 14.530 142.795 17.130 ;
      LAYER pwell ;
        RECT 143.085 15.875 143.995 16.700 ;
        RECT 143.085 15.770 144.185 15.875 ;
        RECT 144.015 15.705 144.185 15.770 ;
        RECT 143.125 14.735 143.910 15.165 ;
        RECT 138.825 14.035 139.610 14.465 ;
        RECT 129.470 8.570 135.980 10.920 ;
        RECT 138.050 6.620 145.150 12.870 ;
        RECT 146.500 10.610 153.600 21.440 ;
      LAYER li1 ;
        RECT 138.230 24.650 144.970 24.820 ;
        RECT 129.650 22.700 135.800 22.870 ;
        RECT 129.650 21.050 129.820 22.700 ;
        RECT 135.630 22.310 135.800 22.700 ;
        RECT 138.230 22.590 138.400 24.650 ;
        RECT 139.080 24.080 144.120 24.250 ;
        RECT 130.300 21.530 132.460 22.220 ;
        RECT 132.990 21.530 135.150 22.220 ;
        RECT 135.530 21.400 135.880 22.310 ;
        RECT 135.630 21.050 135.800 21.400 ;
        RECT 138.200 21.380 138.470 22.590 ;
        RECT 138.740 22.020 138.910 24.020 ;
        RECT 144.290 22.020 144.460 24.020 ;
        RECT 144.800 22.950 144.970 24.650 ;
        RECT 139.080 21.790 144.120 21.960 ;
        RECT 129.650 20.880 135.800 21.050 ;
        RECT 138.230 19.100 138.400 21.380 ;
        RECT 138.740 19.730 138.910 21.730 ;
        RECT 144.290 19.730 144.460 21.730 ;
        RECT 144.730 21.600 145.060 22.950 ;
        RECT 139.080 19.500 144.120 19.670 ;
        RECT 144.800 19.100 144.970 21.600 ;
        RECT 148.210 21.260 151.970 21.350 ;
        RECT 138.230 18.930 144.970 19.100 ;
        RECT 146.680 21.090 153.420 21.260 ;
        RECT 136.995 15.410 137.165 16.240 ;
        RECT 137.335 15.680 139.545 15.910 ;
        RECT 137.335 15.580 138.315 15.680 ;
        RECT 138.915 15.580 139.545 15.680 ;
        RECT 136.995 15.200 138.305 15.410 ;
        RECT 136.995 14.860 137.165 15.200 ;
        RECT 138.485 15.180 138.725 15.510 ;
        RECT 139.715 15.410 139.885 16.240 ;
        RECT 141.295 16.110 141.465 16.940 ;
        RECT 141.635 16.380 143.845 16.610 ;
        RECT 141.635 16.280 142.615 16.380 ;
        RECT 143.215 16.280 143.845 16.380 ;
        RECT 141.295 15.900 142.605 16.110 ;
        RECT 141.295 15.560 141.465 15.900 ;
        RECT 142.785 15.880 143.025 16.210 ;
        RECT 144.015 16.110 144.185 16.940 ;
        RECT 143.195 15.880 144.185 16.110 ;
        RECT 144.015 15.560 144.185 15.880 ;
        RECT 138.895 15.180 139.885 15.410 ;
        RECT 139.715 14.860 139.885 15.180 ;
        RECT 141.295 15.095 141.465 15.180 ;
        RECT 144.015 15.095 144.185 15.180 ;
        RECT 141.295 14.805 142.630 15.095 ;
        RECT 143.290 14.805 144.185 15.095 ;
        RECT 141.295 14.720 141.465 14.805 ;
        RECT 144.015 14.720 144.185 14.805 ;
        RECT 136.995 14.395 137.165 14.480 ;
        RECT 139.715 14.395 139.885 14.480 ;
        RECT 136.995 14.105 138.330 14.395 ;
        RECT 138.990 14.105 139.885 14.395 ;
        RECT 136.995 14.020 137.165 14.105 ;
        RECT 139.715 14.020 139.885 14.105 ;
        RECT 138.230 12.520 144.970 12.690 ;
        RECT 129.650 10.570 135.800 10.740 ;
        RECT 129.650 8.920 129.820 10.570 ;
        RECT 130.300 9.400 132.460 10.090 ;
        RECT 132.990 9.400 135.150 10.090 ;
        RECT 135.630 8.920 135.800 10.570 ;
        RECT 129.650 8.750 135.800 8.920 ;
        RECT 138.230 10.260 138.400 12.520 ;
        RECT 139.080 11.950 144.120 12.120 ;
        RECT 138.230 9.230 138.410 10.260 ;
        RECT 138.740 9.890 138.910 11.890 ;
        RECT 144.290 9.890 144.460 11.890 ;
        RECT 144.800 10.640 144.970 12.520 ;
        RECT 146.680 10.960 146.850 21.090 ;
        RECT 148.210 21.010 151.970 21.090 ;
        RECT 147.530 20.520 152.570 20.690 ;
        RECT 147.190 18.460 147.360 20.460 ;
        RECT 152.740 18.460 152.910 20.460 ;
        RECT 147.530 18.230 152.570 18.400 ;
        RECT 147.190 16.170 147.360 18.170 ;
        RECT 152.740 16.170 152.910 18.170 ;
        RECT 147.530 15.940 152.570 16.110 ;
        RECT 147.190 13.880 147.360 15.880 ;
        RECT 152.740 13.880 152.910 15.880 ;
        RECT 147.530 13.650 152.570 13.820 ;
        RECT 147.190 11.590 147.360 13.590 ;
        RECT 152.740 11.590 152.910 13.590 ;
        RECT 147.530 11.360 152.570 11.530 ;
        RECT 153.250 10.960 153.420 21.090 ;
        RECT 146.680 10.790 153.420 10.960 ;
        RECT 139.080 9.660 144.120 9.830 ;
        RECT 138.230 6.970 138.400 9.230 ;
        RECT 138.740 7.600 138.910 9.600 ;
        RECT 144.290 7.600 144.460 9.600 ;
        RECT 144.700 8.910 145.120 10.640 ;
        RECT 139.080 7.370 144.120 7.540 ;
        RECT 144.800 6.970 144.970 8.910 ;
        RECT 138.230 6.800 144.970 6.970 ;
      LAYER met1 ;
        RECT 132.400 26.630 133.300 26.660 ;
        RECT 136.160 26.630 137.160 26.840 ;
        RECT 132.400 25.730 137.190 26.630 ;
        RECT 132.400 25.700 133.300 25.730 ;
        RECT 136.160 23.500 137.160 25.730 ;
        RECT 154.760 24.990 156.320 26.490 ;
        RECT 139.130 24.280 144.070 24.400 ;
        RECT 139.100 24.050 144.100 24.280 ;
        RECT 128.330 22.240 132.410 22.380 ;
        RECT 128.270 22.170 132.410 22.240 ;
        RECT 133.030 22.170 135.190 22.340 ;
        RECT 128.270 21.600 132.435 22.170 ;
        RECT 128.270 17.750 129.270 21.600 ;
        RECT 130.330 21.580 132.435 21.600 ;
        RECT 133.015 21.580 135.190 22.170 ;
        RECT 133.030 21.390 135.190 21.580 ;
        RECT 135.450 21.290 138.570 22.660 ;
        RECT 138.710 22.040 138.940 24.000 ;
        RECT 139.130 23.940 144.070 24.050 ;
        RECT 138.720 21.710 138.940 22.040 ;
        RECT 139.150 21.990 144.040 22.150 ;
        RECT 144.260 22.040 144.490 24.000 ;
        RECT 154.790 23.230 156.290 24.990 ;
        RECT 139.100 21.760 144.100 21.990 ;
        RECT 138.710 19.750 138.940 21.710 ;
        RECT 139.150 21.610 144.040 21.760 ;
        RECT 144.270 21.710 144.490 22.040 ;
        RECT 138.720 18.320 138.940 19.750 ;
        RECT 139.150 19.700 144.060 19.780 ;
        RECT 144.260 19.750 144.490 21.710 ;
        RECT 144.700 22.940 152.230 23.010 ;
        RECT 155.120 22.940 156.120 23.230 ;
        RECT 144.700 21.740 156.120 22.940 ;
        RECT 144.700 21.530 152.230 21.740 ;
        RECT 139.100 19.470 144.100 19.700 ;
        RECT 139.150 19.330 144.060 19.470 ;
        RECT 144.270 18.320 144.490 19.750 ;
        RECT 138.720 18.020 144.490 18.320 ;
        RECT 128.270 17.470 137.190 17.750 ;
        RECT 143.210 17.700 144.490 18.020 ;
        RECT 143.210 17.690 144.470 17.700 ;
        RECT 143.210 17.670 143.530 17.690 ;
        RECT 128.270 17.110 141.600 17.470 ;
        RECT 128.270 16.750 137.190 17.110 ;
        RECT 141.220 17.100 141.600 17.110 ;
        RECT 141.270 16.940 141.510 17.100 ;
        RECT 128.270 10.130 129.270 16.750 ;
        RECT 136.990 16.380 137.170 16.750 ;
        RECT 138.020 16.690 138.280 16.700 ;
        RECT 138.020 16.465 140.745 16.690 ;
        RECT 136.980 16.240 137.180 16.380 ;
        RECT 136.840 14.860 137.320 16.240 ;
        RECT 138.020 15.590 138.280 16.465 ;
        RECT 136.990 14.480 137.170 14.860 ;
        RECT 132.700 13.810 133.000 13.840 ;
        RECT 135.550 13.810 136.550 14.040 ;
        RECT 136.840 14.020 137.320 14.480 ;
        RECT 132.700 13.680 136.550 13.810 ;
        RECT 138.470 13.680 138.760 15.540 ;
        RECT 132.700 13.510 138.760 13.680 ;
        RECT 132.700 13.480 133.000 13.510 ;
        RECT 135.550 13.390 138.760 13.510 ;
        RECT 135.550 13.040 136.550 13.390 ;
        RECT 139.055 12.920 139.280 16.465 ;
        RECT 139.560 14.860 140.040 16.240 ;
        RECT 139.640 14.480 139.960 14.860 ;
        RECT 139.560 14.020 140.040 14.480 ;
        RECT 140.415 14.285 140.745 16.465 ;
        RECT 141.140 15.560 141.620 16.940 ;
        RECT 143.240 16.270 143.480 17.670 ;
        RECT 145.305 16.940 146.390 21.530 ;
        RECT 147.750 20.950 152.230 21.530 ;
        RECT 147.570 20.720 152.480 20.810 ;
        RECT 147.550 20.490 152.550 20.720 ;
        RECT 147.160 18.480 147.390 20.440 ;
        RECT 147.570 20.430 152.480 20.490 ;
        RECT 147.180 18.150 147.390 18.480 ;
        RECT 147.630 18.430 152.490 18.550 ;
        RECT 152.710 18.480 152.940 20.440 ;
        RECT 147.550 18.200 152.550 18.430 ;
        RECT 141.270 15.180 141.510 15.560 ;
        RECT 141.140 14.720 141.620 15.180 ;
        RECT 142.770 14.285 143.070 16.250 ;
        RECT 143.860 15.560 146.390 16.940 ;
        RECT 147.160 16.190 147.390 18.150 ;
        RECT 147.630 18.050 152.490 18.200 ;
        RECT 152.790 18.150 152.930 18.480 ;
        RECT 147.180 15.860 147.390 16.190 ;
        RECT 147.560 16.140 152.560 16.240 ;
        RECT 152.710 16.190 152.940 18.150 ;
        RECT 147.550 15.910 152.560 16.140 ;
        RECT 143.860 14.720 144.340 15.560 ;
        RECT 139.640 13.580 139.960 14.020 ;
        RECT 140.415 13.955 143.070 14.285 ;
        RECT 139.640 13.570 139.970 13.580 ;
        RECT 145.305 13.570 146.390 15.560 ;
        RECT 147.160 13.900 147.390 15.860 ;
        RECT 147.560 15.780 152.560 15.910 ;
        RECT 152.790 15.860 152.930 16.190 ;
        RECT 147.180 13.570 147.390 13.900 ;
        RECT 147.590 13.850 152.510 14.000 ;
        RECT 152.710 13.900 152.940 15.860 ;
        RECT 147.550 13.620 152.550 13.850 ;
        RECT 139.640 13.160 146.390 13.570 ;
        RECT 139.640 13.150 139.960 13.160 ;
        RECT 144.250 12.920 144.480 12.940 ;
        RECT 138.690 12.685 144.480 12.920 ;
        RECT 128.270 10.040 132.380 10.130 ;
        RECT 128.270 9.450 132.435 10.040 ;
        RECT 128.270 9.350 132.380 9.450 ;
        RECT 133.010 9.350 135.150 10.120 ;
        RECT 122.290 7.190 123.790 7.220 ;
        RECT 128.270 7.190 129.270 9.350 ;
        RECT 135.550 9.180 138.490 10.350 ;
        RECT 122.290 5.690 129.450 7.190 ;
        RECT 136.160 5.790 137.160 8.490 ;
        RECT 138.690 7.620 138.950 12.685 ;
        RECT 139.160 12.150 144.040 12.240 ;
        RECT 139.100 11.920 144.100 12.150 ;
        RECT 139.160 11.840 144.040 11.920 ;
        RECT 144.250 11.870 144.480 12.685 ;
        RECT 139.190 9.860 144.030 9.980 ;
        RECT 144.250 9.910 144.490 11.870 ;
        RECT 145.305 10.830 146.390 13.160 ;
        RECT 147.160 11.610 147.390 13.570 ;
        RECT 147.590 13.500 152.510 13.620 ;
        RECT 152.790 13.570 152.930 13.900 ;
        RECT 139.100 9.630 144.100 9.860 ;
        RECT 139.190 9.470 144.030 9.630 ;
        RECT 144.250 9.580 144.480 9.910 ;
        RECT 139.110 7.570 144.050 7.640 ;
        RECT 144.250 7.630 144.490 9.580 ;
        RECT 144.660 8.760 146.410 10.830 ;
        RECT 147.180 10.400 147.390 11.610 ;
        RECT 147.560 11.560 152.560 11.700 ;
        RECT 152.710 11.610 152.940 13.570 ;
        RECT 155.120 13.210 156.120 21.740 ;
        RECT 147.550 11.330 152.560 11.560 ;
        RECT 147.560 11.240 152.560 11.330 ;
        RECT 152.790 10.400 152.930 11.610 ;
        RECT 147.180 10.260 152.930 10.400 ;
        RECT 145.305 8.740 146.390 8.760 ;
        RECT 147.180 8.150 147.390 10.260 ;
        RECT 146.840 8.120 147.840 8.150 ;
        RECT 153.040 8.120 153.940 8.150 ;
        RECT 144.260 7.620 144.490 7.630 ;
        RECT 139.100 7.340 144.100 7.570 ;
        RECT 139.110 7.260 144.050 7.340 ;
        RECT 146.810 7.220 153.940 8.120 ;
        RECT 146.840 7.150 147.840 7.220 ;
        RECT 153.040 7.190 153.940 7.220 ;
        RECT 147.180 7.100 147.390 7.150 ;
        RECT 122.290 5.660 123.790 5.690 ;
        RECT 134.330 4.890 137.240 5.790 ;
        RECT 134.330 3.800 135.230 4.890 ;
        RECT 136.160 4.830 137.160 4.890 ;
        RECT 134.300 2.900 135.260 3.800 ;
      LAYER met2 ;
        RECT 154.790 27.755 156.290 27.780 ;
        RECT 131.265 26.630 132.115 26.650 ;
        RECT 131.240 25.730 133.330 26.630 ;
        RECT 154.770 26.305 156.310 27.755 ;
        RECT 131.265 25.710 132.115 25.730 ;
        RECT 154.790 24.960 156.290 26.305 ;
        RECT 136.130 23.530 137.190 24.530 ;
        RECT 144.000 24.350 145.840 24.360 ;
        RECT 139.080 24.050 146.040 24.350 ;
        RECT 139.080 23.990 144.120 24.050 ;
        RECT 132.980 22.220 135.240 22.290 ;
        RECT 136.160 22.220 137.160 23.530 ;
        RECT 132.980 22.000 137.900 22.220 ;
        RECT 139.100 22.000 144.090 22.100 ;
        RECT 132.980 21.720 144.090 22.000 ;
        RECT 132.980 21.510 137.900 21.720 ;
        RECT 139.100 21.660 144.090 21.720 ;
        RECT 132.980 21.440 135.240 21.510 ;
        RECT 145.530 20.790 146.040 24.050 ;
        RECT 145.530 20.760 147.920 20.790 ;
        RECT 145.530 20.510 152.530 20.760 ;
        RECT 139.100 19.720 144.110 19.730 ;
        RECT 145.530 19.720 146.040 20.510 ;
        RECT 147.520 20.480 152.530 20.510 ;
        RECT 139.100 19.410 146.040 19.720 ;
        RECT 139.100 19.380 144.110 19.410 ;
        RECT 145.530 16.120 146.040 19.410 ;
        RECT 147.580 18.410 152.540 18.500 ;
        RECT 147.580 18.140 154.360 18.410 ;
        RECT 147.580 18.100 152.540 18.140 ;
        RECT 147.510 16.120 152.610 16.190 ;
        RECT 145.530 15.840 152.610 16.120 ;
        RECT 131.980 13.810 132.260 13.845 ;
        RECT 131.970 13.510 133.030 13.810 ;
        RECT 131.980 13.475 132.260 13.510 ;
        RECT 139.110 12.150 144.090 12.190 ;
        RECT 145.530 12.150 146.040 15.840 ;
        RECT 147.510 15.830 152.610 15.840 ;
        RECT 154.090 14.240 154.360 18.140 ;
        RECT 147.540 13.880 152.560 13.950 ;
        RECT 154.000 13.880 156.150 14.240 ;
        RECT 147.540 13.610 156.150 13.880 ;
        RECT 147.540 13.550 152.560 13.610 ;
        RECT 154.000 13.240 156.150 13.610 ;
        RECT 139.110 11.950 146.040 12.150 ;
        RECT 139.110 11.890 144.090 11.950 ;
        RECT 145.530 11.550 146.040 11.950 ;
        RECT 147.510 11.550 152.610 11.650 ;
        RECT 145.530 11.290 152.610 11.550 ;
        RECT 145.530 11.270 147.920 11.290 ;
        RECT 135.050 10.070 137.870 10.080 ;
        RECT 132.960 9.940 137.870 10.070 ;
        RECT 132.960 9.930 139.200 9.940 ;
        RECT 132.960 9.540 144.080 9.930 ;
        RECT 132.960 9.400 137.870 9.540 ;
        RECT 139.140 9.520 144.080 9.540 ;
        RECT 136.160 8.460 137.160 9.400 ;
        RECT 136.130 7.460 137.190 8.460 ;
        RECT 139.060 7.540 144.100 7.590 ;
        RECT 145.530 7.540 146.040 11.270 ;
        RECT 154.805 8.120 155.655 8.140 ;
        RECT 139.060 7.360 146.040 7.540 ;
        RECT 139.060 7.340 145.810 7.360 ;
        RECT 139.060 7.310 144.100 7.340 ;
        RECT 153.010 7.220 155.680 8.120 ;
        RECT 120.505 7.190 121.955 7.210 ;
        RECT 154.805 7.200 155.655 7.220 ;
        RECT 120.480 5.690 123.820 7.190 ;
        RECT 120.505 5.670 121.955 5.690 ;
        RECT 134.330 2.855 135.230 3.830 ;
        RECT 134.310 2.005 135.250 2.855 ;
        RECT 134.330 1.980 135.230 2.005 ;
      LAYER met3 ;
        RECT 125.220 31.570 125.600 31.890 ;
        RECT 125.260 13.810 125.560 31.570 ;
        RECT 154.790 29.305 156.290 29.310 ;
        RECT 154.765 27.815 156.315 29.305 ;
        RECT 129.505 26.630 130.395 26.655 ;
        RECT 129.500 25.730 132.140 26.630 ;
        RECT 154.790 26.280 156.290 27.815 ;
        RECT 129.505 25.705 130.395 25.730 ;
        RECT 131.955 13.810 132.285 13.825 ;
        RECT 125.260 13.510 132.285 13.810 ;
        RECT 131.955 13.495 132.285 13.510 ;
        RECT 156.415 8.120 157.305 8.145 ;
        RECT 154.780 7.220 157.310 8.120 ;
        RECT 8.225 7.190 9.715 7.215 ;
        RECT 156.415 7.195 157.305 7.220 ;
        RECT 8.220 5.690 121.980 7.190 ;
        RECT 8.225 5.665 9.715 5.690 ;
        RECT 134.330 1.925 135.230 2.880 ;
        RECT 134.305 1.035 135.255 1.925 ;
        RECT 134.330 1.030 135.230 1.035 ;
      LAYER met4 ;
        RECT 3.990 224.150 4.290 224.760 ;
        RECT 7.670 224.150 7.970 224.760 ;
        RECT 11.350 224.150 11.650 224.760 ;
        RECT 15.030 224.150 15.330 224.760 ;
        RECT 18.710 224.150 19.010 224.760 ;
        RECT 22.390 224.150 22.690 224.760 ;
        RECT 26.070 224.150 26.370 224.760 ;
        RECT 29.750 224.150 30.050 224.760 ;
        RECT 33.430 224.150 33.730 224.760 ;
        RECT 37.110 224.150 37.410 224.760 ;
        RECT 40.790 224.150 41.090 224.760 ;
        RECT 44.470 224.150 44.770 224.760 ;
        RECT 48.150 224.150 48.450 224.760 ;
        RECT 51.830 224.150 52.130 224.760 ;
        RECT 55.510 224.150 55.810 224.760 ;
        RECT 59.190 224.150 59.490 224.760 ;
        RECT 62.870 224.150 63.170 224.760 ;
        RECT 66.550 224.150 66.850 224.760 ;
        RECT 70.230 224.150 70.530 224.760 ;
        RECT 73.910 224.150 74.210 224.760 ;
        RECT 77.590 224.150 77.890 224.760 ;
        RECT 81.270 224.150 81.570 224.760 ;
        RECT 84.950 224.150 85.250 224.760 ;
        RECT 88.630 224.150 88.930 224.760 ;
        RECT 3.585 223.700 90.530 224.150 ;
        RECT 3.990 223.680 4.290 223.700 ;
        RECT 7.670 223.670 7.970 223.700 ;
        RECT 63.500 219.770 65.000 223.700 ;
        RECT 50.500 218.270 65.000 219.770 ;
        RECT 147.510 32.570 147.810 224.760 ;
        RECT 125.250 32.270 147.810 32.570 ;
        RECT 125.260 31.895 125.560 32.270 ;
        RECT 125.245 31.565 125.575 31.895 ;
        RECT 50.500 29.030 156.290 30.530 ;
        RECT 154.790 27.810 156.290 29.030 ;
        RECT 112.250 25.730 130.400 26.630 ;
        RECT 2.500 5.690 9.720 7.190 ;
        RECT 112.250 1.000 113.150 25.730 ;
        RECT 134.330 1.000 135.230 1.930 ;
        RECT 156.410 1.000 157.310 8.120 ;
  END
END tt_um_brucemack_sb_mixer
END LIBRARY

