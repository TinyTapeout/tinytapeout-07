VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_ctrl
  CLASS BLOCK ;
  FOREIGN tt_ctrl ;
  ORIGIN 0.000 0.000 ;
  SIZE 184.000 BY 111.520 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 25.450 2.480 27.050 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.710 2.480 90.310 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 151.970 2.480 153.570 109.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.150 2.480 23.750 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 85.410 2.480 87.010 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 148.670 2.480 150.270 109.040 ;
    END
  END VPWR
  PIN ctrl_ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 26.990 0.000 27.290 1.000 ;
    END
  END ctrl_ena
  PIN ctrl_sel_inc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 25.150 0.000 25.450 1.000 ;
    END
  END ctrl_sel_inc
  PIN ctrl_sel_rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 23.310 0.000 23.610 1.000 ;
    END
  END ctrl_sel_rst_n
  PIN k_one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 19.630 0.000 19.930 1.000 ;
    END
  END k_one
  PIN k_zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 21.470 0.000 21.770 1.000 ;
    END
  END k_zero
  PIN pad_ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 163.150 0.000 163.450 1.000 ;
    END
  END pad_ui_in[0]
  PIN pad_ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 164.990 0.000 165.290 1.000 ;
    END
  END pad_ui_in[1]
  PIN pad_ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 178.790 110.520 179.090 111.520 ;
    END
  END pad_ui_in[2]
  PIN pad_ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 176.950 110.520 177.250 111.520 ;
    END
  END pad_ui_in[3]
  PIN pad_ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 175.110 110.520 175.410 111.520 ;
    END
  END pad_ui_in[4]
  PIN pad_ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 173.270 110.520 173.570 111.520 ;
    END
  END pad_ui_in[5]
  PIN pad_ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 171.430 110.520 171.730 111.520 ;
    END
  END pad_ui_in[6]
  PIN pad_ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 169.590 110.520 169.890 111.520 ;
    END
  END pad_ui_in[7]
  PIN pad_ui_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 167.750 110.520 168.050 111.520 ;
    END
  END pad_ui_in[8]
  PIN pad_ui_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 165.910 110.520 166.210 111.520 ;
    END
  END pad_ui_in[9]
  PIN pad_uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 30.670 110.520 30.970 111.520 ;
    END
  END pad_uio_in[0]
  PIN pad_uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 25.150 110.520 25.450 111.520 ;
    END
  END pad_uio_in[1]
  PIN pad_uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 19.630 110.520 19.930 111.520 ;
    END
  END pad_uio_in[2]
  PIN pad_uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 14.110 110.520 14.410 111.520 ;
    END
  END pad_uio_in[3]
  PIN pad_uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 8.590 110.520 8.890 111.520 ;
    END
  END pad_uio_in[4]
  PIN pad_uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 3.070 110.520 3.370 111.520 ;
    END
  END pad_uio_in[5]
  PIN pad_uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 8.590 0.000 8.890 1.000 ;
    END
  END pad_uio_in[6]
  PIN pad_uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 14.110 0.000 14.410 1.000 ;
    END
  END pad_uio_in[7]
  PIN pad_uio_oe_n[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 149.350 110.520 149.650 111.520 ;
    END
  END pad_uio_oe_n[0]
  PIN pad_uio_oe_n[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 28.830 110.520 29.130 111.520 ;
    END
  END pad_uio_oe_n[1]
  PIN pad_uio_oe_n[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 23.310 110.520 23.610 111.520 ;
    END
  END pad_uio_oe_n[2]
  PIN pad_uio_oe_n[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 17.790 110.520 18.090 111.520 ;
    END
  END pad_uio_oe_n[3]
  PIN pad_uio_oe_n[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 12.270 110.520 12.570 111.520 ;
    END
  END pad_uio_oe_n[4]
  PIN pad_uio_oe_n[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 6.750 110.520 7.050 111.520 ;
    END
  END pad_uio_oe_n[5]
  PIN pad_uio_oe_n[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 12.270 0.000 12.570 1.000 ;
    END
  END pad_uio_oe_n[6]
  PIN pad_uio_oe_n[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 17.790 0.000 18.090 1.000 ;
    END
  END pad_uio_oe_n[7]
  PIN pad_uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 32.510 110.520 32.810 111.520 ;
    END
  END pad_uio_out[0]
  PIN pad_uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 26.990 110.520 27.290 111.520 ;
    END
  END pad_uio_out[1]
  PIN pad_uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 21.470 110.520 21.770 111.520 ;
    END
  END pad_uio_out[2]
  PIN pad_uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 15.950 110.520 16.250 111.520 ;
    END
  END pad_uio_out[3]
  PIN pad_uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 10.430 110.520 10.730 111.520 ;
    END
  END pad_uio_out[4]
  PIN pad_uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 4.910 110.520 5.210 111.520 ;
    END
  END pad_uio_out[5]
  PIN pad_uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 10.430 0.000 10.730 1.000 ;
    END
  END pad_uio_out[6]
  PIN pad_uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 15.950 0.000 16.250 1.000 ;
    END
  END pad_uio_out[7]
  PIN pad_uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 164.070 110.520 164.370 111.520 ;
    END
  END pad_uo_out[0]
  PIN pad_uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 162.230 110.520 162.530 111.520 ;
    END
  END pad_uo_out[1]
  PIN pad_uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 160.390 110.520 160.690 111.520 ;
    END
  END pad_uo_out[2]
  PIN pad_uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 158.550 110.520 158.850 111.520 ;
    END
  END pad_uo_out[3]
  PIN pad_uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 156.710 110.520 157.010 111.520 ;
    END
  END pad_uo_out[4]
  PIN pad_uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 110.520 155.170 111.520 ;
    END
  END pad_uo_out[5]
  PIN pad_uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 153.030 110.520 153.330 111.520 ;
    END
  END pad_uo_out[6]
  PIN pad_uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 151.190 110.520 151.490 111.520 ;
    END
  END pad_uo_out[7]
  PIN spine_bot_iw[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 144.750 0.000 145.050 1.000 ;
    END
  END spine_bot_iw[0]
  PIN spine_bot_iw[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 126.350 0.000 126.650 1.000 ;
    END
  END spine_bot_iw[10]
  PIN spine_bot_iw[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 124.510 0.000 124.810 1.000 ;
    END
  END spine_bot_iw[11]
  PIN spine_bot_iw[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 122.670 0.000 122.970 1.000 ;
    END
  END spine_bot_iw[12]
  PIN spine_bot_iw[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 120.830 0.000 121.130 1.000 ;
    END
  END spine_bot_iw[13]
  PIN spine_bot_iw[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 118.990 0.000 119.290 1.000 ;
    END
  END spine_bot_iw[14]
  PIN spine_bot_iw[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 117.150 0.000 117.450 1.000 ;
    END
  END spine_bot_iw[15]
  PIN spine_bot_iw[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 115.310 0.000 115.610 1.000 ;
    END
  END spine_bot_iw[16]
  PIN spine_bot_iw[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 113.470 0.000 113.770 1.000 ;
    END
  END spine_bot_iw[17]
  PIN spine_bot_iw[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 111.630 0.000 111.930 1.000 ;
    END
  END spine_bot_iw[18]
  PIN spine_bot_iw[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 109.790 0.000 110.090 1.000 ;
    END
  END spine_bot_iw[19]
  PIN spine_bot_iw[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 142.910 0.000 143.210 1.000 ;
    END
  END spine_bot_iw[1]
  PIN spine_bot_iw[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 107.950 0.000 108.250 1.000 ;
    END
  END spine_bot_iw[20]
  PIN spine_bot_iw[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 106.110 0.000 106.410 1.000 ;
    END
  END spine_bot_iw[21]
  PIN spine_bot_iw[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 104.270 0.000 104.570 1.000 ;
    END
  END spine_bot_iw[22]
  PIN spine_bot_iw[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 102.430 0.000 102.730 1.000 ;
    END
  END spine_bot_iw[23]
  PIN spine_bot_iw[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 100.590 0.000 100.890 1.000 ;
    END
  END spine_bot_iw[24]
  PIN spine_bot_iw[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 98.750 0.000 99.050 1.000 ;
    END
  END spine_bot_iw[25]
  PIN spine_bot_iw[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 96.910 0.000 97.210 1.000 ;
    END
  END spine_bot_iw[26]
  PIN spine_bot_iw[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 95.070 0.000 95.370 1.000 ;
    END
  END spine_bot_iw[27]
  PIN spine_bot_iw[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 93.230 0.000 93.530 1.000 ;
    END
  END spine_bot_iw[28]
  PIN spine_bot_iw[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 0.000 91.690 1.000 ;
    END
  END spine_bot_iw[29]
  PIN spine_bot_iw[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 141.070 0.000 141.370 1.000 ;
    END
  END spine_bot_iw[2]
  PIN spine_bot_iw[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 139.230 0.000 139.530 1.000 ;
    END
  END spine_bot_iw[3]
  PIN spine_bot_iw[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 137.390 0.000 137.690 1.000 ;
    END
  END spine_bot_iw[4]
  PIN spine_bot_iw[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 0.000 135.850 1.000 ;
    END
  END spine_bot_iw[5]
  PIN spine_bot_iw[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 133.710 0.000 134.010 1.000 ;
    END
  END spine_bot_iw[6]
  PIN spine_bot_iw[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 131.870 0.000 132.170 1.000 ;
    END
  END spine_bot_iw[7]
  PIN spine_bot_iw[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 0.000 130.330 1.000 ;
    END
  END spine_bot_iw[8]
  PIN spine_bot_iw[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 128.190 0.000 128.490 1.000 ;
    END
  END spine_bot_iw[9]
  PIN spine_bot_ow[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 84.030 0.000 84.330 1.000 ;
    END
  END spine_bot_ow[0]
  PIN spine_bot_ow[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 65.630 0.000 65.930 1.000 ;
    END
  END spine_bot_ow[10]
  PIN spine_bot_ow[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 63.790 0.000 64.090 1.000 ;
    END
  END spine_bot_ow[11]
  PIN spine_bot_ow[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 61.950 0.000 62.250 1.000 ;
    END
  END spine_bot_ow[12]
  PIN spine_bot_ow[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 60.110 0.000 60.410 1.000 ;
    END
  END spine_bot_ow[13]
  PIN spine_bot_ow[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 58.270 0.000 58.570 1.000 ;
    END
  END spine_bot_ow[14]
  PIN spine_bot_ow[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 56.430 0.000 56.730 1.000 ;
    END
  END spine_bot_ow[15]
  PIN spine_bot_ow[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 54.590 0.000 54.890 1.000 ;
    END
  END spine_bot_ow[16]
  PIN spine_bot_ow[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 52.750 0.000 53.050 1.000 ;
    END
  END spine_bot_ow[17]
  PIN spine_bot_ow[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 50.910 0.000 51.210 1.000 ;
    END
  END spine_bot_ow[18]
  PIN spine_bot_ow[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 49.070 0.000 49.370 1.000 ;
    END
  END spine_bot_ow[19]
  PIN spine_bot_ow[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 82.190 0.000 82.490 1.000 ;
    END
  END spine_bot_ow[1]
  PIN spine_bot_ow[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 47.230 0.000 47.530 1.000 ;
    END
  END spine_bot_ow[20]
  PIN spine_bot_ow[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.470400 ;
    PORT
      LAYER met4 ;
        RECT 45.390 0.000 45.690 1.000 ;
    END
  END spine_bot_ow[21]
  PIN spine_bot_ow[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 43.550 0.000 43.850 1.000 ;
    END
  END spine_bot_ow[22]
  PIN spine_bot_ow[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 41.710 0.000 42.010 1.000 ;
    END
  END spine_bot_ow[23]
  PIN spine_bot_ow[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 39.870 0.000 40.170 1.000 ;
    END
  END spine_bot_ow[24]
  PIN spine_bot_ow[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 38.030 0.000 38.330 1.000 ;
    END
  END spine_bot_ow[25]
  PIN spine_bot_ow[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 80.350 0.000 80.650 1.000 ;
    END
  END spine_bot_ow[2]
  PIN spine_bot_ow[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 78.510 0.000 78.810 1.000 ;
    END
  END spine_bot_ow[3]
  PIN spine_bot_ow[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 76.670 0.000 76.970 1.000 ;
    END
  END spine_bot_ow[4]
  PIN spine_bot_ow[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 74.830 0.000 75.130 1.000 ;
    END
  END spine_bot_ow[5]
  PIN spine_bot_ow[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 72.990 0.000 73.290 1.000 ;
    END
  END spine_bot_ow[6]
  PIN spine_bot_ow[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 71.150 0.000 71.450 1.000 ;
    END
  END spine_bot_ow[7]
  PIN spine_bot_ow[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 69.310 0.000 69.610 1.000 ;
    END
  END spine_bot_ow[8]
  PIN spine_bot_ow[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 67.470 0.000 67.770 1.000 ;
    END
  END spine_bot_ow[9]
  PIN spine_top_iw[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 144.750 110.520 145.050 111.520 ;
    END
  END spine_top_iw[0]
  PIN spine_top_iw[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 126.350 110.520 126.650 111.520 ;
    END
  END spine_top_iw[10]
  PIN spine_top_iw[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 124.510 110.520 124.810 111.520 ;
    END
  END spine_top_iw[11]
  PIN spine_top_iw[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 122.670 110.520 122.970 111.520 ;
    END
  END spine_top_iw[12]
  PIN spine_top_iw[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 120.830 110.520 121.130 111.520 ;
    END
  END spine_top_iw[13]
  PIN spine_top_iw[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 118.990 110.520 119.290 111.520 ;
    END
  END spine_top_iw[14]
  PIN spine_top_iw[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 117.150 110.520 117.450 111.520 ;
    END
  END spine_top_iw[15]
  PIN spine_top_iw[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 115.310 110.520 115.610 111.520 ;
    END
  END spine_top_iw[16]
  PIN spine_top_iw[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 113.470 110.520 113.770 111.520 ;
    END
  END spine_top_iw[17]
  PIN spine_top_iw[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 111.630 110.520 111.930 111.520 ;
    END
  END spine_top_iw[18]
  PIN spine_top_iw[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 109.790 110.520 110.090 111.520 ;
    END
  END spine_top_iw[19]
  PIN spine_top_iw[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 142.910 110.520 143.210 111.520 ;
    END
  END spine_top_iw[1]
  PIN spine_top_iw[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 107.950 110.520 108.250 111.520 ;
    END
  END spine_top_iw[20]
  PIN spine_top_iw[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 106.110 110.520 106.410 111.520 ;
    END
  END spine_top_iw[21]
  PIN spine_top_iw[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 104.270 110.520 104.570 111.520 ;
    END
  END spine_top_iw[22]
  PIN spine_top_iw[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 102.430 110.520 102.730 111.520 ;
    END
  END spine_top_iw[23]
  PIN spine_top_iw[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 100.590 110.520 100.890 111.520 ;
    END
  END spine_top_iw[24]
  PIN spine_top_iw[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 98.750 110.520 99.050 111.520 ;
    END
  END spine_top_iw[25]
  PIN spine_top_iw[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 96.910 110.520 97.210 111.520 ;
    END
  END spine_top_iw[26]
  PIN spine_top_iw[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 95.070 110.520 95.370 111.520 ;
    END
  END spine_top_iw[27]
  PIN spine_top_iw[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 93.230 110.520 93.530 111.520 ;
    END
  END spine_top_iw[28]
  PIN spine_top_iw[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 110.520 91.690 111.520 ;
    END
  END spine_top_iw[29]
  PIN spine_top_iw[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 141.070 110.520 141.370 111.520 ;
    END
  END spine_top_iw[2]
  PIN spine_top_iw[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 139.230 110.520 139.530 111.520 ;
    END
  END spine_top_iw[3]
  PIN spine_top_iw[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 137.390 110.520 137.690 111.520 ;
    END
  END spine_top_iw[4]
  PIN spine_top_iw[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 110.520 135.850 111.520 ;
    END
  END spine_top_iw[5]
  PIN spine_top_iw[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 133.710 110.520 134.010 111.520 ;
    END
  END spine_top_iw[6]
  PIN spine_top_iw[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 131.870 110.520 132.170 111.520 ;
    END
  END spine_top_iw[7]
  PIN spine_top_iw[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 110.520 130.330 111.520 ;
    END
  END spine_top_iw[8]
  PIN spine_top_iw[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met4 ;
        RECT 128.190 110.520 128.490 111.520 ;
    END
  END spine_top_iw[9]
  PIN spine_top_ow[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 84.030 110.520 84.330 111.520 ;
    END
  END spine_top_ow[0]
  PIN spine_top_ow[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 65.630 110.520 65.930 111.520 ;
    END
  END spine_top_ow[10]
  PIN spine_top_ow[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 63.790 110.520 64.090 111.520 ;
    END
  END spine_top_ow[11]
  PIN spine_top_ow[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 61.950 110.520 62.250 111.520 ;
    END
  END spine_top_ow[12]
  PIN spine_top_ow[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 60.110 110.520 60.410 111.520 ;
    END
  END spine_top_ow[13]
  PIN spine_top_ow[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 58.270 110.520 58.570 111.520 ;
    END
  END spine_top_ow[14]
  PIN spine_top_ow[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 56.430 110.520 56.730 111.520 ;
    END
  END spine_top_ow[15]
  PIN spine_top_ow[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 54.590 110.520 54.890 111.520 ;
    END
  END spine_top_ow[16]
  PIN spine_top_ow[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 52.750 110.520 53.050 111.520 ;
    END
  END spine_top_ow[17]
  PIN spine_top_ow[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 50.910 110.520 51.210 111.520 ;
    END
  END spine_top_ow[18]
  PIN spine_top_ow[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 49.070 110.520 49.370 111.520 ;
    END
  END spine_top_ow[19]
  PIN spine_top_ow[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 82.190 110.520 82.490 111.520 ;
    END
  END spine_top_ow[1]
  PIN spine_top_ow[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 47.230 110.520 47.530 111.520 ;
    END
  END spine_top_ow[20]
  PIN spine_top_ow[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 45.390 110.520 45.690 111.520 ;
    END
  END spine_top_ow[21]
  PIN spine_top_ow[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 43.550 110.520 43.850 111.520 ;
    END
  END spine_top_ow[22]
  PIN spine_top_ow[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 41.710 110.520 42.010 111.520 ;
    END
  END spine_top_ow[23]
  PIN spine_top_ow[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 39.870 110.520 40.170 111.520 ;
    END
  END spine_top_ow[24]
  PIN spine_top_ow[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met4 ;
        RECT 38.030 110.520 38.330 111.520 ;
    END
  END spine_top_ow[25]
  PIN spine_top_ow[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 80.350 110.520 80.650 111.520 ;
    END
  END spine_top_ow[2]
  PIN spine_top_ow[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 78.510 110.520 78.810 111.520 ;
    END
  END spine_top_ow[3]
  PIN spine_top_ow[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 76.670 110.520 76.970 111.520 ;
    END
  END spine_top_ow[4]
  PIN spine_top_ow[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 74.830 110.520 75.130 111.520 ;
    END
  END spine_top_ow[5]
  PIN spine_top_ow[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 72.990 110.520 73.290 111.520 ;
    END
  END spine_top_ow[6]
  PIN spine_top_ow[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 71.150 110.520 71.450 111.520 ;
    END
  END spine_top_ow[7]
  PIN spine_top_ow[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 69.310 110.520 69.610 111.520 ;
    END
  END spine_top_ow[8]
  PIN spine_top_ow[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 1.035700 ;
    PORT
      LAYER met4 ;
        RECT 67.470 110.520 67.770 111.520 ;
    END
  END spine_top_ow[9]
  OBS
      LAYER nwell ;
        RECT 2.570 107.385 181.430 108.990 ;
        RECT 2.570 101.945 181.430 104.775 ;
        RECT 2.570 96.505 181.430 99.335 ;
        RECT 2.570 91.065 181.430 93.895 ;
        RECT 2.570 85.625 181.430 88.455 ;
        RECT 2.570 80.185 181.430 83.015 ;
        RECT 2.570 74.745 181.430 77.575 ;
        RECT 2.570 69.305 181.430 72.135 ;
        RECT 2.570 63.865 181.430 66.695 ;
        RECT 2.570 58.425 181.430 61.255 ;
        RECT 2.570 52.985 181.430 55.815 ;
        RECT 2.570 47.545 181.430 50.375 ;
        RECT 2.570 42.105 181.430 44.935 ;
        RECT 2.570 36.665 181.430 39.495 ;
        RECT 2.570 31.225 181.430 34.055 ;
        RECT 2.570 25.785 181.430 28.615 ;
        RECT 2.570 20.345 181.430 23.175 ;
        RECT 2.570 14.905 181.430 17.735 ;
        RECT 2.570 9.465 181.430 12.295 ;
        RECT 2.570 4.025 181.430 6.855 ;
      LAYER li1 ;
        RECT 2.760 2.635 181.240 108.885 ;
      LAYER met1 ;
        RECT 2.760 0.380 181.240 109.040 ;
      LAYER met2 ;
        RECT 6.070 0.155 174.710 110.005 ;
      LAYER met3 ;
        RECT 3.030 0.175 179.130 109.985 ;
      LAYER met4 ;
        RECT 3.770 110.120 4.510 110.650 ;
        RECT 5.610 110.120 6.350 110.650 ;
        RECT 7.450 110.120 8.190 110.650 ;
        RECT 9.290 110.120 10.030 110.650 ;
        RECT 11.130 110.120 11.870 110.650 ;
        RECT 12.970 110.120 13.710 110.650 ;
        RECT 14.810 110.120 15.550 110.650 ;
        RECT 16.650 110.120 17.390 110.650 ;
        RECT 18.490 110.120 19.230 110.650 ;
        RECT 20.330 110.120 21.070 110.650 ;
        RECT 22.170 110.120 22.910 110.650 ;
        RECT 24.010 110.120 24.750 110.650 ;
        RECT 25.850 110.120 26.590 110.650 ;
        RECT 27.690 110.120 28.430 110.650 ;
        RECT 29.530 110.120 30.270 110.650 ;
        RECT 31.370 110.120 32.110 110.650 ;
        RECT 33.210 110.120 37.630 110.650 ;
        RECT 38.730 110.120 39.470 110.650 ;
        RECT 40.570 110.120 41.310 110.650 ;
        RECT 42.410 110.120 43.150 110.650 ;
        RECT 44.250 110.120 44.990 110.650 ;
        RECT 46.090 110.120 46.830 110.650 ;
        RECT 47.930 110.120 48.670 110.650 ;
        RECT 49.770 110.120 50.510 110.650 ;
        RECT 51.610 110.120 52.350 110.650 ;
        RECT 53.450 110.120 54.190 110.650 ;
        RECT 55.290 110.120 56.030 110.650 ;
        RECT 57.130 110.120 57.870 110.650 ;
        RECT 58.970 110.120 59.710 110.650 ;
        RECT 60.810 110.120 61.550 110.650 ;
        RECT 62.650 110.120 63.390 110.650 ;
        RECT 64.490 110.120 65.230 110.650 ;
        RECT 66.330 110.120 67.070 110.650 ;
        RECT 68.170 110.120 68.910 110.650 ;
        RECT 70.010 110.120 70.750 110.650 ;
        RECT 71.850 110.120 72.590 110.650 ;
        RECT 73.690 110.120 74.430 110.650 ;
        RECT 75.530 110.120 76.270 110.650 ;
        RECT 77.370 110.120 78.110 110.650 ;
        RECT 79.210 110.120 79.950 110.650 ;
        RECT 81.050 110.120 81.790 110.650 ;
        RECT 82.890 110.120 83.630 110.650 ;
        RECT 84.730 110.120 90.990 110.650 ;
        RECT 92.090 110.120 92.830 110.650 ;
        RECT 93.930 110.120 94.670 110.650 ;
        RECT 95.770 110.120 96.510 110.650 ;
        RECT 97.610 110.120 98.350 110.650 ;
        RECT 99.450 110.120 100.190 110.650 ;
        RECT 101.290 110.120 102.030 110.650 ;
        RECT 103.130 110.120 103.870 110.650 ;
        RECT 104.970 110.120 105.710 110.650 ;
        RECT 106.810 110.120 107.550 110.650 ;
        RECT 108.650 110.120 109.390 110.650 ;
        RECT 110.490 110.120 111.230 110.650 ;
        RECT 112.330 110.120 113.070 110.650 ;
        RECT 114.170 110.120 114.910 110.650 ;
        RECT 116.010 110.120 116.750 110.650 ;
        RECT 117.850 110.120 118.590 110.650 ;
        RECT 119.690 110.120 120.430 110.650 ;
        RECT 121.530 110.120 122.270 110.650 ;
        RECT 123.370 110.120 124.110 110.650 ;
        RECT 125.210 110.120 125.950 110.650 ;
        RECT 127.050 110.120 127.790 110.650 ;
        RECT 128.890 110.120 129.630 110.650 ;
        RECT 130.730 110.120 131.470 110.650 ;
        RECT 132.570 110.120 133.310 110.650 ;
        RECT 134.410 110.120 135.150 110.650 ;
        RECT 136.250 110.120 136.990 110.650 ;
        RECT 138.090 110.120 138.830 110.650 ;
        RECT 139.930 110.120 140.670 110.650 ;
        RECT 141.770 110.120 142.510 110.650 ;
        RECT 143.610 110.120 144.350 110.650 ;
        RECT 145.450 110.120 148.950 110.650 ;
        RECT 150.050 110.120 150.790 110.650 ;
        RECT 151.890 110.120 152.630 110.650 ;
        RECT 153.730 110.120 154.470 110.650 ;
        RECT 155.570 110.120 156.310 110.650 ;
        RECT 157.410 110.120 158.150 110.650 ;
        RECT 159.250 110.120 159.990 110.650 ;
        RECT 161.090 110.120 161.830 110.650 ;
        RECT 162.930 110.120 163.670 110.650 ;
        RECT 164.770 110.120 165.510 110.650 ;
        RECT 166.610 110.120 167.350 110.650 ;
        RECT 168.450 110.120 169.190 110.650 ;
        RECT 170.290 110.120 171.030 110.650 ;
        RECT 172.130 110.120 172.870 110.650 ;
        RECT 173.970 110.120 174.710 110.650 ;
        RECT 175.810 110.120 176.550 110.650 ;
        RECT 177.650 110.120 178.390 110.650 ;
        RECT 3.055 109.440 179.105 110.120 ;
        RECT 3.055 2.080 21.750 109.440 ;
        RECT 24.150 2.080 25.050 109.440 ;
        RECT 27.450 2.080 85.010 109.440 ;
        RECT 87.410 2.080 88.310 109.440 ;
        RECT 90.710 2.080 148.270 109.440 ;
        RECT 150.670 2.080 151.570 109.440 ;
        RECT 153.970 2.080 179.105 109.440 ;
        RECT 3.055 1.400 179.105 2.080 ;
        RECT 3.055 0.175 8.190 1.400 ;
        RECT 9.290 0.175 10.030 1.400 ;
        RECT 11.130 0.175 11.870 1.400 ;
        RECT 12.970 0.175 13.710 1.400 ;
        RECT 14.810 0.175 15.550 1.400 ;
        RECT 16.650 0.175 17.390 1.400 ;
        RECT 18.490 0.175 19.230 1.400 ;
        RECT 20.330 0.175 21.070 1.400 ;
        RECT 22.170 0.175 22.910 1.400 ;
        RECT 24.010 0.175 24.750 1.400 ;
        RECT 25.850 0.175 26.590 1.400 ;
        RECT 27.690 0.175 37.630 1.400 ;
        RECT 38.730 0.175 39.470 1.400 ;
        RECT 40.570 0.175 41.310 1.400 ;
        RECT 42.410 0.175 43.150 1.400 ;
        RECT 44.250 0.175 44.990 1.400 ;
        RECT 46.090 0.175 46.830 1.400 ;
        RECT 47.930 0.175 48.670 1.400 ;
        RECT 49.770 0.175 50.510 1.400 ;
        RECT 51.610 0.175 52.350 1.400 ;
        RECT 53.450 0.175 54.190 1.400 ;
        RECT 55.290 0.175 56.030 1.400 ;
        RECT 57.130 0.175 57.870 1.400 ;
        RECT 58.970 0.175 59.710 1.400 ;
        RECT 60.810 0.175 61.550 1.400 ;
        RECT 62.650 0.175 63.390 1.400 ;
        RECT 64.490 0.175 65.230 1.400 ;
        RECT 66.330 0.175 67.070 1.400 ;
        RECT 68.170 0.175 68.910 1.400 ;
        RECT 70.010 0.175 70.750 1.400 ;
        RECT 71.850 0.175 72.590 1.400 ;
        RECT 73.690 0.175 74.430 1.400 ;
        RECT 75.530 0.175 76.270 1.400 ;
        RECT 77.370 0.175 78.110 1.400 ;
        RECT 79.210 0.175 79.950 1.400 ;
        RECT 81.050 0.175 81.790 1.400 ;
        RECT 82.890 0.175 83.630 1.400 ;
        RECT 84.730 0.175 90.990 1.400 ;
        RECT 92.090 0.175 92.830 1.400 ;
        RECT 93.930 0.175 94.670 1.400 ;
        RECT 95.770 0.175 96.510 1.400 ;
        RECT 97.610 0.175 98.350 1.400 ;
        RECT 99.450 0.175 100.190 1.400 ;
        RECT 101.290 0.175 102.030 1.400 ;
        RECT 103.130 0.175 103.870 1.400 ;
        RECT 104.970 0.175 105.710 1.400 ;
        RECT 106.810 0.175 107.550 1.400 ;
        RECT 108.650 0.175 109.390 1.400 ;
        RECT 110.490 0.175 111.230 1.400 ;
        RECT 112.330 0.175 113.070 1.400 ;
        RECT 114.170 0.175 114.910 1.400 ;
        RECT 116.010 0.175 116.750 1.400 ;
        RECT 117.850 0.175 118.590 1.400 ;
        RECT 119.690 0.175 120.430 1.400 ;
        RECT 121.530 0.175 122.270 1.400 ;
        RECT 123.370 0.175 124.110 1.400 ;
        RECT 125.210 0.175 125.950 1.400 ;
        RECT 127.050 0.175 127.790 1.400 ;
        RECT 128.890 0.175 129.630 1.400 ;
        RECT 130.730 0.175 131.470 1.400 ;
        RECT 132.570 0.175 133.310 1.400 ;
        RECT 134.410 0.175 135.150 1.400 ;
        RECT 136.250 0.175 136.990 1.400 ;
        RECT 138.090 0.175 138.830 1.400 ;
        RECT 139.930 0.175 140.670 1.400 ;
        RECT 141.770 0.175 142.510 1.400 ;
        RECT 143.610 0.175 144.350 1.400 ;
        RECT 145.450 0.175 162.750 1.400 ;
        RECT 163.850 0.175 164.590 1.400 ;
        RECT 165.690 0.175 179.105 1.400 ;
  END
END tt_ctrl
END LIBRARY

