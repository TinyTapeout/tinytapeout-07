module tt_mux (k_one,
    k_zero,
    addr,
    spine_iw,
    spine_ow,
    um_ena,
    um_iw,
    um_k_zero,
    um_ow,
    um_pg_vdd);
 output k_one;
 output k_zero;
 input [3:0] addr;
 input [29:0] spine_iw;
 output [25:0] spine_ow;
 output [15:0] um_ena;
 output [287:0] um_iw;
 output [15:0] um_k_zero;
 input [383:0] um_ow;
 output [15:0] um_pg_vdd;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire \block[0].genblk1.grp_sel_buf_I.a ;
 wire \block[0].genblk1.grp_sel_buf_I.z ;
 wire \block[0].genblk1.mux4_I[0].x ;
 wire \block[0].genblk1.mux4_I[10].x ;
 wire \block[0].genblk1.mux4_I[11].x ;
 wire \block[0].genblk1.mux4_I[12].x ;
 wire \block[0].genblk1.mux4_I[13].x ;
 wire \block[0].genblk1.mux4_I[14].x ;
 wire \block[0].genblk1.mux4_I[15].x ;
 wire \block[0].genblk1.mux4_I[16].x ;
 wire \block[0].genblk1.mux4_I[17].x ;
 wire \block[0].genblk1.mux4_I[18].x ;
 wire \block[0].genblk1.mux4_I[19].x ;
 wire \block[0].genblk1.mux4_I[1].x ;
 wire \block[0].genblk1.mux4_I[20].x ;
 wire \block[0].genblk1.mux4_I[21].x ;
 wire \block[0].genblk1.mux4_I[22].x ;
 wire \block[0].genblk1.mux4_I[23].x ;
 wire \block[0].genblk1.mux4_I[2].x ;
 wire \block[0].genblk1.mux4_I[3].x ;
 wire \block[0].genblk1.mux4_I[4].x ;
 wire \block[0].genblk1.mux4_I[5].x ;
 wire \block[0].genblk1.mux4_I[6].x ;
 wire \block[0].genblk1.mux4_I[7].x ;
 wire \block[0].genblk1.mux4_I[8].x ;
 wire \block[0].genblk1.mux4_I[9].x ;
 wire \block[0].genblk1.mux4_sel_buf_I[0].a ;
 wire \block[0].genblk1.mux4_sel_buf_I[0].z ;
 wire \block[0].genblk1.mux4_sel_buf_I[1].a ;
 wire \block[0].genblk1.mux4_sel_buf_I[1].z ;
 wire \block[0].genblk1.tbuf_blk_ena_I.tx ;
 wire \block[0].genblk1.tbuf_spine_ow_I[0].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[10].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[11].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[12].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[13].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[14].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[15].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[16].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[17].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[18].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[19].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[1].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[20].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[21].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[22].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[23].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[2].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[3].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[4].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[5].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[6].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[7].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[8].z ;
 wire \block[0].genblk1.tbuf_spine_ow_I[9].z ;
 wire \block[0].l_ena_0_I.a ;
 wire \block[0].l_ena_0_I.z ;
 wire \block[0].tie_I.hi ;
 wire \block[0].tie_I.lo ;
 wire \block[0].zbuf_bot_iw_I[0].a ;
 wire \block[0].zbuf_bot_iw_I[0].z ;
 wire \block[0].zbuf_bot_iw_I[10].a ;
 wire \block[0].zbuf_bot_iw_I[10].z ;
 wire \block[0].zbuf_bot_iw_I[11].a ;
 wire \block[0].zbuf_bot_iw_I[11].z ;
 wire \block[0].zbuf_bot_iw_I[12].a ;
 wire \block[0].zbuf_bot_iw_I[12].z ;
 wire \block[0].zbuf_bot_iw_I[13].a ;
 wire \block[0].zbuf_bot_iw_I[13].z ;
 wire \block[0].zbuf_bot_iw_I[14].a ;
 wire \block[0].zbuf_bot_iw_I[14].z ;
 wire \block[0].zbuf_bot_iw_I[15].a ;
 wire \block[0].zbuf_bot_iw_I[15].z ;
 wire \block[0].zbuf_bot_iw_I[16].a ;
 wire \block[0].zbuf_bot_iw_I[16].z ;
 wire \block[0].zbuf_bot_iw_I[17].a ;
 wire \block[0].zbuf_bot_iw_I[17].z ;
 wire \block[0].zbuf_bot_iw_I[1].a ;
 wire \block[0].zbuf_bot_iw_I[1].z ;
 wire \block[0].zbuf_bot_iw_I[2].a ;
 wire \block[0].zbuf_bot_iw_I[2].z ;
 wire \block[0].zbuf_bot_iw_I[3].a ;
 wire \block[0].zbuf_bot_iw_I[3].z ;
 wire \block[0].zbuf_bot_iw_I[4].a ;
 wire \block[0].zbuf_bot_iw_I[4].z ;
 wire \block[0].zbuf_bot_iw_I[5].a ;
 wire \block[0].zbuf_bot_iw_I[5].z ;
 wire \block[0].zbuf_bot_iw_I[6].a ;
 wire \block[0].zbuf_bot_iw_I[6].z ;
 wire \block[0].zbuf_bot_iw_I[7].a ;
 wire \block[0].zbuf_bot_iw_I[7].z ;
 wire \block[0].zbuf_bot_iw_I[8].a ;
 wire \block[0].zbuf_bot_iw_I[8].z ;
 wire \block[0].zbuf_bot_iw_I[9].a ;
 wire \block[0].zbuf_bot_iw_I[9].z ;
 wire \block[0].zbuf_ena_I.z ;
 wire \block[0].zbuf_pg_vdd_I.z ;
 wire \block[10].l_ena_0_I.a ;
 wire \block[10].l_ena_0_I.z ;
 wire \block[10].tie_I.hi ;
 wire \block[10].tie_I.lo ;
 wire \block[10].zbuf_bot_iw_I[0].z ;
 wire \block[10].zbuf_bot_iw_I[10].z ;
 wire \block[10].zbuf_bot_iw_I[11].z ;
 wire \block[10].zbuf_bot_iw_I[12].z ;
 wire \block[10].zbuf_bot_iw_I[13].z ;
 wire \block[10].zbuf_bot_iw_I[14].z ;
 wire \block[10].zbuf_bot_iw_I[15].z ;
 wire \block[10].zbuf_bot_iw_I[16].z ;
 wire \block[10].zbuf_bot_iw_I[17].z ;
 wire \block[10].zbuf_bot_iw_I[1].z ;
 wire \block[10].zbuf_bot_iw_I[2].z ;
 wire \block[10].zbuf_bot_iw_I[3].z ;
 wire \block[10].zbuf_bot_iw_I[4].z ;
 wire \block[10].zbuf_bot_iw_I[5].z ;
 wire \block[10].zbuf_bot_iw_I[6].z ;
 wire \block[10].zbuf_bot_iw_I[7].z ;
 wire \block[10].zbuf_bot_iw_I[8].z ;
 wire \block[10].zbuf_bot_iw_I[9].z ;
 wire \block[10].zbuf_ena_I.z ;
 wire \block[10].zbuf_pg_vdd_I.z ;
 wire \block[11].l_ena_0_I.a ;
 wire \block[11].l_ena_0_I.z ;
 wire \block[11].tie_I.hi ;
 wire \block[11].tie_I.lo ;
 wire \block[11].zbuf_bot_iw_I[0].z ;
 wire \block[11].zbuf_bot_iw_I[10].z ;
 wire \block[11].zbuf_bot_iw_I[11].z ;
 wire \block[11].zbuf_bot_iw_I[12].z ;
 wire \block[11].zbuf_bot_iw_I[13].z ;
 wire \block[11].zbuf_bot_iw_I[14].z ;
 wire \block[11].zbuf_bot_iw_I[15].z ;
 wire \block[11].zbuf_bot_iw_I[16].z ;
 wire \block[11].zbuf_bot_iw_I[17].z ;
 wire \block[11].zbuf_bot_iw_I[1].z ;
 wire \block[11].zbuf_bot_iw_I[2].z ;
 wire \block[11].zbuf_bot_iw_I[3].z ;
 wire \block[11].zbuf_bot_iw_I[4].z ;
 wire \block[11].zbuf_bot_iw_I[5].z ;
 wire \block[11].zbuf_bot_iw_I[6].z ;
 wire \block[11].zbuf_bot_iw_I[7].z ;
 wire \block[11].zbuf_bot_iw_I[8].z ;
 wire \block[11].zbuf_bot_iw_I[9].z ;
 wire \block[11].zbuf_ena_I.z ;
 wire \block[11].zbuf_pg_vdd_I.z ;
 wire \block[12].genblk1.grp_sel_buf_I.a ;
 wire \block[12].genblk1.grp_sel_buf_I.z ;
 wire \block[12].genblk1.mux4_I[0].x ;
 wire \block[12].genblk1.mux4_I[10].x ;
 wire \block[12].genblk1.mux4_I[11].x ;
 wire \block[12].genblk1.mux4_I[12].x ;
 wire \block[12].genblk1.mux4_I[13].x ;
 wire \block[12].genblk1.mux4_I[14].x ;
 wire \block[12].genblk1.mux4_I[15].x ;
 wire \block[12].genblk1.mux4_I[16].x ;
 wire \block[12].genblk1.mux4_I[17].x ;
 wire \block[12].genblk1.mux4_I[18].x ;
 wire \block[12].genblk1.mux4_I[19].x ;
 wire \block[12].genblk1.mux4_I[1].x ;
 wire \block[12].genblk1.mux4_I[20].x ;
 wire \block[12].genblk1.mux4_I[21].x ;
 wire \block[12].genblk1.mux4_I[22].x ;
 wire \block[12].genblk1.mux4_I[23].x ;
 wire \block[12].genblk1.mux4_I[2].x ;
 wire \block[12].genblk1.mux4_I[3].x ;
 wire \block[12].genblk1.mux4_I[4].x ;
 wire \block[12].genblk1.mux4_I[5].x ;
 wire \block[12].genblk1.mux4_I[6].x ;
 wire \block[12].genblk1.mux4_I[7].x ;
 wire \block[12].genblk1.mux4_I[8].x ;
 wire \block[12].genblk1.mux4_I[9].x ;
 wire \block[12].genblk1.mux4_sel_buf_I[0].z ;
 wire \block[12].genblk1.mux4_sel_buf_I[1].z ;
 wire \block[12].genblk1.tbuf_blk_ena_I.tx ;
 wire \block[12].l_ena_0_I.a ;
 wire \block[12].l_ena_0_I.z ;
 wire \block[12].tie_I.hi ;
 wire \block[12].tie_I.lo ;
 wire \block[12].zbuf_bot_iw_I[0].z ;
 wire \block[12].zbuf_bot_iw_I[10].z ;
 wire \block[12].zbuf_bot_iw_I[11].z ;
 wire \block[12].zbuf_bot_iw_I[12].z ;
 wire \block[12].zbuf_bot_iw_I[13].z ;
 wire \block[12].zbuf_bot_iw_I[14].z ;
 wire \block[12].zbuf_bot_iw_I[15].z ;
 wire \block[12].zbuf_bot_iw_I[16].z ;
 wire \block[12].zbuf_bot_iw_I[17].z ;
 wire \block[12].zbuf_bot_iw_I[1].z ;
 wire \block[12].zbuf_bot_iw_I[2].z ;
 wire \block[12].zbuf_bot_iw_I[3].z ;
 wire \block[12].zbuf_bot_iw_I[4].z ;
 wire \block[12].zbuf_bot_iw_I[5].z ;
 wire \block[12].zbuf_bot_iw_I[6].z ;
 wire \block[12].zbuf_bot_iw_I[7].z ;
 wire \block[12].zbuf_bot_iw_I[8].z ;
 wire \block[12].zbuf_bot_iw_I[9].z ;
 wire \block[12].zbuf_ena_I.z ;
 wire \block[12].zbuf_pg_vdd_I.z ;
 wire \block[13].l_ena_0_I.a ;
 wire \block[13].l_ena_0_I.z ;
 wire \block[13].tie_I.hi ;
 wire \block[13].tie_I.lo ;
 wire \block[13].zbuf_bot_iw_I[0].z ;
 wire \block[13].zbuf_bot_iw_I[10].z ;
 wire \block[13].zbuf_bot_iw_I[11].z ;
 wire \block[13].zbuf_bot_iw_I[12].z ;
 wire \block[13].zbuf_bot_iw_I[13].z ;
 wire \block[13].zbuf_bot_iw_I[14].z ;
 wire \block[13].zbuf_bot_iw_I[15].z ;
 wire \block[13].zbuf_bot_iw_I[16].z ;
 wire \block[13].zbuf_bot_iw_I[17].z ;
 wire \block[13].zbuf_bot_iw_I[1].z ;
 wire \block[13].zbuf_bot_iw_I[2].z ;
 wire \block[13].zbuf_bot_iw_I[3].z ;
 wire \block[13].zbuf_bot_iw_I[4].z ;
 wire \block[13].zbuf_bot_iw_I[5].z ;
 wire \block[13].zbuf_bot_iw_I[6].z ;
 wire \block[13].zbuf_bot_iw_I[7].z ;
 wire \block[13].zbuf_bot_iw_I[8].z ;
 wire \block[13].zbuf_bot_iw_I[9].z ;
 wire \block[13].zbuf_ena_I.z ;
 wire \block[13].zbuf_pg_vdd_I.z ;
 wire \block[14].l_ena_0_I.a ;
 wire \block[14].l_ena_0_I.z ;
 wire \block[14].tie_I.hi ;
 wire \block[14].tie_I.lo ;
 wire \block[14].zbuf_bot_iw_I[0].z ;
 wire \block[14].zbuf_bot_iw_I[10].z ;
 wire \block[14].zbuf_bot_iw_I[11].z ;
 wire \block[14].zbuf_bot_iw_I[12].z ;
 wire \block[14].zbuf_bot_iw_I[13].z ;
 wire \block[14].zbuf_bot_iw_I[14].z ;
 wire \block[14].zbuf_bot_iw_I[15].z ;
 wire \block[14].zbuf_bot_iw_I[16].z ;
 wire \block[14].zbuf_bot_iw_I[17].z ;
 wire \block[14].zbuf_bot_iw_I[1].z ;
 wire \block[14].zbuf_bot_iw_I[2].z ;
 wire \block[14].zbuf_bot_iw_I[3].z ;
 wire \block[14].zbuf_bot_iw_I[4].z ;
 wire \block[14].zbuf_bot_iw_I[5].z ;
 wire \block[14].zbuf_bot_iw_I[6].z ;
 wire \block[14].zbuf_bot_iw_I[7].z ;
 wire \block[14].zbuf_bot_iw_I[8].z ;
 wire \block[14].zbuf_bot_iw_I[9].z ;
 wire \block[14].zbuf_ena_I.z ;
 wire \block[14].zbuf_pg_vdd_I.z ;
 wire \block[15].l_ena_0_I.a ;
 wire \block[15].l_ena_0_I.z ;
 wire \block[15].tie_I.hi ;
 wire \block[15].tie_I.lo ;
 wire \block[15].zbuf_bot_iw_I[0].z ;
 wire \block[15].zbuf_bot_iw_I[10].z ;
 wire \block[15].zbuf_bot_iw_I[11].z ;
 wire \block[15].zbuf_bot_iw_I[12].z ;
 wire \block[15].zbuf_bot_iw_I[13].z ;
 wire \block[15].zbuf_bot_iw_I[14].z ;
 wire \block[15].zbuf_bot_iw_I[15].z ;
 wire \block[15].zbuf_bot_iw_I[16].z ;
 wire \block[15].zbuf_bot_iw_I[17].z ;
 wire \block[15].zbuf_bot_iw_I[1].z ;
 wire \block[15].zbuf_bot_iw_I[2].z ;
 wire \block[15].zbuf_bot_iw_I[3].z ;
 wire \block[15].zbuf_bot_iw_I[4].z ;
 wire \block[15].zbuf_bot_iw_I[5].z ;
 wire \block[15].zbuf_bot_iw_I[6].z ;
 wire \block[15].zbuf_bot_iw_I[7].z ;
 wire \block[15].zbuf_bot_iw_I[8].z ;
 wire \block[15].zbuf_bot_iw_I[9].z ;
 wire \block[15].zbuf_ena_I.z ;
 wire \block[15].zbuf_pg_vdd_I.z ;
 wire \block[1].l_ena_0_I.a ;
 wire \block[1].l_ena_0_I.z ;
 wire \block[1].tie_I.hi ;
 wire \block[1].tie_I.lo ;
 wire \block[1].zbuf_bot_iw_I[0].z ;
 wire \block[1].zbuf_bot_iw_I[10].z ;
 wire \block[1].zbuf_bot_iw_I[11].z ;
 wire \block[1].zbuf_bot_iw_I[12].z ;
 wire \block[1].zbuf_bot_iw_I[13].z ;
 wire \block[1].zbuf_bot_iw_I[14].z ;
 wire \block[1].zbuf_bot_iw_I[15].z ;
 wire \block[1].zbuf_bot_iw_I[16].z ;
 wire \block[1].zbuf_bot_iw_I[17].z ;
 wire \block[1].zbuf_bot_iw_I[1].z ;
 wire \block[1].zbuf_bot_iw_I[2].z ;
 wire \block[1].zbuf_bot_iw_I[3].z ;
 wire \block[1].zbuf_bot_iw_I[4].z ;
 wire \block[1].zbuf_bot_iw_I[5].z ;
 wire \block[1].zbuf_bot_iw_I[6].z ;
 wire \block[1].zbuf_bot_iw_I[7].z ;
 wire \block[1].zbuf_bot_iw_I[8].z ;
 wire \block[1].zbuf_bot_iw_I[9].z ;
 wire \block[1].zbuf_ena_I.z ;
 wire \block[1].zbuf_pg_vdd_I.z ;
 wire \block[2].l_ena_0_I.a ;
 wire \block[2].l_ena_0_I.z ;
 wire \block[2].tie_I.hi ;
 wire \block[2].tie_I.lo ;
 wire \block[2].zbuf_bot_iw_I[0].z ;
 wire \block[2].zbuf_bot_iw_I[10].z ;
 wire \block[2].zbuf_bot_iw_I[11].z ;
 wire \block[2].zbuf_bot_iw_I[12].z ;
 wire \block[2].zbuf_bot_iw_I[13].z ;
 wire \block[2].zbuf_bot_iw_I[14].z ;
 wire \block[2].zbuf_bot_iw_I[15].z ;
 wire \block[2].zbuf_bot_iw_I[16].z ;
 wire \block[2].zbuf_bot_iw_I[17].z ;
 wire \block[2].zbuf_bot_iw_I[1].z ;
 wire \block[2].zbuf_bot_iw_I[2].z ;
 wire \block[2].zbuf_bot_iw_I[3].z ;
 wire \block[2].zbuf_bot_iw_I[4].z ;
 wire \block[2].zbuf_bot_iw_I[5].z ;
 wire \block[2].zbuf_bot_iw_I[6].z ;
 wire \block[2].zbuf_bot_iw_I[7].z ;
 wire \block[2].zbuf_bot_iw_I[8].z ;
 wire \block[2].zbuf_bot_iw_I[9].z ;
 wire \block[2].zbuf_ena_I.z ;
 wire \block[2].zbuf_pg_vdd_I.z ;
 wire \block[3].l_ena_0_I.a ;
 wire \block[3].l_ena_0_I.z ;
 wire \block[3].tie_I.hi ;
 wire \block[3].tie_I.lo ;
 wire \block[3].zbuf_bot_iw_I[0].z ;
 wire \block[3].zbuf_bot_iw_I[10].z ;
 wire \block[3].zbuf_bot_iw_I[11].z ;
 wire \block[3].zbuf_bot_iw_I[12].z ;
 wire \block[3].zbuf_bot_iw_I[13].z ;
 wire \block[3].zbuf_bot_iw_I[14].z ;
 wire \block[3].zbuf_bot_iw_I[15].z ;
 wire \block[3].zbuf_bot_iw_I[16].z ;
 wire \block[3].zbuf_bot_iw_I[17].z ;
 wire \block[3].zbuf_bot_iw_I[1].z ;
 wire \block[3].zbuf_bot_iw_I[2].z ;
 wire \block[3].zbuf_bot_iw_I[3].z ;
 wire \block[3].zbuf_bot_iw_I[4].z ;
 wire \block[3].zbuf_bot_iw_I[5].z ;
 wire \block[3].zbuf_bot_iw_I[6].z ;
 wire \block[3].zbuf_bot_iw_I[7].z ;
 wire \block[3].zbuf_bot_iw_I[8].z ;
 wire \block[3].zbuf_bot_iw_I[9].z ;
 wire \block[3].zbuf_ena_I.z ;
 wire \block[3].zbuf_pg_vdd_I.z ;
 wire \block[4].genblk1.grp_sel_buf_I.a ;
 wire \block[4].genblk1.grp_sel_buf_I.z ;
 wire \block[4].genblk1.mux4_I[0].x ;
 wire \block[4].genblk1.mux4_I[10].x ;
 wire \block[4].genblk1.mux4_I[11].x ;
 wire \block[4].genblk1.mux4_I[12].x ;
 wire \block[4].genblk1.mux4_I[13].x ;
 wire \block[4].genblk1.mux4_I[14].x ;
 wire \block[4].genblk1.mux4_I[15].x ;
 wire \block[4].genblk1.mux4_I[16].x ;
 wire \block[4].genblk1.mux4_I[17].x ;
 wire \block[4].genblk1.mux4_I[18].x ;
 wire \block[4].genblk1.mux4_I[19].x ;
 wire \block[4].genblk1.mux4_I[1].x ;
 wire \block[4].genblk1.mux4_I[20].x ;
 wire \block[4].genblk1.mux4_I[21].x ;
 wire \block[4].genblk1.mux4_I[22].x ;
 wire \block[4].genblk1.mux4_I[23].x ;
 wire \block[4].genblk1.mux4_I[2].x ;
 wire \block[4].genblk1.mux4_I[3].x ;
 wire \block[4].genblk1.mux4_I[4].x ;
 wire \block[4].genblk1.mux4_I[5].x ;
 wire \block[4].genblk1.mux4_I[6].x ;
 wire \block[4].genblk1.mux4_I[7].x ;
 wire \block[4].genblk1.mux4_I[8].x ;
 wire \block[4].genblk1.mux4_I[9].x ;
 wire \block[4].genblk1.mux4_sel_buf_I[0].z ;
 wire \block[4].genblk1.mux4_sel_buf_I[1].z ;
 wire \block[4].genblk1.tbuf_blk_ena_I.tx ;
 wire \block[4].l_ena_0_I.a ;
 wire \block[4].l_ena_0_I.z ;
 wire \block[4].tie_I.hi ;
 wire \block[4].tie_I.lo ;
 wire \block[4].zbuf_bot_iw_I[0].z ;
 wire \block[4].zbuf_bot_iw_I[10].z ;
 wire \block[4].zbuf_bot_iw_I[11].z ;
 wire \block[4].zbuf_bot_iw_I[12].z ;
 wire \block[4].zbuf_bot_iw_I[13].z ;
 wire \block[4].zbuf_bot_iw_I[14].z ;
 wire \block[4].zbuf_bot_iw_I[15].z ;
 wire \block[4].zbuf_bot_iw_I[16].z ;
 wire \block[4].zbuf_bot_iw_I[17].z ;
 wire \block[4].zbuf_bot_iw_I[1].z ;
 wire \block[4].zbuf_bot_iw_I[2].z ;
 wire \block[4].zbuf_bot_iw_I[3].z ;
 wire \block[4].zbuf_bot_iw_I[4].z ;
 wire \block[4].zbuf_bot_iw_I[5].z ;
 wire \block[4].zbuf_bot_iw_I[6].z ;
 wire \block[4].zbuf_bot_iw_I[7].z ;
 wire \block[4].zbuf_bot_iw_I[8].z ;
 wire \block[4].zbuf_bot_iw_I[9].z ;
 wire \block[4].zbuf_ena_I.z ;
 wire \block[4].zbuf_pg_vdd_I.z ;
 wire \block[5].l_ena_0_I.a ;
 wire \block[5].l_ena_0_I.z ;
 wire \block[5].tie_I.hi ;
 wire \block[5].tie_I.lo ;
 wire \block[5].zbuf_bot_iw_I[0].z ;
 wire \block[5].zbuf_bot_iw_I[10].z ;
 wire \block[5].zbuf_bot_iw_I[11].z ;
 wire \block[5].zbuf_bot_iw_I[12].z ;
 wire \block[5].zbuf_bot_iw_I[13].z ;
 wire \block[5].zbuf_bot_iw_I[14].z ;
 wire \block[5].zbuf_bot_iw_I[15].z ;
 wire \block[5].zbuf_bot_iw_I[16].z ;
 wire \block[5].zbuf_bot_iw_I[17].z ;
 wire \block[5].zbuf_bot_iw_I[1].z ;
 wire \block[5].zbuf_bot_iw_I[2].z ;
 wire \block[5].zbuf_bot_iw_I[3].z ;
 wire \block[5].zbuf_bot_iw_I[4].z ;
 wire \block[5].zbuf_bot_iw_I[5].z ;
 wire \block[5].zbuf_bot_iw_I[6].z ;
 wire \block[5].zbuf_bot_iw_I[7].z ;
 wire \block[5].zbuf_bot_iw_I[8].z ;
 wire \block[5].zbuf_bot_iw_I[9].z ;
 wire \block[5].zbuf_ena_I.z ;
 wire \block[5].zbuf_pg_vdd_I.z ;
 wire \block[6].l_ena_0_I.a ;
 wire \block[6].l_ena_0_I.z ;
 wire \block[6].tie_I.hi ;
 wire \block[6].tie_I.lo ;
 wire \block[6].zbuf_bot_iw_I[0].z ;
 wire \block[6].zbuf_bot_iw_I[10].z ;
 wire \block[6].zbuf_bot_iw_I[11].z ;
 wire \block[6].zbuf_bot_iw_I[12].z ;
 wire \block[6].zbuf_bot_iw_I[13].z ;
 wire \block[6].zbuf_bot_iw_I[14].z ;
 wire \block[6].zbuf_bot_iw_I[15].z ;
 wire \block[6].zbuf_bot_iw_I[16].z ;
 wire \block[6].zbuf_bot_iw_I[17].z ;
 wire \block[6].zbuf_bot_iw_I[1].z ;
 wire \block[6].zbuf_bot_iw_I[2].z ;
 wire \block[6].zbuf_bot_iw_I[3].z ;
 wire \block[6].zbuf_bot_iw_I[4].z ;
 wire \block[6].zbuf_bot_iw_I[5].z ;
 wire \block[6].zbuf_bot_iw_I[6].z ;
 wire \block[6].zbuf_bot_iw_I[7].z ;
 wire \block[6].zbuf_bot_iw_I[8].z ;
 wire \block[6].zbuf_bot_iw_I[9].z ;
 wire \block[6].zbuf_ena_I.z ;
 wire \block[6].zbuf_pg_vdd_I.z ;
 wire \block[7].l_ena_0_I.a ;
 wire \block[7].l_ena_0_I.z ;
 wire \block[7].tie_I.hi ;
 wire \block[7].tie_I.lo ;
 wire \block[7].zbuf_bot_iw_I[0].z ;
 wire \block[7].zbuf_bot_iw_I[10].z ;
 wire \block[7].zbuf_bot_iw_I[11].z ;
 wire \block[7].zbuf_bot_iw_I[12].z ;
 wire \block[7].zbuf_bot_iw_I[13].z ;
 wire \block[7].zbuf_bot_iw_I[14].z ;
 wire \block[7].zbuf_bot_iw_I[15].z ;
 wire \block[7].zbuf_bot_iw_I[16].z ;
 wire \block[7].zbuf_bot_iw_I[17].z ;
 wire \block[7].zbuf_bot_iw_I[1].z ;
 wire \block[7].zbuf_bot_iw_I[2].z ;
 wire \block[7].zbuf_bot_iw_I[3].z ;
 wire \block[7].zbuf_bot_iw_I[4].z ;
 wire \block[7].zbuf_bot_iw_I[5].z ;
 wire \block[7].zbuf_bot_iw_I[6].z ;
 wire \block[7].zbuf_bot_iw_I[7].z ;
 wire \block[7].zbuf_bot_iw_I[8].z ;
 wire \block[7].zbuf_bot_iw_I[9].z ;
 wire \block[7].zbuf_ena_I.z ;
 wire \block[7].zbuf_pg_vdd_I.z ;
 wire \block[8].genblk1.grp_sel_buf_I.a ;
 wire \block[8].genblk1.grp_sel_buf_I.z ;
 wire \block[8].genblk1.mux4_I[0].x ;
 wire \block[8].genblk1.mux4_I[10].x ;
 wire \block[8].genblk1.mux4_I[11].x ;
 wire \block[8].genblk1.mux4_I[12].x ;
 wire \block[8].genblk1.mux4_I[13].x ;
 wire \block[8].genblk1.mux4_I[14].x ;
 wire \block[8].genblk1.mux4_I[15].x ;
 wire \block[8].genblk1.mux4_I[16].x ;
 wire \block[8].genblk1.mux4_I[17].x ;
 wire \block[8].genblk1.mux4_I[18].x ;
 wire \block[8].genblk1.mux4_I[19].x ;
 wire \block[8].genblk1.mux4_I[1].x ;
 wire \block[8].genblk1.mux4_I[20].x ;
 wire \block[8].genblk1.mux4_I[21].x ;
 wire \block[8].genblk1.mux4_I[22].x ;
 wire \block[8].genblk1.mux4_I[23].x ;
 wire \block[8].genblk1.mux4_I[2].x ;
 wire \block[8].genblk1.mux4_I[3].x ;
 wire \block[8].genblk1.mux4_I[4].x ;
 wire \block[8].genblk1.mux4_I[5].x ;
 wire \block[8].genblk1.mux4_I[6].x ;
 wire \block[8].genblk1.mux4_I[7].x ;
 wire \block[8].genblk1.mux4_I[8].x ;
 wire \block[8].genblk1.mux4_I[9].x ;
 wire \block[8].genblk1.mux4_sel_buf_I[0].z ;
 wire \block[8].genblk1.mux4_sel_buf_I[1].z ;
 wire \block[8].genblk1.tbuf_blk_ena_I.tx ;
 wire \block[8].l_ena_0_I.a ;
 wire \block[8].l_ena_0_I.z ;
 wire \block[8].tie_I.hi ;
 wire \block[8].tie_I.lo ;
 wire \block[8].zbuf_bot_iw_I[0].z ;
 wire \block[8].zbuf_bot_iw_I[10].z ;
 wire \block[8].zbuf_bot_iw_I[11].z ;
 wire \block[8].zbuf_bot_iw_I[12].z ;
 wire \block[8].zbuf_bot_iw_I[13].z ;
 wire \block[8].zbuf_bot_iw_I[14].z ;
 wire \block[8].zbuf_bot_iw_I[15].z ;
 wire \block[8].zbuf_bot_iw_I[16].z ;
 wire \block[8].zbuf_bot_iw_I[17].z ;
 wire \block[8].zbuf_bot_iw_I[1].z ;
 wire \block[8].zbuf_bot_iw_I[2].z ;
 wire \block[8].zbuf_bot_iw_I[3].z ;
 wire \block[8].zbuf_bot_iw_I[4].z ;
 wire \block[8].zbuf_bot_iw_I[5].z ;
 wire \block[8].zbuf_bot_iw_I[6].z ;
 wire \block[8].zbuf_bot_iw_I[7].z ;
 wire \block[8].zbuf_bot_iw_I[8].z ;
 wire \block[8].zbuf_bot_iw_I[9].z ;
 wire \block[8].zbuf_ena_I.z ;
 wire \block[8].zbuf_pg_vdd_I.z ;
 wire \block[9].l_ena_0_I.a ;
 wire \block[9].l_ena_0_I.z ;
 wire \block[9].tie_I.hi ;
 wire \block[9].tie_I.lo ;
 wire \block[9].zbuf_bot_iw_I[0].z ;
 wire \block[9].zbuf_bot_iw_I[10].z ;
 wire \block[9].zbuf_bot_iw_I[11].z ;
 wire \block[9].zbuf_bot_iw_I[12].z ;
 wire \block[9].zbuf_bot_iw_I[13].z ;
 wire \block[9].zbuf_bot_iw_I[14].z ;
 wire \block[9].zbuf_bot_iw_I[15].z ;
 wire \block[9].zbuf_bot_iw_I[16].z ;
 wire \block[9].zbuf_bot_iw_I[17].z ;
 wire \block[9].zbuf_bot_iw_I[1].z ;
 wire \block[9].zbuf_bot_iw_I[2].z ;
 wire \block[9].zbuf_bot_iw_I[3].z ;
 wire \block[9].zbuf_bot_iw_I[4].z ;
 wire \block[9].zbuf_bot_iw_I[5].z ;
 wire \block[9].zbuf_bot_iw_I[6].z ;
 wire \block[9].zbuf_bot_iw_I[7].z ;
 wire \block[9].zbuf_bot_iw_I[8].z ;
 wire \block[9].zbuf_bot_iw_I[9].z ;
 wire \block[9].zbuf_ena_I.z ;
 wire \block[9].zbuf_pg_vdd_I.z ;
 wire \branch_addr_match_buf_I[0].z ;
 wire \branch_addr_match_buf_I[1].z ;
 wire \branch_addr_match_buf_I[2].z ;
 wire \branch_addr_match_buf_I[3].z ;
 wire \branch_ena_buf_I.z ;
 wire \branch_sel_buf_I.a ;
 wire \branch_sel_buf_I.z ;
 wire \branch_sel_n_buf_I.z ;
 wire \buf_bus_ena_I.z ;
 wire \buf_spine_ow_I[0].z ;
 wire \buf_spine_ow_I[10].z ;
 wire \buf_spine_ow_I[11].z ;
 wire \buf_spine_ow_I[12].z ;
 wire \buf_spine_ow_I[13].z ;
 wire \buf_spine_ow_I[14].z ;
 wire \buf_spine_ow_I[15].z ;
 wire \buf_spine_ow_I[16].z ;
 wire \buf_spine_ow_I[17].z ;
 wire \buf_spine_ow_I[18].z ;
 wire \buf_spine_ow_I[19].z ;
 wire \buf_spine_ow_I[1].z ;
 wire \buf_spine_ow_I[20].z ;
 wire \buf_spine_ow_I[21].z ;
 wire \buf_spine_ow_I[22].z ;
 wire \buf_spine_ow_I[23].z ;
 wire \buf_spine_ow_I[2].z ;
 wire \buf_spine_ow_I[3].z ;
 wire \buf_spine_ow_I[4].z ;
 wire \buf_spine_ow_I[5].z ;
 wire \buf_spine_ow_I[6].z ;
 wire \buf_spine_ow_I[7].z ;
 wire \buf_spine_ow_I[8].z ;
 wire \buf_spine_ow_I[9].z ;
 wire \bus_pull_ow_I[0].a ;
 wire \bus_pull_ow_I[0].tx ;
 wire \bus_pull_tie_I.hi ;
 wire one_;
 wire \tbuf_row_ena_I.tx ;
 wire \tbuf_spine_ow_I[0].z ;
 wire \tbuf_spine_ow_I[10].z ;
 wire \tbuf_spine_ow_I[11].z ;
 wire \tbuf_spine_ow_I[12].z ;
 wire \tbuf_spine_ow_I[13].z ;
 wire \tbuf_spine_ow_I[14].z ;
 wire \tbuf_spine_ow_I[15].z ;
 wire \tbuf_spine_ow_I[16].z ;
 wire \tbuf_spine_ow_I[17].z ;
 wire \tbuf_spine_ow_I[18].z ;
 wire \tbuf_spine_ow_I[19].z ;
 wire \tbuf_spine_ow_I[1].z ;
 wire \tbuf_spine_ow_I[20].z ;
 wire \tbuf_spine_ow_I[21].z ;
 wire \tbuf_spine_ow_I[22].z ;
 wire \tbuf_spine_ow_I[23].z ;
 wire \tbuf_spine_ow_I[2].z ;
 wire \tbuf_spine_ow_I[3].z ;
 wire \tbuf_spine_ow_I[4].z ;
 wire \tbuf_spine_ow_I[5].z ;
 wire \tbuf_spine_ow_I[6].z ;
 wire \tbuf_spine_ow_I[7].z ;
 wire \tbuf_spine_ow_I[8].z ;
 wire \tbuf_spine_ow_I[9].z ;
 wire \tie_spine_guard_I[0].hi ;
 wire \tie_spine_guard_I[0].lo ;
 wire \tie_spine_guard_I[1].hi ;
 wire \tie_spine_guard_I[1].lo ;
 wire \zbuf_bus_iw_I[0].genblk1.l ;
 wire \zbuf_bus_iw_I[10].genblk1.l ;
 wire \zbuf_bus_iw_I[11].genblk1.l ;
 wire \zbuf_bus_iw_I[12].genblk1.l ;
 wire \zbuf_bus_iw_I[13].genblk1.l ;
 wire \zbuf_bus_iw_I[14].genblk1.l ;
 wire \zbuf_bus_iw_I[15].genblk1.l ;
 wire \zbuf_bus_iw_I[16].genblk1.l ;
 wire \zbuf_bus_iw_I[17].genblk1.l ;
 wire \zbuf_bus_iw_I[1].genblk1.l ;
 wire \zbuf_bus_iw_I[2].genblk1.l ;
 wire \zbuf_bus_iw_I[3].genblk1.l ;
 wire \zbuf_bus_iw_I[4].genblk1.l ;
 wire \zbuf_bus_iw_I[5].genblk1.l ;
 wire \zbuf_bus_iw_I[6].genblk1.l ;
 wire \zbuf_bus_iw_I[7].genblk1.l ;
 wire \zbuf_bus_iw_I[8].genblk1.l ;
 wire \zbuf_bus_iw_I[9].genblk1.l ;
 wire \zbuf_bus_sel_I[0].genblk1.l ;
 wire \zbuf_bus_sel_I[1].genblk1.l ;
 wire \zbuf_bus_sel_I[2].genblk1.l ;
 wire \zbuf_bus_sel_I[2].z ;
 wire \zbuf_bus_sel_I[3].genblk1.l ;
 wire \zbuf_bus_sel_I[3].z ;
 wire \zbuf_bus_sel_I[4].genblk1.l ;
 wire \zbuf_bus_sel_I[4].z ;

 sky130_fd_sc_hd__clkinv_1 _09_ (.A(\branch_addr_match_buf_I[0].z ),
    .Y(_00_));
 sky130_fd_sc_hd__clkinv_1 _10_ (.A(\branch_addr_match_buf_I[1].z ),
    .Y(_01_));
 sky130_fd_sc_hd__xnor2_1 _11_ (.A(\branch_addr_match_buf_I[3].z ),
    .B(addr[3]),
    .Y(_02_));
 sky130_fd_sc_hd__xnor2_1 _12_ (.A(\branch_addr_match_buf_I[2].z ),
    .B(addr[2]),
    .Y(_03_));
 sky130_fd_sc_hd__o2bb2ai_1 _13_ (.A1_N(_01_),
    .A2_N(addr[1]),
    .B1(_00_),
    .B2(addr[0]),
    .Y(_04_));
 sky130_fd_sc_hd__o2111ai_1 _14_ (.A1(_01_),
    .A2(addr[1]),
    .B1(\branch_ena_buf_I.z ),
    .C1(_02_),
    .D1(_03_),
    .Y(_05_));
 sky130_fd_sc_hd__a211oi_1 _15_ (.A1(_00_),
    .A2(addr[0]),
    .B1(_04_),
    .C1(_05_),
    .Y(\branch_sel_buf_I.a ));
 sky130_fd_sc_hd__nor4b_1 _16_ (.A(\zbuf_bus_sel_I[2].z ),
    .B(\zbuf_bus_sel_I[3].z ),
    .C(\zbuf_bus_sel_I[4].z ),
    .D_N(\buf_bus_ena_I.z ),
    .Y(\block[0].genblk1.grp_sel_buf_I.a ));
 sky130_fd_sc_hd__nor2_1 _17_ (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .B(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .Y(_06_));
 sky130_fd_sc_hd__and2_1 _18_ (.A(\block[0].genblk1.grp_sel_buf_I.z ),
    .B(_06_),
    .X(\block[0].l_ena_0_I.a ));
 sky130_fd_sc_hd__nor2b_1 _19_ (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .B_N(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .Y(_07_));
 sky130_fd_sc_hd__and2_1 _20_ (.A(\block[0].genblk1.grp_sel_buf_I.z ),
    .B(_07_),
    .X(\block[1].l_ena_0_I.a ));
 sky130_fd_sc_hd__nor2b_1 _21_ (.A(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .B_N(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .Y(_08_));
 sky130_fd_sc_hd__and2_1 _22_ (.A(\block[0].genblk1.grp_sel_buf_I.z ),
    .B(_08_),
    .X(\block[2].l_ena_0_I.a ));
 sky130_fd_sc_hd__and3_1 _23_ (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .B(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .C(\block[0].genblk1.grp_sel_buf_I.z ),
    .X(\block[3].l_ena_0_I.a ));
 sky130_fd_sc_hd__nor4bb_1 _24_ (.A(\zbuf_bus_sel_I[3].z ),
    .B(\zbuf_bus_sel_I[4].z ),
    .C_N(\buf_bus_ena_I.z ),
    .D_N(\zbuf_bus_sel_I[2].z ),
    .Y(\block[4].genblk1.grp_sel_buf_I.a ));
 sky130_fd_sc_hd__and2_1 _25_ (.A(\block[4].genblk1.grp_sel_buf_I.z ),
    .B(_06_),
    .X(\block[4].l_ena_0_I.a ));
 sky130_fd_sc_hd__and2_1 _26_ (.A(\block[4].genblk1.grp_sel_buf_I.z ),
    .B(_07_),
    .X(\block[5].l_ena_0_I.a ));
 sky130_fd_sc_hd__and2_1 _27_ (.A(\block[4].genblk1.grp_sel_buf_I.z ),
    .B(_08_),
    .X(\block[6].l_ena_0_I.a ));
 sky130_fd_sc_hd__and3_1 _28_ (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .B(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .C(\block[4].genblk1.grp_sel_buf_I.z ),
    .X(\block[7].l_ena_0_I.a ));
 sky130_fd_sc_hd__nor4bb_1 _29_ (.A(\zbuf_bus_sel_I[2].z ),
    .B(\zbuf_bus_sel_I[4].z ),
    .C_N(\buf_bus_ena_I.z ),
    .D_N(\zbuf_bus_sel_I[3].z ),
    .Y(\block[8].genblk1.grp_sel_buf_I.a ));
 sky130_fd_sc_hd__and2_1 _30_ (.A(\block[8].genblk1.grp_sel_buf_I.z ),
    .B(_06_),
    .X(\block[8].l_ena_0_I.a ));
 sky130_fd_sc_hd__and2_1 _31_ (.A(\block[8].genblk1.grp_sel_buf_I.z ),
    .B(_07_),
    .X(\block[9].l_ena_0_I.a ));
 sky130_fd_sc_hd__and2_1 _32_ (.A(\block[8].genblk1.grp_sel_buf_I.z ),
    .B(_08_),
    .X(\block[10].l_ena_0_I.a ));
 sky130_fd_sc_hd__and3_1 _33_ (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .B(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .C(\block[8].genblk1.grp_sel_buf_I.z ),
    .X(\block[11].l_ena_0_I.a ));
 sky130_fd_sc_hd__and4b_1 _34_ (.A_N(\zbuf_bus_sel_I[4].z ),
    .B(\buf_bus_ena_I.z ),
    .C(\zbuf_bus_sel_I[2].z ),
    .D(\zbuf_bus_sel_I[3].z ),
    .X(\block[12].genblk1.grp_sel_buf_I.a ));
 sky130_fd_sc_hd__and2_1 _35_ (.A(\block[12].genblk1.grp_sel_buf_I.z ),
    .B(_06_),
    .X(\block[12].l_ena_0_I.a ));
 sky130_fd_sc_hd__and2_1 _36_ (.A(\block[12].genblk1.grp_sel_buf_I.z ),
    .B(_07_),
    .X(\block[13].l_ena_0_I.a ));
 sky130_fd_sc_hd__and2_1 _37_ (.A(\block[12].genblk1.grp_sel_buf_I.z ),
    .B(_08_),
    .X(\block[14].l_ena_0_I.a ));
 sky130_fd_sc_hd__and3_1 _38_ (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .B(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .C(\block[12].genblk1.grp_sel_buf_I.z ),
    .X(\block[15].l_ena_0_I.a ));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[0].cell0_I  (.DIODE(um_ow[0]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[10].cell0_I  (.DIODE(um_ow[10]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[11].cell0_I  (.DIODE(um_ow[11]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[12].cell0_I  (.DIODE(um_ow[12]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[13].cell0_I  (.DIODE(um_ow[13]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[14].cell0_I  (.DIODE(um_ow[14]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[15].cell0_I  (.DIODE(um_ow[15]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[16].cell0_I  (.DIODE(um_ow[16]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[17].cell0_I  (.DIODE(um_ow[17]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[18].cell0_I  (.DIODE(um_ow[18]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[19].cell0_I  (.DIODE(um_ow[19]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[1].cell0_I  (.DIODE(um_ow[1]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[20].cell0_I  (.DIODE(um_ow[20]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[21].cell0_I  (.DIODE(um_ow[21]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[22].cell0_I  (.DIODE(um_ow[22]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[23].cell0_I  (.DIODE(um_ow[23]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[2].cell0_I  (.DIODE(um_ow[2]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[3].cell0_I  (.DIODE(um_ow[3]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[4].cell0_I  (.DIODE(um_ow[4]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[5].cell0_I  (.DIODE(um_ow[5]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[6].cell0_I  (.DIODE(um_ow[6]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[7].cell0_I  (.DIODE(um_ow[7]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[8].cell0_I  (.DIODE(um_ow[8]));
 sky130_fd_sc_hd__diode_2 \block[0].diode_I[9].cell0_I  (.DIODE(um_ow[9]));
 sky130_fd_sc_hd__buf_2 \block[0].genblk1.grp_sel_buf_I.genblk1.cell0_I  (.A(\block[0].genblk1.grp_sel_buf_I.a ),
    .X(\block[0].genblk1.grp_sel_buf_I.z ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[0].cell0_I  (.A0(um_ow[0]),
    .A1(um_ow[24]),
    .A2(um_ow[48]),
    .A3(um_ow[72]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[10].cell0_I  (.A0(um_ow[10]),
    .A1(um_ow[34]),
    .A2(um_ow[58]),
    .A3(um_ow[82]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[11].cell0_I  (.A0(um_ow[11]),
    .A1(um_ow[35]),
    .A2(um_ow[59]),
    .A3(um_ow[83]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[12].cell0_I  (.A0(um_ow[12]),
    .A1(um_ow[36]),
    .A2(um_ow[60]),
    .A3(um_ow[84]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[13].cell0_I  (.A0(um_ow[13]),
    .A1(um_ow[37]),
    .A2(um_ow[61]),
    .A3(um_ow[85]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[14].cell0_I  (.A0(um_ow[14]),
    .A1(um_ow[38]),
    .A2(um_ow[62]),
    .A3(um_ow[86]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[15].cell0_I  (.A0(um_ow[15]),
    .A1(um_ow[39]),
    .A2(um_ow[63]),
    .A3(um_ow[87]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[16].cell0_I  (.A0(um_ow[16]),
    .A1(um_ow[40]),
    .A2(um_ow[64]),
    .A3(um_ow[88]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[17].cell0_I  (.A0(um_ow[17]),
    .A1(um_ow[41]),
    .A2(um_ow[65]),
    .A3(um_ow[89]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[18].cell0_I  (.A0(um_ow[18]),
    .A1(um_ow[42]),
    .A2(um_ow[66]),
    .A3(um_ow[90]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[19].cell0_I  (.A0(um_ow[19]),
    .A1(um_ow[43]),
    .A2(um_ow[67]),
    .A3(um_ow[91]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[1].cell0_I  (.A0(um_ow[1]),
    .A1(um_ow[25]),
    .A2(um_ow[49]),
    .A3(um_ow[73]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[20].cell0_I  (.A0(um_ow[20]),
    .A1(um_ow[44]),
    .A2(um_ow[68]),
    .A3(um_ow[92]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[21].cell0_I  (.A0(um_ow[21]),
    .A1(um_ow[45]),
    .A2(um_ow[69]),
    .A3(um_ow[93]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[22].cell0_I  (.A0(um_ow[22]),
    .A1(um_ow[46]),
    .A2(um_ow[70]),
    .A3(um_ow[94]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[23].cell0_I  (.A0(um_ow[23]),
    .A1(um_ow[47]),
    .A2(um_ow[71]),
    .A3(um_ow[95]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[2].cell0_I  (.A0(um_ow[2]),
    .A1(um_ow[26]),
    .A2(um_ow[50]),
    .A3(um_ow[74]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[3].cell0_I  (.A0(um_ow[3]),
    .A1(um_ow[27]),
    .A2(um_ow[51]),
    .A3(um_ow[75]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[4].cell0_I  (.A0(um_ow[4]),
    .A1(um_ow[28]),
    .A2(um_ow[52]),
    .A3(um_ow[76]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[5].cell0_I  (.A0(um_ow[5]),
    .A1(um_ow[29]),
    .A2(um_ow[53]),
    .A3(um_ow[77]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[6].cell0_I  (.A0(um_ow[6]),
    .A1(um_ow[30]),
    .A2(um_ow[54]),
    .A3(um_ow[78]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[7].cell0_I  (.A0(um_ow[7]),
    .A1(um_ow[31]),
    .A2(um_ow[55]),
    .A3(um_ow[79]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[8].cell0_I  (.A0(um_ow[8]),
    .A1(um_ow[32]),
    .A2(um_ow[56]),
    .A3(um_ow[80]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_2 \block[0].genblk1.mux4_I[9].cell0_I  (.A0(um_ow[9]),
    .A1(um_ow[33]),
    .A2(um_ow[57]),
    .A3(um_ow[81]),
    .S0(\block[0].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[0].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[0].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__buf_2 \block[0].genblk1.mux4_sel_buf_I[0].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .X(\block[0].genblk1.mux4_sel_buf_I[0].z ));
 sky130_fd_sc_hd__buf_2 \block[0].genblk1.mux4_sel_buf_I[1].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .X(\block[0].genblk1.mux4_sel_buf_I[1].z ));
 sky130_fd_sc_hd__bufinv_8 \block[0].genblk1.tbuf_blk_ena_I.cell0_I  (.A(\block[0].genblk1.grp_sel_buf_I.z ),
    .Y(\block[0].genblk1.tbuf_blk_ena_I.tx ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[0].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[0].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[10].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[10].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[11].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[11].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[12].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[12].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[13].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[13].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[14].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[14].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[15].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[15].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[16].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[16].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[17].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[17].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[18].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[18].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[19].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[19].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[1].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[1].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[20].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[20].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[21].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[21].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[22].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[22].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[23].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[23].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[2].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[2].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[3].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[3].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[4].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[4].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[5].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[5].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[6].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[6].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[7].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[7].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[8].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[8].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__ebufn_8 \block[0].genblk1.tbuf_spine_ow_I[9].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_I[9].x ),
    .TE_B(\block[0].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__buf_8 \block[0].l_ena_0_I.genblk1.cell0_I  (.A(\block[0].l_ena_0_I.a ),
    .X(\block[0].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[0].tie_I.cell_I  (.HI(\block[0].tie_I.hi ),
    .LO(\block[0].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[0].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[0].l_ena_0_I.z ),
    .X(\block[0].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[0].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[0].l_ena_0_I.z ),
    .Y(\block[0].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[0].cell0_I  (.DIODE(um_ow[240]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[10].cell0_I  (.DIODE(um_ow[250]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[11].cell0_I  (.DIODE(um_ow[251]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[12].cell0_I  (.DIODE(um_ow[252]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[13].cell0_I  (.DIODE(um_ow[253]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[14].cell0_I  (.DIODE(um_ow[254]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[15].cell0_I  (.DIODE(um_ow[255]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[16].cell0_I  (.DIODE(um_ow[256]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[17].cell0_I  (.DIODE(um_ow[257]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[18].cell0_I  (.DIODE(um_ow[258]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[19].cell0_I  (.DIODE(um_ow[259]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[1].cell0_I  (.DIODE(um_ow[241]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[20].cell0_I  (.DIODE(um_ow[260]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[21].cell0_I  (.DIODE(um_ow[261]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[22].cell0_I  (.DIODE(um_ow[262]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[23].cell0_I  (.DIODE(um_ow[263]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[2].cell0_I  (.DIODE(um_ow[242]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[3].cell0_I  (.DIODE(um_ow[243]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[4].cell0_I  (.DIODE(um_ow[244]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[5].cell0_I  (.DIODE(um_ow[245]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[6].cell0_I  (.DIODE(um_ow[246]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[7].cell0_I  (.DIODE(um_ow[247]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[8].cell0_I  (.DIODE(um_ow[248]));
 sky130_fd_sc_hd__diode_2 \block[10].diode_I[9].cell0_I  (.DIODE(um_ow[249]));
 sky130_fd_sc_hd__buf_8 \block[10].l_ena_0_I.genblk1.cell0_I  (.A(\block[10].l_ena_0_I.a ),
    .X(\block[10].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[10].tie_I.cell_I  (.HI(\block[10].tie_I.hi ),
    .LO(\block[10].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[10].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[10].l_ena_0_I.z ),
    .X(\block[10].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[10].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[10].l_ena_0_I.z ),
    .Y(\block[10].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[0].cell0_I  (.DIODE(um_ow[264]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[10].cell0_I  (.DIODE(um_ow[274]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[11].cell0_I  (.DIODE(um_ow[275]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[12].cell0_I  (.DIODE(um_ow[276]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[13].cell0_I  (.DIODE(um_ow[277]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[14].cell0_I  (.DIODE(um_ow[278]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[15].cell0_I  (.DIODE(um_ow[279]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[16].cell0_I  (.DIODE(um_ow[280]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[17].cell0_I  (.DIODE(um_ow[281]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[18].cell0_I  (.DIODE(um_ow[282]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[19].cell0_I  (.DIODE(um_ow[283]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[1].cell0_I  (.DIODE(um_ow[265]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[20].cell0_I  (.DIODE(um_ow[284]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[21].cell0_I  (.DIODE(um_ow[285]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[22].cell0_I  (.DIODE(um_ow[286]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[23].cell0_I  (.DIODE(um_ow[287]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[2].cell0_I  (.DIODE(um_ow[266]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[3].cell0_I  (.DIODE(um_ow[267]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[4].cell0_I  (.DIODE(um_ow[268]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[5].cell0_I  (.DIODE(um_ow[269]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[6].cell0_I  (.DIODE(um_ow[270]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[7].cell0_I  (.DIODE(um_ow[271]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[8].cell0_I  (.DIODE(um_ow[272]));
 sky130_fd_sc_hd__diode_2 \block[11].diode_I[9].cell0_I  (.DIODE(um_ow[273]));
 sky130_fd_sc_hd__buf_8 \block[11].l_ena_0_I.genblk1.cell0_I  (.A(\block[11].l_ena_0_I.a ),
    .X(\block[11].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[11].tie_I.cell_I  (.HI(\block[11].tie_I.hi ),
    .LO(\block[11].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[11].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[11].l_ena_0_I.z ),
    .X(\block[11].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[11].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[11].l_ena_0_I.z ),
    .Y(\block[11].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[0].cell0_I  (.DIODE(um_ow[288]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[10].cell0_I  (.DIODE(um_ow[298]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[11].cell0_I  (.DIODE(um_ow[299]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[12].cell0_I  (.DIODE(um_ow[300]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[13].cell0_I  (.DIODE(um_ow[301]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[14].cell0_I  (.DIODE(um_ow[302]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[15].cell0_I  (.DIODE(um_ow[303]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[16].cell0_I  (.DIODE(um_ow[304]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[17].cell0_I  (.DIODE(um_ow[305]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[18].cell0_I  (.DIODE(um_ow[306]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[19].cell0_I  (.DIODE(um_ow[307]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[1].cell0_I  (.DIODE(um_ow[289]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[20].cell0_I  (.DIODE(um_ow[308]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[21].cell0_I  (.DIODE(um_ow[309]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[22].cell0_I  (.DIODE(um_ow[310]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[23].cell0_I  (.DIODE(um_ow[311]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[2].cell0_I  (.DIODE(um_ow[290]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[3].cell0_I  (.DIODE(um_ow[291]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[4].cell0_I  (.DIODE(um_ow[292]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[5].cell0_I  (.DIODE(um_ow[293]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[6].cell0_I  (.DIODE(um_ow[294]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[7].cell0_I  (.DIODE(um_ow[295]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[8].cell0_I  (.DIODE(um_ow[296]));
 sky130_fd_sc_hd__diode_2 \block[12].diode_I[9].cell0_I  (.DIODE(um_ow[297]));
 sky130_fd_sc_hd__buf_2 \block[12].genblk1.grp_sel_buf_I.genblk1.cell0_I  (.A(\block[12].genblk1.grp_sel_buf_I.a ),
    .X(\block[12].genblk1.grp_sel_buf_I.z ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[0].cell0_I  (.A0(um_ow[288]),
    .A1(um_ow[312]),
    .A2(um_ow[336]),
    .A3(um_ow[360]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[10].cell0_I  (.A0(um_ow[298]),
    .A1(um_ow[322]),
    .A2(um_ow[346]),
    .A3(um_ow[370]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[11].cell0_I  (.A0(um_ow[299]),
    .A1(um_ow[323]),
    .A2(um_ow[347]),
    .A3(um_ow[371]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[12].cell0_I  (.A0(um_ow[300]),
    .A1(um_ow[324]),
    .A2(um_ow[348]),
    .A3(um_ow[372]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[13].cell0_I  (.A0(um_ow[301]),
    .A1(um_ow[325]),
    .A2(um_ow[349]),
    .A3(um_ow[373]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[14].cell0_I  (.A0(um_ow[302]),
    .A1(um_ow[326]),
    .A2(um_ow[350]),
    .A3(um_ow[374]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[15].cell0_I  (.A0(um_ow[303]),
    .A1(um_ow[327]),
    .A2(um_ow[351]),
    .A3(um_ow[375]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[16].cell0_I  (.A0(um_ow[304]),
    .A1(um_ow[328]),
    .A2(um_ow[352]),
    .A3(um_ow[376]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[17].cell0_I  (.A0(um_ow[305]),
    .A1(um_ow[329]),
    .A2(um_ow[353]),
    .A3(um_ow[377]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[18].cell0_I  (.A0(um_ow[306]),
    .A1(um_ow[330]),
    .A2(um_ow[354]),
    .A3(um_ow[378]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[19].cell0_I  (.A0(um_ow[307]),
    .A1(um_ow[331]),
    .A2(um_ow[355]),
    .A3(um_ow[379]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[1].cell0_I  (.A0(um_ow[289]),
    .A1(um_ow[313]),
    .A2(um_ow[337]),
    .A3(um_ow[361]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[20].cell0_I  (.A0(um_ow[308]),
    .A1(um_ow[332]),
    .A2(um_ow[356]),
    .A3(um_ow[380]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[21].cell0_I  (.A0(um_ow[309]),
    .A1(um_ow[333]),
    .A2(um_ow[357]),
    .A3(um_ow[381]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[22].cell0_I  (.A0(um_ow[310]),
    .A1(um_ow[334]),
    .A2(um_ow[358]),
    .A3(um_ow[382]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[23].cell0_I  (.A0(um_ow[311]),
    .A1(um_ow[335]),
    .A2(um_ow[359]),
    .A3(um_ow[383]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[2].cell0_I  (.A0(um_ow[290]),
    .A1(um_ow[314]),
    .A2(um_ow[338]),
    .A3(um_ow[362]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[3].cell0_I  (.A0(um_ow[291]),
    .A1(um_ow[315]),
    .A2(um_ow[339]),
    .A3(um_ow[363]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[4].cell0_I  (.A0(um_ow[292]),
    .A1(um_ow[316]),
    .A2(um_ow[340]),
    .A3(um_ow[364]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[5].cell0_I  (.A0(um_ow[293]),
    .A1(um_ow[317]),
    .A2(um_ow[341]),
    .A3(um_ow[365]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[6].cell0_I  (.A0(um_ow[294]),
    .A1(um_ow[318]),
    .A2(um_ow[342]),
    .A3(um_ow[366]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[7].cell0_I  (.A0(um_ow[295]),
    .A1(um_ow[319]),
    .A2(um_ow[343]),
    .A3(um_ow[367]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[8].cell0_I  (.A0(um_ow[296]),
    .A1(um_ow[320]),
    .A2(um_ow[344]),
    .A3(um_ow[368]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_2 \block[12].genblk1.mux4_I[9].cell0_I  (.A0(um_ow[297]),
    .A1(um_ow[321]),
    .A2(um_ow[345]),
    .A3(um_ow[369]),
    .S0(\block[12].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[12].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[12].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__buf_2 \block[12].genblk1.mux4_sel_buf_I[0].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .X(\block[12].genblk1.mux4_sel_buf_I[0].z ));
 sky130_fd_sc_hd__buf_2 \block[12].genblk1.mux4_sel_buf_I[1].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .X(\block[12].genblk1.mux4_sel_buf_I[1].z ));
 sky130_fd_sc_hd__bufinv_8 \block[12].genblk1.tbuf_blk_ena_I.cell0_I  (.A(\block[12].genblk1.grp_sel_buf_I.z ),
    .Y(\block[12].genblk1.tbuf_blk_ena_I.tx ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[0].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[0].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[10].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[10].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[11].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[11].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[12].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[12].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[13].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[13].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[14].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[14].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[15].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[15].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[16].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[16].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[17].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[17].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[18].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[18].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[19].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[19].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[1].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[1].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[20].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[20].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[21].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[21].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[22].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[22].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[23].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[23].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[2].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[2].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[3].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[3].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[4].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[4].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[5].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[5].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[6].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[6].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[7].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[7].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[8].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[8].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__ebufn_8 \block[12].genblk1.tbuf_spine_ow_I[9].genblk1.cell0_I  (.A(\block[12].genblk1.mux4_I[9].x ),
    .TE_B(\block[12].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__buf_8 \block[12].l_ena_0_I.genblk1.cell0_I  (.A(\block[12].l_ena_0_I.a ),
    .X(\block[12].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[12].tie_I.cell_I  (.HI(\block[12].tie_I.hi ),
    .LO(\block[12].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[12].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[12].l_ena_0_I.z ),
    .X(\block[12].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[12].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[12].l_ena_0_I.z ),
    .Y(\block[12].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[0].cell0_I  (.DIODE(um_ow[312]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[10].cell0_I  (.DIODE(um_ow[322]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[11].cell0_I  (.DIODE(um_ow[323]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[12].cell0_I  (.DIODE(um_ow[324]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[13].cell0_I  (.DIODE(um_ow[325]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[14].cell0_I  (.DIODE(um_ow[326]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[15].cell0_I  (.DIODE(um_ow[327]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[16].cell0_I  (.DIODE(um_ow[328]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[17].cell0_I  (.DIODE(um_ow[329]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[18].cell0_I  (.DIODE(um_ow[330]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[19].cell0_I  (.DIODE(um_ow[331]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[1].cell0_I  (.DIODE(um_ow[313]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[20].cell0_I  (.DIODE(um_ow[332]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[21].cell0_I  (.DIODE(um_ow[333]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[22].cell0_I  (.DIODE(um_ow[334]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[23].cell0_I  (.DIODE(um_ow[335]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[2].cell0_I  (.DIODE(um_ow[314]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[3].cell0_I  (.DIODE(um_ow[315]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[4].cell0_I  (.DIODE(um_ow[316]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[5].cell0_I  (.DIODE(um_ow[317]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[6].cell0_I  (.DIODE(um_ow[318]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[7].cell0_I  (.DIODE(um_ow[319]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[8].cell0_I  (.DIODE(um_ow[320]));
 sky130_fd_sc_hd__diode_2 \block[13].diode_I[9].cell0_I  (.DIODE(um_ow[321]));
 sky130_fd_sc_hd__buf_8 \block[13].l_ena_0_I.genblk1.cell0_I  (.A(\block[13].l_ena_0_I.a ),
    .X(\block[13].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[13].tie_I.cell_I  (.HI(\block[13].tie_I.hi ),
    .LO(\block[13].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[13].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[13].l_ena_0_I.z ),
    .X(\block[13].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[13].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[13].l_ena_0_I.z ),
    .Y(\block[13].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[0].cell0_I  (.DIODE(um_ow[336]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[10].cell0_I  (.DIODE(um_ow[346]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[11].cell0_I  (.DIODE(um_ow[347]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[12].cell0_I  (.DIODE(um_ow[348]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[13].cell0_I  (.DIODE(um_ow[349]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[14].cell0_I  (.DIODE(um_ow[350]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[15].cell0_I  (.DIODE(um_ow[351]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[16].cell0_I  (.DIODE(um_ow[352]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[17].cell0_I  (.DIODE(um_ow[353]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[18].cell0_I  (.DIODE(um_ow[354]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[19].cell0_I  (.DIODE(um_ow[355]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[1].cell0_I  (.DIODE(um_ow[337]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[20].cell0_I  (.DIODE(um_ow[356]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[21].cell0_I  (.DIODE(um_ow[357]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[22].cell0_I  (.DIODE(um_ow[358]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[23].cell0_I  (.DIODE(um_ow[359]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[2].cell0_I  (.DIODE(um_ow[338]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[3].cell0_I  (.DIODE(um_ow[339]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[4].cell0_I  (.DIODE(um_ow[340]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[5].cell0_I  (.DIODE(um_ow[341]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[6].cell0_I  (.DIODE(um_ow[342]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[7].cell0_I  (.DIODE(um_ow[343]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[8].cell0_I  (.DIODE(um_ow[344]));
 sky130_fd_sc_hd__diode_2 \block[14].diode_I[9].cell0_I  (.DIODE(um_ow[345]));
 sky130_fd_sc_hd__buf_8 \block[14].l_ena_0_I.genblk1.cell0_I  (.A(\block[14].l_ena_0_I.a ),
    .X(\block[14].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[14].tie_I.cell_I  (.HI(\block[14].tie_I.hi ),
    .LO(\block[14].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[14].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[14].l_ena_0_I.z ),
    .X(\block[14].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[14].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[14].l_ena_0_I.z ),
    .Y(\block[14].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[0].cell0_I  (.DIODE(um_ow[360]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[10].cell0_I  (.DIODE(um_ow[370]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[11].cell0_I  (.DIODE(um_ow[371]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[12].cell0_I  (.DIODE(um_ow[372]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[13].cell0_I  (.DIODE(um_ow[373]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[14].cell0_I  (.DIODE(um_ow[374]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[15].cell0_I  (.DIODE(um_ow[375]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[16].cell0_I  (.DIODE(um_ow[376]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[17].cell0_I  (.DIODE(um_ow[377]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[18].cell0_I  (.DIODE(um_ow[378]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[19].cell0_I  (.DIODE(um_ow[379]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[1].cell0_I  (.DIODE(um_ow[361]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[20].cell0_I  (.DIODE(um_ow[380]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[21].cell0_I  (.DIODE(um_ow[381]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[22].cell0_I  (.DIODE(um_ow[382]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[23].cell0_I  (.DIODE(um_ow[383]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[2].cell0_I  (.DIODE(um_ow[362]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[3].cell0_I  (.DIODE(um_ow[363]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[4].cell0_I  (.DIODE(um_ow[364]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[5].cell0_I  (.DIODE(um_ow[365]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[6].cell0_I  (.DIODE(um_ow[366]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[7].cell0_I  (.DIODE(um_ow[367]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[8].cell0_I  (.DIODE(um_ow[368]));
 sky130_fd_sc_hd__diode_2 \block[15].diode_I[9].cell0_I  (.DIODE(um_ow[369]));
 sky130_fd_sc_hd__buf_8 \block[15].l_ena_0_I.genblk1.cell0_I  (.A(\block[15].l_ena_0_I.a ),
    .X(\block[15].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[15].tie_I.cell_I  (.HI(\block[15].tie_I.hi ),
    .LO(\block[15].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[15].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[15].l_ena_0_I.z ),
    .X(\block[15].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[15].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[15].l_ena_0_I.z ),
    .Y(\block[15].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[0].cell0_I  (.DIODE(um_ow[24]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[10].cell0_I  (.DIODE(um_ow[34]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[11].cell0_I  (.DIODE(um_ow[35]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[12].cell0_I  (.DIODE(um_ow[36]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[13].cell0_I  (.DIODE(um_ow[37]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[14].cell0_I  (.DIODE(um_ow[38]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[15].cell0_I  (.DIODE(um_ow[39]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[16].cell0_I  (.DIODE(um_ow[40]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[17].cell0_I  (.DIODE(um_ow[41]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[18].cell0_I  (.DIODE(um_ow[42]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[19].cell0_I  (.DIODE(um_ow[43]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[1].cell0_I  (.DIODE(um_ow[25]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[20].cell0_I  (.DIODE(um_ow[44]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[21].cell0_I  (.DIODE(um_ow[45]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[22].cell0_I  (.DIODE(um_ow[46]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[23].cell0_I  (.DIODE(um_ow[47]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[2].cell0_I  (.DIODE(um_ow[26]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[3].cell0_I  (.DIODE(um_ow[27]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[4].cell0_I  (.DIODE(um_ow[28]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[5].cell0_I  (.DIODE(um_ow[29]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[6].cell0_I  (.DIODE(um_ow[30]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[7].cell0_I  (.DIODE(um_ow[31]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[8].cell0_I  (.DIODE(um_ow[32]));
 sky130_fd_sc_hd__diode_2 \block[1].diode_I[9].cell0_I  (.DIODE(um_ow[33]));
 sky130_fd_sc_hd__buf_8 \block[1].l_ena_0_I.genblk1.cell0_I  (.A(\block[1].l_ena_0_I.a ),
    .X(\block[1].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[1].tie_I.cell_I  (.HI(\block[1].tie_I.hi ),
    .LO(\block[1].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[1].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[1].l_ena_0_I.z ),
    .X(\block[1].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[1].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[1].l_ena_0_I.z ),
    .Y(\block[1].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[0].cell0_I  (.DIODE(um_ow[48]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[10].cell0_I  (.DIODE(um_ow[58]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[11].cell0_I  (.DIODE(um_ow[59]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[12].cell0_I  (.DIODE(um_ow[60]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[13].cell0_I  (.DIODE(um_ow[61]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[14].cell0_I  (.DIODE(um_ow[62]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[15].cell0_I  (.DIODE(um_ow[63]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[16].cell0_I  (.DIODE(um_ow[64]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[17].cell0_I  (.DIODE(um_ow[65]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[18].cell0_I  (.DIODE(um_ow[66]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[19].cell0_I  (.DIODE(um_ow[67]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[1].cell0_I  (.DIODE(um_ow[49]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[20].cell0_I  (.DIODE(um_ow[68]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[21].cell0_I  (.DIODE(um_ow[69]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[22].cell0_I  (.DIODE(um_ow[70]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[23].cell0_I  (.DIODE(um_ow[71]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[2].cell0_I  (.DIODE(um_ow[50]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[3].cell0_I  (.DIODE(um_ow[51]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[4].cell0_I  (.DIODE(um_ow[52]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[5].cell0_I  (.DIODE(um_ow[53]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[6].cell0_I  (.DIODE(um_ow[54]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[7].cell0_I  (.DIODE(um_ow[55]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[8].cell0_I  (.DIODE(um_ow[56]));
 sky130_fd_sc_hd__diode_2 \block[2].diode_I[9].cell0_I  (.DIODE(um_ow[57]));
 sky130_fd_sc_hd__buf_8 \block[2].l_ena_0_I.genblk1.cell0_I  (.A(\block[2].l_ena_0_I.a ),
    .X(\block[2].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[2].tie_I.cell_I  (.HI(\block[2].tie_I.hi ),
    .LO(\block[2].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[2].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[2].l_ena_0_I.z ),
    .X(\block[2].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[2].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[2].l_ena_0_I.z ),
    .Y(\block[2].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[0].cell0_I  (.DIODE(um_ow[72]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[10].cell0_I  (.DIODE(um_ow[82]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[11].cell0_I  (.DIODE(um_ow[83]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[12].cell0_I  (.DIODE(um_ow[84]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[13].cell0_I  (.DIODE(um_ow[85]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[14].cell0_I  (.DIODE(um_ow[86]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[15].cell0_I  (.DIODE(um_ow[87]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[16].cell0_I  (.DIODE(um_ow[88]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[17].cell0_I  (.DIODE(um_ow[89]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[18].cell0_I  (.DIODE(um_ow[90]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[19].cell0_I  (.DIODE(um_ow[91]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[1].cell0_I  (.DIODE(um_ow[73]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[20].cell0_I  (.DIODE(um_ow[92]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[21].cell0_I  (.DIODE(um_ow[93]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[22].cell0_I  (.DIODE(um_ow[94]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[23].cell0_I  (.DIODE(um_ow[95]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[2].cell0_I  (.DIODE(um_ow[74]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[3].cell0_I  (.DIODE(um_ow[75]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[4].cell0_I  (.DIODE(um_ow[76]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[5].cell0_I  (.DIODE(um_ow[77]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[6].cell0_I  (.DIODE(um_ow[78]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[7].cell0_I  (.DIODE(um_ow[79]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[8].cell0_I  (.DIODE(um_ow[80]));
 sky130_fd_sc_hd__diode_2 \block[3].diode_I[9].cell0_I  (.DIODE(um_ow[81]));
 sky130_fd_sc_hd__buf_8 \block[3].l_ena_0_I.genblk1.cell0_I  (.A(\block[3].l_ena_0_I.a ),
    .X(\block[3].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[3].tie_I.cell_I  (.HI(\block[3].tie_I.hi ),
    .LO(\block[3].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[3].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[3].l_ena_0_I.z ),
    .X(\block[3].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[3].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[3].l_ena_0_I.z ),
    .Y(\block[3].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[0].cell0_I  (.DIODE(um_ow[96]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[10].cell0_I  (.DIODE(um_ow[106]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[11].cell0_I  (.DIODE(um_ow[107]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[12].cell0_I  (.DIODE(um_ow[108]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[13].cell0_I  (.DIODE(um_ow[109]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[14].cell0_I  (.DIODE(um_ow[110]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[15].cell0_I  (.DIODE(um_ow[111]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[16].cell0_I  (.DIODE(um_ow[112]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[17].cell0_I  (.DIODE(um_ow[113]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[18].cell0_I  (.DIODE(um_ow[114]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[19].cell0_I  (.DIODE(um_ow[115]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[1].cell0_I  (.DIODE(um_ow[97]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[20].cell0_I  (.DIODE(um_ow[116]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[21].cell0_I  (.DIODE(um_ow[117]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[22].cell0_I  (.DIODE(um_ow[118]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[23].cell0_I  (.DIODE(um_ow[119]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[2].cell0_I  (.DIODE(um_ow[98]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[3].cell0_I  (.DIODE(um_ow[99]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[4].cell0_I  (.DIODE(um_ow[100]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[5].cell0_I  (.DIODE(um_ow[101]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[6].cell0_I  (.DIODE(um_ow[102]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[7].cell0_I  (.DIODE(um_ow[103]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[8].cell0_I  (.DIODE(um_ow[104]));
 sky130_fd_sc_hd__diode_2 \block[4].diode_I[9].cell0_I  (.DIODE(um_ow[105]));
 sky130_fd_sc_hd__buf_2 \block[4].genblk1.grp_sel_buf_I.genblk1.cell0_I  (.A(\block[4].genblk1.grp_sel_buf_I.a ),
    .X(\block[4].genblk1.grp_sel_buf_I.z ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[0].cell0_I  (.A0(um_ow[96]),
    .A1(um_ow[120]),
    .A2(um_ow[144]),
    .A3(um_ow[168]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[10].cell0_I  (.A0(um_ow[106]),
    .A1(um_ow[130]),
    .A2(um_ow[154]),
    .A3(um_ow[178]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[11].cell0_I  (.A0(um_ow[107]),
    .A1(um_ow[131]),
    .A2(um_ow[155]),
    .A3(um_ow[179]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[12].cell0_I  (.A0(um_ow[108]),
    .A1(um_ow[132]),
    .A2(um_ow[156]),
    .A3(um_ow[180]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[13].cell0_I  (.A0(um_ow[109]),
    .A1(um_ow[133]),
    .A2(um_ow[157]),
    .A3(um_ow[181]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[14].cell0_I  (.A0(um_ow[110]),
    .A1(um_ow[134]),
    .A2(um_ow[158]),
    .A3(um_ow[182]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[15].cell0_I  (.A0(um_ow[111]),
    .A1(um_ow[135]),
    .A2(um_ow[159]),
    .A3(um_ow[183]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[16].cell0_I  (.A0(um_ow[112]),
    .A1(um_ow[136]),
    .A2(um_ow[160]),
    .A3(um_ow[184]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[17].cell0_I  (.A0(um_ow[113]),
    .A1(um_ow[137]),
    .A2(um_ow[161]),
    .A3(um_ow[185]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[18].cell0_I  (.A0(um_ow[114]),
    .A1(um_ow[138]),
    .A2(um_ow[162]),
    .A3(um_ow[186]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[19].cell0_I  (.A0(um_ow[115]),
    .A1(um_ow[139]),
    .A2(um_ow[163]),
    .A3(um_ow[187]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[1].cell0_I  (.A0(um_ow[97]),
    .A1(um_ow[121]),
    .A2(um_ow[145]),
    .A3(um_ow[169]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[20].cell0_I  (.A0(um_ow[116]),
    .A1(um_ow[140]),
    .A2(um_ow[164]),
    .A3(um_ow[188]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[21].cell0_I  (.A0(um_ow[117]),
    .A1(um_ow[141]),
    .A2(um_ow[165]),
    .A3(um_ow[189]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[22].cell0_I  (.A0(um_ow[118]),
    .A1(um_ow[142]),
    .A2(um_ow[166]),
    .A3(um_ow[190]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[23].cell0_I  (.A0(um_ow[119]),
    .A1(um_ow[143]),
    .A2(um_ow[167]),
    .A3(um_ow[191]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[2].cell0_I  (.A0(um_ow[98]),
    .A1(um_ow[122]),
    .A2(um_ow[146]),
    .A3(um_ow[170]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[3].cell0_I  (.A0(um_ow[99]),
    .A1(um_ow[123]),
    .A2(um_ow[147]),
    .A3(um_ow[171]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[4].cell0_I  (.A0(um_ow[100]),
    .A1(um_ow[124]),
    .A2(um_ow[148]),
    .A3(um_ow[172]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[5].cell0_I  (.A0(um_ow[101]),
    .A1(um_ow[125]),
    .A2(um_ow[149]),
    .A3(um_ow[173]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[6].cell0_I  (.A0(um_ow[102]),
    .A1(um_ow[126]),
    .A2(um_ow[150]),
    .A3(um_ow[174]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[7].cell0_I  (.A0(um_ow[103]),
    .A1(um_ow[127]),
    .A2(um_ow[151]),
    .A3(um_ow[175]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[8].cell0_I  (.A0(um_ow[104]),
    .A1(um_ow[128]),
    .A2(um_ow[152]),
    .A3(um_ow[176]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_2 \block[4].genblk1.mux4_I[9].cell0_I  (.A0(um_ow[105]),
    .A1(um_ow[129]),
    .A2(um_ow[153]),
    .A3(um_ow[177]),
    .S0(\block[4].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[4].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[4].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__buf_2 \block[4].genblk1.mux4_sel_buf_I[0].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .X(\block[4].genblk1.mux4_sel_buf_I[0].z ));
 sky130_fd_sc_hd__buf_2 \block[4].genblk1.mux4_sel_buf_I[1].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .X(\block[4].genblk1.mux4_sel_buf_I[1].z ));
 sky130_fd_sc_hd__bufinv_8 \block[4].genblk1.tbuf_blk_ena_I.cell0_I  (.A(\block[4].genblk1.grp_sel_buf_I.z ),
    .Y(\block[4].genblk1.tbuf_blk_ena_I.tx ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[0].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[0].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[10].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[10].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[11].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[11].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[12].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[12].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[13].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[13].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[14].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[14].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[15].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[15].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[16].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[16].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[17].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[17].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[18].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[18].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[19].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[19].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[1].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[1].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[20].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[20].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[21].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[21].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[22].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[22].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[23].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[23].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[2].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[2].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[3].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[3].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[4].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[4].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[5].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[5].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[6].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[6].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[7].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[7].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[8].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[8].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__ebufn_8 \block[4].genblk1.tbuf_spine_ow_I[9].genblk1.cell0_I  (.A(\block[4].genblk1.mux4_I[9].x ),
    .TE_B(\block[4].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__buf_8 \block[4].l_ena_0_I.genblk1.cell0_I  (.A(\block[4].l_ena_0_I.a ),
    .X(\block[4].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[4].tie_I.cell_I  (.HI(\block[4].tie_I.hi ),
    .LO(\block[4].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[4].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[4].l_ena_0_I.z ),
    .X(\block[4].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[4].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[4].l_ena_0_I.z ),
    .Y(\block[4].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[0].cell0_I  (.DIODE(um_ow[120]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[10].cell0_I  (.DIODE(um_ow[130]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[11].cell0_I  (.DIODE(um_ow[131]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[12].cell0_I  (.DIODE(um_ow[132]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[13].cell0_I  (.DIODE(um_ow[133]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[14].cell0_I  (.DIODE(um_ow[134]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[15].cell0_I  (.DIODE(um_ow[135]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[16].cell0_I  (.DIODE(um_ow[136]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[17].cell0_I  (.DIODE(um_ow[137]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[18].cell0_I  (.DIODE(um_ow[138]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[19].cell0_I  (.DIODE(um_ow[139]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[1].cell0_I  (.DIODE(um_ow[121]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[20].cell0_I  (.DIODE(um_ow[140]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[21].cell0_I  (.DIODE(um_ow[141]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[22].cell0_I  (.DIODE(um_ow[142]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[23].cell0_I  (.DIODE(um_ow[143]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[2].cell0_I  (.DIODE(um_ow[122]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[3].cell0_I  (.DIODE(um_ow[123]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[4].cell0_I  (.DIODE(um_ow[124]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[5].cell0_I  (.DIODE(um_ow[125]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[6].cell0_I  (.DIODE(um_ow[126]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[7].cell0_I  (.DIODE(um_ow[127]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[8].cell0_I  (.DIODE(um_ow[128]));
 sky130_fd_sc_hd__diode_2 \block[5].diode_I[9].cell0_I  (.DIODE(um_ow[129]));
 sky130_fd_sc_hd__buf_8 \block[5].l_ena_0_I.genblk1.cell0_I  (.A(\block[5].l_ena_0_I.a ),
    .X(\block[5].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[5].tie_I.cell_I  (.HI(\block[5].tie_I.hi ),
    .LO(\block[5].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[5].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[5].l_ena_0_I.z ),
    .X(\block[5].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[5].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[5].l_ena_0_I.z ),
    .Y(\block[5].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[0].cell0_I  (.DIODE(um_ow[144]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[10].cell0_I  (.DIODE(um_ow[154]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[11].cell0_I  (.DIODE(um_ow[155]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[12].cell0_I  (.DIODE(um_ow[156]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[13].cell0_I  (.DIODE(um_ow[157]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[14].cell0_I  (.DIODE(um_ow[158]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[15].cell0_I  (.DIODE(um_ow[159]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[16].cell0_I  (.DIODE(um_ow[160]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[17].cell0_I  (.DIODE(um_ow[161]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[18].cell0_I  (.DIODE(um_ow[162]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[19].cell0_I  (.DIODE(um_ow[163]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[1].cell0_I  (.DIODE(um_ow[145]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[20].cell0_I  (.DIODE(um_ow[164]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[21].cell0_I  (.DIODE(um_ow[165]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[22].cell0_I  (.DIODE(um_ow[166]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[23].cell0_I  (.DIODE(um_ow[167]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[2].cell0_I  (.DIODE(um_ow[146]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[3].cell0_I  (.DIODE(um_ow[147]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[4].cell0_I  (.DIODE(um_ow[148]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[5].cell0_I  (.DIODE(um_ow[149]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[6].cell0_I  (.DIODE(um_ow[150]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[7].cell0_I  (.DIODE(um_ow[151]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[8].cell0_I  (.DIODE(um_ow[152]));
 sky130_fd_sc_hd__diode_2 \block[6].diode_I[9].cell0_I  (.DIODE(um_ow[153]));
 sky130_fd_sc_hd__buf_8 \block[6].l_ena_0_I.genblk1.cell0_I  (.A(\block[6].l_ena_0_I.a ),
    .X(\block[6].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[6].tie_I.cell_I  (.HI(\block[6].tie_I.hi ),
    .LO(\block[6].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[6].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[6].l_ena_0_I.z ),
    .X(\block[6].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[6].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[6].l_ena_0_I.z ),
    .Y(\block[6].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[0].cell0_I  (.DIODE(um_ow[168]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[10].cell0_I  (.DIODE(um_ow[178]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[11].cell0_I  (.DIODE(um_ow[179]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[12].cell0_I  (.DIODE(um_ow[180]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[13].cell0_I  (.DIODE(um_ow[181]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[14].cell0_I  (.DIODE(um_ow[182]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[15].cell0_I  (.DIODE(um_ow[183]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[16].cell0_I  (.DIODE(um_ow[184]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[17].cell0_I  (.DIODE(um_ow[185]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[18].cell0_I  (.DIODE(um_ow[186]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[19].cell0_I  (.DIODE(um_ow[187]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[1].cell0_I  (.DIODE(um_ow[169]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[20].cell0_I  (.DIODE(um_ow[188]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[21].cell0_I  (.DIODE(um_ow[189]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[22].cell0_I  (.DIODE(um_ow[190]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[23].cell0_I  (.DIODE(um_ow[191]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[2].cell0_I  (.DIODE(um_ow[170]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[3].cell0_I  (.DIODE(um_ow[171]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[4].cell0_I  (.DIODE(um_ow[172]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[5].cell0_I  (.DIODE(um_ow[173]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[6].cell0_I  (.DIODE(um_ow[174]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[7].cell0_I  (.DIODE(um_ow[175]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[8].cell0_I  (.DIODE(um_ow[176]));
 sky130_fd_sc_hd__diode_2 \block[7].diode_I[9].cell0_I  (.DIODE(um_ow[177]));
 sky130_fd_sc_hd__buf_8 \block[7].l_ena_0_I.genblk1.cell0_I  (.A(\block[7].l_ena_0_I.a ),
    .X(\block[7].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[7].tie_I.cell_I  (.HI(\block[7].tie_I.hi ),
    .LO(\block[7].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[7].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[7].l_ena_0_I.z ),
    .X(\block[7].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[7].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[7].l_ena_0_I.z ),
    .Y(\block[7].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[0].cell0_I  (.DIODE(um_ow[192]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[10].cell0_I  (.DIODE(um_ow[202]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[11].cell0_I  (.DIODE(um_ow[203]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[12].cell0_I  (.DIODE(um_ow[204]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[13].cell0_I  (.DIODE(um_ow[205]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[14].cell0_I  (.DIODE(um_ow[206]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[15].cell0_I  (.DIODE(um_ow[207]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[16].cell0_I  (.DIODE(um_ow[208]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[17].cell0_I  (.DIODE(um_ow[209]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[18].cell0_I  (.DIODE(um_ow[210]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[19].cell0_I  (.DIODE(um_ow[211]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[1].cell0_I  (.DIODE(um_ow[193]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[20].cell0_I  (.DIODE(um_ow[212]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[21].cell0_I  (.DIODE(um_ow[213]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[22].cell0_I  (.DIODE(um_ow[214]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[23].cell0_I  (.DIODE(um_ow[215]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[2].cell0_I  (.DIODE(um_ow[194]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[3].cell0_I  (.DIODE(um_ow[195]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[4].cell0_I  (.DIODE(um_ow[196]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[5].cell0_I  (.DIODE(um_ow[197]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[6].cell0_I  (.DIODE(um_ow[198]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[7].cell0_I  (.DIODE(um_ow[199]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[8].cell0_I  (.DIODE(um_ow[200]));
 sky130_fd_sc_hd__diode_2 \block[8].diode_I[9].cell0_I  (.DIODE(um_ow[201]));
 sky130_fd_sc_hd__buf_2 \block[8].genblk1.grp_sel_buf_I.genblk1.cell0_I  (.A(\block[8].genblk1.grp_sel_buf_I.a ),
    .X(\block[8].genblk1.grp_sel_buf_I.z ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[0].cell0_I  (.A0(um_ow[192]),
    .A1(um_ow[216]),
    .A2(um_ow[240]),
    .A3(um_ow[264]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[0].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[10].cell0_I  (.A0(um_ow[202]),
    .A1(um_ow[226]),
    .A2(um_ow[250]),
    .A3(um_ow[274]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[10].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[11].cell0_I  (.A0(um_ow[203]),
    .A1(um_ow[227]),
    .A2(um_ow[251]),
    .A3(um_ow[275]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[11].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[12].cell0_I  (.A0(um_ow[204]),
    .A1(um_ow[228]),
    .A2(um_ow[252]),
    .A3(um_ow[276]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[12].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[13].cell0_I  (.A0(um_ow[205]),
    .A1(um_ow[229]),
    .A2(um_ow[253]),
    .A3(um_ow[277]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[13].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[14].cell0_I  (.A0(um_ow[206]),
    .A1(um_ow[230]),
    .A2(um_ow[254]),
    .A3(um_ow[278]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[14].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[15].cell0_I  (.A0(um_ow[207]),
    .A1(um_ow[231]),
    .A2(um_ow[255]),
    .A3(um_ow[279]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[15].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[16].cell0_I  (.A0(um_ow[208]),
    .A1(um_ow[232]),
    .A2(um_ow[256]),
    .A3(um_ow[280]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[16].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[17].cell0_I  (.A0(um_ow[209]),
    .A1(um_ow[233]),
    .A2(um_ow[257]),
    .A3(um_ow[281]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[17].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[18].cell0_I  (.A0(um_ow[210]),
    .A1(um_ow[234]),
    .A2(um_ow[258]),
    .A3(um_ow[282]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[18].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[19].cell0_I  (.A0(um_ow[211]),
    .A1(um_ow[235]),
    .A2(um_ow[259]),
    .A3(um_ow[283]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[19].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[1].cell0_I  (.A0(um_ow[193]),
    .A1(um_ow[217]),
    .A2(um_ow[241]),
    .A3(um_ow[265]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[1].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[20].cell0_I  (.A0(um_ow[212]),
    .A1(um_ow[236]),
    .A2(um_ow[260]),
    .A3(um_ow[284]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[20].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[21].cell0_I  (.A0(um_ow[213]),
    .A1(um_ow[237]),
    .A2(um_ow[261]),
    .A3(um_ow[285]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[21].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[22].cell0_I  (.A0(um_ow[214]),
    .A1(um_ow[238]),
    .A2(um_ow[262]),
    .A3(um_ow[286]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[22].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[23].cell0_I  (.A0(um_ow[215]),
    .A1(um_ow[239]),
    .A2(um_ow[263]),
    .A3(um_ow[287]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[23].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[2].cell0_I  (.A0(um_ow[194]),
    .A1(um_ow[218]),
    .A2(um_ow[242]),
    .A3(um_ow[266]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[2].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[3].cell0_I  (.A0(um_ow[195]),
    .A1(um_ow[219]),
    .A2(um_ow[243]),
    .A3(um_ow[267]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[3].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[4].cell0_I  (.A0(um_ow[196]),
    .A1(um_ow[220]),
    .A2(um_ow[244]),
    .A3(um_ow[268]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[4].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[5].cell0_I  (.A0(um_ow[197]),
    .A1(um_ow[221]),
    .A2(um_ow[245]),
    .A3(um_ow[269]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[5].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[6].cell0_I  (.A0(um_ow[198]),
    .A1(um_ow[222]),
    .A2(um_ow[246]),
    .A3(um_ow[270]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[6].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[7].cell0_I  (.A0(um_ow[199]),
    .A1(um_ow[223]),
    .A2(um_ow[247]),
    .A3(um_ow[271]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[7].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[8].cell0_I  (.A0(um_ow[200]),
    .A1(um_ow[224]),
    .A2(um_ow[248]),
    .A3(um_ow[272]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[8].x ));
 sky130_fd_sc_hd__mux4_2 \block[8].genblk1.mux4_I[9].cell0_I  (.A0(um_ow[201]),
    .A1(um_ow[225]),
    .A2(um_ow[249]),
    .A3(um_ow[273]),
    .S0(\block[8].genblk1.mux4_sel_buf_I[0].z ),
    .S1(\block[8].genblk1.mux4_sel_buf_I[1].z ),
    .X(\block[8].genblk1.mux4_I[9].x ));
 sky130_fd_sc_hd__buf_2 \block[8].genblk1.mux4_sel_buf_I[0].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[0].a ),
    .X(\block[8].genblk1.mux4_sel_buf_I[0].z ));
 sky130_fd_sc_hd__buf_2 \block[8].genblk1.mux4_sel_buf_I[1].genblk1.cell0_I  (.A(\block[0].genblk1.mux4_sel_buf_I[1].a ),
    .X(\block[8].genblk1.mux4_sel_buf_I[1].z ));
 sky130_fd_sc_hd__bufinv_8 \block[8].genblk1.tbuf_blk_ena_I.cell0_I  (.A(\block[8].genblk1.grp_sel_buf_I.z ),
    .Y(\block[8].genblk1.tbuf_blk_ena_I.tx ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[0].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[0].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[10].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[10].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[11].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[11].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[12].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[12].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[13].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[13].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[14].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[14].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[15].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[15].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[16].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[16].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[17].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[17].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[18].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[18].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[19].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[19].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[1].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[1].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[20].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[20].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[21].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[21].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[22].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[22].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[23].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[23].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[2].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[2].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[3].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[3].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[4].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[4].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[5].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[5].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[6].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[6].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[7].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[7].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[8].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[8].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__ebufn_8 \block[8].genblk1.tbuf_spine_ow_I[9].genblk1.cell0_I  (.A(\block[8].genblk1.mux4_I[9].x ),
    .TE_B(\block[8].genblk1.tbuf_blk_ena_I.tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__buf_8 \block[8].l_ena_0_I.genblk1.cell0_I  (.A(\block[8].l_ena_0_I.a ),
    .X(\block[8].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[8].tie_I.cell_I  (.HI(\block[8].tie_I.hi ),
    .LO(\block[8].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[8].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[8].l_ena_0_I.z ),
    .X(\block[8].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[8].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[8].l_ena_0_I.z ),
    .Y(\block[8].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[0].cell0_I  (.DIODE(um_ow[216]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[10].cell0_I  (.DIODE(um_ow[226]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[11].cell0_I  (.DIODE(um_ow[227]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[12].cell0_I  (.DIODE(um_ow[228]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[13].cell0_I  (.DIODE(um_ow[229]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[14].cell0_I  (.DIODE(um_ow[230]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[15].cell0_I  (.DIODE(um_ow[231]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[16].cell0_I  (.DIODE(um_ow[232]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[17].cell0_I  (.DIODE(um_ow[233]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[18].cell0_I  (.DIODE(um_ow[234]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[19].cell0_I  (.DIODE(um_ow[235]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[1].cell0_I  (.DIODE(um_ow[217]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[20].cell0_I  (.DIODE(um_ow[236]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[21].cell0_I  (.DIODE(um_ow[237]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[22].cell0_I  (.DIODE(um_ow[238]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[23].cell0_I  (.DIODE(um_ow[239]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[2].cell0_I  (.DIODE(um_ow[218]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[3].cell0_I  (.DIODE(um_ow[219]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[4].cell0_I  (.DIODE(um_ow[220]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[5].cell0_I  (.DIODE(um_ow[221]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[6].cell0_I  (.DIODE(um_ow[222]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[7].cell0_I  (.DIODE(um_ow[223]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[8].cell0_I  (.DIODE(um_ow[224]));
 sky130_fd_sc_hd__diode_2 \block[9].diode_I[9].cell0_I  (.DIODE(um_ow[225]));
 sky130_fd_sc_hd__buf_8 \block[9].l_ena_0_I.genblk1.cell0_I  (.A(\block[9].l_ena_0_I.a ),
    .X(\block[9].l_ena_0_I.z ));
 sky130_fd_sc_hd__conb_1 \block[9].tie_I.cell_I  (.HI(\block[9].tie_I.hi ),
    .LO(\block[9].tie_I.lo ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[0].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[0].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[0].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[10].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[10].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[10].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[11].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[11].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[11].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[12].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[12].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[12].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[13].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[13].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[13].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[14].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[14].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[14].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[15].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[15].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[15].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[16].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[16].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[16].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[17].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[17].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[17].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[1].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[1].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[1].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[2].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[2].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[2].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[3].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[3].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[3].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[4].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[4].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[4].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[5].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[5].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[5].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[6].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[6].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[6].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[7].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[7].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[7].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[8].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[8].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[8].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_bot_iw_I[9].genblk1.cell0_I  (.A(\block[0].zbuf_bot_iw_I[9].a ),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_bot_iw_I[9].z ));
 sky130_fd_sc_hd__and2_2 \block[9].zbuf_ena_I.genblk1.cell0_I  (.A(one_),
    .B(\block[9].l_ena_0_I.z ),
    .X(\block[9].zbuf_ena_I.z ));
 sky130_fd_sc_hd__bufinv_8 \block[9].zbuf_pg_vdd_I.genblk1.cell0_I  (.A(\block[9].l_ena_0_I.z ),
    .Y(\block[9].zbuf_pg_vdd_I.z ));
 sky130_fd_sc_hd__buf_2 \branch_addr_match_buf_I[0].genblk1.cell0_I  (.A(spine_iw[7]),
    .X(\branch_addr_match_buf_I[0].z ));
 sky130_fd_sc_hd__buf_2 \branch_addr_match_buf_I[1].genblk1.cell0_I  (.A(spine_iw[8]),
    .X(\branch_addr_match_buf_I[1].z ));
 sky130_fd_sc_hd__buf_2 \branch_addr_match_buf_I[2].genblk1.cell0_I  (.A(spine_iw[9]),
    .X(\branch_addr_match_buf_I[2].z ));
 sky130_fd_sc_hd__buf_2 \branch_addr_match_buf_I[3].genblk1.cell0_I  (.A(spine_iw[10]),
    .X(\branch_addr_match_buf_I[3].z ));
 sky130_fd_sc_hd__buf_2 \branch_ena_buf_I.genblk1.cell0_I  (.A(spine_iw[1]),
    .X(\branch_ena_buf_I.z ));
 sky130_fd_sc_hd__buf_8 \branch_sel_buf_I.genblk1.cell0_I  (.A(\branch_sel_buf_I.a ),
    .X(\branch_sel_buf_I.z ));
 sky130_fd_sc_hd__inv_2 \branch_sel_n_buf_I.genblk1.cell0_I  (.A(\branch_sel_buf_I.z ),
    .Y(\branch_sel_n_buf_I.z ));
 sky130_fd_sc_hd__buf_8 \buf_bus_ena_I.genblk1.cell0_I  (.A(\branch_sel_buf_I.z ),
    .X(\buf_bus_ena_I.z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[0].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[0].z ),
    .X(\buf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[10].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[10].z ),
    .X(\buf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[11].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[11].z ),
    .X(\buf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[12].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[12].z ),
    .X(\buf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[13].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[13].z ),
    .X(\buf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[14].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[14].z ),
    .X(\buf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[15].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[15].z ),
    .X(\buf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[16].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[16].z ),
    .X(\buf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[17].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[17].z ),
    .X(\buf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[18].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[18].z ),
    .X(\buf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[19].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[19].z ),
    .X(\buf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[1].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[1].z ),
    .X(\buf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[20].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[20].z ),
    .X(\buf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[21].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[21].z ),
    .X(\buf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[22].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[22].z ),
    .X(\buf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[23].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[23].z ),
    .X(\buf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[2].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[2].z ),
    .X(\buf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[3].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[3].z ),
    .X(\buf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[4].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[4].z ),
    .X(\buf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[5].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[5].z ),
    .X(\buf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[6].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[6].z ),
    .X(\buf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[7].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[7].z ),
    .X(\buf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[8].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[8].z ),
    .X(\buf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__buf_2 \buf_spine_ow_I[9].genblk1.cell0_I  (.A(\block[0].genblk1.tbuf_spine_ow_I[9].z ),
    .X(\buf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[0].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[10].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[11].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[12].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[13].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[14].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[15].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[16].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[17].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[18].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[19].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[1].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[20].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[21].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[22].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[23].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[2].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[3].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[4].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[5].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[6].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[7].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[8].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__ebufn_1 \bus_pull_ow_I[9].genblk1.cell0_I  (.A(\bus_pull_ow_I[0].a ),
    .TE_B(\bus_pull_ow_I[0].tx ),
    .Z(\block[0].genblk1.tbuf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__conb_1 \bus_pull_tie_I.cell_I  (.HI(\bus_pull_tie_I.hi ),
    .LO(\bus_pull_ow_I[0].a ));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[0].cell0_I  (.DIODE(spine_iw[0]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[10].cell0_I  (.DIODE(spine_iw[10]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[11].cell0_I  (.DIODE(spine_iw[11]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[12].cell0_I  (.DIODE(spine_iw[12]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[13].cell0_I  (.DIODE(spine_iw[13]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[14].cell0_I  (.DIODE(spine_iw[14]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[15].cell0_I  (.DIODE(spine_iw[15]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[16].cell0_I  (.DIODE(spine_iw[16]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[17].cell0_I  (.DIODE(spine_iw[17]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[18].cell0_I  (.DIODE(spine_iw[18]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[19].cell0_I  (.DIODE(spine_iw[19]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[1].cell0_I  (.DIODE(spine_iw[1]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[20].cell0_I  (.DIODE(spine_iw[20]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[21].cell0_I  (.DIODE(spine_iw[21]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[22].cell0_I  (.DIODE(spine_iw[22]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[23].cell0_I  (.DIODE(spine_iw[23]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[24].cell0_I  (.DIODE(spine_iw[24]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[25].cell0_I  (.DIODE(spine_iw[25]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[26].cell0_I  (.DIODE(spine_iw[26]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[27].cell0_I  (.DIODE(spine_iw[27]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[28].cell0_I  (.DIODE(spine_iw[28]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[29].cell0_I  (.DIODE(spine_iw[29]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[2].cell0_I  (.DIODE(spine_iw[2]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[3].cell0_I  (.DIODE(spine_iw[3]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[4].cell0_I  (.DIODE(spine_iw[4]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[5].cell0_I  (.DIODE(spine_iw[5]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[6].cell0_I  (.DIODE(spine_iw[6]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[7].cell0_I  (.DIODE(spine_iw[7]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[8].cell0_I  (.DIODE(spine_iw[8]));
 sky130_fd_sc_hd__diode_2 \diode_spine_I[9].cell0_I  (.DIODE(spine_iw[9]));
 sky130_fd_sc_hd__bufinv_8 \tbuf_row_ena_I.cell0_I  (.A(\branch_sel_buf_I.z ),
    .Y(\tbuf_row_ena_I.tx ));
 sky130_fd_sc_hd__bufinv_8 \tbuf_row_ena_n_I.cell0_I  (.A(\branch_sel_n_buf_I.z ),
    .Y(\bus_pull_ow_I[0].tx ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[0].genblk1.cell0_I  (.A(\buf_spine_ow_I[0].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[0].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[10].genblk1.cell0_I  (.A(\buf_spine_ow_I[10].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[10].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[11].genblk1.cell0_I  (.A(\buf_spine_ow_I[11].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[11].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[12].genblk1.cell0_I  (.A(\buf_spine_ow_I[12].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[12].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[13].genblk1.cell0_I  (.A(\buf_spine_ow_I[13].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[13].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[14].genblk1.cell0_I  (.A(\buf_spine_ow_I[14].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[14].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[15].genblk1.cell0_I  (.A(\buf_spine_ow_I[15].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[15].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[16].genblk1.cell0_I  (.A(\buf_spine_ow_I[16].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[16].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[17].genblk1.cell0_I  (.A(\buf_spine_ow_I[17].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[17].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[18].genblk1.cell0_I  (.A(\buf_spine_ow_I[18].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[18].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[19].genblk1.cell0_I  (.A(\buf_spine_ow_I[19].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[19].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[1].genblk1.cell0_I  (.A(\buf_spine_ow_I[1].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[1].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[20].genblk1.cell0_I  (.A(\buf_spine_ow_I[20].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[20].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[21].genblk1.cell0_I  (.A(\buf_spine_ow_I[21].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[21].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[22].genblk1.cell0_I  (.A(\buf_spine_ow_I[22].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[22].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[23].genblk1.cell0_I  (.A(\buf_spine_ow_I[23].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[23].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[2].genblk1.cell0_I  (.A(\buf_spine_ow_I[2].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[2].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[3].genblk1.cell0_I  (.A(\buf_spine_ow_I[3].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[3].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[4].genblk1.cell0_I  (.A(\buf_spine_ow_I[4].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[4].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[5].genblk1.cell0_I  (.A(\buf_spine_ow_I[5].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[5].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[6].genblk1.cell0_I  (.A(\buf_spine_ow_I[6].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[6].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[7].genblk1.cell0_I  (.A(\buf_spine_ow_I[7].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[7].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[8].genblk1.cell0_I  (.A(\buf_spine_ow_I[8].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[8].z ));
 sky130_fd_sc_hd__ebufn_8 \tbuf_spine_ow_I[9].genblk1.cell0_I  (.A(\buf_spine_ow_I[9].z ),
    .TE_B(\tbuf_row_ena_I.tx ),
    .Z(\tbuf_spine_ow_I[9].z ));
 sky130_fd_sc_hd__conb_1 \tie_I.cell_I  (.HI(k_one),
    .LO(k_zero));
 sky130_fd_sc_hd__conb_1 \tie_spine_guard_I[0].cell_I  (.HI(\tie_spine_guard_I[0].hi ),
    .LO(\tie_spine_guard_I[0].lo ));
 sky130_fd_sc_hd__conb_1 \tie_spine_guard_I[1].cell_I  (.HI(\tie_spine_guard_I[1].hi ),
    .LO(\tie_spine_guard_I[1].lo ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[0].genblk1.cell0_I  (.A(spine_iw[11]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[0].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[0].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[0].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[10].genblk1.cell0_I  (.A(spine_iw[21]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[10].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[10].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[10].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[10].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[11].genblk1.cell0_I  (.A(spine_iw[22]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[11].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[11].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[11].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[11].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[12].genblk1.cell0_I  (.A(spine_iw[23]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[12].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[12].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[12].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[12].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[13].genblk1.cell0_I  (.A(spine_iw[24]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[13].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[13].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[13].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[13].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[14].genblk1.cell0_I  (.A(spine_iw[25]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[14].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[14].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[14].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[15].genblk1.cell0_I  (.A(spine_iw[26]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[15].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[15].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[15].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[15].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[16].genblk1.cell0_I  (.A(spine_iw[27]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[16].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[16].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[16].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[16].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[17].genblk1.cell0_I  (.A(spine_iw[28]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[17].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[17].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[17].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[17].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[1].genblk1.cell0_I  (.A(spine_iw[12]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[1].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[1].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[1].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[1].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[2].genblk1.cell0_I  (.A(spine_iw[13]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[2].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[2].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[2].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[3].genblk1.cell0_I  (.A(spine_iw[14]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[3].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[3].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[4].genblk1.cell0_I  (.A(spine_iw[15]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[4].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[4].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[4].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[5].genblk1.cell0_I  (.A(spine_iw[16]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[5].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[5].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[5].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[5].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[6].genblk1.cell0_I  (.A(spine_iw[17]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[6].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[6].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[6].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[6].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[7].genblk1.cell0_I  (.A(spine_iw[18]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[7].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[7].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[7].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[7].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[8].genblk1.cell0_I  (.A(spine_iw[19]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[8].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[8].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[8].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[8].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_iw_I[9].genblk1.cell0_I  (.A(spine_iw[20]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_iw_I[9].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_iw_I[9].genblk1.cell1_I  (.A(\zbuf_bus_iw_I[9].genblk1.l ),
    .X(\block[0].zbuf_bot_iw_I[9].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_sel_I[0].genblk1.cell0_I  (.A(spine_iw[2]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_sel_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[0].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[0].genblk1.l ),
    .X(\block[0].genblk1.mux4_sel_buf_I[0].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_sel_I[1].genblk1.cell0_I  (.A(spine_iw[3]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_sel_I[1].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[1].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[1].genblk1.l ),
    .X(\block[0].genblk1.mux4_sel_buf_I[1].a ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_sel_I[2].genblk1.cell0_I  (.A(spine_iw[4]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_sel_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[2].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[2].genblk1.l ),
    .X(\zbuf_bus_sel_I[2].z ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_sel_I[3].genblk1.cell0_I  (.A(spine_iw[5]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_sel_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[3].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[3].genblk1.l ),
    .X(\zbuf_bus_sel_I[3].z ));
 sky130_fd_sc_hd__and2_2 \zbuf_bus_sel_I[4].genblk1.cell0_I  (.A(spine_iw[6]),
    .B(\branch_sel_buf_I.z ),
    .X(\zbuf_bus_sel_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \zbuf_bus_sel_I[4].genblk1.cell1_I  (.A(\zbuf_bus_sel_I[4].genblk1.l ),
    .X(\zbuf_bus_sel_I[4].z ));
 sky130_fd_sc_hd__conb_1 TIE_ONE_one_ (.HI(one_));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1085 ();
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\block[0].genblk1.mux4_sel_buf_I[1].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\block[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\block[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(um_ow[114]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(um_ow[118]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(um_ow[119]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(um_ow[139]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(um_ow[140]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(um_ow[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(um_ow[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(um_ow[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(um_ow[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(um_ow[42]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\block[0].zbuf_bot_iw_I[14].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\block[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\block[0].zbuf_bot_iw_I[3].a ));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2071 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_2658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_2781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_2789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_2913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_2181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_2237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_2809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_2844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2863 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_2907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1858 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_2293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_2402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_2466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_2769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2899 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_2937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1760 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2226 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_2356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2590 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2812 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_2809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2842 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2891 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2899 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2940 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2880 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_2937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2807 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_2869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_2843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2868 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2927 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_2937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1618 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2803 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2842 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2886 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2924 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_2932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_2937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_2841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_2892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_2359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2450 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_2321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_2901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2801 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2917 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1619 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_2097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_2141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_2151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_2421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_2428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_2471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_2893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1918 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_2067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2071 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_2325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_2387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_2789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2937 ();
 assign um_k_zero[0] = \block[0].tie_I.lo ;
 assign um_iw[0] = \block[0].zbuf_bot_iw_I[0].z ;
 assign um_iw[10] = \block[0].zbuf_bot_iw_I[10].z ;
 assign um_iw[11] = \block[0].zbuf_bot_iw_I[11].z ;
 assign um_iw[12] = \block[0].zbuf_bot_iw_I[12].z ;
 assign um_iw[13] = \block[0].zbuf_bot_iw_I[13].z ;
 assign um_iw[14] = \block[0].zbuf_bot_iw_I[14].z ;
 assign um_iw[15] = \block[0].zbuf_bot_iw_I[15].z ;
 assign um_iw[16] = \block[0].zbuf_bot_iw_I[16].z ;
 assign um_iw[17] = \block[0].zbuf_bot_iw_I[17].z ;
 assign um_iw[1] = \block[0].zbuf_bot_iw_I[1].z ;
 assign um_iw[2] = \block[0].zbuf_bot_iw_I[2].z ;
 assign um_iw[3] = \block[0].zbuf_bot_iw_I[3].z ;
 assign um_iw[4] = \block[0].zbuf_bot_iw_I[4].z ;
 assign um_iw[5] = \block[0].zbuf_bot_iw_I[5].z ;
 assign um_iw[6] = \block[0].zbuf_bot_iw_I[6].z ;
 assign um_iw[7] = \block[0].zbuf_bot_iw_I[7].z ;
 assign um_iw[8] = \block[0].zbuf_bot_iw_I[8].z ;
 assign um_iw[9] = \block[0].zbuf_bot_iw_I[9].z ;
 assign um_ena[0] = \block[0].zbuf_ena_I.z ;
 assign um_pg_vdd[0] = \block[0].zbuf_pg_vdd_I.z ;
 assign um_k_zero[10] = \block[10].tie_I.lo ;
 assign um_iw[180] = \block[10].zbuf_bot_iw_I[0].z ;
 assign um_iw[190] = \block[10].zbuf_bot_iw_I[10].z ;
 assign um_iw[191] = \block[10].zbuf_bot_iw_I[11].z ;
 assign um_iw[192] = \block[10].zbuf_bot_iw_I[12].z ;
 assign um_iw[193] = \block[10].zbuf_bot_iw_I[13].z ;
 assign um_iw[194] = \block[10].zbuf_bot_iw_I[14].z ;
 assign um_iw[195] = \block[10].zbuf_bot_iw_I[15].z ;
 assign um_iw[196] = \block[10].zbuf_bot_iw_I[16].z ;
 assign um_iw[197] = \block[10].zbuf_bot_iw_I[17].z ;
 assign um_iw[181] = \block[10].zbuf_bot_iw_I[1].z ;
 assign um_iw[182] = \block[10].zbuf_bot_iw_I[2].z ;
 assign um_iw[183] = \block[10].zbuf_bot_iw_I[3].z ;
 assign um_iw[184] = \block[10].zbuf_bot_iw_I[4].z ;
 assign um_iw[185] = \block[10].zbuf_bot_iw_I[5].z ;
 assign um_iw[186] = \block[10].zbuf_bot_iw_I[6].z ;
 assign um_iw[187] = \block[10].zbuf_bot_iw_I[7].z ;
 assign um_iw[188] = \block[10].zbuf_bot_iw_I[8].z ;
 assign um_iw[189] = \block[10].zbuf_bot_iw_I[9].z ;
 assign um_ena[10] = \block[10].zbuf_ena_I.z ;
 assign um_pg_vdd[10] = \block[10].zbuf_pg_vdd_I.z ;
 assign um_k_zero[11] = \block[11].tie_I.lo ;
 assign um_iw[198] = \block[11].zbuf_bot_iw_I[0].z ;
 assign um_iw[208] = \block[11].zbuf_bot_iw_I[10].z ;
 assign um_iw[209] = \block[11].zbuf_bot_iw_I[11].z ;
 assign um_iw[210] = \block[11].zbuf_bot_iw_I[12].z ;
 assign um_iw[211] = \block[11].zbuf_bot_iw_I[13].z ;
 assign um_iw[212] = \block[11].zbuf_bot_iw_I[14].z ;
 assign um_iw[213] = \block[11].zbuf_bot_iw_I[15].z ;
 assign um_iw[214] = \block[11].zbuf_bot_iw_I[16].z ;
 assign um_iw[215] = \block[11].zbuf_bot_iw_I[17].z ;
 assign um_iw[199] = \block[11].zbuf_bot_iw_I[1].z ;
 assign um_iw[200] = \block[11].zbuf_bot_iw_I[2].z ;
 assign um_iw[201] = \block[11].zbuf_bot_iw_I[3].z ;
 assign um_iw[202] = \block[11].zbuf_bot_iw_I[4].z ;
 assign um_iw[203] = \block[11].zbuf_bot_iw_I[5].z ;
 assign um_iw[204] = \block[11].zbuf_bot_iw_I[6].z ;
 assign um_iw[205] = \block[11].zbuf_bot_iw_I[7].z ;
 assign um_iw[206] = \block[11].zbuf_bot_iw_I[8].z ;
 assign um_iw[207] = \block[11].zbuf_bot_iw_I[9].z ;
 assign um_ena[11] = \block[11].zbuf_ena_I.z ;
 assign um_pg_vdd[11] = \block[11].zbuf_pg_vdd_I.z ;
 assign um_k_zero[12] = \block[12].tie_I.lo ;
 assign um_iw[216] = \block[12].zbuf_bot_iw_I[0].z ;
 assign um_iw[226] = \block[12].zbuf_bot_iw_I[10].z ;
 assign um_iw[227] = \block[12].zbuf_bot_iw_I[11].z ;
 assign um_iw[228] = \block[12].zbuf_bot_iw_I[12].z ;
 assign um_iw[229] = \block[12].zbuf_bot_iw_I[13].z ;
 assign um_iw[230] = \block[12].zbuf_bot_iw_I[14].z ;
 assign um_iw[231] = \block[12].zbuf_bot_iw_I[15].z ;
 assign um_iw[232] = \block[12].zbuf_bot_iw_I[16].z ;
 assign um_iw[233] = \block[12].zbuf_bot_iw_I[17].z ;
 assign um_iw[217] = \block[12].zbuf_bot_iw_I[1].z ;
 assign um_iw[218] = \block[12].zbuf_bot_iw_I[2].z ;
 assign um_iw[219] = \block[12].zbuf_bot_iw_I[3].z ;
 assign um_iw[220] = \block[12].zbuf_bot_iw_I[4].z ;
 assign um_iw[221] = \block[12].zbuf_bot_iw_I[5].z ;
 assign um_iw[222] = \block[12].zbuf_bot_iw_I[6].z ;
 assign um_iw[223] = \block[12].zbuf_bot_iw_I[7].z ;
 assign um_iw[224] = \block[12].zbuf_bot_iw_I[8].z ;
 assign um_iw[225] = \block[12].zbuf_bot_iw_I[9].z ;
 assign um_ena[12] = \block[12].zbuf_ena_I.z ;
 assign um_pg_vdd[12] = \block[12].zbuf_pg_vdd_I.z ;
 assign um_k_zero[13] = \block[13].tie_I.lo ;
 assign um_iw[234] = \block[13].zbuf_bot_iw_I[0].z ;
 assign um_iw[244] = \block[13].zbuf_bot_iw_I[10].z ;
 assign um_iw[245] = \block[13].zbuf_bot_iw_I[11].z ;
 assign um_iw[246] = \block[13].zbuf_bot_iw_I[12].z ;
 assign um_iw[247] = \block[13].zbuf_bot_iw_I[13].z ;
 assign um_iw[248] = \block[13].zbuf_bot_iw_I[14].z ;
 assign um_iw[249] = \block[13].zbuf_bot_iw_I[15].z ;
 assign um_iw[250] = \block[13].zbuf_bot_iw_I[16].z ;
 assign um_iw[251] = \block[13].zbuf_bot_iw_I[17].z ;
 assign um_iw[235] = \block[13].zbuf_bot_iw_I[1].z ;
 assign um_iw[236] = \block[13].zbuf_bot_iw_I[2].z ;
 assign um_iw[237] = \block[13].zbuf_bot_iw_I[3].z ;
 assign um_iw[238] = \block[13].zbuf_bot_iw_I[4].z ;
 assign um_iw[239] = \block[13].zbuf_bot_iw_I[5].z ;
 assign um_iw[240] = \block[13].zbuf_bot_iw_I[6].z ;
 assign um_iw[241] = \block[13].zbuf_bot_iw_I[7].z ;
 assign um_iw[242] = \block[13].zbuf_bot_iw_I[8].z ;
 assign um_iw[243] = \block[13].zbuf_bot_iw_I[9].z ;
 assign um_ena[13] = \block[13].zbuf_ena_I.z ;
 assign um_pg_vdd[13] = \block[13].zbuf_pg_vdd_I.z ;
 assign um_k_zero[14] = \block[14].tie_I.lo ;
 assign um_iw[252] = \block[14].zbuf_bot_iw_I[0].z ;
 assign um_iw[262] = \block[14].zbuf_bot_iw_I[10].z ;
 assign um_iw[263] = \block[14].zbuf_bot_iw_I[11].z ;
 assign um_iw[264] = \block[14].zbuf_bot_iw_I[12].z ;
 assign um_iw[265] = \block[14].zbuf_bot_iw_I[13].z ;
 assign um_iw[266] = \block[14].zbuf_bot_iw_I[14].z ;
 assign um_iw[267] = \block[14].zbuf_bot_iw_I[15].z ;
 assign um_iw[268] = \block[14].zbuf_bot_iw_I[16].z ;
 assign um_iw[269] = \block[14].zbuf_bot_iw_I[17].z ;
 assign um_iw[253] = \block[14].zbuf_bot_iw_I[1].z ;
 assign um_iw[254] = \block[14].zbuf_bot_iw_I[2].z ;
 assign um_iw[255] = \block[14].zbuf_bot_iw_I[3].z ;
 assign um_iw[256] = \block[14].zbuf_bot_iw_I[4].z ;
 assign um_iw[257] = \block[14].zbuf_bot_iw_I[5].z ;
 assign um_iw[258] = \block[14].zbuf_bot_iw_I[6].z ;
 assign um_iw[259] = \block[14].zbuf_bot_iw_I[7].z ;
 assign um_iw[260] = \block[14].zbuf_bot_iw_I[8].z ;
 assign um_iw[261] = \block[14].zbuf_bot_iw_I[9].z ;
 assign um_ena[14] = \block[14].zbuf_ena_I.z ;
 assign um_pg_vdd[14] = \block[14].zbuf_pg_vdd_I.z ;
 assign um_k_zero[15] = \block[15].tie_I.lo ;
 assign um_iw[270] = \block[15].zbuf_bot_iw_I[0].z ;
 assign um_iw[280] = \block[15].zbuf_bot_iw_I[10].z ;
 assign um_iw[281] = \block[15].zbuf_bot_iw_I[11].z ;
 assign um_iw[282] = \block[15].zbuf_bot_iw_I[12].z ;
 assign um_iw[283] = \block[15].zbuf_bot_iw_I[13].z ;
 assign um_iw[284] = \block[15].zbuf_bot_iw_I[14].z ;
 assign um_iw[285] = \block[15].zbuf_bot_iw_I[15].z ;
 assign um_iw[286] = \block[15].zbuf_bot_iw_I[16].z ;
 assign um_iw[287] = \block[15].zbuf_bot_iw_I[17].z ;
 assign um_iw[271] = \block[15].zbuf_bot_iw_I[1].z ;
 assign um_iw[272] = \block[15].zbuf_bot_iw_I[2].z ;
 assign um_iw[273] = \block[15].zbuf_bot_iw_I[3].z ;
 assign um_iw[274] = \block[15].zbuf_bot_iw_I[4].z ;
 assign um_iw[275] = \block[15].zbuf_bot_iw_I[5].z ;
 assign um_iw[276] = \block[15].zbuf_bot_iw_I[6].z ;
 assign um_iw[277] = \block[15].zbuf_bot_iw_I[7].z ;
 assign um_iw[278] = \block[15].zbuf_bot_iw_I[8].z ;
 assign um_iw[279] = \block[15].zbuf_bot_iw_I[9].z ;
 assign um_ena[15] = \block[15].zbuf_ena_I.z ;
 assign um_pg_vdd[15] = \block[15].zbuf_pg_vdd_I.z ;
 assign um_k_zero[1] = \block[1].tie_I.lo ;
 assign um_iw[18] = \block[1].zbuf_bot_iw_I[0].z ;
 assign um_iw[28] = \block[1].zbuf_bot_iw_I[10].z ;
 assign um_iw[29] = \block[1].zbuf_bot_iw_I[11].z ;
 assign um_iw[30] = \block[1].zbuf_bot_iw_I[12].z ;
 assign um_iw[31] = \block[1].zbuf_bot_iw_I[13].z ;
 assign um_iw[32] = \block[1].zbuf_bot_iw_I[14].z ;
 assign um_iw[33] = \block[1].zbuf_bot_iw_I[15].z ;
 assign um_iw[34] = \block[1].zbuf_bot_iw_I[16].z ;
 assign um_iw[35] = \block[1].zbuf_bot_iw_I[17].z ;
 assign um_iw[19] = \block[1].zbuf_bot_iw_I[1].z ;
 assign um_iw[20] = \block[1].zbuf_bot_iw_I[2].z ;
 assign um_iw[21] = \block[1].zbuf_bot_iw_I[3].z ;
 assign um_iw[22] = \block[1].zbuf_bot_iw_I[4].z ;
 assign um_iw[23] = \block[1].zbuf_bot_iw_I[5].z ;
 assign um_iw[24] = \block[1].zbuf_bot_iw_I[6].z ;
 assign um_iw[25] = \block[1].zbuf_bot_iw_I[7].z ;
 assign um_iw[26] = \block[1].zbuf_bot_iw_I[8].z ;
 assign um_iw[27] = \block[1].zbuf_bot_iw_I[9].z ;
 assign um_ena[1] = \block[1].zbuf_ena_I.z ;
 assign um_pg_vdd[1] = \block[1].zbuf_pg_vdd_I.z ;
 assign um_k_zero[2] = \block[2].tie_I.lo ;
 assign um_iw[36] = \block[2].zbuf_bot_iw_I[0].z ;
 assign um_iw[46] = \block[2].zbuf_bot_iw_I[10].z ;
 assign um_iw[47] = \block[2].zbuf_bot_iw_I[11].z ;
 assign um_iw[48] = \block[2].zbuf_bot_iw_I[12].z ;
 assign um_iw[49] = \block[2].zbuf_bot_iw_I[13].z ;
 assign um_iw[50] = \block[2].zbuf_bot_iw_I[14].z ;
 assign um_iw[51] = \block[2].zbuf_bot_iw_I[15].z ;
 assign um_iw[52] = \block[2].zbuf_bot_iw_I[16].z ;
 assign um_iw[53] = \block[2].zbuf_bot_iw_I[17].z ;
 assign um_iw[37] = \block[2].zbuf_bot_iw_I[1].z ;
 assign um_iw[38] = \block[2].zbuf_bot_iw_I[2].z ;
 assign um_iw[39] = \block[2].zbuf_bot_iw_I[3].z ;
 assign um_iw[40] = \block[2].zbuf_bot_iw_I[4].z ;
 assign um_iw[41] = \block[2].zbuf_bot_iw_I[5].z ;
 assign um_iw[42] = \block[2].zbuf_bot_iw_I[6].z ;
 assign um_iw[43] = \block[2].zbuf_bot_iw_I[7].z ;
 assign um_iw[44] = \block[2].zbuf_bot_iw_I[8].z ;
 assign um_iw[45] = \block[2].zbuf_bot_iw_I[9].z ;
 assign um_ena[2] = \block[2].zbuf_ena_I.z ;
 assign um_pg_vdd[2] = \block[2].zbuf_pg_vdd_I.z ;
 assign um_k_zero[3] = \block[3].tie_I.lo ;
 assign um_iw[54] = \block[3].zbuf_bot_iw_I[0].z ;
 assign um_iw[64] = \block[3].zbuf_bot_iw_I[10].z ;
 assign um_iw[65] = \block[3].zbuf_bot_iw_I[11].z ;
 assign um_iw[66] = \block[3].zbuf_bot_iw_I[12].z ;
 assign um_iw[67] = \block[3].zbuf_bot_iw_I[13].z ;
 assign um_iw[68] = \block[3].zbuf_bot_iw_I[14].z ;
 assign um_iw[69] = \block[3].zbuf_bot_iw_I[15].z ;
 assign um_iw[70] = \block[3].zbuf_bot_iw_I[16].z ;
 assign um_iw[71] = \block[3].zbuf_bot_iw_I[17].z ;
 assign um_iw[55] = \block[3].zbuf_bot_iw_I[1].z ;
 assign um_iw[56] = \block[3].zbuf_bot_iw_I[2].z ;
 assign um_iw[57] = \block[3].zbuf_bot_iw_I[3].z ;
 assign um_iw[58] = \block[3].zbuf_bot_iw_I[4].z ;
 assign um_iw[59] = \block[3].zbuf_bot_iw_I[5].z ;
 assign um_iw[60] = \block[3].zbuf_bot_iw_I[6].z ;
 assign um_iw[61] = \block[3].zbuf_bot_iw_I[7].z ;
 assign um_iw[62] = \block[3].zbuf_bot_iw_I[8].z ;
 assign um_iw[63] = \block[3].zbuf_bot_iw_I[9].z ;
 assign um_ena[3] = \block[3].zbuf_ena_I.z ;
 assign um_pg_vdd[3] = \block[3].zbuf_pg_vdd_I.z ;
 assign um_k_zero[4] = \block[4].tie_I.lo ;
 assign um_iw[72] = \block[4].zbuf_bot_iw_I[0].z ;
 assign um_iw[82] = \block[4].zbuf_bot_iw_I[10].z ;
 assign um_iw[83] = \block[4].zbuf_bot_iw_I[11].z ;
 assign um_iw[84] = \block[4].zbuf_bot_iw_I[12].z ;
 assign um_iw[85] = \block[4].zbuf_bot_iw_I[13].z ;
 assign um_iw[86] = \block[4].zbuf_bot_iw_I[14].z ;
 assign um_iw[87] = \block[4].zbuf_bot_iw_I[15].z ;
 assign um_iw[88] = \block[4].zbuf_bot_iw_I[16].z ;
 assign um_iw[89] = \block[4].zbuf_bot_iw_I[17].z ;
 assign um_iw[73] = \block[4].zbuf_bot_iw_I[1].z ;
 assign um_iw[74] = \block[4].zbuf_bot_iw_I[2].z ;
 assign um_iw[75] = \block[4].zbuf_bot_iw_I[3].z ;
 assign um_iw[76] = \block[4].zbuf_bot_iw_I[4].z ;
 assign um_iw[77] = \block[4].zbuf_bot_iw_I[5].z ;
 assign um_iw[78] = \block[4].zbuf_bot_iw_I[6].z ;
 assign um_iw[79] = \block[4].zbuf_bot_iw_I[7].z ;
 assign um_iw[80] = \block[4].zbuf_bot_iw_I[8].z ;
 assign um_iw[81] = \block[4].zbuf_bot_iw_I[9].z ;
 assign um_ena[4] = \block[4].zbuf_ena_I.z ;
 assign um_pg_vdd[4] = \block[4].zbuf_pg_vdd_I.z ;
 assign um_k_zero[5] = \block[5].tie_I.lo ;
 assign um_iw[90] = \block[5].zbuf_bot_iw_I[0].z ;
 assign um_iw[100] = \block[5].zbuf_bot_iw_I[10].z ;
 assign um_iw[101] = \block[5].zbuf_bot_iw_I[11].z ;
 assign um_iw[102] = \block[5].zbuf_bot_iw_I[12].z ;
 assign um_iw[103] = \block[5].zbuf_bot_iw_I[13].z ;
 assign um_iw[104] = \block[5].zbuf_bot_iw_I[14].z ;
 assign um_iw[105] = \block[5].zbuf_bot_iw_I[15].z ;
 assign um_iw[106] = \block[5].zbuf_bot_iw_I[16].z ;
 assign um_iw[107] = \block[5].zbuf_bot_iw_I[17].z ;
 assign um_iw[91] = \block[5].zbuf_bot_iw_I[1].z ;
 assign um_iw[92] = \block[5].zbuf_bot_iw_I[2].z ;
 assign um_iw[93] = \block[5].zbuf_bot_iw_I[3].z ;
 assign um_iw[94] = \block[5].zbuf_bot_iw_I[4].z ;
 assign um_iw[95] = \block[5].zbuf_bot_iw_I[5].z ;
 assign um_iw[96] = \block[5].zbuf_bot_iw_I[6].z ;
 assign um_iw[97] = \block[5].zbuf_bot_iw_I[7].z ;
 assign um_iw[98] = \block[5].zbuf_bot_iw_I[8].z ;
 assign um_iw[99] = \block[5].zbuf_bot_iw_I[9].z ;
 assign um_ena[5] = \block[5].zbuf_ena_I.z ;
 assign um_pg_vdd[5] = \block[5].zbuf_pg_vdd_I.z ;
 assign um_k_zero[6] = \block[6].tie_I.lo ;
 assign um_iw[108] = \block[6].zbuf_bot_iw_I[0].z ;
 assign um_iw[118] = \block[6].zbuf_bot_iw_I[10].z ;
 assign um_iw[119] = \block[6].zbuf_bot_iw_I[11].z ;
 assign um_iw[120] = \block[6].zbuf_bot_iw_I[12].z ;
 assign um_iw[121] = \block[6].zbuf_bot_iw_I[13].z ;
 assign um_iw[122] = \block[6].zbuf_bot_iw_I[14].z ;
 assign um_iw[123] = \block[6].zbuf_bot_iw_I[15].z ;
 assign um_iw[124] = \block[6].zbuf_bot_iw_I[16].z ;
 assign um_iw[125] = \block[6].zbuf_bot_iw_I[17].z ;
 assign um_iw[109] = \block[6].zbuf_bot_iw_I[1].z ;
 assign um_iw[110] = \block[6].zbuf_bot_iw_I[2].z ;
 assign um_iw[111] = \block[6].zbuf_bot_iw_I[3].z ;
 assign um_iw[112] = \block[6].zbuf_bot_iw_I[4].z ;
 assign um_iw[113] = \block[6].zbuf_bot_iw_I[5].z ;
 assign um_iw[114] = \block[6].zbuf_bot_iw_I[6].z ;
 assign um_iw[115] = \block[6].zbuf_bot_iw_I[7].z ;
 assign um_iw[116] = \block[6].zbuf_bot_iw_I[8].z ;
 assign um_iw[117] = \block[6].zbuf_bot_iw_I[9].z ;
 assign um_ena[6] = \block[6].zbuf_ena_I.z ;
 assign um_pg_vdd[6] = \block[6].zbuf_pg_vdd_I.z ;
 assign um_k_zero[7] = \block[7].tie_I.lo ;
 assign um_iw[126] = \block[7].zbuf_bot_iw_I[0].z ;
 assign um_iw[136] = \block[7].zbuf_bot_iw_I[10].z ;
 assign um_iw[137] = \block[7].zbuf_bot_iw_I[11].z ;
 assign um_iw[138] = \block[7].zbuf_bot_iw_I[12].z ;
 assign um_iw[139] = \block[7].zbuf_bot_iw_I[13].z ;
 assign um_iw[140] = \block[7].zbuf_bot_iw_I[14].z ;
 assign um_iw[141] = \block[7].zbuf_bot_iw_I[15].z ;
 assign um_iw[142] = \block[7].zbuf_bot_iw_I[16].z ;
 assign um_iw[143] = \block[7].zbuf_bot_iw_I[17].z ;
 assign um_iw[127] = \block[7].zbuf_bot_iw_I[1].z ;
 assign um_iw[128] = \block[7].zbuf_bot_iw_I[2].z ;
 assign um_iw[129] = \block[7].zbuf_bot_iw_I[3].z ;
 assign um_iw[130] = \block[7].zbuf_bot_iw_I[4].z ;
 assign um_iw[131] = \block[7].zbuf_bot_iw_I[5].z ;
 assign um_iw[132] = \block[7].zbuf_bot_iw_I[6].z ;
 assign um_iw[133] = \block[7].zbuf_bot_iw_I[7].z ;
 assign um_iw[134] = \block[7].zbuf_bot_iw_I[8].z ;
 assign um_iw[135] = \block[7].zbuf_bot_iw_I[9].z ;
 assign um_ena[7] = \block[7].zbuf_ena_I.z ;
 assign um_pg_vdd[7] = \block[7].zbuf_pg_vdd_I.z ;
 assign um_k_zero[8] = \block[8].tie_I.lo ;
 assign um_iw[144] = \block[8].zbuf_bot_iw_I[0].z ;
 assign um_iw[154] = \block[8].zbuf_bot_iw_I[10].z ;
 assign um_iw[155] = \block[8].zbuf_bot_iw_I[11].z ;
 assign um_iw[156] = \block[8].zbuf_bot_iw_I[12].z ;
 assign um_iw[157] = \block[8].zbuf_bot_iw_I[13].z ;
 assign um_iw[158] = \block[8].zbuf_bot_iw_I[14].z ;
 assign um_iw[159] = \block[8].zbuf_bot_iw_I[15].z ;
 assign um_iw[160] = \block[8].zbuf_bot_iw_I[16].z ;
 assign um_iw[161] = \block[8].zbuf_bot_iw_I[17].z ;
 assign um_iw[145] = \block[8].zbuf_bot_iw_I[1].z ;
 assign um_iw[146] = \block[8].zbuf_bot_iw_I[2].z ;
 assign um_iw[147] = \block[8].zbuf_bot_iw_I[3].z ;
 assign um_iw[148] = \block[8].zbuf_bot_iw_I[4].z ;
 assign um_iw[149] = \block[8].zbuf_bot_iw_I[5].z ;
 assign um_iw[150] = \block[8].zbuf_bot_iw_I[6].z ;
 assign um_iw[151] = \block[8].zbuf_bot_iw_I[7].z ;
 assign um_iw[152] = \block[8].zbuf_bot_iw_I[8].z ;
 assign um_iw[153] = \block[8].zbuf_bot_iw_I[9].z ;
 assign um_ena[8] = \block[8].zbuf_ena_I.z ;
 assign um_pg_vdd[8] = \block[8].zbuf_pg_vdd_I.z ;
 assign um_k_zero[9] = \block[9].tie_I.lo ;
 assign um_iw[162] = \block[9].zbuf_bot_iw_I[0].z ;
 assign um_iw[172] = \block[9].zbuf_bot_iw_I[10].z ;
 assign um_iw[173] = \block[9].zbuf_bot_iw_I[11].z ;
 assign um_iw[174] = \block[9].zbuf_bot_iw_I[12].z ;
 assign um_iw[175] = \block[9].zbuf_bot_iw_I[13].z ;
 assign um_iw[176] = \block[9].zbuf_bot_iw_I[14].z ;
 assign um_iw[177] = \block[9].zbuf_bot_iw_I[15].z ;
 assign um_iw[178] = \block[9].zbuf_bot_iw_I[16].z ;
 assign um_iw[179] = \block[9].zbuf_bot_iw_I[17].z ;
 assign um_iw[163] = \block[9].zbuf_bot_iw_I[1].z ;
 assign um_iw[164] = \block[9].zbuf_bot_iw_I[2].z ;
 assign um_iw[165] = \block[9].zbuf_bot_iw_I[3].z ;
 assign um_iw[166] = \block[9].zbuf_bot_iw_I[4].z ;
 assign um_iw[167] = \block[9].zbuf_bot_iw_I[5].z ;
 assign um_iw[168] = \block[9].zbuf_bot_iw_I[6].z ;
 assign um_iw[169] = \block[9].zbuf_bot_iw_I[7].z ;
 assign um_iw[170] = \block[9].zbuf_bot_iw_I[8].z ;
 assign um_iw[171] = \block[9].zbuf_bot_iw_I[9].z ;
 assign um_ena[9] = \block[9].zbuf_ena_I.z ;
 assign um_pg_vdd[9] = \block[9].zbuf_pg_vdd_I.z ;
 assign spine_ow[1] = \tbuf_spine_ow_I[0].z ;
 assign spine_ow[11] = \tbuf_spine_ow_I[10].z ;
 assign spine_ow[12] = \tbuf_spine_ow_I[11].z ;
 assign spine_ow[13] = \tbuf_spine_ow_I[12].z ;
 assign spine_ow[14] = \tbuf_spine_ow_I[13].z ;
 assign spine_ow[15] = \tbuf_spine_ow_I[14].z ;
 assign spine_ow[16] = \tbuf_spine_ow_I[15].z ;
 assign spine_ow[17] = \tbuf_spine_ow_I[16].z ;
 assign spine_ow[18] = \tbuf_spine_ow_I[17].z ;
 assign spine_ow[19] = \tbuf_spine_ow_I[18].z ;
 assign spine_ow[20] = \tbuf_spine_ow_I[19].z ;
 assign spine_ow[2] = \tbuf_spine_ow_I[1].z ;
 assign spine_ow[21] = \tbuf_spine_ow_I[20].z ;
 assign spine_ow[22] = \tbuf_spine_ow_I[21].z ;
 assign spine_ow[23] = \tbuf_spine_ow_I[22].z ;
 assign spine_ow[24] = \tbuf_spine_ow_I[23].z ;
 assign spine_ow[3] = \tbuf_spine_ow_I[2].z ;
 assign spine_ow[4] = \tbuf_spine_ow_I[3].z ;
 assign spine_ow[5] = \tbuf_spine_ow_I[4].z ;
 assign spine_ow[6] = \tbuf_spine_ow_I[5].z ;
 assign spine_ow[7] = \tbuf_spine_ow_I[6].z ;
 assign spine_ow[8] = \tbuf_spine_ow_I[7].z ;
 assign spine_ow[9] = \tbuf_spine_ow_I[8].z ;
 assign spine_ow[10] = \tbuf_spine_ow_I[9].z ;
 assign spine_ow[0] = \tie_spine_guard_I[0].lo ;
 assign spine_ow[25] = \tie_spine_guard_I[1].lo ;
endmodule
